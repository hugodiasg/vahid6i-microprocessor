* NGSPICE file created from vahid6i.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

.subckt vahid6i D_R_data[0] D_R_data[10] D_R_data[11] D_R_data[12] D_R_data[13] D_R_data[14]
+ D_R_data[15] D_R_data[1] D_R_data[2] D_R_data[3] D_R_data[4] D_R_data[5] D_R_data[6]
+ D_R_data[7] D_R_data[8] D_R_data[9] D_W_data[0] D_W_data[10] D_W_data[11] D_W_data[12]
+ D_W_data[13] D_W_data[14] D_W_data[15] D_W_data[1] D_W_data[2] D_W_data[3] D_W_data[4]
+ D_W_data[5] D_W_data[6] D_W_data[7] D_W_data[8] D_W_data[9] D_addr[0] D_addr[1]
+ D_addr[2] D_addr[3] D_addr[4] D_addr[5] D_addr[6] D_addr[7] D_rd D_wr I_addr[0]
+ I_addr[10] I_addr[11] I_addr[12] I_addr[13] I_addr[14] I_addr[15] I_addr[1] I_addr[2]
+ I_addr[3] I_addr[4] I_addr[5] I_addr[6] I_addr[7] I_addr[8] I_addr[9] I_data[0]
+ I_data[10] I_data[11] I_data[12] I_data[13] I_data[14] I_data[15] I_data[1] I_data[2]
+ I_data[3] I_data[4] I_data[5] I_data[6] I_data[7] I_data[8] I_data[9] I_rd VGND
+ VPWR clock led_clock leds[0] leds[1] leds[2] leds[3] reset
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3155_ uc_0._20_\[9\] _0724_ _0562_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__mux2_1
X_3086_ po_0.regf_0.rf\[3\]\[13\] _0858_ _1331_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__mux2_1
X_2106_ po_0._1_\[8\] _0637_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__and2b_1
X_2037_ _0581_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__nor2_1
XFILLER_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2939_ _1171_ _1247_ _1250_ _1251_ _1252_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__a32o_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2724_ po_0.regf_0.rf\[10\]\[7\] _0944_ _1086_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__mux2_1
X_2655_ _1050_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
X_1606_ _1422_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__clkbuf_1
X_2586_ _1012_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
Xfanout127 net133 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout138 net139 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout105 net106 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
Xfanout116 net118 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xfanout149 net183 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
X_3207_ net126 _0031_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_3138_ po_0.regf_0.rq_addr\[1\] _0566_ _0563_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__mux2_1
XFILLER_15_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3069_ po_0.regf_0.rf\[3\]\[5\] _0772_ _1332_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__mux2_1
XFILLER_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2440_ po_0.regf_0.rf\[5\]\[14\] _0871_ _0908_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__mux2_1
X_2371_ po_0.regf_0.w_addr\[2\] VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2707_ po_0.regf_0.w_addr\[2\] _0882_ po_0.regf_0.w_wr _0885_ VGND VGND VPWR VPWR
+ _1078_ sky130_fd_sc_hd__and4b_2
X_2638_ _1040_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__buf_2
X_2569_ _1003_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1940_ _0423_ _0501_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__and2b_1
X_1871_ po_0.regf_0.rf\[8\]\[2\] po_0.regf_0.rf\[9\]\[2\] po_0.regf_0.rf\[10\]\[2\]
+ po_0.regf_0.rf\[11\]\[2\] _0411_ _0412_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__mux4_1
X_3541_ net180 _0325_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfxtp_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3472_ net168 _0256_ VGND VGND VPWR VPWR uc_0._00_ sky130_fd_sc_hd__dfxtp_1
X_2423_ _0908_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__buf_2
X_2354_ _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2285_ _0775_ po_0.alu_0._11_\[8\] _0706_ _0637_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__a22o_1
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2070_ _0612_ VGND VGND VPWR VPWR po_0.alu_0._10_\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2972_ uc_0._01_ _1139_ _1144_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__o21ba_1
X_1923_ po_0.regf_0.rf\[12\]\[7\] po_0.regf_0.rf\[13\]\[7\] po_0.regf_0.rf\[14\]\[7\]
+ po_0.regf_0.rf\[15\]\[7\] _0419_ _0420_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux4_1
X_1854_ _0422_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__buf_2
X_1785_ po_0.regf_0.rf\[0\]\[11\] po_0.regf_0.rf\[1\]\[11\] po_0.regf_0.rf\[2\]\[11\]
+ po_0.regf_0.rf\[3\]\[11\] _1488_ _1489_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__mux4_1
X_3524_ net160 _0308_ VGND VGND VPWR VPWR po_0.regf_0.rp_rd sky130_fd_sc_hd__dfxtp_1
X_3455_ net153 _0015_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__dfxtp_1
X_2406_ _0905_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
X_3386_ net157 _0174_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2337_ _0853_ _0675_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__nand2_1
X_2268_ net85 _0775_ _1401_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__or3_1
XFILLER_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2199_ _0711_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__clkbuf_2
XFILLER_52_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_5 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ po_0.regf_0._3_\[0\] net89 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlxtp_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _1391_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2122_ _0656_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__nor2_2
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2053_ _0587_ _0589_ _0585_ _0586_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__o211ai_1
X_2955_ _1237_ _1249_ _1256_ _1243_ net63 VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__a41oi_1
X_1906_ _0469_ _0470_ _0399_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__mux2_1
X_2886_ _1200_ _0566_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__or2_1
X_1837_ _0406_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__buf_2
X_1768_ po_0.regf_0.rf\[12\]\[9\] po_0.regf_0.rf\[13\]\[9\] po_0.regf_0.rf\[14\]\[9\]
+ po_0.regf_0.rf\[15\]\[9\] _1461_ _1463_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__mux4_1
X_3507_ net143 _0291_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1699_ _1502_ _1484_ _1485_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__a21bo_1
X_3438_ net167 _0226_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfxtp_2
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ net124 _0157_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput42 net42 VGND VGND VPWR VPWR D_W_data[1] sky130_fd_sc_hd__buf_2
Xoutput75 net75 VGND VGND VPWR VPWR I_addr[8] sky130_fd_sc_hd__clkbuf_4
Xoutput53 net53 VGND VGND VPWR VPWR D_addr[2] sky130_fd_sc_hd__buf_2
Xoutput64 net64 VGND VGND VPWR VPWR I_addr[12] sky130_fd_sc_hd__buf_2
XFILLER_0_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2740_ po_0.regf_0.rf\[10\]\[15\] _0960_ _1078_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__mux2_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2671_ _1058_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
X_1622_ _1431_ uc_0.bc_0._55_\[1\] uc_0.bc_0._55_\[0\] uc_0.bc_0._55_\[2\] uc_0.bc_0._55_\[3\]
+ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__a311oi_2
X_3223_ net126 _0047_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3154_ _1382_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__clkbuf_1
X_3085_ _1346_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__clkbuf_1
X_2105_ net50 po_0._1_\[9\] VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__xor2_2
XFILLER_54_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2036_ net86 po_0._1_\[1\] VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__nor2_1
XFILLER_35_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2938_ _1241_ net97 _1226_ _1246_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__a31o_1
XFILLER_10_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2869_ _1185_ _0557_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__nor2_1
XFILLER_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2723_ _1087_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
X_2654_ po_0.regf_0.rf\[12\]\[7\] _0944_ _1048_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__mux2_1
X_2585_ _0811_ po_0.regf_0.rf\[14\]\[8\] _1009_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__mux2_1
X_1605_ _1414_ _1416_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__or2b_1
Xfanout128 net132 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout106 net107 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout117 net118 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_1
Xfanout139 net149 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3206_ net109 _0030_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_3137_ _1373_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3068_ _1337_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2019_ po_0.muxf_0.rf_w_data\[7\] VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2370_ _0883_ _0884_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__and2b_1
XFILLER_68_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2706_ _1077_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_1
X_2637_ _0718_ _0715_ _0716_ _1039_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__and4_2
X_2568_ _0714_ po_0.regf_0.rf\[14\]\[0\] _1002_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__mux2_1
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2499_ po_0.regf_0.rf\[1\]\[1\] _0931_ _0963_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__mux2_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1870_ _0425_ _0427_ _0433_ _0438_ VGND VGND VPWR VPWR po_0.regf_0._3_\[1\] sky130_fd_sc_hd__o22a_1
X_3540_ net179 _0324_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfxtp_1
X_3471_ net168 _0255_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_2
X_2422_ _0915_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2353_ net6 _0701_ _0869_ _0793_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__a22o_2
XFILLER_69_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2284_ _0805_ _0668_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__nand2_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1999_ _0403_ _0553_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__and2b_1
XFILLER_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2971_ net65 _1215_ _1280_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__o21ba_1
X_1922_ _0417_ _0484_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__and2b_1
X_1853_ _0002_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__clkbuf_2
X_1784_ _0358_ _1550_ _1485_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__a21bo_1
X_3523_ net166 _0307_ VGND VGND VPWR VPWR po_0.regf_0.rq_rd sky130_fd_sc_hd__dfxtp_1
X_3454_ net153 _0014_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__dfxtp_1
X_2405_ po_0.regf_0.rf\[6\]\[15\] _0880_ _0887_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__mux2_1
X_3385_ net157 _0173_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2336_ _0675_ _0853_ _0758_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__o21a_1
XFILLER_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2267_ _0786_ _0789_ _0758_ _0790_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__a31o_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2198_ _1405_ po_0.alu_0._11_\[1\] _0705_ net86 _0727_ VGND VGND VPWR VPWR _0728_
+ sky130_fd_sc_hd__a221o_1
XFILLER_4_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_6 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3170_ _0704_ net51 _1389_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__mux2_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2121_ net84 po_0._1_\[11\] VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__and2_1
XFILLER_66_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2052_ po_0._1_\[2\] _0588_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__or2b_1
XFILLER_66_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2954_ _1262_ _1265_ _1145_ _1207_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__a31o_1
X_1905_ po_0.regf_0.rf\[4\]\[5\] po_0.regf_0.rf\[5\]\[5\] po_0.regf_0.rf\[6\]\[5\]
+ po_0.regf_0.rf\[7\]\[5\] _0404_ _0406_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__mux4_1
X_2885_ net72 po_0.muxf_0.rf_w_data\[5\] VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__nand2_1
X_1836_ _0001_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__buf_2
X_1767_ _1511_ _0343_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__and2b_1
X_3506_ net144 _0290_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1698_ po_0.regf_0.rf\[12\]\[2\] po_0.regf_0.rf\[13\]\[2\] po_0.regf_0.rf\[14\]\[2\]
+ po_0.regf_0.rf\[15\]\[2\] _1481_ _1482_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__mux4_1
X_3437_ net167 _0225_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfxtp_2
X_3368_ net129 _0156_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _0838_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3299_ net123 _0087_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput43 net43 VGND VGND VPWR VPWR D_W_data[2] sky130_fd_sc_hd__buf_2
Xoutput76 net76 VGND VGND VPWR VPWR I_addr[9] sky130_fd_sc_hd__buf_2
Xoutput65 net65 VGND VGND VPWR VPWR I_addr[13] sky130_fd_sc_hd__buf_2
Xoutput54 net54 VGND VGND VPWR VPWR D_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2670_ po_0.regf_0.rf\[12\]\[15\] _0960_ _1040_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__mux2_1
X_1621_ net82 net81 net80 VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__or3b_1
X_3222_ net109 _0046_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3153_ _0883_ _1381_ _1372_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__mux2_1
X_2104_ _0640_ _0642_ VGND VGND VPWR VPWR po_0.alu_0._10_\[8\] sky130_fd_sc_hd__xor2_1
X_3084_ po_0.regf_0.rf\[3\]\[12\] _0848_ _1331_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__mux2_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2035_ net86 po_0._1_\[1\] VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__and2_1
XFILLER_35_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2937_ _1248_ _1246_ _1242_ _1144_ _1139_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__a311oi_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2868_ _1186_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__clkbuf_2
X_1819_ _1453_ _0389_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__and2b_1
X_2799_ _1128_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__clkbuf_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2722_ po_0.regf_0.rf\[10\]\[6\] _0941_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__mux2_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2653_ _1049_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
X_2584_ _1011_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
X_1604_ _1421_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__clkbuf_1
Xfanout129 net132 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
Xfanout107 net115 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
Xfanout118 net121 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
X_3205_ net113 _0029_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3136_ po_0.regf_0.rq_addr\[0\] _0557_ _0563_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__mux2_1
X_3067_ po_0.regf_0.rf\[3\]\[4\] _0762_ _1332_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__mux2_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2018_ _0569_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2705_ po_0.regf_0.rf\[11\]\[15\] _0960_ _1059_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__mux2_1
X_2636_ _0884_ _0883_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__nor2_1
X_2567_ _1001_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__buf_2
X_2498_ _0964_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3119_ po_0.regf_0.rf\[2\]\[12\] _0848_ _1350_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__mux2_1
XFILLER_82_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3470_ net151 _0254_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfxtp_2
X_2421_ po_0.regf_0.rf\[5\]\[5\] _0773_ _0909_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__mux2_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2352_ _0866_ _0867_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__o21ai_1
X_2283_ _0638_ _0639_ _0805_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__a21o_1
XFILLER_56_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1998_ po_0.regf_0.rf\[0\]\[15\] po_0.regf_0.rf\[1\]\[15\] po_0.regf_0.rf\[2\]\[15\]
+ po_0.regf_0.rf\[3\]\[15\] _0405_ _0407_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__mux4_1
X_2619_ _1030_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2970_ _1275_ _1186_ _1276_ _1279_ _1214_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__o311a_1
X_1921_ po_0.regf_0.rf\[8\]\[7\] po_0.regf_0.rf\[9\]\[7\] po_0.regf_0.rf\[10\]\[7\]
+ po_0.regf_0.rf\[11\]\[7\] _0411_ _0412_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__mux4_1
XFILLER_61_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1852_ po_0.regf_0.rf\[4\]\[1\] po_0.regf_0.rf\[5\]\[1\] po_0.regf_0.rf\[6\]\[1\]
+ po_0.regf_0.rf\[7\]\[1\] _0419_ _0420_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux4_1
X_1783_ po_0.regf_0.rf\[12\]\[11\] po_0.regf_0.rf\[13\]\[11\] po_0.regf_0.rf\[14\]\[11\]
+ po_0.regf_0.rf\[15\]\[11\] _1542_ _1543_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__mux4_1
X_3522_ net180 _0306_ VGND VGND VPWR VPWR po_0.alu_0.s0 sky130_fd_sc_hd__dfxtp_1
X_3453_ net153 _0013_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__dfxtp_1
X_2404_ _0904_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
X_3384_ net170 _0172_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2335_ _0664_ _0844_ _0852_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2266_ _0775_ po_0.alu_0._11_\[7\] _0706_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__a21o_1
X_2197_ _1429_ _0581_ _0582_ _0725_ _0726_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__o311a_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_7 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2120_ net84 po_0._1_\[11\] VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__nor2_1
X_2051_ _0595_ VGND VGND VPWR VPWR po_0.alu_0._10_\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2953_ _1234_ _1264_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__nand2_1
X_1904_ po_0.regf_0.rf\[0\]\[5\] po_0.regf_0.rf\[1\]\[5\] po_0.regf_0.rf\[2\]\[5\]
+ po_0.regf_0.rf\[3\]\[5\] _0404_ _0406_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__mux4_1
XFILLER_30_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2884_ _1189_ _1190_ _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__o21ai_1
X_1835_ _0404_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__clkbuf_4
X_1766_ po_0.regf_0.rf\[0\]\[9\] po_0.regf_0.rf\[1\]\[9\] po_0.regf_0.rf\[2\]\[9\]
+ po_0.regf_0.rf\[3\]\[9\] _1512_ _1513_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__mux4_1
X_3505_ net147 _0289_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1697_ _1486_ _1491_ _1493_ _1501_ VGND VGND VPWR VPWR po_0.regf_0._5_\[1\] sky130_fd_sc_hd__o22a_1
X_3436_ net167 _0224_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfxtp_2
X_3367_ net106 _0155_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2318_ _0722_ _0723_ net3 _0836_ _0837_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__a32o_4
X_3298_ net122 _0086_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2249_ _0774_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput66 net96 VGND VGND VPWR VPWR I_addr[14] sky130_fd_sc_hd__clkbuf_4
Xoutput44 net44 VGND VGND VPWR VPWR D_W_data[3] sky130_fd_sc_hd__clkbuf_4
Xoutput55 net55 VGND VGND VPWR VPWR D_addr[4] sky130_fd_sc_hd__buf_2
Xoutput77 net77 VGND VGND VPWR VPWR I_rd sky130_fd_sc_hd__buf_2
XFILLER_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1620_ _1430_ VGND VGND VPWR VPWR po_0.alu_0._10_\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3221_ net109 _0045_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3152_ uc_0._20_\[8\] _0704_ _0563_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__mux2_1
X_2103_ _0634_ _0641_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__nand2_1
X_3083_ _1345_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__clkbuf_1
X_2034_ net87 po_0._1_\[0\] VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__and2b_1
XFILLER_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2936_ _1248_ _1249_ _1234_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__nand3_1
XFILLER_50_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2867_ _1146_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__clkbuf_2
XFILLER_30_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1818_ po_0.regf_0.rf\[8\]\[15\] po_0.regf_0.rf\[9\]\[15\] po_0.regf_0.rf\[10\]\[15\]
+ po_0.regf_0.rf\[11\]\[15\] _1455_ _1457_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__mux4_1
X_2798_ po_0.regf_0.rf\[8\]\[9\] _0819_ _1124_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__mux2_1
X_1749_ po_0.regf_0.rf\[12\]\[7\] po_0.regf_0.rf\[13\]\[7\] po_0.regf_0.rf\[14\]\[7\]
+ po_0.regf_0.rf\[15\]\[7\] _1475_ _1476_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__mux4_1
X_3419_ net128 _0207_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2721_ _1078_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__buf_2
X_2652_ po_0.regf_0.rf\[12\]\[6\] _0941_ _1048_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__mux2_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2583_ _0796_ po_0.regf_0.rf\[14\]\[7\] _1009_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__mux2_1
X_1603_ _1414_ _1416_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__or2b_1
Xfanout108 net111 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout119 net121 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlymetal6s2s_1
X_3204_ net109 _0028_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3135_ _0716_ _1311_ _1372_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__a21o_1
X_3066_ _1336_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__clkbuf_1
X_2017_ po_0.regf_0.rq_addr\[2\] _0568_ _0564_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__mux2_1
XFILLER_82_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2919_ _1232_ _1234_ _1171_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__or3b_1
XFILLER_5_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2704_ _1076_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__clkbuf_1
X_2635_ _1038_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
X_2566_ _0883_ _1000_ _0884_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__or3b_4
X_2497_ po_0.regf_0.rf\[1\]\[0\] _0927_ _0963_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__mux2_1
X_3118_ _1364_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3049_ po_0.regf_0.rf\[4\]\[12\] _0848_ _1312_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__mux2_1
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout90 net91 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dlymetal6s2s_1
X_2420_ _0914_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
X_2351_ _0745_ po_0.alu_0._11_\[14\] _0815_ _0680_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__a22oi_1
X_2282_ _0600_ _0799_ _0800_ _0804_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__o31ai_4
XFILLER_69_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1997_ _0551_ _0434_ _0401_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__a21bo_1
X_2618_ _0796_ po_0.regf_0.rf\[13\]\[7\] _1028_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__mux2_1
X_2549_ po_0.regf_0.rf\[15\]\[8\] _0946_ _0989_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__mux2_1
XFILLER_85_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1920_ _0477_ _0479_ _0481_ _0483_ VGND VGND VPWR VPWR po_0.regf_0._3_\[6\] sky130_fd_sc_hd__o22a_1
X_1851_ _0396_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__clkbuf_4
X_1782_ _1500_ _0356_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__and2b_1
X_3521_ net179 _0305_ VGND VGND VPWR VPWR po_0.alu_0.s1 sky130_fd_sc_hd__dfxtp_1
X_3452_ net166 _0012_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__dfxtp_1
X_2403_ po_0.regf_0.rf\[6\]\[14\] _0871_ _0887_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__mux2_1
X_3383_ net120 _0171_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_2334_ net38 po_0._1_\[12\] VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__nand2_1
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2265_ _0622_ _0788_ _0633_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__o21ai_1
X_2196_ _0581_ _0582_ po_0._1_\[0\] net87 VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_8 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2050_ _0591_ _0594_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__or2b_1
XFILLER_47_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2952_ _1263_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__clkbuf_2
X_1903_ _0462_ _0464_ _0466_ _0468_ VGND VGND VPWR VPWR po_0.regf_0._3_\[4\] sky130_fd_sc_hd__o22a_1
X_2883_ net70 po_0.muxf_0.rf_w_data\[3\] net71 po_0.muxf_0.rf_w_data\[4\] _1192_ VGND
+ VGND VPWR VPWR _1201_ sky130_fd_sc_hd__o221ai_4
X_1834_ _0000_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__clkbuf_4
X_1765_ _0341_ _1484_ _1492_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__a21o_1
X_3504_ net140 _0288_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_1696_ _1496_ _1499_ _1500_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__mux2_1
X_3435_ net172 _0223_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_3366_ net116 _0154_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ net144 _0085_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2317_ net84 _1406_ _1402_ _0729_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__o31a_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _0773_ po_0.regf_0.rf\[7\]\[5\] _0720_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__mux2_1
X_2179_ net87 _1404_ _1401_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__or3_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput56 net56 VGND VGND VPWR VPWR D_addr[5] sky130_fd_sc_hd__buf_2
Xoutput45 net45 VGND VGND VPWR VPWR D_W_data[4] sky130_fd_sc_hd__buf_2
Xoutput67 net67 VGND VGND VPWR VPWR I_addr[15] sky130_fd_sc_hd__buf_2
Xoutput78 net78 VGND VGND VPWR VPWR led_clock sky130_fd_sc_hd__clkbuf_4
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3220_ net109 _0044_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3151_ _1380_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2102_ po_0._1_\[7\] net85 VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__or2b_1
XFILLER_82_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3082_ po_0.regf_0.rf\[3\]\[11\] _0838_ _1339_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__mux2_1
XFILLER_54_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2033_ _0579_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2935_ _1246_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__clkbuf_2
X_2866_ net71 VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1817_ _0387_ _1470_ _1467_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a21bo_1
X_2797_ _1127_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__clkbuf_1
X_1748_ _1511_ _1546_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__and2b_1
X_1679_ _1452_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__buf_2
X_3418_ net128 _0206_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_3349_ net103 _0137_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2720_ _1085_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2651_ _1040_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__buf_2
X_1602_ _1420_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__clkbuf_1
X_2582_ _1010_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout109 net111 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlymetal6s2s_1
X_3203_ net100 _0027_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3134_ uc_0.bc_0._54_\[0\] _1369_ _1370_ _1371_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__o211ai_4
XFILLER_82_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3065_ po_0.regf_0.rf\[3\]\[3\] _0752_ _1332_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__mux2_1
X_2016_ po_0.muxf_0.rf_w_data\[6\] VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__clkbuf_2
XFILLER_23_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2918_ _1233_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__clkbuf_2
X_2849_ _1169_ _1161_ _1148_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__mux2_1
XFILLER_2_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2703_ po_0.regf_0.rf\[11\]\[14\] _0958_ _1059_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__mux2_1
X_2634_ _0880_ po_0.regf_0.rf\[13\]\[15\] _1020_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__mux2_1
X_2565_ po_0.regf_0.w_addr\[2\] po_0.regf_0.w_addr\[3\] po_0.regf_0.w_wr VGND VGND
+ VPWR VPWR _1000_ sky130_fd_sc_hd__nand3_1
X_2496_ _0962_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__buf_2
XFILLER_67_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3117_ po_0.regf_0.rf\[2\]\[11\] _0838_ _1358_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__mux2_1
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3048_ _1326_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout91 po_0.regf_0.rp_rd VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
X_2350_ _0865_ _0863_ _0864_ _0708_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__a31o_1
X_2281_ _0801_ _0803_ _0632_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__a21oi_2
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1996_ po_0.regf_0.rf\[12\]\[15\] po_0.regf_0.rf\[13\]\[15\] po_0.regf_0.rf\[14\]\[15\]
+ po_0.regf_0.rf\[15\]\[15\] _0419_ _0420_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__mux4_1
X_2617_ _1029_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
X_2548_ _0991_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
X_2479_ _0951_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1850_ _0394_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__clkbuf_4
X_1781_ po_0.regf_0.rf\[8\]\[11\] po_0.regf_0.rf\[9\]\[11\] po_0.regf_0.rf\[10\]\[11\]
+ po_0.regf_0.rf\[11\]\[11\] _1494_ _1495_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux4_1
X_3520_ net140 _0304_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_3451_ net166 _0239_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfxtp_2
X_2402_ _0903_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3382_ net150 _0170_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_2333_ _0683_ _0815_ _0703_ _0700_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__a211o_1
XFILLER_69_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2264_ _0757_ _0777_ _0614_ _0787_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__a211oi_1
X_2195_ po_0.alu_0.s1 po_0.alu_0.s0 VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__and2b_1
XFILLER_65_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1979_ po_0.regf_0.rf\[0\]\[13\] po_0.regf_0.rf\[1\]\[13\] po_0.regf_0.rf\[2\]\[13\]
+ po_0.regf_0.rf\[3\]\[13\] _0495_ _0496_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__mux4_1
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2951_ net97 net76 net62 net63 VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__and4_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1902_ _0434_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__and2b_1
XFILLER_30_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2882_ net72 VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__clkbuf_2
X_1833_ _0399_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__clkbuf_2
X_1764_ po_0.regf_0.rf\[4\]\[9\] po_0.regf_0.rf\[5\]\[9\] po_0.regf_0.rf\[6\]\[9\]
+ po_0.regf_0.rf\[7\]\[9\] _1542_ _1543_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__mux4_1
X_3503_ net114 _0287_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_1695_ _1452_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__buf_2
X_3434_ net161 _0222_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_3365_ net116 _0153_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ net146 _0084_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2316_ _0832_ _0758_ _0834_ _0835_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__a31o_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _0772_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2178_ po_0.alu_0._10_\[0\] po_0.alu_0._11_\[0\] _0708_ VGND VGND VPWR VPWR _0709_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput35 net35 VGND VGND VPWR VPWR D_W_data[0] sky130_fd_sc_hd__buf_2
Xoutput46 net46 VGND VGND VPWR VPWR D_W_data[5] sky130_fd_sc_hd__clkbuf_4
Xoutput57 net57 VGND VGND VPWR VPWR D_addr[6] sky130_fd_sc_hd__buf_2
Xoutput79 net79 VGND VGND VPWR VPWR leds[0] sky130_fd_sc_hd__clkbuf_4
Xoutput68 net68 VGND VGND VPWR VPWR I_addr[1] sky130_fd_sc_hd__buf_2
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3150_ uc_0._20_\[11\] po_0.regf_0.rp_addr\[3\] _0574_ VGND VGND VPWR VPWR _1380_
+ sky130_fd_sc_hd__mux2_1
X_3081_ _1344_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__clkbuf_1
X_2101_ _0638_ _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__nand2_1
X_2032_ uc_0._20_\[11\] po_0.regf_0.rp_addr\[3\] _0575_ VGND VGND VPWR VPWR _0579_
+ sky130_fd_sc_hd__mux2_1
X_2934_ net97 VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__clkbuf_2
X_2865_ _1184_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__clkbuf_1
X_1816_ po_0.regf_0.rf\[12\]\[15\] po_0.regf_0.rf\[13\]\[15\] po_0.regf_0.rf\[14\]\[15\]
+ po_0.regf_0.rf\[15\]\[15\] _1471_ _1472_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__mux4_1
X_2796_ po_0.regf_0.rf\[8\]\[8\] _0810_ _1124_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__mux2_1
X_1747_ po_0.regf_0.rf\[0\]\[7\] po_0.regf_0.rf\[1\]\[7\] po_0.regf_0.rf\[2\]\[7\]
+ po_0.regf_0.rf\[3\]\[7\] _1512_ _1513_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__mux4_1
X_1678_ po_0.regf_0.rf\[12\]\[1\] po_0.regf_0.rf\[13\]\[1\] po_0.regf_0.rf\[14\]\[1\]
+ po_0.regf_0.rf\[15\]\[1\] _1481_ _1482_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__mux4_1
X_3417_ net113 _0205_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3348_ net104 _0136_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3279_ net171 _0067_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2650_ _1047_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
X_1601_ _1414_ _1416_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__or2b_1
X_2581_ _0783_ po_0.regf_0.rf\[14\]\[6\] _1009_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__mux2_1
X_3202_ net100 _0026_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_3133_ _0558_ _0561_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__and2_1
XFILLER_82_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3064_ _1335_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__clkbuf_1
X_2015_ _0567_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2917_ net98 net74 _1208_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__and3_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2848_ _1164_ _1141_ _1165_ _1168_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__a31o_1
X_2779_ po_0.regf_0.rf\[8\]\[0\] _0713_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__mux2_1
XFILLER_85_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2702_ _1075_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2633_ _1037_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
X_2564_ _0999_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
X_2495_ _0718_ po_0.regf_0.w_addr\[3\] _0906_ _0907_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__and4bb_2
XFILLER_59_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3116_ _1363_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3047_ po_0.regf_0.rf\[4\]\[11\] _0838_ _1320_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__mux2_1
XFILLER_82_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout92 net93 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2280_ _0614_ _0623_ _0777_ _0802_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__o31ai_1
XFILLER_49_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1995_ _0417_ _0549_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__and2b_1
X_2616_ _0783_ po_0.regf_0.rf\[13\]\[6\] _1028_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__mux2_1
X_2547_ po_0.regf_0.rf\[15\]\[7\] _0944_ _0989_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__mux2_1
X_2478_ po_0.regf_0.rf\[9\]\[10\] _0950_ _0942_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__mux2_1
XFILLER_28_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1780_ _0350_ _0352_ _1493_ _0355_ VGND VGND VPWR VPWR po_0.regf_0._5_\[10\] sky130_fd_sc_hd__o22a_1
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3450_ net166 _0238_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfxtp_1
X_2401_ po_0.regf_0.rf\[6\]\[13\] _0859_ _0887_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__mux2_1
X_3381_ net150 _0169_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_2332_ _0850_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2263_ _0622_ _0623_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__or2_1
X_2194_ po_0.muxf_0.rf_w_data\[1\] VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__buf_2
XFILLER_37_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1978_ _0534_ _0400_ _0432_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__a21o_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2950_ _1248_ _1249_ _1256_ _1234_ net63 VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__a41o_1
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2881_ _1135_ _1185_ _1187_ _1199_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__o31a_1
X_1901_ po_0.regf_0.rf\[8\]\[4\] po_0.regf_0.rf\[9\]\[4\] po_0.regf_0.rf\[10\]\[4\]
+ po_0.regf_0.rf\[11\]\[4\] _0435_ _0436_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux4_1
X_1832_ _0398_ _0400_ _0401_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__a21bo_1
X_1763_ _1554_ _1556_ _0338_ _0340_ VGND VGND VPWR VPWR po_0.regf_0._5_\[8\] sky130_fd_sc_hd__o22a_1
X_1694_ po_0.regf_0.rf\[4\]\[1\] po_0.regf_0.rf\[5\]\[1\] po_0.regf_0.rf\[6\]\[1\]
+ po_0.regf_0.rf\[7\]\[1\] _1497_ _1498_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__mux4_1
X_3502_ net124 _0286_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3433_ net157 _0221_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ net104 _0152_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ net142 _0083_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2315_ _0775_ po_0.alu_0._11_\[11\] _0706_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__a21o_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ net12 _0700_ _0703_ _0566_ _0771_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__a221o_4
XFILLER_38_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2177_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__buf_2
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput36 net36 VGND VGND VPWR VPWR D_W_data[10] sky130_fd_sc_hd__clkbuf_4
Xoutput58 net58 VGND VGND VPWR VPWR D_addr[7] sky130_fd_sc_hd__buf_2
Xoutput47 net47 VGND VGND VPWR VPWR D_W_data[6] sky130_fd_sc_hd__buf_2
Xoutput69 net69 VGND VGND VPWR VPWR I_addr[2] sky130_fd_sc_hd__buf_2
XFILLER_56_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3080_ po_0.regf_0.rf\[3\]\[10\] _0829_ _1339_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__mux2_1
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2100_ _0637_ po_0._1_\[8\] VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__or2_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2031_ _0578_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2933_ net73 _1225_ net97 _1209_ _1246_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__a41o_1
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2864_ _1183_ _1172_ _1148_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__mux2_1
X_1815_ _0381_ _0383_ _1493_ _0386_ VGND VGND VPWR VPWR po_0.regf_0._5_\[14\] sky130_fd_sc_hd__o22a_1
X_2795_ _1126_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__clkbuf_1
X_1746_ _1544_ _1484_ _1492_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__a21o_1
X_1677_ _1456_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__buf_2
X_3416_ net141 _0204_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3347_ net112 _0135_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ net173 _0066_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2229_ _0598_ po_0._1_\[3\] _0755_ _0746_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__o22a_1
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1600_ _1419_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__clkbuf_1
X_2580_ _1001_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__buf_2
XFILLER_4_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3201_ net102 _0025_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_3132_ _1441_ _0559_ _1451_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__or3_2
XFILLER_82_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3063_ po_0.regf_0.rf\[3\]\[2\] _0741_ _1332_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__mux2_1
XFILLER_82_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2014_ po_0.regf_0.rq_addr\[1\] _0566_ _0564_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__mux2_1
XFILLER_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2916_ _1213_ _1209_ _1225_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__a21oi_1
X_2847_ _1166_ _1167_ _1140_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__and3b_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2778_ _1116_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__buf_2
X_1729_ _1529_ _1466_ _1468_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__a21bo_1
XFILLER_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2701_ po_0.regf_0.rf\[11\]\[13\] _0956_ _1059_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__mux2_1
X_2632_ _0871_ po_0.regf_0.rf\[13\]\[14\] _1020_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2563_ po_0.regf_0.rf\[15\]\[15\] _0960_ _0981_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__mux2_1
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2494_ _0961_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3115_ po_0.regf_0.rf\[2\]\[10\] _0829_ _1358_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__mux2_1
XFILLER_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3046_ _1325_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout93 net95 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1994_ po_0.regf_0.rf\[8\]\[15\] po_0.regf_0.rf\[9\]\[15\] po_0.regf_0.rf\[10\]\[15\]
+ po_0.regf_0.rf\[11\]\[15\] _0411_ _0412_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__mux4_1
X_2615_ _1020_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__buf_2
X_2546_ _0990_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
X_2477_ _0829_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__clkbuf_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3029_ _1316_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2400_ _0902_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
X_3380_ net119 _0168_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_2331_ _0849_ po_0.regf_0.rf\[7\]\[12\] _0719_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__mux2_1
X_2262_ _0620_ _0621_ _0778_ _0628_ _0633_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__a221o_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2193_ _0698_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__clkbuf_2
XFILLER_37_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1977_ po_0.regf_0.rf\[4\]\[13\] po_0.regf_0.rf\[5\]\[13\] po_0.regf_0.rf\[6\]\[13\]
+ po_0.regf_0.rf\[7\]\[13\] _0395_ _0397_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__mux4_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2529_ _0980_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2880_ _1194_ _1142_ _1195_ _1198_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__a31o_1
X_1900_ _0465_ _0431_ _0432_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__a21bo_1
X_1831_ _0003_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__clkbuf_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1762_ _1550_ _0339_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__and2b_1
X_1693_ _0005_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__buf_2
X_3501_ net123 _0285_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3432_ net172 _0220_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3363_ net114 _0151_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ net141 _0082_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2314_ _0833_ _0824_ _0658_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__o21ai_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2245_ _0613_ _0745_ _1401_ _0711_ _0770_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__o311a_1
X_2176_ _1404_ po_0.alu_0.s0 VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__or2b_1
XFILLER_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput37 net37 VGND VGND VPWR VPWR D_W_data[11] sky130_fd_sc_hd__buf_2
Xoutput48 net85 VGND VGND VPWR VPWR D_W_data[7] sky130_fd_sc_hd__buf_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput59 net59 VGND VGND VPWR VPWR D_rd sky130_fd_sc_hd__buf_2
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2030_ uc_0._20_\[10\] po_0.regf_0.rp_addr\[2\] _0575_ VGND VGND VPWR VPWR _0578_
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2932_ net76 VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__clkbuf_2
X_2863_ _1171_ _1173_ _1174_ _1182_ _1142_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__a32o_1
X_1814_ _0384_ _0385_ _1465_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__mux2_1
X_2794_ po_0.regf_0.rf\[8\]\[7\] _0795_ _1124_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__mux2_1
X_1745_ po_0.regf_0.rf\[4\]\[7\] po_0.regf_0.rf\[5\]\[7\] po_0.regf_0.rf\[6\]\[7\]
+ po_0.regf_0.rf\[7\]\[7\] _1542_ _1543_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__mux4_1
X_1676_ _1454_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__clkbuf_4
X_3415_ net105 _0203_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_3346_ net112 _0134_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ net174 _0065_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2228_ _0588_ po_0._1_\[2\] po_0._1_\[3\] net44 VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__a22o_1
X_2159_ _0689_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__nor2_1
XFILLER_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3200_ net102 _0024_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3131_ _1440_ _1432_ _1439_ _1451_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__or4_2
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3062_ _1334_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__clkbuf_1
X_2013_ po_0.muxf_0.rf_w_data\[5\] VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__buf_2
XFILLER_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2915_ _1229_ _1226_ _1227_ _1186_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__a31o_1
X_2846_ _1136_ _1151_ _1161_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__a21o_1
X_2777_ po_0.regf_0.w_addr\[2\] _0882_ po_0.regf_0.w_wr _1039_ VGND VGND VPWR VPWR
+ _1116_ sky130_fd_sc_hd__and4b_2
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1728_ po_0.regf_0.rf\[12\]\[5\] po_0.regf_0.rf\[13\]\[5\] po_0.regf_0.rf\[14\]\[5\]
+ po_0.regf_0.rf\[15\]\[5\] _1461_ _1463_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__mux4_1
X_1659_ _0006_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__buf_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ net137 _0117_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2700_ _1074_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__clkbuf_1
X_2631_ _1036_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
X_2562_ _0998_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2493_ po_0.regf_0.rf\[9\]\[15\] _0960_ _0928_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__mux2_1
XFILLER_4_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3114_ _1362_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__clkbuf_1
X_3045_ po_0.regf_0.rf\[4\]\[10\] _0829_ _1320_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__mux2_1
XFILLER_55_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2829_ net68 VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__clkbuf_2
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout83 net38 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout94 net95 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1993_ _0543_ _0545_ _0410_ _0548_ VGND VGND VPWR VPWR po_0.regf_0._3_\[14\] sky130_fd_sc_hd__o22a_1
X_2614_ _1027_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
X_2545_ po_0.regf_0.rf\[15\]\[6\] _0941_ _0989_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__mux2_1
X_2476_ _0949_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3028_ po_0.regf_0.rf\[4\]\[2\] _0741_ _1313_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__mux2_1
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2330_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__clkbuf_2
XFILLER_69_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2261_ _0785_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
X_2192_ po_0.muxf_0.s0 VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__clkbuf_2
XFILLER_65_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1976_ _0527_ _0529_ _0531_ _0533_ VGND VGND VPWR VPWR po_0.regf_0._3_\[12\] sky130_fd_sc_hd__o22a_1
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2528_ po_0.regf_0.rf\[1\]\[15\] _0960_ _0962_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2459_ po_0.regf_0.rf\[9\]\[4\] _0937_ _0929_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__mux2_1
XFILLER_56_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1830_ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__buf_2
X_3500_ net120 _0284_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_1761_ po_0.regf_0.rf\[8\]\[8\] po_0.regf_0.rf\[9\]\[8\] po_0.regf_0.rf\[10\]\[8\]
+ po_0.regf_0.rf\[11\]\[8\] _1471_ _1472_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__mux4_1
X_1692_ _0004_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__clkbuf_4
X_3431_ net156 _0219_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_3362_ net122 _0150_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _0646_ po_0._1_\[10\] VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__and2_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ net146 _0081_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ po_0.alu_0._11_\[5\] _0708_ _0705_ _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__a211o_1
X_2175_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__clkbuf_2
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1959_ po_0.regf_0.rf\[4\]\[11\] po_0.regf_0.rf\[5\]\[11\] po_0.regf_0.rf\[6\]\[11\]
+ po_0.regf_0.rf\[7\]\[11\] _0395_ _0397_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__mux4_1
Xoutput49 net49 VGND VGND VPWR VPWR D_W_data[8] sky130_fd_sc_hd__buf_2
Xoutput38 net83 VGND VGND VPWR VPWR D_W_data[12] sky130_fd_sc_hd__buf_2
XFILLER_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2931_ _1237_ _1215_ _1240_ _1245_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__o22a_1
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2862_ _1180_ _1181_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__or2_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1813_ po_0.regf_0.rf\[4\]\[14\] po_0.regf_0.rf\[5\]\[14\] po_0.regf_0.rf\[6\]\[14\]
+ po_0.regf_0.rf\[7\]\[14\] _1460_ _1462_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__mux4_1
X_2793_ _1125_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1744_ _1456_ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__buf_2
XFILLER_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3414_ net105 _0202_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_1675_ _1459_ _1469_ _1474_ _1480_ VGND VGND VPWR VPWR po_0.regf_0._5_\[0\] sky130_fd_sc_hd__o22a_1
X_3345_ net138 _0133_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ net173 _0064_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _0754_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2158_ net41 po_0._1_\[15\] VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__and2b_1
X_2089_ _0625_ _0629_ VGND VGND VPWR VPWR po_0.alu_0._10_\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3130_ net88 _1311_ _0575_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__a21bo_1
X_3061_ po_0.regf_0.rf\[3\]\[1\] _0731_ _1332_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__mux2_1
XFILLER_35_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2012_ _0565_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2914_ _1226_ _1227_ _1229_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__a21oi_1
X_2845_ _1136_ _1151_ _1161_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__and3_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2776_ _1115_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__clkbuf_1
X_1727_ _1453_ _1527_ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__and2b_1
X_1658_ po_0.regf_0.rf\[12\]\[0\] po_0.regf_0.rf\[13\]\[0\] po_0.regf_0.rf\[14\]\[0\]
+ po_0.regf_0.rf\[15\]\[0\] _1461_ _1463_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__mux4_1
X_3328_ net137 _0116_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ _1403_ _1407_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__or2b_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ net133 _0051_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2630_ _0859_ po_0.regf_0.rf\[13\]\[13\] _1020_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__mux2_1
X_2561_ po_0.regf_0.rf\[15\]\[14\] _0958_ _0981_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__mux2_1
X_2492_ _0879_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3113_ po_0.regf_0.rf\[2\]\[9\] _0819_ _1358_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__mux2_1
X_3044_ _1324_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2828_ net68 po_0.muxf_0.rf_w_data\[1\] VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__nor2_2
X_2759_ _0796_ po_0.regf_0.rf\[0\]\[7\] _1105_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__mux2_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout84 net37 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
Xfanout95 po_0.regf_0.rq_rd VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1992_ _0546_ _0547_ _0422_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__mux2_1
XFILLER_60_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2613_ _0773_ po_0.regf_0.rf\[13\]\[5\] _1021_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__mux2_1
X_2544_ _0981_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__buf_2
X_2475_ po_0.regf_0.rf\[9\]\[9\] _0948_ _0942_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__mux2_1
XFILLER_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3027_ _1315_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2260_ _0783_ po_0.regf_0.rf\[7\]\[6\] _0784_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__mux2_1
XFILLER_69_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2191_ _0721_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1975_ _0532_ _0431_ _0424_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__a21o_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2527_ _0979_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
X_2458_ _0762_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__clkbuf_2
XFILLER_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2389_ po_0.regf_0.rf\[6\]\[7\] _0796_ _0895_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__mux2_1
XFILLER_68_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1760_ _1557_ _1466_ _1468_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__a21bo_1
X_1691_ po_0.regf_0.rf\[0\]\[1\] po_0.regf_0.rf\[1\]\[1\] po_0.regf_0.rf\[2\]\[1\]
+ po_0.regf_0.rf\[3\]\[1\] _1494_ _1495_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__mux4_1
X_3430_ net151 _0218_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_3361_ net145 _0149_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2312_ _0646_ po_0._1_\[10\] _0658_ _0824_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__a211o_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ net147 _0080_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _0767_ _0768_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__nor2_1
X_2174_ _1404_ _1401_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__nor2_2
XFILLER_65_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1958_ _0511_ _0513_ _0515_ _0517_ VGND VGND VPWR VPWR po_0.regf_0._3_\[10\] sky130_fd_sc_hd__o22a_1
X_1889_ po_0.regf_0.rf\[8\]\[3\] po_0.regf_0.rf\[9\]\[3\] po_0.regf_0.rf\[10\]\[3\]
+ po_0.regf_0.rf\[11\]\[3\] _0405_ _0407_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__mux4_1
Xoutput39 net39 VGND VGND VPWR VPWR D_W_data[13] sky130_fd_sc_hd__buf_2
X_3559_ po_0.alu_0._10_\[0\] _1558_ VGND VGND VPWR VPWR po_0.alu_0._11_\[0\] sky130_fd_sc_hd__ebufn_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2930_ _1237_ _1243_ _1244_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__o21ba_1
XFILLER_62_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2861_ _1175_ _1176_ _1179_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__and3_1
X_1812_ po_0.regf_0.rf\[0\]\[14\] po_0.regf_0.rf\[1\]\[14\] po_0.regf_0.rf\[2\]\[14\]
+ po_0.regf_0.rf\[3\]\[14\] _1497_ _1498_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__mux4_1
X_2792_ po_0.regf_0.rf\[8\]\[6\] _0782_ _1124_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__mux2_1
X_1743_ _1454_ VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__clkbuf_4
X_1674_ _1477_ _1478_ _1479_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__a21o_1
X_3413_ net103 _0201_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_3344_ net137 _0132_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ net159 _0011_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__dfxtp_2
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2226_ _0753_ po_0.regf_0.rf\[7\]\[3\] _0720_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__mux2_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2157_ po_0._1_\[15\] net41 VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__and2b_1
X_2088_ _0617_ _0628_ _0624_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__and3_1
XFILLER_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3060_ _1333_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2011_ po_0.regf_0.rq_addr\[0\] _0557_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__mux2_1
XFILLER_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2913_ _1204_ _1221_ _1228_ net98 _0568_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__a32o_1
X_2844_ _1152_ _1163_ _1160_ _1162_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__o211ai_1
X_2775_ _0880_ po_0.regf_0.rf\[0\]\[15\] _1097_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__mux2_1
X_1726_ po_0.regf_0.rf\[8\]\[5\] po_0.regf_0.rf\[9\]\[5\] po_0.regf_0.rf\[10\]\[5\]
+ po_0.regf_0.rf\[11\]\[5\] _1455_ _1457_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__mux4_1
X_1657_ _1462_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__clkbuf_4
X_1588_ _1411_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__clkbuf_1
X_3327_ net130 _0115_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3258_ net133 _0050_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3189_ _1289_ _1309_ _1400_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o21a_1
X_2209_ _0592_ _0593_ _0736_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__o31a_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2560_ _0997_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
X_2491_ _0959_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3112_ _1361_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3043_ po_0.regf_0.rf\[4\]\[9\] _0819_ _1320_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__mux2_1
XFILLER_63_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2827_ _1135_ _1137_ _1143_ _1149_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a31o_1
X_2758_ _1106_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__clkbuf_1
X_1709_ _1454_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__clkbuf_4
X_2689_ po_0.regf_0.rf\[11\]\[7\] _0944_ _1067_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__mux2_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout96 net66 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_4
Xfanout85 net48 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
XFILLER_10_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1991_ po_0.regf_0.rf\[4\]\[14\] po_0.regf_0.rf\[5\]\[14\] po_0.regf_0.rf\[6\]\[14\]
+ po_0.regf_0.rf\[7\]\[14\] _0414_ _0415_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__mux4_1
XFILLER_9_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2612_ _1026_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2543_ _0988_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
X_2474_ _0819_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__clkbuf_2
XFILLER_68_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3026_ po_0.regf_0.rf\[4\]\[1\] _0731_ _1313_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__mux2_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2190_ _0714_ po_0.regf_0.rf\[7\]\[0\] _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__mux2_1
XFILLER_1_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1974_ po_0.regf_0.rf\[4\]\[12\] po_0.regf_0.rf\[5\]\[12\] po_0.regf_0.rf\[6\]\[12\]
+ po_0.regf_0.rf\[7\]\[12\] _0428_ _0429_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__mux4_1
XFILLER_60_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2526_ po_0.regf_0.rf\[1\]\[14\] _0958_ _0962_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__mux2_1
X_2457_ _0936_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
X_2388_ _0896_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3009_ net79 net20 _1295_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__mux2_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1690_ _0005_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__buf_2
XFILLER_51_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3360_ net145 _0148_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2311_ _0831_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ net170 _0079_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2242_ _0765_ _0766_ _0757_ _0707_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__a31o_1
X_2173_ po_0.muxf_0.rf_w_data\[0\] VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__buf_2
XFILLER_53_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1957_ _0423_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__and2b_1
X_1888_ _0454_ _0447_ _0401_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__a21bo_1
X_3558_ net164 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
X_2509_ _0962_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__buf_2
X_3489_ net147 _0273_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2860_ _1175_ _1176_ _1179_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__a21oi_1
XFILLER_70_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1811_ _1453_ _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__and2b_1
X_2791_ _1116_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__buf_2
X_1742_ _1536_ _1538_ _1493_ _1541_ VGND VGND VPWR VPWR po_0.regf_0._5_\[6\] sky130_fd_sc_hd__o22a_1
X_1673_ _1467_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__buf_2
X_3412_ net104 _0200_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ net131 _0131_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ net153 _0010_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__dfxtp_1
X_2225_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2156_ _0680_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__inv_2
X_2087_ _0626_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__nand2_2
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2989_ _0744_ net26 _1289_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__mux2_1
XFILLER_21_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2010_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__buf_2
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2912_ _1219_ _1220_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__and2_1
X_2843_ _1155_ _0724_ _1160_ _1162_ _1163_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__a221o_1
X_2774_ _1114_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__clkbuf_1
X_1725_ _1520_ _1522_ _1524_ _1526_ VGND VGND VPWR VPWR po_0.regf_0._5_\[4\] sky130_fd_sc_hd__o22a_1
X_1656_ _0005_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__buf_2
X_1587_ _1403_ _1407_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__or2b_1
X_3326_ net130 _0114_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3257_ net134 _0049_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ net77 _1308_ _1309_ _1400_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__o31a_1
X_2208_ _0590_ _0736_ _0707_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__a21oi_1
XFILLER_66_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2139_ net39 po_0._1_\[13\] VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__nor2_1
XFILLER_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2490_ po_0.regf_0.rf\[9\]\[14\] _0958_ _0928_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__mux2_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3111_ po_0.regf_0.rf\[2\]\[8\] _0810_ _1358_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__mux2_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3042_ _1323_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2826_ _1145_ _1148_ _1138_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__mux2_1
X_2757_ _0783_ po_0.regf_0.rf\[0\]\[6\] _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__mux2_1
X_1708_ _1452_ VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__clkbuf_2
X_2688_ _1068_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
X_1639_ _1447_ VGND VGND VPWR VPWR uc_0.bc_0._54_\[0\] sky130_fd_sc_hd__buf_2
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ net144 _0097_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout97 net75 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout86 net42 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1990_ po_0.regf_0.rf\[0\]\[14\] po_0.regf_0.rf\[1\]\[14\] po_0.regf_0.rf\[2\]\[14\]
+ po_0.regf_0.rf\[3\]\[14\] _0414_ _0415_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__mux4_1
XFILLER_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2611_ _0763_ po_0.regf_0.rf\[13\]\[4\] _1021_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__mux2_1
X_2542_ po_0.regf_0.rf\[15\]\[5\] _0939_ _0982_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__mux2_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2473_ _0947_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3025_ _1314_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2809_ _1133_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1973_ _0447_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__and2b_1
X_3574_ po_0.alu_0._10_\[15\] _1573_ VGND VGND VPWR VPWR po_0.alu_0._11_\[15\] sky130_fd_sc_hd__ebufn_1
X_2525_ _0978_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
X_2456_ po_0.regf_0.rf\[9\]\[3\] _0935_ _0929_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__mux2_1
XFILLER_29_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2387_ po_0.regf_0.rf\[6\]\[6\] _0783_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__mux2_1
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3008_ _1303_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2310_ _0830_ po_0.regf_0.rf\[7\]\[10\] _0784_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__mux2_1
X_3290_ net157 _0078_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2241_ _0765_ _0757_ _0766_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__a21oi_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2172_ _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__buf_2
XFILLER_80_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1956_ po_0.regf_0.rf\[8\]\[10\] po_0.regf_0.rf\[9\]\[10\] po_0.regf_0.rf\[10\]\[10\]
+ po_0.regf_0.rf\[11\]\[10\] _0448_ _0449_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__mux4_1
X_1887_ po_0.regf_0.rf\[12\]\[3\] po_0.regf_0.rf\[13\]\[3\] po_0.regf_0.rf\[14\]\[3\]
+ po_0.regf_0.rf\[15\]\[3\] _0395_ _0397_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__mux4_1
X_3557_ net181 uc_0.bc_0._54_\[3\] VGND VGND VPWR VPWR uc_0.bc_0._55_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2508_ _0969_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
X_3488_ net127 _0272_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_2439_ _0924_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1810_ po_0.regf_0.rf\[8\]\[14\] po_0.regf_0.rf\[9\]\[14\] po_0.regf_0.rf\[10\]\[14\]
+ po_0.regf_0.rf\[11\]\[14\] _1455_ _1457_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux4_1
X_2790_ _1123_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1741_ _1539_ _1540_ _1500_ VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__mux2_1
X_1672_ _1465_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__buf_2
X_3411_ net112 _0199_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3342_ net131 _0130_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ net171 _0009_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__dfxtp_2
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ net10 _0700_ _0703_ _0744_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__a221o_4
X_2155_ _0686_ _0687_ VGND VGND VPWR VPWR po_0.alu_0._10_\[14\] sky130_fd_sc_hd__nor2_1
XFILLER_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2086_ net47 _0621_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__or2b_1
XFILLER_34_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2988_ _1292_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1939_ po_0.regf_0.rf\[8\]\[8\] po_0.regf_0.rf\[9\]\[8\] po_0.regf_0.rf\[10\]\[8\]
+ po_0.regf_0.rf\[11\]\[8\] _0435_ _0436_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__mux4_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2911_ net74 po_0.muxf_0.rf_w_data\[7\] VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__nand2_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2842_ _1151_ _0724_ _1136_ po_0.muxf_0.rf_w_data\[0\] VGND VGND VPWR VPWR _1163_
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2773_ _0871_ po_0.regf_0.rf\[0\]\[14\] _1097_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__mux2_1
X_1724_ _1525_ _1478_ _1479_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__a21o_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1655_ _1460_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__clkbuf_4
X_1586_ _1410_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__clkbuf_1
X_3325_ net136 _0113_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ net134 _0048_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2207_ _1429_ _0582_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__o21ai_2
XFILLER_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3187_ _0572_ _0559_ _0573_ _1389_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__o31a_1
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2138_ net83 VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__inv_2
X_2069_ _0609_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__and2b_1
XFILLER_81_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3110_ _1360_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3041_ po_0.regf_0.rf\[4\]\[8\] _0810_ _1320_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__mux2_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2825_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__buf_2
XFILLER_31_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2756_ _1097_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__buf_2
X_1707_ _1509_ _1470_ _1485_ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__a21bo_1
X_2687_ po_0.regf_0.rf\[11\]\[6\] _0941_ _1067_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__mux2_1
X_1638_ _1446_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__inv_2
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ net144 _0096_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ po_0.regf_0._5_\[15\] net93 VGND VGND VPWR VPWR po_0._1_\[15\] sky130_fd_sc_hd__dlxtp_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout87 net35 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout98 net73 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_2
XFILLER_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2610_ _1025_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
X_2541_ _0987_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
X_2472_ po_0.regf_0.rf\[9\]\[8\] _0946_ _0942_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__mux2_1
XFILLER_5_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3024_ po_0.regf_0.rf\[4\]\[0\] _0713_ _1313_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__mux2_1
XFILLER_24_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2808_ po_0.regf_0.rf\[8\]\[14\] _0870_ _1116_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__mux2_1
X_2739_ _1095_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1972_ po_0.regf_0.rf\[0\]\[12\] po_0.regf_0.rf\[1\]\[12\] po_0.regf_0.rf\[2\]\[12\]
+ po_0.regf_0.rf\[3\]\[12\] _0448_ _0449_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__mux4_1
X_3573_ po_0.alu_0._10_\[14\] _1572_ VGND VGND VPWR VPWR po_0.alu_0._11_\[14\] sky130_fd_sc_hd__ebufn_1
X_2524_ po_0.regf_0.rf\[1\]\[13\] _0956_ _0962_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__mux2_1
X_2455_ _0752_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__clkbuf_2
X_2386_ _0887_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__buf_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3007_ uc_0._20_\[11\] net19 _1295_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__mux2_1
XFILLER_24_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _0614_ _0615_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__or2_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2171_ po_0.muxf_0.s0 _0698_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__nor2_1
XFILLER_65_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1955_ _0514_ _0444_ _0445_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__a21bo_1
X_1886_ _0440_ _0446_ _0451_ _0453_ VGND VGND VPWR VPWR po_0.regf_0._3_\[2\] sky130_fd_sc_hd__o22a_1
X_3556_ net181 uc_0.bc_0._54_\[2\] VGND VGND VPWR VPWR uc_0.bc_0._55_\[2\] sky130_fd_sc_hd__dfxtp_1
X_2507_ po_0.regf_0.rf\[1\]\[5\] _0939_ _0963_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__mux2_1
X_3487_ net126 _0271_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_2438_ po_0.regf_0.rf\[5\]\[13\] _0859_ _0908_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__mux2_1
X_2369_ po_0.regf_0.w_addr\[1\] VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1740_ po_0.regf_0.rf\[4\]\[6\] po_0.regf_0.rf\[5\]\[6\] po_0.regf_0.rf\[6\]\[6\]
+ po_0.regf_0.rf\[7\]\[6\] _1460_ _1462_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__mux4_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1671_ po_0.regf_0.rf\[4\]\[0\] po_0.regf_0.rf\[5\]\[0\] po_0.regf_0.rf\[6\]\[0\]
+ po_0.regf_0.rf\[7\]\[0\] _1475_ _1476_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__mux4_1
X_3410_ net114 _0198_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3341_ net138 _0129_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ net160 _0008_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__dfxtp_2
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _0598_ _0745_ _1402_ _0711_ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__o311a_1
X_2154_ _0679_ _0681_ _0682_ _0685_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__and4_1
X_2085_ po_0._1_\[6\] net47 VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__or2b_1
XFILLER_61_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2987_ _0734_ net25 _1289_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__mux2_1
X_1938_ _0499_ _0444_ _0445_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__a21bo_1
X_1869_ _0434_ _0437_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__and2b_1
X_3539_ net180 _0323_ VGND VGND VPWR VPWR po_0.muxf_0.s1 sky130_fd_sc_hd__dfxtp_1
XFILLER_67_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2910_ _1225_ _0570_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__or2_2
X_2841_ _1161_ _0734_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__or2_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2772_ _1113_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__clkbuf_1
X_1723_ po_0.regf_0.rf\[4\]\[4\] po_0.regf_0.rf\[5\]\[4\] po_0.regf_0.rf\[6\]\[4\]
+ po_0.regf_0.rf\[7\]\[4\] _1475_ _1476_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__mux4_1
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1654_ _0004_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__clkbuf_4
X_1585_ _1403_ _1407_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__or2b_1
X_3324_ net136 _0112_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ po_0.regf_0._3_\[15\] net89 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlxtp_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ net86 po_0._1_\[1\] VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__nand2_1
X_3186_ _1399_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__clkbuf_1
X_2137_ _0664_ _0671_ VGND VGND VPWR VPWR po_0.alu_0._10_\[12\] sky130_fd_sc_hd__xnor2_1
X_2068_ _0601_ _0610_ _0608_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__nand3_1
XFILLER_81_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3040_ _1322_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2824_ uc_0._01_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__nor2_1
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2755_ _1104_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__clkbuf_1
X_1706_ po_0.regf_0.rf\[12\]\[3\] po_0.regf_0.rf\[13\]\[3\] po_0.regf_0.rf\[14\]\[3\]
+ po_0.regf_0.rf\[15\]\[3\] _1481_ _1482_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__mux4_1
X_2686_ _1059_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__buf_2
X_1637_ _1436_ _1437_ _1438_ _1445_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__o31ai_2
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ net141 _0095_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3238_ po_0.regf_0._5_\[14\] net93 VGND VGND VPWR VPWR po_0._1_\[14\] sky130_fd_sc_hd__dlxtp_1
X_3169_ _1389_ uc_0.bc_0._54_\[0\] net59 _1311_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout99 net70 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
Xfanout88 net91 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2540_ po_0.regf_0.rf\[15\]\[4\] _0937_ _0982_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__mux2_1
XFILLER_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2471_ _0810_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__clkbuf_2
XFILLER_68_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3023_ _1312_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__buf_2
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2807_ _1132_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__clkbuf_1
X_2738_ po_0.regf_0.rf\[10\]\[14\] _0958_ _1078_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__mux2_1
X_2669_ _1057_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1971_ _0528_ _0434_ _0401_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__a21bo_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3572_ po_0.alu_0._10_\[13\] _1571_ VGND VGND VPWR VPWR po_0.alu_0._11_\[13\] sky130_fd_sc_hd__ebufn_1
X_2523_ _0977_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_2454_ _0934_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
X_2385_ _0894_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput1 D_R_data[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3006_ _1302_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2170_ _0700_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__buf_2
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1954_ po_0.regf_0.rf\[12\]\[10\] po_0.regf_0.rf\[13\]\[10\] po_0.regf_0.rf\[14\]\[10\]
+ po_0.regf_0.rf\[15\]\[10\] _0441_ _0442_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__mux4_1
X_1885_ _0452_ _0431_ _0410_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__a21o_1
X_3555_ net177 uc_0.bc_0._54_\[1\] VGND VGND VPWR VPWR uc_0.bc_0._55_\[1\] sky130_fd_sc_hd__dfxtp_1
X_3486_ net113 _0270_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2506_ _0968_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
X_2437_ _0923_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2368_ po_0.regf_0.w_addr\[0\] VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2299_ _0820_ po_0.regf_0.rf\[7\]\[9\] _0784_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__mux2_1
XFILLER_56_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1670_ _1462_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__buf_2
X_3340_ net138 _0128_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ net126 _0063_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _1405_ po_0.alu_0._11_\[3\] _0706_ _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__a211o_1
X_2153_ _0681_ _0682_ _0679_ _0685_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__a22oi_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2084_ _0622_ _0623_ _0624_ _0617_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__a2bb2oi_1
X_2986_ _1291_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1937_ po_0.regf_0.rf\[12\]\[8\] po_0.regf_0.rf\[13\]\[8\] po_0.regf_0.rf\[14\]\[8\]
+ po_0.regf_0.rf\[15\]\[8\] _0441_ _0442_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__mux4_1
X_1868_ po_0.regf_0.rf\[8\]\[1\] po_0.regf_0.rf\[9\]\[1\] po_0.regf_0.rf\[10\]\[1\]
+ po_0.regf_0.rf\[11\]\[1\] _0435_ _0436_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__mux4_1
X_1799_ po_0.regf_0.rf\[8\]\[13\] po_0.regf_0.rf\[9\]\[13\] po_0.regf_0.rf\[10\]\[13\]
+ po_0.regf_0.rf\[11\]\[13\] _1494_ _1495_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__mux4_1
X_3538_ net180 _0322_ VGND VGND VPWR VPWR po_0.muxf_0.s0 sky130_fd_sc_hd__dfxtp_1
X_3469_ net179 _0253_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfxtp_2
XFILLER_67_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2840_ net69 VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2771_ _0859_ po_0.regf_0.rf\[0\]\[13\] _1097_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__mux2_1
X_1722_ _1487_ _1523_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__and2b_1
X_1653_ _1453_ _1458_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__and2b_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1584_ _1409_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__clkbuf_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ net141 _0111_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ po_0.regf_0._3_\[14\] net89 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlxtp_1
X_2205_ po_0.muxf_0.rf_w_data\[2\] VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__clkbuf_4
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _0570_ net58 _1393_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__mux2_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2136_ _0667_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__nor2_1
XFILLER_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2067_ _0606_ _0607_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__nor2_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2969_ _1277_ _1171_ _1278_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__nand3b_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2823_ uc_0._00_ uc_0._02_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__or2_1
X_2754_ _0773_ po_0.regf_0.rf\[0\]\[5\] _1098_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__mux2_1
X_1705_ _1503_ _1505_ _1493_ _1508_ VGND VGND VPWR VPWR po_0.regf_0._5_\[2\] sky130_fd_sc_hd__o22a_1
X_2685_ _1066_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
X_1636_ net34 _1444_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__nor2_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ net122 _0094_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ po_0.regf_0._5_\[13\] net92 VGND VGND VPWR VPWR po_0._1_\[13\] sky130_fd_sc_hd__dlxtp_1
X_3168_ _0572_ uc_0.bc_0._54_\[0\] uc_0.bc_0._54_\[2\] _1311_ net60 VGND VGND VPWR
+ VPWR _0324_ sky130_fd_sc_hd__a32o_1
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2119_ _0649_ _0655_ VGND VGND VPWR VPWR po_0.alu_0._10_\[10\] sky130_fd_sc_hd__xnor2_1
X_3099_ _1354_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout89 net91 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2470_ _0945_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3022_ _0882_ _0906_ _1039_ _0886_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__and4b_4
XFILLER_36_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2806_ po_0.regf_0.rf\[8\]\[13\] _0858_ _1116_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__mux2_1
X_2737_ _1094_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__clkbuf_1
X_2668_ po_0.regf_0.rf\[12\]\[14\] _0958_ _1040_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__mux2_1
X_1619_ _1428_ _1429_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__and2_1
X_2599_ _0880_ po_0.regf_0.rf\[14\]\[15\] _1001_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__mux2_1
XFILLER_59_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1970_ po_0.regf_0.rf\[12\]\[12\] po_0.regf_0.rf\[13\]\[12\] po_0.regf_0.rf\[14\]\[12\]
+ po_0.regf_0.rf\[15\]\[12\] _0419_ _0420_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__mux4_1
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3571_ po_0.alu_0._10_\[12\] _1570_ VGND VGND VPWR VPWR po_0.alu_0._11_\[12\] sky130_fd_sc_hd__ebufn_1
X_2522_ po_0.regf_0.rf\[1\]\[12\] _0954_ _0962_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__mux2_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2453_ po_0.regf_0.rf\[9\]\[2\] _0933_ _0929_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__mux2_1
X_2384_ po_0.regf_0.rf\[6\]\[5\] _0773_ _0888_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__mux2_1
XFILLER_68_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 D_R_data[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3005_ uc_0._20_\[10\] net18 _1296_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__mux2_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1953_ _0494_ _0512_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__and2b_1
X_1884_ po_0.regf_0.rf\[4\]\[2\] po_0.regf_0.rf\[5\]\[2\] po_0.regf_0.rf\[6\]\[2\]
+ po_0.regf_0.rf\[7\]\[2\] _0428_ _0429_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__mux4_1
X_3554_ net179 uc_0.bc_0._54_\[0\] VGND VGND VPWR VPWR uc_0.bc_0._55_\[0\] sky130_fd_sc_hd__dfxtp_1
X_3485_ net110 _0269_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_2505_ po_0.regf_0.rf\[1\]\[4\] _0937_ _0963_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__mux2_1
X_2436_ po_0.regf_0.rf\[5\]\[12\] _0849_ _0908_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__mux2_1
X_2367_ po_0.regf_0.w_addr\[3\] VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2298_ _0819_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3270_ net126 _0062_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _0747_ _0725_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__and3_1
XFILLER_85_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2152_ _0683_ po_0._1_\[13\] _0684_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__o21a_1
XFILLER_38_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2083_ po_0._1_\[5\] _0613_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__or2b_1
XFILLER_53_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2985_ _0724_ net24 _1289_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__mux2_1
XFILLER_21_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1936_ _0494_ _0497_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__and2b_1
X_1867_ _0396_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__clkbuf_4
X_1798_ _0365_ _0367_ _0369_ _0371_ VGND VGND VPWR VPWR po_0.regf_0._5_\[12\] sky130_fd_sc_hd__o22a_1
X_3537_ net159 _0321_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[3\] sky130_fd_sc_hd__dfxtp_1
X_3468_ net164 _0252_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dfxtp_1
X_2419_ po_0.regf_0.rf\[5\]\[4\] _0763_ _0909_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__mux2_1
X_3399_ net120 _0187_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2770_ _1112_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__clkbuf_1
X_1721_ po_0.regf_0.rf\[0\]\[4\] po_0.regf_0.rf\[1\]\[4\] po_0.regf_0.rf\[2\]\[4\]
+ po_0.regf_0.rf\[3\]\[4\] _1488_ _1489_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__mux4_1
X_1652_ po_0.regf_0.rf\[8\]\[0\] po_0.regf_0.rf\[9\]\[0\] po_0.regf_0.rf\[10\]\[0\]
+ po_0.regf_0.rf\[11\]\[0\] _1455_ _1457_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__mux4_1
X_1583_ _1403_ _1407_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__or2b_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ net122 _0110_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ po_0.regf_0._3_\[13\] net91 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlxtp_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2204_ _0733_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _1398_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2135_ _0634_ _0641_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__a21oi_2
XFILLER_66_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2066_ _0606_ _0607_ _0608_ _0601_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2968_ net64 _1233_ _1263_ net65 VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__a31o_1
X_1919_ _0434_ _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__and2b_1
X_2899_ _1213_ _1209_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__nand2_1
XFILLER_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2822_ _1144_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__clkbuf_2
X_2753_ _1103_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__clkbuf_1
X_1704_ _1506_ _1507_ _1500_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__mux2_1
X_2684_ po_0.regf_0.rf\[11\]\[5\] _0939_ _1060_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__mux2_1
X_1635_ _1443_ uc_0.bc_0._55_\[1\] uc_0.bc_0._55_\[2\] uc_0.bc_0._55_\[3\] VGND VGND
+ VPWR VPWR _1444_ sky130_fd_sc_hd__a211oi_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ net123 _0093_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ po_0.regf_0._5_\[12\] net93 VGND VGND VPWR VPWR po_0._1_\[12\] sky130_fd_sc_hd__dlxtp_1
XFILLER_39_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3167_ _0723_ _1370_ _1390_ _0564_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__a211oi_1
X_3098_ po_0.regf_0.rf\[2\]\[2\] _0741_ _1351_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__mux2_1
X_2118_ _0651_ _0652_ _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__nand3_1
XFILLER_81_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2049_ _0592_ _0593_ _0585_ _0586_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__o211ai_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3021_ _1440_ _1139_ _1311_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__o21a_1
XFILLER_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2805_ _1131_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__clkbuf_1
X_2736_ po_0.regf_0.rf\[10\]\[13\] _0956_ _1078_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__mux2_1
X_2667_ _1056_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
X_1618_ po_0._1_\[0\] net87 VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__nand2_1
X_2598_ _1018_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
X_3219_ net100 _0043_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3570_ po_0.alu_0._10_\[11\] _1569_ VGND VGND VPWR VPWR po_0.alu_0._11_\[11\] sky130_fd_sc_hd__ebufn_1
X_2521_ _0976_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2452_ _0741_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__clkbuf_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2383_ _0893_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput3 D_R_data[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_3004_ _1301_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2719_ po_0.regf_0.rf\[10\]\[5\] _0939_ _1079_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__mux2_1
XFILLER_10_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1952_ po_0.regf_0.rf\[0\]\[10\] po_0.regf_0.rf\[1\]\[10\] po_0.regf_0.rf\[2\]\[10\]
+ po_0.regf_0.rf\[3\]\[10\] _0495_ _0496_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__mux4_1
X_1883_ _0447_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__and2b_1
X_3553_ net177 _0337_ VGND VGND VPWR VPWR uc_0._01_ sky130_fd_sc_hd__dfxtp_1
X_3484_ net101 _0268_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_2504_ _0967_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
X_2435_ _0922_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
X_2366_ _0881_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__clkbuf_1
X_2297_ _0722_ _0723_ net16 _0817_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__a32o_4
XFILLER_64_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _0587_ _0746_ _0602_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__o21ai_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2151_ _0672_ po_0._1_\[12\] _0675_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__or3_1
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2082_ _0620_ _0621_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__nor2_1
XFILLER_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2984_ _1290_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__clkbuf_1
X_1935_ po_0.regf_0.rf\[0\]\[8\] po_0.regf_0.rf\[1\]\[8\] po_0.regf_0.rf\[2\]\[8\]
+ po_0.regf_0.rf\[3\]\[8\] _0495_ _0496_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__mux4_1
X_1866_ _0394_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__buf_4
X_1797_ _1550_ _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__and2b_1
X_3536_ net158 _0320_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[2\] sky130_fd_sc_hd__dfxtp_1
X_3467_ net155 _0251_ VGND VGND VPWR VPWR uc_0._20_\[11\] sky130_fd_sc_hd__dfxtp_1
X_2418_ _0913_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
X_3398_ net150 _0186_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_2349_ _0863_ _0864_ _0865_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1720_ _1521_ _1466_ _1468_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__a21bo_1
X_1651_ _1456_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__buf_2
X_3321_ net122 _0109_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_1582_ _1408_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__clkbuf_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ po_0.regf_0._3_\[12\] net89 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlxtp_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _0732_ po_0.regf_0.rf\[7\]\[1\] _0720_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__mux2_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _0568_ net57 _1393_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__mux2_1
X_2134_ _0668_ _0643_ _0649_ _0658_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__or4_1
XFILLER_26_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2065_ po_0._1_\[3\] _0598_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__or2b_1
X_2967_ net64 net65 _1233_ _1263_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__and4_1
X_1918_ po_0.regf_0.rf\[8\]\[6\] po_0.regf_0.rf\[9\]\[6\] po_0.regf_0.rf\[10\]\[6\]
+ po_0.regf_0.rf\[11\]\[6\] _0435_ _0436_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__mux4_1
X_2898_ _1214_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__clkbuf_2
X_1849_ _0402_ _0409_ _0410_ _0418_ VGND VGND VPWR VPWR po_0.regf_0._3_\[0\] sky130_fd_sc_hd__o22a_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3519_ net114 _0303_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2821_ _1140_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2752_ _0763_ po_0.regf_0.rf\[0\]\[4\] _1098_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__mux2_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1703_ po_0.regf_0.rf\[4\]\[2\] po_0.regf_0.rf\[5\]\[2\] po_0.regf_0.rf\[6\]\[2\]
+ po_0.regf_0.rf\[7\]\[2\] _1497_ _1498_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__mux4_1
X_2683_ _1065_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
X_1634_ net80 net81 net82 net79 _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__a2111o_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ net141 _0092_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ po_0.regf_0._5_\[11\] net93 VGND VGND VPWR VPWR po_0._1_\[11\] sky130_fd_sc_hd__dlxtp_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3166_ _0722_ _1390_ _1370_ _1371_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__o211a_1
X_3097_ _1353_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__clkbuf_1
X_2117_ _0640_ _0642_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__nand3_1
XFILLER_81_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2048_ po_0._1_\[2\] _0588_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__and2b_1
XFILLER_22_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3020_ _1310_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__buf_2
XFILLER_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2804_ po_0.regf_0.rf\[8\]\[12\] _0848_ _1116_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__mux2_1
X_2735_ _1093_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__clkbuf_1
X_2666_ po_0.regf_0.rf\[12\]\[13\] _0956_ _1040_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__mux2_1
X_1617_ po_0._1_\[0\] net87 VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__or2_1
X_2597_ _0871_ po_0.regf_0.rf\[14\]\[14\] _1001_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__mux2_1
XFILLER_75_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3218_ net100 _0042_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3149_ _1379_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2520_ po_0.regf_0.rf\[1\]\[11\] _0952_ _0970_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__mux2_1
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2451_ _0932_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
X_2382_ po_0.regf_0.rf\[6\]\[4\] _0763_ _0888_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__mux2_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput4 D_R_data[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
X_3003_ uc_0._20_\[9\] net32 _1296_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__mux2_1
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2718_ _1084_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
X_2649_ po_0.regf_0.rf\[12\]\[5\] _0939_ _1041_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__mux2_1
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1951_ _0510_ _0400_ _0432_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__a21o_1
XFILLER_14_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1882_ po_0.regf_0.rf\[0\]\[2\] po_0.regf_0.rf\[1\]\[2\] po_0.regf_0.rf\[2\]\[2\]
+ po_0.regf_0.rf\[3\]\[2\] _0448_ _0449_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__mux4_1
X_3552_ net177 _0336_ VGND VGND VPWR VPWR uc_0._02_ sky130_fd_sc_hd__dfxtp_1
X_2503_ po_0.regf_0.rf\[1\]\[3\] _0935_ _0963_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__mux2_1
X_3483_ net101 _0267_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_2434_ po_0.regf_0.rf\[5\]\[11\] _0839_ _0916_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__mux2_1
X_2365_ _0880_ po_0.regf_0.rf\[7\]\[15\] _0719_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__mux2_1
X_2296_ _0650_ _1406_ _1402_ _0793_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__o31a_1
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_20 _1500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2150_ net39 VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__inv_2
X_2081_ _0620_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__and2_1
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2983_ _0704_ net17 _1289_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__mux2_1
X_1934_ _0406_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__buf_2
X_1865_ _0422_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__clkbuf_2
X_1796_ po_0.regf_0.rf\[8\]\[12\] po_0.regf_0.rf\[9\]\[12\] po_0.regf_0.rf\[10\]\[12\]
+ po_0.regf_0.rf\[11\]\[12\] _1471_ _1472_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__mux4_1
X_3535_ net159 _0319_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[1\] sky130_fd_sc_hd__dfxtp_1
X_3466_ net155 _0250_ VGND VGND VPWR VPWR uc_0._20_\[10\] sky130_fd_sc_hd__dfxtp_1
X_2417_ po_0.regf_0.rf\[5\]\[3\] _0753_ _0909_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__mux2_1
X_3397_ net150 _0185_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2348_ _0681_ _0682_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__nand2_1
X_2279_ _0620_ _0621_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__nand2_1
XFILLER_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1650_ _0005_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1581_ _1403_ _1407_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__or2b_1
X_3320_ net129 _0108_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ po_0.regf_0._3_\[11\] net88 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlxtp_1
XFILLER_85_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2202_ _0731_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ _1397_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2133_ _0638_ _0639_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__and2_1
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2064_ _0605_ po_0._1_\[4\] VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__nor2_1
X_2966_ net64 net65 _1242_ _1263_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__and4_1
X_1917_ _0480_ _0444_ _0432_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a21bo_1
X_2897_ uc_0._01_ _1139_ _1144_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__or3_1
X_1848_ _0413_ _0416_ _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux2_1
X_1779_ _0353_ _0354_ _1465_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux2_1
X_3518_ net124 _0302_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3449_ net165 _0237_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfxtp_1
XFILLER_76_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2820_ _1138_ _0704_ _1142_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__o21a_1
X_2751_ _1102_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__clkbuf_1
X_1702_ po_0.regf_0.rf\[0\]\[2\] po_0.regf_0.rf\[1\]\[2\] po_0.regf_0.rf\[2\]\[2\]
+ po_0.regf_0.rf\[3\]\[2\] _1494_ _1495_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__mux4_1
X_2682_ po_0.regf_0.rf\[11\]\[4\] _0937_ _1060_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__mux2_1
X_1633_ uc_0.bc_0._55_\[0\] VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__inv_2
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3303_ net120 _0091_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ po_0.regf_0._5_\[10\] net92 VGND VGND VPWR VPWR po_0._1_\[10\] sky130_fd_sc_hd__dlxtp_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3165_ uc_0.bc_0._54_\[0\] _1389_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__nor2_1
X_3096_ po_0.regf_0.rf\[2\]\[1\] _0731_ _1351_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__mux2_1
XFILLER_66_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2116_ _0650_ po_0._1_\[9\] VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__xnor2_1
X_2047_ _0588_ po_0._1_\[2\] VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__and2b_1
X_2949_ _1261_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2803_ _1130_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__clkbuf_1
X_2734_ po_0.regf_0.rf\[10\]\[12\] _0954_ _1078_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__mux2_1
X_2665_ _1055_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
X_2596_ _1017_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
X_1616_ _1427_ VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__clkbuf_1
X_3217_ net102 _0041_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_3148_ uc_0._20_\[10\] po_0.regf_0.rp_addr\[2\] _0574_ VGND VGND VPWR VPWR _1379_
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3079_ _1343_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2450_ po_0.regf_0.rf\[9\]\[1\] _0931_ _0929_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__mux2_1
X_2381_ _0892_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
Xinput5 D_R_data[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3002_ _1300_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2717_ po_0.regf_0.rf\[10\]\[4\] _0937_ _1079_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__mux2_1
X_2648_ _1046_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
X_2579_ _1008_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1950_ po_0.regf_0.rf\[4\]\[10\] po_0.regf_0.rf\[5\]\[10\] po_0.regf_0.rf\[6\]\[10\]
+ po_0.regf_0.rf\[7\]\[10\] _0395_ _0397_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__mux4_1
X_1881_ _0396_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__buf_2
X_3551_ net178 _0335_ VGND VGND VPWR VPWR uc_0._03_ sky130_fd_sc_hd__dfxtp_1
X_2502_ _0966_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
X_3482_ net105 _0266_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_2433_ _0921_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
X_2364_ _0879_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2295_ _0813_ _0708_ _0814_ _0816_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__o31ai_1
XFILLER_24_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_10 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 po_0.regf_0._5_\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2080_ po_0._1_\[6\] VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2982_ uc_0._03_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__buf_2
X_1933_ _0404_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__clkbuf_4
X_1864_ _0430_ _0431_ _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__a21bo_1
Xinput30 I_data[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
X_1795_ _0368_ _1466_ _1468_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__a21bo_1
X_3534_ net159 _0318_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[0\] sky130_fd_sc_hd__dfxtp_1
X_3465_ net160 _0249_ VGND VGND VPWR VPWR uc_0._20_\[9\] sky130_fd_sc_hd__dfxtp_1
X_2416_ _0912_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
X_3396_ net119 _0184_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_2347_ _0852_ _0673_ _0674_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__o21ba_1
X_2278_ net48 po_0._1_\[7\] VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__or2_1
XFILLER_84_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1580_ _1406_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3250_ po_0.regf_0._3_\[10\] net88 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlxtp_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _0722_ _0723_ net8 _0730_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__a31o_2
X_3181_ _0566_ net56 _1393_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__mux2_1
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2132_ net84 _0665_ _0666_ _0647_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__a22o_1
XFILLER_66_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2063_ _0605_ po_0._1_\[4\] VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__and2_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2965_ _1269_ _1243_ _1264_ net65 VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__a31oi_1
X_1916_ po_0.regf_0.rf\[12\]\[6\] po_0.regf_0.rf\[13\]\[6\] po_0.regf_0.rf\[14\]\[6\]
+ po_0.regf_0.rf\[15\]\[6\] _0441_ _0442_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__mux4_1
X_2896_ net98 VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__clkbuf_2
X_1847_ _0002_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__clkbuf_2
X_1778_ po_0.regf_0.rf\[4\]\[10\] po_0.regf_0.rf\[5\]\[10\] po_0.regf_0.rf\[6\]\[10\]
+ po_0.regf_0.rf\[7\]\[10\] _1460_ _1462_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux4_1
X_3517_ net124 _0301_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3448_ net163 _0236_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfxtp_4
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ net158 _0167_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2750_ _0753_ po_0.regf_0.rf\[0\]\[3\] _1098_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__mux2_1
X_1701_ _1487_ _1504_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__and2b_1
X_2681_ _1064_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
X_1632_ _1441_ VGND VGND VPWR VPWR uc_0.bc_0._54_\[1\] sky130_fd_sc_hd__inv_2
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ net117 _0090_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ po_0.regf_0._5_\[9\] net92 VGND VGND VPWR VPWR po_0._1_\[9\] sky130_fd_sc_hd__dlxtp_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3164_ _1369_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__clkbuf_2
X_3095_ _1352_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__clkbuf_1
X_2115_ po_0._1_\[8\] _0643_ _0637_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or3b_1
X_2046_ _0585_ _0586_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2948_ _1260_ _1256_ _1148_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__mux2_1
X_2879_ _1196_ _1197_ _1171_ _1147_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__a31o_1
XFILLER_77_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2802_ po_0.regf_0.rf\[8\]\[11\] _0838_ _1124_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__mux2_1
X_2733_ _1092_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__clkbuf_1
X_2664_ po_0.regf_0.rf\[12\]\[12\] _0954_ _1040_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__mux2_1
X_2595_ _0859_ po_0.regf_0.rf\[14\]\[13\] _1001_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__mux2_1
X_1615_ _1413_ _1415_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__or2b_1
X_3216_ net102 _0040_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3147_ _1378_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3078_ po_0.regf_0.rf\[3\]\[9\] _0819_ _1339_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__mux2_1
X_2029_ _0577_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2380_ po_0.regf_0.rf\[6\]\[3\] _0753_ _0888_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__mux2_1
Xinput6 D_R_data[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3001_ uc_0._20_\[8\] net31 _1296_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__mux2_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2716_ _1083_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2647_ po_0.regf_0.rf\[12\]\[4\] _0937_ _1041_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__mux2_1
X_2578_ _0773_ po_0.regf_0.rf\[14\]\[5\] _1002_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__mux2_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _0394_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__clkbuf_4
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3550_ net178 _0334_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfxtp_1
X_2501_ po_0.regf_0.rf\[1\]\[2\] _0933_ _0963_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__mux2_1
X_3481_ net101 _0265_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_2432_ po_0.regf_0.rf\[5\]\[10\] _0830_ _0916_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__mux2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2363_ po_0.muxf_0.s0 _0698_ net7 _0876_ _0878_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__a32o_2
XFILLER_56_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2294_ _1406_ po_0.alu_0._11_\[9\] _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_11 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2981_ net67 _1207_ _1287_ _1288_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__o31ai_1
X_1932_ _0399_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__clkbuf_2
XFILLER_61_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1863_ _0003_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__buf_2
Xinput20 I_data[12] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
Xinput31 I_data[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
X_1794_ po_0.regf_0.rf\[12\]\[12\] po_0.regf_0.rf\[13\]\[12\] po_0.regf_0.rf\[14\]\[12\]
+ po_0.regf_0.rf\[15\]\[12\] _1461_ _1463_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__mux4_1
X_3533_ net153 _0317_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[3\] sky130_fd_sc_hd__dfxtp_1
X_3464_ net159 _0248_ VGND VGND VPWR VPWR uc_0._20_\[8\] sky130_fd_sc_hd__dfxtp_1
X_2415_ po_0.regf_0.rf\[5\]\[2\] _0742_ _0909_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__mux2_1
X_3395_ net158 _0183_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2346_ _0861_ _0862_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__nand2_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2277_ _0590_ _0736_ _0755_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _0724_ _0702_ _0728_ _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__a22o_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3180_ _1396_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2131_ _0658_ _0659_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__nor2_1
X_2062_ net45 VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__clkbuf_2
XFILLER_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2964_ _1269_ _1215_ _1272_ _1274_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__o22a_1
X_1915_ _0403_ _0478_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__and2b_1
X_2895_ _1135_ _1200_ _1187_ _1212_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__o31a_1
X_1846_ po_0.regf_0.rf\[4\]\[0\] po_0.regf_0.rf\[5\]\[0\] po_0.regf_0.rf\[6\]\[0\]
+ po_0.regf_0.rf\[7\]\[0\] _0414_ _0415_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux4_1
X_1777_ po_0.regf_0.rf\[0\]\[10\] po_0.regf_0.rf\[1\]\[10\] po_0.regf_0.rf\[2\]\[10\]
+ po_0.regf_0.rf\[3\]\[10\] _1497_ _1498_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__mux4_1
X_3516_ net120 _0300_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_3447_ net164 _0235_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfxtp_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ net152 _0166_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2329_ net4 _0701_ _0847_ _0793_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__a22o_2
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1700_ po_0.regf_0.rf\[8\]\[2\] po_0.regf_0.rf\[9\]\[2\] po_0.regf_0.rf\[10\]\[2\]
+ po_0.regf_0.rf\[11\]\[2\] _1488_ _1489_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__mux4_1
X_2680_ po_0.regf_0.rf\[11\]\[3\] _0935_ _1060_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__mux2_1
XFILLER_8_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1631_ _1432_ _1439_ _1440_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__o21bai_2
X_3301_ net116 _0089_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ po_0.regf_0._5_\[8\] net92 VGND VGND VPWR VPWR po_0._1_\[8\] sky130_fd_sc_hd__dlxtp_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _1388_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2114_ po_0._1_\[9\] _0650_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__or2b_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3094_ po_0.regf_0.rf\[2\]\[0\] _0713_ _1351_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__mux2_1
XFILLER_66_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2045_ _0587_ _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__nor2_1
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2947_ _1144_ _1255_ _1257_ _1258_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__a32o_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2878_ _1138_ _1155_ _1161_ _1172_ _1185_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__a41o_1
X_1829_ _0002_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__buf_2
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2801_ _1129_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__clkbuf_1
X_2732_ po_0.regf_0.rf\[10\]\[11\] _0952_ _1086_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__mux2_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2663_ _1054_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
X_2594_ _1016_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
X_1614_ _1426_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__clkbuf_1
X_3215_ net108 _0039_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3146_ uc_0._20_\[9\] po_0.regf_0.rp_addr\[1\] _0574_ VGND VGND VPWR VPWR _1378_
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3077_ _1342_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2028_ uc_0._20_\[9\] po_0.regf_0.rp_addr\[1\] _0575_ VGND VGND VPWR VPWR _0577_
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput7 D_R_data[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3000_ _1299_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2715_ po_0.regf_0.rf\[10\]\[3\] _0935_ _1079_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__mux2_1
X_2646_ _1045_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
X_2577_ _1007_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3129_ net92 _1311_ _0564_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__a21o_1
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3480_ net110 _0264_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2500_ _0965_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
X_2431_ _0920_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
X_2362_ net41 _0745_ _1402_ _0877_ _0729_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__o311a_1
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2293_ _0705_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__clkbuf_2
XFILLER_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_23 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2629_ _1035_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2980_ _1285_ _1283_ net67 VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__o21ai_1
X_1931_ _0492_ _0400_ _0424_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__a21o_1
X_1862_ _0422_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__clkbuf_2
Xinput10 D_R_data[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 I_data[13] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 I_data[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
X_1793_ _1453_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__and2b_1
X_3532_ net154 _0316_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[2\] sky130_fd_sc_hd__dfxtp_1
X_3463_ net162 _0247_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[7\] sky130_fd_sc_hd__dfxtp_1
X_2414_ _0911_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
X_3394_ net152 _0182_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2345_ _0661_ _0662_ _0673_ _0674_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__nor4_1
X_2276_ _0610_ _0798_ _0628_ _0633_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__nand4_2
XFILLER_37_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2130_ po_0._1_\[11\] VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__inv_2
X_2061_ _0604_ VGND VGND VPWR VPWR po_0.alu_0._10_\[3\] sky130_fd_sc_hd__clkbuf_1
X_2963_ _1269_ _1243_ _1264_ _1187_ _1273_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__a311oi_1
X_1914_ po_0.regf_0.rf\[0\]\[6\] po_0.regf_0.rf\[1\]\[6\] po_0.regf_0.rf\[2\]\[6\]
+ po_0.regf_0.rf\[3\]\[6\] _0405_ _0407_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__mux4_1
X_2894_ _1205_ _1206_ _1207_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__a211o_1
X_1845_ _0406_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__clkbuf_4
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1776_ _1511_ _0351_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__and2b_1
X_3515_ net116 _0299_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_3446_ net164 _0234_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfxtp_2
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ net174 _0165_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2328_ _0745_ po_0.alu_0._11_\[12\] _0815_ net83 _0846_ VGND VGND VPWR VPWR _0847_
+ sky130_fd_sc_hd__a221o_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2259_ _0719_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__buf_2
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1630_ net34 VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__clkbuf_2
X_3300_ net119 _0088_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ po_0.regf_0._5_\[7\] net92 VGND VGND VPWR VPWR po_0._1_\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _0715_ _1387_ _1372_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__mux2_1
XFILLER_66_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2113_ net50 VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__clkbuf_2
X_3093_ _1350_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__buf_2
XFILLER_66_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2044_ _0588_ po_0._1_\[2\] VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__nor2_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2946_ _1248_ _1246_ _1242_ _1256_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__a31o_1
X_2877_ _1189_ _1174_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__or2_1
X_1828_ po_0.regf_0.rf\[12\]\[0\] po_0.regf_0.rf\[13\]\[0\] po_0.regf_0.rf\[14\]\[0\]
+ po_0.regf_0.rf\[15\]\[0\] _0395_ _0397_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__mux4_1
X_1759_ po_0.regf_0.rf\[12\]\[8\] po_0.regf_0.rf\[13\]\[8\] po_0.regf_0.rf\[14\]\[8\]
+ po_0.regf_0.rf\[15\]\[8\] _1461_ _1463_ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__mux4_1
X_3429_ net151 _0217_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2800_ po_0.regf_0.rf\[8\]\[10\] _0829_ _1124_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__mux2_1
X_2731_ _1091_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2662_ po_0.regf_0.rf\[12\]\[11\] _0952_ _1048_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__mux2_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2593_ _0849_ po_0.regf_0.rf\[14\]\[12\] _1001_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__mux2_1
X_1613_ _1413_ _1415_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__or2b_1
X_3214_ net111 _0038_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3145_ _1377_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3076_ po_0.regf_0.rf\[3\]\[8\] _0810_ _1339_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__mux2_1
X_2027_ _0576_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2929_ _1241_ _1237_ _1226_ _1186_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__a31o_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 D_R_data[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2714_ _1082_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
X_2645_ po_0.regf_0.rf\[12\]\[3\] _0935_ _1041_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__mux2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2576_ _0763_ po_0.regf_0.rf\[14\]\[4\] _1002_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__mux2_1
XFILLER_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3128_ _1403_ _0561_ _0558_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a21bo_1
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3059_ po_0.regf_0.rf\[3\]\[0\] _0713_ _1332_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__mux2_1
XFILLER_42_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2430_ po_0.regf_0.rf\[5\]\[9\] _0820_ _0916_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__mux2_1
X_2361_ po_0.alu_0._11_\[15\] _0775_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__or2b_1
X_2292_ _0638_ _0653_ _0807_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__and3_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_13 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_24 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2628_ _0849_ po_0.regf_0.rf\[13\]\[12\] _1020_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__mux2_1
X_2559_ po_0.regf_0.rf\[15\]\[13\] _0956_ _0981_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__mux2_1
XFILLER_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1930_ po_0.regf_0.rf\[4\]\[8\] po_0.regf_0.rf\[5\]\[8\] po_0.regf_0.rf\[6\]\[8\]
+ po_0.regf_0.rf\[7\]\[8\] _0395_ _0397_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__mux4_1
X_1861_ po_0.regf_0.rf\[12\]\[1\] po_0.regf_0.rf\[13\]\[1\] po_0.regf_0.rf\[14\]\[1\]
+ po_0.regf_0.rf\[15\]\[1\] _0428_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux4_1
Xinput22 I_data[14] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 D_R_data[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput33 clock VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
X_1792_ po_0.regf_0.rf\[0\]\[12\] po_0.regf_0.rf\[1\]\[12\] po_0.regf_0.rf\[2\]\[12\]
+ po_0.regf_0.rf\[3\]\[12\] _1455_ _1457_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__mux4_1
X_3531_ net160 _0315_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[1\] sky130_fd_sc_hd__dfxtp_1
X_3462_ net162 _0246_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[6\] sky130_fd_sc_hd__dfxtp_1
X_2413_ po_0.regf_0.rf\[5\]\[1\] _0732_ _0909_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__mux2_1
X_3393_ net175 _0181_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2344_ _0843_ _0805_ _0656_ _0842_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2275_ _0614_ _0615_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__nor2_1
XFILLER_52_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2060_ _0601_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__and2_1
XFILLER_81_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2962_ _1243_ _1264_ _1269_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__a21oi_1
X_1913_ _0476_ _0400_ _0424_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__a21o_1
X_2893_ _1209_ _1210_ _1144_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__and3b_1
X_1844_ _0404_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__buf_4
X_1775_ po_0.regf_0.rf\[8\]\[10\] po_0.regf_0.rf\[9\]\[10\] po_0.regf_0.rf\[10\]\[10\]
+ po_0.regf_0.rf\[11\]\[10\] _1512_ _1513_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__mux4_1
X_3514_ net117 _0298_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_3445_ net164 _0233_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfxtp_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ net148 _0164_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2327_ _0661_ _0662_ _0844_ _0845_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__o31a_1
XFILLER_57_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2258_ _0782_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2189_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__buf_2
XFILLER_25_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ po_0.regf_0._5_\[6\] net94 VGND VGND VPWR VPWR po_0._1_\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ uc_0._20_\[11\] _0744_ _0562_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__mux2_1
XFILLER_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2112_ _0647_ _0648_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__nand2_1
X_3092_ _0886_ po_0.regf_0.w_addr\[3\] _0906_ _0885_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__and4bb_4
X_2043_ net43 VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2945_ _1248_ _1249_ _1256_ _1243_ _1186_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__a41oi_1
X_2876_ _1188_ _1191_ _1192_ _1175_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__a2bb2o_1
X_1827_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__buf_2
X_1758_ _1511_ _1555_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__and2b_1
X_1689_ _0004_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__clkbuf_4
X_3428_ net150 _0216_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_3359_ net140 _0147_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2730_ po_0.regf_0.rf\[10\]\[10\] _0950_ _1086_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__mux2_1
XFILLER_8_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2661_ _1053_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
X_1612_ _1425_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__clkbuf_1
X_2592_ _1015_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3213_ net135 _0037_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3144_ uc_0._20_\[8\] po_0.regf_0.rp_addr\[0\] _0575_ VGND VGND VPWR VPWR _1377_
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3075_ _1341_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2026_ uc_0._20_\[8\] po_0.regf_0.rp_addr\[0\] _0575_ VGND VGND VPWR VPWR _0576_
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2928_ _1242_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__clkbuf_2
X_2859_ _1150_ _1177_ _1178_ _1160_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__o31a_1
XFILLER_85_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput9 D_R_data[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2713_ po_0.regf_0.rf\[10\]\[2\] _0933_ _1079_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__mux2_1
X_2644_ _1044_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
X_2575_ _1006_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3127_ _0572_ _0559_ uc_0.bc_0._54_\[3\] _0558_ _1407_ VGND VGND VPWR VPWR _0305_
+ sky130_fd_sc_hd__a32o_1
X_3058_ _1331_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__buf_2
XFILLER_70_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2009_ _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__buf_2
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2360_ _0873_ _0758_ _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__nand3_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2291_ _0638_ _0807_ _0653_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_14 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2627_ _1034_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
X_2558_ _0996_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
X_2489_ _0870_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__clkbuf_2
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1860_ _0396_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__buf_2
Xinput12 D_R_data[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
X_1791_ _0364_ _1484_ _1492_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__a21o_1
Xinput23 I_data[15] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xinput34 reset VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
X_3530_ net160 _0314_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[0\] sky130_fd_sc_hd__dfxtp_1
X_3461_ net162 _0245_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[5\] sky130_fd_sc_hd__dfxtp_1
X_2412_ _0910_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
X_3392_ net148 _0180_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2343_ _0860_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
X_2274_ _0797_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1989_ _0494_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__and2b_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2961_ _1270_ _1145_ _1271_ _1207_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__a31o_1
X_1912_ po_0.regf_0.rf\[4\]\[6\] po_0.regf_0.rf\[5\]\[6\] po_0.regf_0.rf\[6\]\[6\]
+ po_0.regf_0.rf\[7\]\[6\] _0419_ _0420_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__mux4_1
X_2892_ _1172_ _1185_ _1166_ _1200_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__a31o_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1843_ po_0.regf_0.rf\[0\]\[0\] po_0.regf_0.rf\[1\]\[0\] po_0.regf_0.rf\[2\]\[0\]
+ po_0.regf_0.rf\[3\]\[0\] _0411_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux4_1
X_1774_ _0349_ _1470_ _1467_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__a21bo_1
X_3513_ net119 _0297_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_3444_ net164 _0232_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ net171 _0163_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2326_ _0844_ _0664_ _0708_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__a21oi_1
X_2257_ net13 _0700_ _0703_ _0568_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__a221o_4
XFILLER_84_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2188_ _0715_ _0716_ _0717_ _0718_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__nand4b_4
XFILLER_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _1386_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkbuf_1
X_3091_ _1349_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkbuf_1
X_2111_ po_0._1_\[10\] _0646_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__or2b_1
X_2042_ net43 po_0._1_\[2\] VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__and2_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2944_ _1248_ _1249_ _1256_ _1233_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__nand4_1
X_2875_ _1188_ _1191_ _1193_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__or3_1
X_1826_ _0001_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1757_ po_0.regf_0.rf\[0\]\[8\] po_0.regf_0.rf\[1\]\[8\] po_0.regf_0.rf\[2\]\[8\]
+ po_0.regf_0.rf\[3\]\[8\] _1512_ _1513_ VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__mux4_1
X_1688_ _1492_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__buf_2
X_3427_ net158 _0215_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3358_ net131 _0146_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _0829_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ net157 _0077_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2660_ po_0.regf_0.rf\[12\]\[10\] _0950_ _1048_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__mux2_1
XFILLER_8_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1611_ _1413_ _1415_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__or2b_1
X_2591_ _0839_ po_0.regf_0.rf\[14\]\[11\] _1009_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__mux2_1
XFILLER_5_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3212_ net135 _0036_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3143_ _1376_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3074_ po_0.regf_0.rf\[3\]\[7\] _0795_ _1339_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__mux2_1
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2025_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__buf_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2927_ net74 po_0.muxf_0.rf_w_data\[7\] _1241_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__o21a_1
X_2858_ net61 po_0.muxf_0.rf_w_data\[0\] _1151_ po_0.muxf_0.rf_w_data\[1\] VGND VGND
+ VPWR VPWR _1178_ sky130_fd_sc_hd__a22oi_4
X_1809_ _0380_ _1470_ _1467_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__a21bo_1
X_2789_ po_0.regf_0.rf\[8\]\[5\] _0772_ _1117_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__mux2_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2712_ _1081_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2643_ po_0.regf_0.rf\[12\]\[2\] _0933_ _1041_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__mux2_1
X_2574_ _0753_ po_0.regf_0.rf\[14\]\[3\] _1002_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__mux2_1
XFILLER_67_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3126_ _1368_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3057_ _0886_ po_0.regf_0.w_addr\[3\] _0906_ _0717_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__and4bb_4
XFILLER_63_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2008_ _0558_ _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__nand2_4
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2290_ _0812_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_15 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2626_ _0839_ po_0.regf_0.rf\[13\]\[11\] _1028_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__mux2_1
X_2557_ po_0.regf_0.rf\[15\]\[12\] _0954_ _0981_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__mux2_1
X_2488_ _0957_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3109_ po_0.regf_0.rf\[2\]\[7\] _0795_ _1358_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__mux2_1
XFILLER_43_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1790_ po_0.regf_0.rf\[4\]\[12\] po_0.regf_0.rf\[5\]\[12\] po_0.regf_0.rf\[6\]\[12\]
+ po_0.regf_0.rf\[7\]\[12\] _1542_ _1543_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__mux4_1
Xinput13 D_R_data[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput24 I_data[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
X_3460_ net177 _0244_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2411_ po_0.regf_0.rf\[5\]\[0\] _0714_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__mux2_1
X_3391_ net171 _0179_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2342_ _0859_ po_0.regf_0.rf\[7\]\[13\] _0719_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__mux2_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2273_ _0796_ po_0.regf_0.rf\[7\]\[7\] _0784_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__mux2_1
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1988_ po_0.regf_0.rf\[8\]\[14\] po_0.regf_0.rf\[9\]\[14\] po_0.regf_0.rf\[10\]\[14\]
+ po_0.regf_0.rf\[11\]\[14\] _0495_ _0496_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__mux4_1
X_2609_ _0753_ po_0.regf_0.rf\[13\]\[3\] _1021_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2960_ _1213_ _1225_ _1209_ _1263_ _1269_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__a41o_1
X_2891_ _1208_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__clkbuf_2
X_1911_ _0475_ VGND VGND VPWR VPWR po_0.regf_0._3_\[5\] sky130_fd_sc_hd__clkbuf_1
X_1842_ _0406_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__buf_2
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1773_ po_0.regf_0.rf\[12\]\[10\] po_0.regf_0.rf\[13\]\[10\] po_0.regf_0.rf\[14\]\[10\]
+ po_0.regf_0.rf\[15\]\[10\] _1481_ _1482_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__mux4_1
X_3512_ net123 _0296_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3443_ net163 _0231_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfxtp_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ net173 _0162_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ _0656_ _0842_ _0843_ _0805_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__a2bb2oi_1
X_2256_ _0776_ _0780_ _0729_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__o21a_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2187_ po_0.regf_0.w_addr\[2\] VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__clkbuf_2
XFILLER_65_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3090_ po_0.regf_0.rf\[3\]\[15\] _0879_ _1331_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__mux2_1
XFILLER_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2110_ _0646_ po_0._1_\[10\] VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__or2b_1
X_2041_ po_0._1_\[1\] _0584_ _0580_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2943_ net62 VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__clkbuf_2
XFILLER_62_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2874_ _1172_ _0744_ _1192_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__o21ai_1
X_1825_ _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__clkbuf_4
X_1756_ _1553_ _1484_ _1492_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__a21o_1
X_1687_ _0007_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__clkbuf_2
X_3426_ net156 _0214_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3357_ net145 _0145_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ net2 _0701_ _0828_ _0793_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__a22o_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3288_ net170 _0076_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2239_ _0605_ po_0._1_\[4\] VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__nand2_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1610_ _1424_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__clkbuf_1
X_2590_ _1014_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3211_ net127 _0035_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3142_ po_0.regf_0.rq_addr\[3\] _0570_ _0563_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__mux2_1
XFILLER_39_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3073_ _1340_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2024_ _0572_ _1447_ _0573_ _0562_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__a31oi_4
XFILLER_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2926_ _1219_ _1223_ _1227_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__nand3_2
X_2857_ net69 po_0.muxf_0.rf_w_data\[2\] VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__nor2_1
X_1808_ po_0.regf_0.rf\[12\]\[14\] po_0.regf_0.rf\[13\]\[14\] po_0.regf_0.rf\[14\]\[14\]
+ po_0.regf_0.rf\[15\]\[14\] _1481_ _1482_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__mux4_1
X_2788_ _1122_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1739_ po_0.regf_0.rf\[0\]\[6\] po_0.regf_0.rf\[1\]\[6\] po_0.regf_0.rf\[2\]\[6\]
+ po_0.regf_0.rf\[3\]\[6\] _1494_ _1495_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__mux4_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3409_ net138 _0197_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2711_ po_0.regf_0.rf\[10\]\[1\] _0931_ _1079_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__mux2_1
X_2642_ _1043_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
X_2573_ _1005_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3125_ po_0.regf_0.rf\[2\]\[15\] _0879_ _1350_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__mux2_1
XFILLER_67_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3056_ _1330_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2007_ _1440_ uc_0.bc_0._54_\[1\] _0559_ _0560_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__or4bb_2
XFILLER_23_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2909_ net74 VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__clkbuf_2
XFILLER_58_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_16 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2625_ _1033_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
X_2556_ _0995_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
X_2487_ po_0.regf_0.rf\[9\]\[13\] _0956_ _0928_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__mux2_1
X_3108_ _1359_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3039_ po_0.regf_0.rf\[4\]\[7\] _0795_ _1320_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__mux2_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput14 D_R_data[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
Xinput25 I_data[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
XFILLER_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2410_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__buf_2
X_3390_ net171 _0178_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2341_ _0858_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2272_ _0795_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1987_ _0542_ _0447_ _0003_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__a21bo_1
X_2608_ _1024_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
X_2539_ _0986_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout180 net181 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2890_ net99 _1185_ _1200_ _1166_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__and4_1
X_1910_ _0471_ _0474_ _0445_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__mux2_1
XFILLER_30_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1841_ _0404_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__clkbuf_4
X_1772_ _0342_ _0344_ _0346_ _0348_ VGND VGND VPWR VPWR po_0.regf_0._5_\[9\] sky130_fd_sc_hd__o22a_1
X_3511_ net122 _0295_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3442_ net162 _0230_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfxtp_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ net174 _0161_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _0668_ _0643_ _0649_ _0658_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__and4_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ _0778_ _0628_ _1401_ _0779_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__o211a_1
X_2186_ po_0.regf_0.w_addr\[1\] po_0.regf_0.w_addr\[0\] VGND VGND VPWR VPWR _0717_
+ sky130_fd_sc_hd__and2_1
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2040_ _0584_ po_0._1_\[1\] VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__nand2_1
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2942_ net97 _1246_ _1233_ net62 VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__a31o_1
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2873_ _1150_ _1177_ _1178_ _1176_ _1160_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__o311ai_4
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1824_ _0000_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__clkbuf_2
X_1755_ po_0.regf_0.rf\[4\]\[8\] po_0.regf_0.rf\[5\]\[8\] po_0.regf_0.rf\[6\]\[8\]
+ po_0.regf_0.rf\[7\]\[8\] _1542_ _1543_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__mux4_1
X_1686_ _1487_ _1490_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__and2b_1
X_3425_ net175 _0213_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3356_ net144 _0144_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3287_ net120 _0075_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _0824_ _0708_ _0826_ _0827_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__o31ai_1
X_2238_ _0764_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2169_ _0699_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__buf_2
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3210_ net127 _0034_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3141_ _1375_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__clkbuf_1
X_3072_ po_0.regf_0.rf\[3\]\[6\] _0782_ _1339_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__mux2_1
XFILLER_54_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2023_ uc_0.bc_0._54_\[3\] uc_0.bc_0._54_\[2\] VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__or2_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2925_ _1238_ _1145_ _1239_ _1207_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__a31o_1
X_2856_ net99 po_0.muxf_0.rf_w_data\[3\] VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__nand2_1
X_1807_ _0373_ _0375_ _0377_ _0379_ VGND VGND VPWR VPWR po_0.regf_0._5_\[13\] sky130_fd_sc_hd__o22a_1
X_2787_ po_0.regf_0.rf\[8\]\[4\] _0762_ _1117_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__mux2_1
X_1738_ _1511_ _1537_ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__and2b_1
X_1669_ _1460_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__clkbuf_4
X_3408_ net137 _0196_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3339_ net128 _0127_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2710_ _1080_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__clkbuf_1
X_2641_ po_0.regf_0.rf\[12\]\[1\] _0931_ _1041_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__mux2_1
X_2572_ _0742_ po_0.regf_0.rf\[14\]\[2\] _1002_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__mux2_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3124_ _1367_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3055_ po_0.regf_0.rf\[4\]\[15\] _0879_ _1312_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__mux2_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2006_ _1439_ _1449_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__or2_1
X_2908_ _1213_ _1215_ _1218_ _1224_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__o22a_1
X_2839_ net69 _0734_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__nand2_2
XFILLER_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_17 _0423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2624_ _0830_ po_0.regf_0.rf\[13\]\[10\] _1028_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__mux2_1
X_2555_ po_0.regf_0.rf\[15\]\[11\] _0952_ _0989_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__mux2_1
X_2486_ _0858_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__clkbuf_2
XFILLER_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3107_ po_0.regf_0.rf\[2\]\[6\] _0782_ _1358_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__mux2_1
X_3038_ _1321_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 I_data[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput15 D_R_data[8] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2340_ net5 _0701_ _0851_ _0857_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__o2bb2ai_4
X_2271_ _0791_ _0792_ _0793_ _0794_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a31o_2
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1986_ po_0.regf_0.rf\[12\]\[14\] po_0.regf_0.rf\[13\]\[14\] po_0.regf_0.rf\[14\]\[14\]
+ po_0.regf_0.rf\[15\]\[14\] _0435_ _0436_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__mux4_1
X_2607_ _0742_ po_0.regf_0.rf\[13\]\[2\] _1021_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__mux2_1
X_2538_ po_0.regf_0.rf\[15\]\[3\] _0935_ _0982_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__mux2_1
X_2469_ po_0.regf_0.rf\[9\]\[7\] _0944_ _0942_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__mux2_1
XFILLER_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout181 net182 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
Xfanout170 net172 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1840_ _0003_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__buf_2
XFILLER_30_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3510_ net146 _0294_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1771_ _1550_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__and2b_1
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3441_ net162 _0229_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfxtp_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3372_ net173 _0160_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _0822_ _0823_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__o21ba_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _0778_ _0628_ _1404_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__a21oi_1
X_2185_ po_0.regf_0.w_wr VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__clkbuf_2
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1969_ _0417_ _0526_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__and2b_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2941_ _1254_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__clkbuf_1
X_2872_ _1189_ _1190_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__nor2_1
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1823_ _0388_ _0390_ _1479_ _0393_ VGND VGND VPWR VPWR po_0.regf_0._5_\[15\] sky130_fd_sc_hd__o22a_1
X_1754_ _1545_ _1547_ _1549_ _1552_ VGND VGND VPWR VPWR po_0.regf_0._5_\[7\] sky130_fd_sc_hd__o22a_1
X_1685_ po_0.regf_0.rf\[8\]\[1\] po_0.regf_0.rf\[9\]\[1\] po_0.regf_0.rf\[10\]\[1\]
+ po_0.regf_0.rf\[11\]\[1\] _1488_ _1489_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__mux4_1
X_3424_ net174 _0212_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3355_ net128 _0143_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ net152 _0074_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _0745_ po_0.alu_0._11_\[10\] _0815_ _0646_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__a22oi_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ _0763_ po_0.regf_0.rf\[7\]\[4\] _0720_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__mux2_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2168_ _0698_ po_0.muxf_0.s0 VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__and2_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2099_ _0637_ po_0._1_\[8\] VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__nand2_1
XFILLER_80_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3140_ po_0.regf_0.rq_addr\[2\] _0568_ _0563_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__mux2_1
XFILLER_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3071_ _1331_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__buf_2
X_2022_ _1441_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__buf_2
X_2924_ _1213_ _1225_ _1209_ _1237_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__a31o_1
X_2855_ net99 _0744_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__or2_1
X_1806_ _0378_ _1478_ _1479_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__a21o_1
X_2786_ _1121_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__clkbuf_1
X_1737_ po_0.regf_0.rf\[8\]\[6\] po_0.regf_0.rf\[9\]\[6\] po_0.regf_0.rf\[10\]\[6\]
+ po_0.regf_0.rf\[11\]\[6\] _1512_ _1513_ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__mux4_1
X_1668_ _1470_ _1473_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__and2b_1
X_3407_ net130 _0195_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3338_ net113 _0126_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1599_ _1414_ _1416_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__or2b_1
XFILLER_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ net110 _0061_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2640_ _1042_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2571_ _1004_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3123_ po_0.regf_0.rf\[2\]\[14\] _0870_ _1350_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__mux2_1
X_3054_ _1329_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2005_ _1446_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__clkbuf_2
XFILLER_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2907_ _1222_ _1142_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__and3_1
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2838_ _1159_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__clkbuf_1
X_2769_ _0849_ po_0.regf_0.rf\[0\]\[12\] _1097_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__mux2_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 _0704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2623_ _1032_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
X_2554_ _0994_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
X_2485_ _0955_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
X_3106_ _1350_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__buf_2
X_3037_ po_0.regf_0.rf\[4\]\[6\] _0782_ _1320_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__mux2_1
XFILLER_23_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput16 D_R_data[9] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 I_data[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2270_ net14 _0700_ _0703_ _0570_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__a22o_1
XFILLER_77_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1985_ _0535_ _0537_ _0539_ _0541_ VGND VGND VPWR VPWR po_0.regf_0._3_\[13\] sky130_fd_sc_hd__o22a_1
X_2606_ _1023_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
X_2537_ _0985_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
X_2468_ _0795_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__clkbuf_2
X_2399_ po_0.regf_0.rf\[6\]\[12\] _0849_ _0887_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__mux2_1
XFILLER_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout182 net183 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout171 net172 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout160 net161 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1770_ po_0.regf_0.rf\[8\]\[9\] po_0.regf_0.rf\[9\]\[9\] po_0.regf_0.rf\[10\]\[9\]
+ po_0.regf_0.rf\[11\]\[9\] _1471_ _1472_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__mux4_1
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3440_ net167 _0228_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfxtp_2
X_3371_ net141 _0159_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2322_ _0646_ po_0._1_\[10\] po_0._1_\[11\] net84 VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__a22o_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2253_ _0777_ _0757_ po_0._1_\[5\] _0613_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_77_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2184_ po_0.regf_0.w_addr\[3\] VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1968_ po_0.regf_0.rf\[8\]\[12\] po_0.regf_0.rf\[9\]\[12\] po_0.regf_0.rf\[10\]\[12\]
+ po_0.regf_0.rf\[11\]\[12\] _0411_ _0412_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__mux4_1
X_1899_ po_0.regf_0.rf\[12\]\[4\] po_0.regf_0.rf\[13\]\[4\] po_0.regf_0.rf\[14\]\[4\]
+ po_0.regf_0.rf\[15\]\[4\] _0428_ _0429_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__mux4_1
X_3569_ po_0.alu_0._10_\[10\] _1568_ VGND VGND VPWR VPWR po_0.alu_0._11_\[10\] sky130_fd_sc_hd__ebufn_1
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2940_ _1253_ _1249_ _1148_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__mux2_1
XFILLER_15_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2871_ po_0.muxf_0.rf_w_data\[4\] VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__inv_2
X_1822_ _0391_ _0392_ _1465_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__mux2_1
X_1753_ _1550_ _1551_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__and2b_1
X_1684_ _1456_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__buf_2
X_3423_ net171 _0211_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ net128 _0142_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3285_ net150 _0073_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _0825_ _0648_ _0647_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__and3_1
X_2236_ _0762_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2167_ po_0.muxf_0.s1 VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__inv_2
X_2098_ net49 VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__clkbuf_2
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3070_ _1338_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2021_ _0571_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2923_ _1237_ _1234_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__nand2_1
X_2854_ net99 _1166_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nand2_1
X_1805_ po_0.regf_0.rf\[4\]\[13\] po_0.regf_0.rf\[5\]\[13\] po_0.regf_0.rf\[6\]\[13\]
+ po_0.regf_0.rf\[7\]\[13\] _1475_ _1476_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__mux4_1
X_2785_ po_0.regf_0.rf\[8\]\[3\] _0752_ _1117_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__mux2_1
X_1736_ _1535_ _1470_ _1485_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__a21bo_1
X_1667_ po_0.regf_0.rf\[0\]\[0\] po_0.regf_0.rf\[1\]\[0\] po_0.regf_0.rf\[2\]\[0\]
+ po_0.regf_0.rf\[3\]\[0\] _1471_ _1472_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__mux4_1
X_3406_ net130 _0194_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_1598_ _1418_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__clkbuf_1
X_3337_ net113 _0125_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ net109 _0060_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3199_ net108 _0023_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2219_ _0587_ _0602_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__or3_1
XFILLER_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2570_ _0732_ po_0.regf_0.rf\[14\]\[1\] _1002_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__mux2_1
X_3122_ _1366_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3053_ po_0.regf_0.rf\[4\]\[14\] _0870_ _1312_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__mux2_1
XFILLER_48_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2004_ _1441_ _1451_ _1447_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__or3_2
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2906_ _1200_ po_0.muxf_0.rf_w_data\[5\] _1219_ _1220_ _1221_ VGND VGND VPWR VPWR
+ _1223_ sky130_fd_sc_hd__o2111ai_2
X_2837_ _1158_ _1155_ _1148_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__mux2_1
X_2768_ _1111_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__clkbuf_1
X_1719_ po_0.regf_0.rf\[12\]\[4\] po_0.regf_0.rf\[13\]\[4\] po_0.regf_0.rf\[14\]\[4\]
+ po_0.regf_0.rf\[15\]\[4\] _1461_ _1463_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__mux4_1
X_2699_ po_0.regf_0.rf\[11\]\[12\] _0954_ _1059_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__mux2_1
XFILLER_58_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 _0795_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2622_ _0820_ po_0.regf_0.rf\[13\]\[9\] _1028_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__mux2_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2553_ po_0.regf_0.rf\[15\]\[10\] _0950_ _0989_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__mux2_1
X_2484_ po_0.regf_0.rf\[9\]\[12\] _0954_ _0928_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__mux2_1
XFILLER_28_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3105_ _1357_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__clkbuf_1
X_3036_ _1312_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__buf_2
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput17 I_data[0] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 I_data[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1984_ _0423_ _0540_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__and2b_1
X_2605_ _0732_ po_0.regf_0.rf\[13\]\[1\] _1021_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__mux2_1
X_2536_ po_0.regf_0.rf\[15\]\[2\] _0933_ _0982_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__mux2_1
X_2467_ _0943_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
X_2398_ _0901_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3019_ _1308_ _1309_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__nor2_1
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout183 net33 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_2
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout150 net152 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout172 net182 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout161 net169 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3370_ net140 _0158_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _0840_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2252_ _0605_ po_0._1_\[4\] po_0._1_\[5\] _0613_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__a22oi_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2183_ _0713_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1967_ _0519_ _0521_ _0523_ _0525_ VGND VGND VPWR VPWR po_0.regf_0._3_\[11\] sky130_fd_sc_hd__o22a_1
X_1898_ _0403_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__and2b_1
X_3568_ po_0.alu_0._10_\[9\] _1567_ VGND VGND VPWR VPWR po_0.alu_0._11_\[9\] sky130_fd_sc_hd__ebufn_1
X_2519_ _0975_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3499_ net118 _0283_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2870_ net71 VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__inv_2
X_1821_ po_0.regf_0.rf\[4\]\[15\] po_0.regf_0.rf\[5\]\[15\] po_0.regf_0.rf\[6\]\[15\]
+ po_0.regf_0.rf\[7\]\[15\] _1460_ _1462_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__mux4_1
X_1752_ po_0.regf_0.rf\[8\]\[7\] po_0.regf_0.rf\[9\]\[7\] po_0.regf_0.rf\[10\]\[7\]
+ po_0.regf_0.rf\[11\]\[7\] _1471_ _1472_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__mux4_1
X_1683_ _1454_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__clkbuf_4
X_3422_ net176 _0210_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ net113 _0141_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ net119 _0072_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _0650_ po_0._1_\[9\] _0822_ _0807_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2235_ _0722_ _0723_ net11 _0761_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__a31o_2
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2166_ _0695_ _0697_ VGND VGND VPWR VPWR po_0.alu_0._10_\[15\] sky130_fd_sc_hd__nand2_1
XFILLER_65_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2097_ _0636_ VGND VGND VPWR VPWR po_0.alu_0._10_\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_80_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2999_ _0570_ net30 _1296_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__mux2_1
XFILLER_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2020_ po_0.regf_0.rq_addr\[3\] _0570_ _0564_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__mux2_1
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2922_ net97 VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__clkbuf_2
X_2853_ _1138_ _1155_ _1161_ _1172_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__a31o_1
X_1804_ _1487_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__and2b_1
X_2784_ _1120_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__clkbuf_1
X_1735_ po_0.regf_0.rf\[12\]\[6\] po_0.regf_0.rf\[13\]\[6\] po_0.regf_0.rf\[14\]\[6\]
+ po_0.regf_0.rf\[15\]\[6\] _1481_ _1482_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__mux4_1
X_1666_ _1456_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__clkbuf_4
X_3405_ net136 _0193_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1597_ _1414_ _1416_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__or2b_1
X_3336_ net129 _0124_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3267_ net101 _0059_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3198_ net108 _0022_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2218_ _0592_ _0593_ _0736_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__o21a_1
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2149_ _0680_ po_0._1_\[14\] VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__or2_1
XFILLER_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3121_ po_0.regf_0.rf\[2\]\[13\] _0858_ _1350_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__mux2_1
X_3052_ _1328_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__clkbuf_1
X_2003_ po_0.muxf_0.rf_w_data\[4\] VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__buf_2
XFILLER_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2905_ _1219_ _1220_ _1221_ _1204_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__a22o_1
X_2836_ _1153_ _1142_ _1154_ _1157_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__a31o_1
X_2767_ _0839_ po_0.regf_0.rf\[0\]\[11\] _1105_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__mux2_1
X_1718_ _1453_ _1519_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__and2b_1
X_2698_ _1073_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__clkbuf_1
X_1649_ _1454_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__clkbuf_4
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3319_ net105 _0107_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2621_ _1031_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
X_2552_ _0993_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
X_2483_ _0848_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__clkbuf_2
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3104_ po_0.regf_0.rf\[2\]\[5\] _0772_ _1351_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__mux2_1
X_3035_ _1319_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2819_ _1141_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__clkbuf_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 I_data[10] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 I_data[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1983_ po_0.regf_0.rf\[8\]\[13\] po_0.regf_0.rf\[9\]\[13\] po_0.regf_0.rf\[10\]\[13\]
+ po_0.regf_0.rf\[11\]\[13\] _0448_ _0449_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__mux4_1
X_2604_ _1022_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
X_2535_ _0984_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
X_2466_ po_0.regf_0.rf\[9\]\[6\] _0941_ _0942_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__mux2_1
X_2397_ po_0.regf_0.rf\[6\]\[11\] _0839_ _0895_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__mux2_1
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3018_ _0572_ uc_0.bc_0._54_\[0\] uc_0.bc_0._54_\[3\] uc_0.bc_0._54_\[2\] VGND VGND
+ VPWR VPWR _1309_ sky130_fd_sc_hd__nor4_1
XFILLER_43_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout140 net143 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout173 net176 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout151 net152 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
Xfanout162 net163 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _0839_ po_0.regf_0.rf\[7\]\[11\] _0784_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__mux2_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ _0775_ po_0.alu_0._11_\[6\] _0706_ _0620_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__a22o_1
X_2182_ net1 _0701_ _0703_ _0704_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__a221o_2
XFILLER_65_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1966_ _0423_ _0524_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__and2b_1
X_1897_ po_0.regf_0.rf\[0\]\[4\] po_0.regf_0.rf\[1\]\[4\] po_0.regf_0.rf\[2\]\[4\]
+ po_0.regf_0.rf\[3\]\[4\] _0405_ _0407_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__mux4_1
X_3567_ po_0.alu_0._10_\[8\] _1566_ VGND VGND VPWR VPWR po_0.alu_0._11_\[8\] sky130_fd_sc_hd__ebufn_1
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2518_ po_0.regf_0.rf\[1\]\[10\] _0950_ _0970_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3498_ net117 _0282_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_2449_ _0731_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__clkbuf_2
XFILLER_83_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1820_ po_0.regf_0.rf\[0\]\[15\] po_0.regf_0.rf\[1\]\[15\] po_0.regf_0.rf\[2\]\[15\]
+ po_0.regf_0.rf\[3\]\[15\] _1497_ _1498_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__mux4_1
XFILLER_30_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1751_ _1465_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__clkbuf_2
X_1682_ _1452_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__clkbuf_2
X_3421_ net174 _0209_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3352_ net128 _0140_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _0807_ _0822_ _0823_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__a21oi_1
X_3283_ net158 _0071_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _0557_ _0702_ _0760_ _0729_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__a22o_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ _0689_ _0690_ _0696_ _0686_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__o22ai_1
XFILLER_80_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2096_ _0634_ _0635_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__and2_1
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2998_ _1298_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__clkbuf_1
X_1949_ _0504_ _0506_ _0410_ _0509_ VGND VGND VPWR VPWR po_0.regf_0._3_\[9\] sky130_fd_sc_hd__o22a_1
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2921_ _1135_ _1225_ _1187_ _1236_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__o31a_1
X_2852_ net99 VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__clkbuf_2
X_1803_ po_0.regf_0.rf\[0\]\[13\] po_0.regf_0.rf\[1\]\[13\] po_0.regf_0.rf\[2\]\[13\]
+ po_0.regf_0.rf\[3\]\[13\] _1488_ _1489_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__mux4_1
X_2783_ po_0.regf_0.rf\[8\]\[2\] _0741_ _1117_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__mux2_1
X_1734_ _1528_ _1530_ _1532_ _1534_ VGND VGND VPWR VPWR po_0.regf_0._5_\[5\] sky130_fd_sc_hd__o22a_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3404_ net136 _0192_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1665_ _1454_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__clkbuf_4
X_1596_ _1417_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__clkbuf_1
X_3335_ net105 _0123_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3266_ net100 _0058_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _1405_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__clkbuf_2
X_3197_ net135 _0021_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2148_ _0680_ po_0._1_\[14\] VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__nand2_1
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2079_ net47 VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3120_ _1365_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__clkbuf_1
X_3051_ po_0.regf_0.rf\[4\]\[13\] _0858_ _1312_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__mux2_1
X_2002_ _0550_ _0552_ _0554_ _0556_ VGND VGND VPWR VPWR po_0.regf_0._3_\[15\] sky130_fd_sc_hd__o22a_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2904_ _1189_ _1190_ _1203_ _1201_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__o211ai_2
X_2835_ _1138_ _1155_ _1156_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__a21oi_1
X_2766_ _1110_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__clkbuf_1
X_2697_ po_0.regf_0.rf\[11\]\[11\] _0952_ _1067_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__mux2_1
X_1717_ po_0.regf_0.rf\[8\]\[4\] po_0.regf_0.rf\[9\]\[4\] po_0.regf_0.rf\[10\]\[4\]
+ po_0.regf_0.rf\[11\]\[4\] _1455_ _1457_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__mux4_1
X_1648_ _0004_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__clkbuf_2
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ net116 _0106_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_1579_ _1405_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__clkbuf_2
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3249_ po_0.regf_0._3_\[9\] net88 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlxtp_1
XFILLER_73_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2620_ _0811_ po_0.regf_0.rf\[13\]\[8\] _1028_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__mux2_1
X_2551_ po_0.regf_0.rf\[15\]\[9\] _0948_ _0989_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__mux2_1
X_2482_ _0953_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3103_ _1356_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3034_ po_0.regf_0.rf\[4\]\[5\] _0772_ _1313_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__mux2_1
XFILLER_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2818_ _1139_ _1140_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__nor2_1
X_2749_ _1101_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__clkbuf_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput19 I_data[11] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1982_ _0538_ _0444_ _0445_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__a21bo_1
X_2603_ _0714_ po_0.regf_0.rf\[13\]\[0\] _1021_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__mux2_1
X_2534_ po_0.regf_0.rf\[15\]\[1\] _0931_ _0982_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__mux2_1
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2465_ _0928_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__buf_2
X_2396_ _0900_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3017_ _0559_ uc_0.bc_0._54_\[3\] uc_0.bc_0._54_\[2\] uc_0.bc_0._54_\[1\] VGND VGND
+ VPWR VPWR _1308_ sky130_fd_sc_hd__nor4_1
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout130 net132 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
Xfanout141 net143 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
Xfanout152 net156 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout174 net175 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
Xfanout163 net165 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _1404_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__clkbuf_2
X_2181_ _0706_ _0709_ _0710_ _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__o211a_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1965_ po_0.regf_0.rf\[8\]\[11\] po_0.regf_0.rf\[9\]\[11\] po_0.regf_0.rf\[10\]\[11\]
+ po_0.regf_0.rf\[11\]\[11\] _0448_ _0449_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__mux4_1
X_1896_ _0461_ _0423_ _0424_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__a21o_1
X_3566_ po_0.alu_0._10_\[7\] _1565_ VGND VGND VPWR VPWR po_0.alu_0._11_\[7\] sky130_fd_sc_hd__ebufn_1
X_2517_ _0974_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
X_3497_ net119 _0281_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_2448_ _0930_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2379_ _0891_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1750_ _1548_ _1478_ _1492_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__a21bo_1
XFILLER_11_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1681_ _1483_ _1484_ _1485_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__a21bo_1
X_3420_ net176 _0208_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3351_ net105 _0139_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2302_ _0650_ po_0._1_\[9\] _0647_ _0648_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__a2bb2o_1
X_3282_ net152 _0070_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _1405_ po_0.alu_0._11_\[4\] _0705_ _0605_ _0759_ VGND VGND VPWR VPWR _0760_
+ sky130_fd_sc_hd__a221o_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2164_ po_0._1_\[14\] _0688_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__nor2_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2095_ _0630_ _0625_ _0631_ _0632_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__or4_1
X_2997_ _0568_ net29 _1296_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__mux2_1
X_1948_ _0507_ _0508_ _0422_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__mux2_1
X_1879_ _0399_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__buf_2
X_3549_ net100 _0333_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2920_ _1230_ _1231_ _1235_ _1215_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__o211ai_1
X_2851_ _1140_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1802_ _0374_ _1550_ _1485_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__a21bo_1
X_2782_ _1119_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__clkbuf_1
X_1733_ _1533_ _1478_ _1479_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__a21o_1
X_1664_ _1452_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__buf_2
X_3403_ net170 _0191_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_1595_ _1414_ _1416_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__or2b_1
X_3334_ net103 _0122_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3265_ net102 _0057_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ po_0.muxf_0.rf_w_data\[3\] VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ net135 _0020_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2147_ net40 VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__clkbuf_2
X_2078_ _0619_ VGND VGND VPWR VPWR po_0.alu_0._10_\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3050_ _1327_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__clkbuf_1
X_2001_ _0555_ _0431_ _0424_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__a21o_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2903_ net98 po_0.muxf_0.rf_w_data\[6\] VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__or2_1
X_2834_ _1138_ _1155_ _1140_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__o21ai_1
X_2765_ _0830_ po_0.regf_0.rf\[0\]\[10\] _1105_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__mux2_1
X_1716_ _1510_ _1515_ _1493_ _1518_ VGND VGND VPWR VPWR po_0.regf_0._5_\[3\] sky130_fd_sc_hd__o22a_1
X_2696_ _1072_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__clkbuf_1
X_1647_ _1452_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__clkbuf_2
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ net116 _0105_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_1578_ _1404_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__clkbuf_2
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ po_0.regf_0._3_\[8\] net88 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlxtp_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3179_ _0557_ net55 _1393_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__mux2_1
XFILLER_73_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2550_ _0992_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_2481_ po_0.regf_0.rf\[9\]\[11\] _0952_ _0942_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__mux2_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3102_ po_0.regf_0.rf\[2\]\[4\] _0762_ _1351_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__mux2_1
X_3033_ _1318_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2817_ uc_0._02_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__clkbuf_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2748_ _0742_ po_0.regf_0.rf\[0\]\[2\] _1098_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__mux2_1
X_2679_ _1063_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1981_ po_0.regf_0.rf\[12\]\[13\] po_0.regf_0.rf\[13\]\[13\] po_0.regf_0.rf\[14\]\[13\]
+ po_0.regf_0.rf\[15\]\[13\] _0441_ _0442_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__mux4_1
XFILLER_9_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2602_ _1020_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__buf_2
X_2533_ _0983_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
X_2464_ _0782_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__clkbuf_2
X_2395_ po_0.regf_0.rf\[6\]\[10\] _0830_ _0895_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__mux2_1
XFILLER_56_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3016_ _1307_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout131 net132 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
Xfanout120 net121 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout164 net165 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
Xfanout142 net143 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout153 net155 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout175 net176 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
XFILLER_74_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2180_ _0699_ _0702_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__nor2_1
XFILLER_38_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1964_ _0522_ _0444_ _0445_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__a21bo_1
X_1895_ po_0.regf_0.rf\[4\]\[4\] po_0.regf_0.rf\[5\]\[4\] po_0.regf_0.rf\[6\]\[4\]
+ po_0.regf_0.rf\[7\]\[4\] _0419_ _0420_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__mux4_1
X_3565_ po_0.alu_0._10_\[6\] _1564_ VGND VGND VPWR VPWR po_0.alu_0._11_\[6\] sky130_fd_sc_hd__ebufn_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2516_ po_0.regf_0.rf\[1\]\[9\] _0948_ _0970_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__mux2_1
X_3496_ net123 _0280_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2447_ po_0.regf_0.rf\[9\]\[0\] _0927_ _0929_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__mux2_1
X_2378_ po_0.regf_0.rf\[6\]\[2\] _0742_ _0888_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__mux2_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1680_ _1467_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__clkbuf_2
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3350_ net106 _0138_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ _0637_ po_0._1_\[8\] po_0._1_\[9\] _0650_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__a22oi_2
X_3281_ net174 _0069_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ _0610_ _0756_ _0757_ _0758_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__o211a_1
X_2163_ _0688_ po_0._1_\[14\] _0691_ _0694_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__o211ai_1
XFILLER_65_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2094_ _0630_ _0625_ _0633_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__o21bai_2
XFILLER_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2996_ _1297_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__clkbuf_1
X_1947_ po_0.regf_0.rf\[4\]\[9\] po_0.regf_0.rf\[5\]\[9\] po_0.regf_0.rf\[6\]\[9\]
+ po_0.regf_0.rf\[7\]\[9\] _0414_ _0415_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__mux4_1
X_1878_ _0443_ _0444_ _0445_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__a21bo_1
X_3548_ net153 _0332_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfxtp_1
X_3479_ net111 _0263_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2850_ _1170_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1801_ po_0.regf_0.rf\[12\]\[13\] po_0.regf_0.rf\[13\]\[13\] po_0.regf_0.rf\[14\]\[13\]
+ po_0.regf_0.rf\[15\]\[13\] _1542_ _1543_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__mux4_1
X_2781_ po_0.regf_0.rf\[8\]\[1\] _0731_ _1117_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__mux2_1
X_1732_ po_0.regf_0.rf\[4\]\[5\] po_0.regf_0.rf\[5\]\[5\] po_0.regf_0.rf\[6\]\[5\]
+ po_0.regf_0.rf\[7\]\[5\] _1475_ _1476_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__mux4_1
X_1663_ _1464_ _1466_ _1468_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__a21bo_1
X_3402_ net157 _0190_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _1415_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__dlymetal6s2s_1
X_3333_ net103 _0121_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ net102 _0056_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2215_ _0743_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ net127 _0019_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2146_ _0672_ po_0._1_\[12\] _0675_ _0677_ _0679_ VGND VGND VPWR VPWR po_0.alu_0._10_\[13\]
+ sky130_fd_sc_hd__o311a_1
XFILLER_66_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2077_ _0617_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__and2_1
X_2979_ net66 _1142_ _1276_ _1282_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__a31oi_1
XFILLER_57_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2000_ po_0.regf_0.rf\[4\]\[15\] po_0.regf_0.rf\[5\]\[15\] po_0.regf_0.rf\[6\]\[15\]
+ po_0.regf_0.rf\[7\]\[15\] _0428_ _0429_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__mux4_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2902_ net98 po_0.muxf_0.rf_w_data\[6\] VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__nand2_1
X_2833_ _1151_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__clkbuf_2
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2764_ _1109_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__clkbuf_1
X_1715_ _1516_ _1517_ _1500_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__mux2_1
X_2695_ po_0.regf_0.rf\[11\]\[10\] _0950_ _1067_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__mux2_1
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1646_ _0006_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1577_ po_0.alu_0.s1 VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__clkbuf_2
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ net103 _0104_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ po_0.regf_0._3_\[7\] net88 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlxtp_1
X_3178_ _1395_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2129_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2480_ _0838_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__clkbuf_2
X_3101_ _1355_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_1
X_3032_ po_0.regf_0.rf\[4\]\[4\] _0762_ _1313_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__mux2_1
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2816_ uc_0._00_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__clkbuf_2
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2747_ _1100_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2678_ po_0.regf_0.rf\[11\]\[2\] _0933_ _1060_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__mux2_1
X_1629_ _1436_ _1437_ _1438_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__nor3_2
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1980_ _0494_ _0536_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__and2b_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2601_ _1000_ _0884_ _0883_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__or3b_4
X_2532_ po_0.regf_0.rf\[15\]\[0\] _0927_ _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2463_ _0940_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
X_2394_ _0899_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3015_ net82 net23 _1295_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__mux2_1
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout110 net111 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_1
Xfanout121 net125 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout165 net169 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_1
Xfanout132 net133 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout143 net149 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout154 net155 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_1
Xfanout176 net182 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1963_ po_0.regf_0.rf\[12\]\[11\] po_0.regf_0.rf\[13\]\[11\] po_0.regf_0.rf\[14\]\[11\]
+ po_0.regf_0.rf\[15\]\[11\] _0441_ _0442_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__mux4_1
XFILLER_21_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1894_ _0455_ _0457_ _0410_ _0460_ VGND VGND VPWR VPWR po_0.regf_0._3_\[3\] sky130_fd_sc_hd__o22a_1
X_3564_ po_0.alu_0._10_\[5\] _1563_ VGND VGND VPWR VPWR po_0.alu_0._11_\[5\] sky130_fd_sc_hd__ebufn_1
X_3495_ net118 _0279_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2515_ _0973_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
X_2446_ _0928_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__buf_2
X_2377_ _0890_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2300_ _0821_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
X_3280_ net146 _0068_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _0725_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__buf_2
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2162_ _0685_ _0679_ _0692_ _0693_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2093_ _0631_ _0632_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__nor2_1
XFILLER_80_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2995_ _0566_ net28 _1296_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__mux2_1
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1946_ po_0.regf_0.rf\[0\]\[9\] po_0.regf_0.rf\[1\]\[9\] po_0.regf_0.rf\[2\]\[9\]
+ po_0.regf_0.rf\[3\]\[9\] _0414_ _0415_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__mux4_1
X_1877_ _0003_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__buf_2
X_3547_ net168 _0331_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3478_ net137 _0262_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2429_ _0919_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1800_ _1500_ _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__and2b_1
X_2780_ _1118_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__clkbuf_1
X_1731_ _1487_ _1531_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__and2b_1
X_1662_ _1467_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__buf_2
X_3401_ net123 _0189_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3332_ net103 _0120_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_1593_ _1406_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__clkbuf_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ net108 _0055_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _0742_ po_0.regf_0.rf\[7\]\[2\] _0720_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__mux2_1
X_3194_ net127 _0018_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ _0667_ _0670_ _0678_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__o21bai_2
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2076_ _0609_ _0614_ _0615_ _0616_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__or4_1
XFILLER_34_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2978_ _1135_ _1187_ net96 _1284_ _1286_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__o32a_1
X_1929_ _0485_ _0487_ _0489_ _0491_ VGND VGND VPWR VPWR po_0.regf_0._3_\[7\] sky130_fd_sc_hd__o22a_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2901_ _1216_ _1145_ _1217_ _1207_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__a31o_1
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2832_ _1152_ _1150_ _1136_ _0704_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__a2bb2o_1
X_2763_ _0820_ po_0.regf_0.rf\[0\]\[9\] _1105_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__mux2_1
X_1714_ po_0.regf_0.rf\[4\]\[3\] po_0.regf_0.rf\[5\]\[3\] po_0.regf_0.rf\[6\]\[3\]
+ po_0.regf_0.rf\[7\]\[3\] _1497_ _1498_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__mux4_1
X_2694_ _1071_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_1
X_1645_ _1440_ _1451_ VGND VGND VPWR VPWR uc_0.bc_0._54_\[2\] sky130_fd_sc_hd__nor2_1
X_1576_ _1402_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__clkbuf_2
X_3315_ net112 _0103_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ po_0.regf_0._3_\[6\] net89 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlxtp_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _0744_ net54 _1393_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__mux2_1
XFILLER_39_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2128_ _0661_ _0662_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__or2_1
XFILLER_66_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2059_ _0596_ _0597_ _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__nand3_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput80 net80 VGND VGND VPWR VPWR leds[1] sky130_fd_sc_hd__buf_2
X_3100_ po_0.regf_0.rf\[2\]\[3\] _0752_ _1351_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__mux2_1
X_3031_ _1317_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2815_ _1136_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__clkbuf_2
X_2746_ _0732_ po_0.regf_0.rf\[0\]\[1\] _1098_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__mux2_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2677_ _1062_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
X_1628_ net46 net45 net85 net47 VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__or4_2
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3229_ po_0.regf_0._5_\[5\] net95 VGND VGND VPWR VPWR po_0._1_\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2600_ _1019_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
X_2531_ _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__buf_2
XFILLER_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2462_ po_0.regf_0.rf\[9\]\[5\] _0939_ _0929_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__mux2_1
X_2393_ po_0.regf_0.rf\[6\]\[9\] _0820_ _0895_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__mux2_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3014_ _1306_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2729_ _1090_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__clkbuf_1
Xfanout111 net115 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
Xfanout100 net101 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
Xfanout122 net124 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
Xfanout133 net149 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
Xfanout144 net148 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
Xfanout155 net156 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout177 net179 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout166 net168 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1962_ _0494_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__and2b_1
X_1893_ _0458_ _0459_ _0417_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__mux2_1
X_3563_ po_0.alu_0._10_\[4\] _1562_ VGND VGND VPWR VPWR po_0.alu_0._11_\[4\] sky130_fd_sc_hd__ebufn_1
X_3494_ net146 _0278_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2514_ po_0.regf_0.rf\[1\]\[8\] _0946_ _0970_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__mux2_1
X_2445_ _0886_ _0715_ _0906_ _0907_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__and4b_2
X_2376_ po_0.regf_0.rf\[6\]\[1\] _0732_ _0888_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__mux2_1
XFILLER_17_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _0598_ po_0._1_\[3\] _0755_ _0746_ _0610_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__o221ai_4
XFILLER_38_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2161_ _0680_ po_0._1_\[14\] VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__nor2_1
XFILLER_65_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2092_ net85 po_0._1_\[7\] VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__and2_1
XFILLER_53_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2994_ _1295_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__buf_2
X_1945_ _0494_ _0505_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__and2b_1
X_1876_ _0422_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__buf_2
X_3546_ net180 _0330_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dfxtp_1
X_3477_ net137 _0261_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2428_ po_0.regf_0.rf\[5\]\[8\] _0811_ _0916_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__mux2_1
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2359_ _0689_ _0690_ _0865_ _0874_ _0681_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__o221ai_1
XFILLER_69_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1730_ po_0.regf_0.rf\[0\]\[5\] po_0.regf_0.rf\[1\]\[5\] po_0.regf_0.rf\[2\]\[5\]
+ po_0.regf_0.rf\[3\]\[5\] _1488_ _1489_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__mux4_1
X_1661_ _0007_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__clkbuf_2
X_3400_ net170 _0188_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3331_ net112 _0119_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1592_ _1413_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__clkbuf_2
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ net108 _0054_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2213_ _0741_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__dlymetal6s2s_1
X_3193_ net134 _0017_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _0673_ _0674_ _0664_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__o21ai_1
XFILLER_26_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2075_ _0614_ _0615_ _0616_ _0609_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__o22ai_2
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2977_ net96 _1276_ _1285_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__o21a_1
X_1928_ _0490_ _0431_ _0410_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__a21o_1
X_1859_ _0394_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3529_ net154 _0313_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2900_ _1172_ _1185_ _1200_ _1166_ _1213_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__a41o_1
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2831_ _1150_ _1137_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__or3_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2762_ _1108_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__clkbuf_1
X_1713_ po_0.regf_0.rf\[0\]\[3\] po_0.regf_0.rf\[1\]\[3\] po_0.regf_0.rf\[2\]\[3\]
+ po_0.regf_0.rf\[3\]\[3\] _1494_ _1495_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__mux4_1
X_2693_ po_0.regf_0.rf\[11\]\[9\] _0948_ _1067_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__mux2_1
X_1644_ net82 net81 _1448_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__or3b_1
X_1575_ _1401_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__clkbuf_2
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ net118 _0102_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ po_0.regf_0._3_\[5\] net90 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlxtp_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _1394_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2127_ net83 po_0._1_\[12\] VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__nor2_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2058_ _0599_ _0600_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__nor2_1
XFILLER_81_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput70 net99 VGND VGND VPWR VPWR I_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_68_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput81 net81 VGND VGND VPWR VPWR leds[2] sky130_fd_sc_hd__clkbuf_4
X_3030_ po_0.regf_0.rf\[4\]\[3\] _0752_ _1313_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__mux2_1
XFILLER_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2814_ _1136_ po_0.muxf_0.rf_w_data\[0\] VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__nand2_1
X_2745_ _1099_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__clkbuf_1
X_2676_ po_0.regf_0.rf\[11\]\[1\] _0931_ _1060_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__mux2_1
X_1627_ net87 net86 net44 net43 VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__or4_2
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3228_ po_0.regf_0._5_\[4\] net94 VGND VGND VPWR VPWR po_0._1_\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_27_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3159_ _0718_ _1385_ _1372_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__mux2_1
XFILLER_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2530_ _0718_ _0715_ _0716_ _0717_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__and4_2
X_2461_ _0772_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__clkbuf_2
X_2392_ _0898_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3013_ net81 net22 _1295_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__mux2_1
XFILLER_36_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2728_ po_0.regf_0.rf\[10\]\[9\] _0948_ _1086_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__mux2_1
X_2659_ _1052_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
Xfanout101 net107 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout112 net114 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
Xfanout134 net139 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
Xfanout145 net148 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
Xfanout123 net124 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
Xfanout156 net169 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout167 net168 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
Xfanout178 net179 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1961_ po_0.regf_0.rf\[0\]\[11\] po_0.regf_0.rf\[1\]\[11\] po_0.regf_0.rf\[2\]\[11\]
+ po_0.regf_0.rf\[3\]\[11\] _0495_ _0496_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__mux4_1
XFILLER_53_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1892_ po_0.regf_0.rf\[4\]\[3\] po_0.regf_0.rf\[5\]\[3\] po_0.regf_0.rf\[6\]\[3\]
+ po_0.regf_0.rf\[7\]\[3\] _0414_ _0415_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__mux4_1
X_3562_ po_0.alu_0._10_\[3\] _1561_ VGND VGND VPWR VPWR po_0.alu_0._11_\[3\] sky130_fd_sc_hd__ebufn_1
X_2513_ _0972_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
X_3493_ net146 _0277_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2444_ _0713_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__clkbuf_2
X_2375_ _0889_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _0680_ po_0._1_\[14\] VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__and2_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2091_ net85 po_0._1_\[7\] VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2993_ uc_0._03_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__clkbuf_4
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1944_ po_0.regf_0.rf\[8\]\[9\] po_0.regf_0.rf\[9\]\[9\] po_0.regf_0.rf\[10\]\[9\]
+ po_0.regf_0.rf\[11\]\[9\] _0495_ _0496_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__mux4_1
X_1875_ po_0.regf_0.rf\[12\]\[2\] po_0.regf_0.rf\[13\]\[2\] po_0.regf_0.rf\[14\]\[2\]
+ po_0.regf_0.rf\[15\]\[2\] _0441_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__mux4_1
X_3545_ net126 _0329_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dfxtp_1
X_3476_ net130 _0260_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2427_ _0918_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2358_ _0861_ _0862_ _0864_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__a21boi_1
XFILLER_84_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2289_ _0811_ po_0.regf_0.rf\[7\]\[8\] _0784_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__mux2_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1660_ _1465_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__buf_2
X_1591_ _1402_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__dlymetal6s2s_1
X_3330_ net112 _0118_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ net135 _0053_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3192_ net134 _0016_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _0722_ _0723_ net9 _0740_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__a31o_2
XFILLER_78_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2143_ _0672_ po_0._1_\[12\] _0675_ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__o211ai_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2074_ po_0._1_\[4\] _0605_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__and2b_1
XFILLER_53_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2976_ net96 _1276_ _1186_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__a21oi_1
X_1927_ po_0.regf_0.rf\[4\]\[7\] po_0.regf_0.rf\[5\]\[7\] po_0.regf_0.rf\[6\]\[7\]
+ po_0.regf_0.rf\[7\]\[7\] _0428_ _0429_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__mux4_1
X_1858_ _0403_ _0426_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__and2b_1
X_1789_ _0357_ _0359_ _0361_ _0363_ VGND VGND VPWR VPWR po_0.regf_0._5_\[11\] sky130_fd_sc_hd__o22a_1
XFILLER_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3528_ net154 _0312_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[2\] sky130_fd_sc_hd__dfxtp_1
X_3459_ net167 _0243_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2830_ _1151_ po_0.muxf_0.rf_w_data\[1\] VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__and2_1
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2761_ _0811_ po_0.regf_0.rf\[0\]\[8\] _1105_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__mux2_1
XFILLER_31_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2692_ _1070_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
X_1712_ _1511_ _1514_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__and2b_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 _0744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1643_ _1450_ VGND VGND VPWR VPWR uc_0.bc_0._54_\[3\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1574_ po_0.alu_0.s0 VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__clkbuf_2
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ net145 _0101_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ po_0.regf_0._3_\[4\] net90 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlxtp_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ _0734_ net53 _1393_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__mux2_1
XFILLER_66_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2126_ net83 po_0._1_\[12\] VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__and2_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2057_ _0596_ _0597_ _0599_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__o2bb2ai_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2959_ _1269_ _1234_ _1264_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__nand3_1
XFILLER_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput60 net60 VGND VGND VPWR VPWR D_wr sky130_fd_sc_hd__buf_2
Xoutput71 net71 VGND VGND VPWR VPWR I_addr[4] sky130_fd_sc_hd__buf_2
Xoutput82 net82 VGND VGND VPWR VPWR leds[3] sky130_fd_sc_hd__buf_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2813_ net61 VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2744_ _0714_ po_0.regf_0.rf\[0\]\[0\] _1098_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__mux2_1
X_2675_ _1061_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
X_1626_ _1433_ _1434_ _1435_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__nand3_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ po_0.regf_0._5_\[3\] net94 VGND VGND VPWR VPWR po_0._1_\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_27_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3158_ uc_0._20_\[10\] _0734_ _0562_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__mux2_1
XFILLER_36_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2109_ net36 VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__dlymetal6s2s_1
X_3089_ _1348_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2460_ _0938_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_2391_ po_0.regf_0.rf\[6\]\[8\] _0811_ _0895_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__mux2_1
X_3012_ _1305_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2727_ _1089_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__clkbuf_1
X_2658_ po_0.regf_0.rf\[12\]\[9\] _0948_ _1048_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__mux2_1
X_2589_ _0830_ po_0.regf_0.rf\[14\]\[10\] _1009_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__mux2_1
Xfanout113 net114 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout102 net107 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlymetal6s2s_1
X_1609_ _1413_ _1415_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__or2b_1
Xfanout135 net139 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout124 net125 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xfanout146 net147 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
Xfanout168 net169 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
Xfanout179 net180 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
Xfanout157 net158 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1960_ _0518_ _0400_ _0432_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__a21o_1
XFILLER_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1891_ po_0.regf_0.rf\[0\]\[3\] po_0.regf_0.rf\[1\]\[3\] po_0.regf_0.rf\[2\]\[3\]
+ po_0.regf_0.rf\[3\]\[3\] _0411_ _0412_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__mux4_1
X_3561_ po_0.alu_0._10_\[2\] _1560_ VGND VGND VPWR VPWR po_0.alu_0._11_\[2\] sky130_fd_sc_hd__ebufn_1
X_2512_ po_0.regf_0.rf\[1\]\[7\] _0944_ _0970_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__mux2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3492_ net142 _0276_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2443_ _0926_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2374_ po_0.regf_0.rf\[6\]\[0\] _0714_ _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__mux2_1
XFILLER_68_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2090_ _0621_ _0620_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__and2b_1
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2992_ _1294_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__clkbuf_1
X_1943_ _0503_ _0447_ _0401_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__a21bo_1
X_1874_ _0396_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__buf_2
X_3544_ net108 _0328_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dfxtp_1
X_3475_ net130 _0259_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2426_ po_0.regf_0.rf\[5\]\[7\] _0796_ _0916_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__mux2_1
XFILLER_69_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2357_ _0692_ _0866_ _0691_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2288_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__clkbuf_2
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1590_ _1412_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__clkbuf_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ net135 _0052_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3191_ uc_0.bc_0._54_\[1\] _0559_ _0560_ _1310_ _1135_ VGND VGND VPWR VPWR _0337_
+ sky130_fd_sc_hd__a32o_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _0734_ _0702_ _0739_ _0729_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__a22o_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2142_ _0667_ _0670_ _0664_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__o21ai_1
X_2073_ _0613_ po_0._1_\[5\] VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__and2_1
XFILLER_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2975_ net96 _1147_ _1277_ _1283_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__o31a_1
X_1926_ _0447_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__and2b_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1857_ po_0.regf_0.rf\[0\]\[1\] po_0.regf_0.rf\[1\]\[1\] po_0.regf_0.rf\[2\]\[1\]
+ po_0.regf_0.rf\[3\]\[1\] _0405_ _0407_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux4_1
X_1788_ _0362_ _1478_ _1479_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__a21o_1
X_3527_ net162 _0311_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[1\] sky130_fd_sc_hd__dfxtp_1
X_3458_ net178 _0242_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[2\] sky130_fd_sc_hd__dfxtp_1
X_3389_ net173 _0177_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2409_ _0882_ _0906_ _0907_ _0886_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__and4b_4
XFILLER_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2760_ _1107_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__clkbuf_1
X_2691_ po_0.regf_0.rf\[11\]\[8\] _0946_ _1067_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__mux2_1
X_1711_ po_0.regf_0.rf\[8\]\[3\] po_0.regf_0.rf\[9\]\[3\] po_0.regf_0.rf\[10\]\[3\]
+ po_0.regf_0.rf\[11\]\[3\] _1512_ _1513_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__mux4_1
XANTENNA_2 _0810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1642_ _1439_ _1449_ _1440_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__o21ba_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ net144 _0100_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ po_0.regf_0._3_\[3\] net90 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlxtp_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _1369_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__buf_4
XFILLER_66_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2125_ _0658_ _0660_ VGND VGND VPWR VPWR po_0.alu_0._10_\[11\] sky130_fd_sc_hd__xnor2_1
XFILLER_19_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2056_ _0598_ po_0._1_\[3\] VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__nor2_2
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2958_ net64 VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1909_ _0472_ _0473_ _0399_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__mux2_1
X_2889_ _1147_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__clkbuf_2
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput50 net50 VGND VGND VPWR VPWR D_W_data[9] sky130_fd_sc_hd__clkbuf_4
Xoutput61 net61 VGND VGND VPWR VPWR I_addr[0] sky130_fd_sc_hd__buf_2
Xoutput72 net72 VGND VGND VPWR VPWR I_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_51_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2812_ uc_0._01_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__buf_2
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2743_ _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__buf_2
X_2674_ po_0.regf_0.rf\[11\]\[0\] _0927_ _1060_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__mux2_1
X_1625_ net50 net49 net84 net36 VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__nor4_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3226_ po_0.regf_0._5_\[2\] net94 VGND VGND VPWR VPWR po_0._1_\[2\] sky130_fd_sc_hd__dlxtp_1
X_3157_ _1384_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__clkbuf_1
X_2108_ _0643_ _0645_ VGND VGND VPWR VPWR po_0.alu_0._10_\[9\] sky130_fd_sc_hd__xor2_1
X_3088_ po_0.regf_0.rf\[3\]\[14\] _0870_ _1331_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__mux2_1
X_2039_ net86 VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__inv_2
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2390_ _0897_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3011_ net80 net21 _1295_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__mux2_1
XFILLER_36_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2726_ po_0.regf_0.rf\[10\]\[8\] _0946_ _1086_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__mux2_1
X_2657_ _1051_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
X_1608_ _1423_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__clkbuf_1
Xfanout103 net106 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
X_2588_ _1013_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout136 net138 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout114 net115 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
Xfanout147 net148 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
Xfanout125 net183 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
Xfanout169 net183 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
Xfanout158 net161 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
X_3209_ net134 _0033_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1890_ _0403_ _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__and2b_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3560_ po_0.alu_0._10_\[1\] _1559_ VGND VGND VPWR VPWR po_0.alu_0._11_\[1\] sky130_fd_sc_hd__ebufn_1
X_2511_ _0971_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
X_3491_ net142 _0275_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2442_ po_0.regf_0.rf\[5\]\[15\] _0880_ _0908_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__mux2_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2373_ _0887_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__buf_2
XFILLER_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2709_ po_0.regf_0.rf\[10\]\[0\] _0927_ _1079_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__mux2_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2991_ _0557_ net27 _1289_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__mux2_1
X_1942_ po_0.regf_0.rf\[12\]\[9\] po_0.regf_0.rf\[13\]\[9\] po_0.regf_0.rf\[14\]\[9\]
+ po_0.regf_0.rf\[15\]\[9\] _0435_ _0436_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__mux4_1
X_1873_ _0394_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__clkbuf_4
X_3543_ net178 _0327_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dfxtp_1
X_3474_ net136 _0258_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2425_ _0917_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2356_ _0872_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2287_ net15 _0701_ _0809_ _0793_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__a22o_2
XFILLER_84_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _1405_ po_0.alu_0._11_\[2\] _0705_ _0588_ _0738_ VGND VGND VPWR VPWR _0739_
+ sky130_fd_sc_hd__a221o_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3190_ _0572_ _0573_ _1308_ _1145_ _1389_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__o221a_1
XFILLER_38_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2141_ _0673_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__nor2_1
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2072_ _0613_ po_0._1_\[5\] VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__nor2_2
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2974_ _1281_ _1282_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__nor2_1
X_1925_ po_0.regf_0.rf\[0\]\[7\] po_0.regf_0.rf\[1\]\[7\] po_0.regf_0.rf\[2\]\[7\]
+ po_0.regf_0.rf\[3\]\[7\] _0448_ _0449_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux4_1
X_1856_ _0421_ _0423_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__a21o_1
X_1787_ po_0.regf_0.rf\[4\]\[11\] po_0.regf_0.rf\[5\]\[11\] po_0.regf_0.rf\[6\]\[11\]
+ po_0.regf_0.rf\[7\]\[11\] _1475_ _1476_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__mux4_1
X_3526_ net166 _0310_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[0\] sky130_fd_sc_hd__dfxtp_1
X_3457_ net177 _0241_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3388_ net173 _0176_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2408_ _0884_ _0883_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__and2b_1
XFILLER_69_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2339_ _0854_ _0855_ _0856_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1710_ _1456_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__buf_2
X_2690_ _1069_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 _0819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1641_ net80 net82 net81 _1448_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__and4bb_1
X_3311_ net140 _0099_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ po_0.regf_0._3_\[2\] net90 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlxtp_1
X_3173_ _1392_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__clkbuf_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2124_ _0654_ _0659_ _0647_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__a21boi_1
XFILLER_19_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2055_ _0598_ po_0._1_\[3\] VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__and2_1
XFILLER_22_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2957_ net63 _1215_ _1266_ _1268_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__o22a_1
X_1908_ po_0.regf_0.rf\[12\]\[5\] po_0.regf_0.rf\[13\]\[5\] po_0.regf_0.rf\[14\]\[5\]
+ po_0.regf_0.rf\[15\]\[5\] _0000_ _0001_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux4_1
X_2888_ _1204_ _1203_ _1202_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__a21o_1
X_1839_ _0403_ _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__and2b_1
X_3509_ net147 _0293_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput51 net51 VGND VGND VPWR VPWR D_addr[0] sky130_fd_sc_hd__buf_2
Xoutput40 net40 VGND VGND VPWR VPWR D_W_data[14] sky130_fd_sc_hd__buf_2
Xoutput73 net98 VGND VGND VPWR VPWR I_addr[6] sky130_fd_sc_hd__clkbuf_4
Xoutput62 net62 VGND VGND VPWR VPWR I_addr[10] sky130_fd_sc_hd__buf_2
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2811_ _1134_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__clkbuf_1
X_2742_ _0718_ _0882_ _0716_ _1039_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__or4bb_4
X_2673_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__buf_2
X_1624_ net39 net83 net41 net40 VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__nor4_1
X_3225_ po_0.regf_0._5_\[1\] net94 VGND VGND VPWR VPWR po_0._1_\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3156_ _0884_ _1383_ _1372_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__mux2_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3087_ _1347_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__clkbuf_1
X_2107_ _0640_ _0642_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__a21oi_1
X_2038_ _0580_ _0583_ VGND VGND VPWR VPWR po_0.alu_0._10_\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3010_ _1304_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2725_ _1088_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2656_ po_0.regf_0.rf\[12\]\[8\] _0946_ _1048_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__mux2_1
X_1607_ _1413_ _1415_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__or2b_1
Xfanout104 net106 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
X_2587_ _0820_ po_0.regf_0.rf\[14\]\[9\] _1009_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__mux2_1
Xfanout126 net127 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout137 net138 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
Xfanout115 net125 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout148 net149 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
Xfanout159 net160 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
X_3208_ net134 _0032_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3139_ _1374_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2510_ po_0.regf_0.rf\[1\]\[6\] _0941_ _0970_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__mux2_1
X_3490_ net147 _0274_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2441_ _0925_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2372_ _0882_ _0716_ _0885_ _0886_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__and4b_4
XFILLER_68_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2708_ _1078_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__buf_2
X_2639_ po_0.regf_0.rf\[12\]\[0\] _0927_ _1041_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__mux2_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2990_ _1293_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1941_ _0493_ _0498_ _0500_ _0502_ VGND VGND VPWR VPWR po_0.regf_0._3_\[8\] sky130_fd_sc_hd__o22a_1
XFILLER_61_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1872_ _0417_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__and2b_1
X_3542_ net166 _0326_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfxtp_2
X_3473_ net136 _0257_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2424_ po_0.regf_0.rf\[5\]\[6\] _0783_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__mux2_1
XFILLER_69_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2355_ _0871_ po_0.regf_0.rf\[7\]\[14\] _0719_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__mux2_1
X_2286_ _0806_ _0807_ _0758_ _0808_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__a31o_1
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ net39 po_0._1_\[13\] VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__and2_1
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2071_ net46 VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__clkbuf_2
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2973_ _1140_ net96 _1277_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__and3_1
X_1924_ _0486_ _0434_ _0401_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__a21bo_1
X_1855_ _0003_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__buf_2
X_1786_ _1487_ _0360_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__and2b_1
X_3525_ net159 _0309_ VGND VGND VPWR VPWR po_0.regf_0.w_wr sky130_fd_sc_hd__dfxtp_1
X_3456_ net177 _0240_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[0\] sky130_fd_sc_hd__dfxtp_1
X_2407_ po_0.regf_0.w_wr VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__dlymetal6s2s_1
X_3387_ net170 _0175_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2338_ _1406_ po_0.alu_0._11_\[13\] _0815_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__a21o_1
X_2269_ _0711_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__buf_2
XFILLER_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1640_ uc_0.bc_0._55_\[2\] uc_0.bc_0._55_\[3\] uc_0.bc_0._55_\[0\] uc_0.bc_0._55_\[1\]
+ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__and4bb_1
XANTENNA_4 _1511_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3310_ net140 _0098_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ po_0.regf_0._3_\[1\] net89 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlxtp_1
X_3172_ _0724_ net52 _1389_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__mux2_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2123_ _0648_ _0651_ _0652_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__and3_1
XFILLER_54_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2054_ net44 VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__buf_2
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2956_ _1226_ _1241_ _1264_ _1187_ _1267_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__a311oi_1
X_1907_ po_0.regf_0.rf\[8\]\[5\] po_0.regf_0.rf\[9\]\[5\] po_0.regf_0.rf\[10\]\[5\]
+ po_0.regf_0.rf\[11\]\[5\] _0000_ _0001_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__mux4_1
X_2887_ _1202_ _1203_ _1204_ _1139_ _1171_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__a311oi_1
X_1838_ po_0.regf_0.rf\[8\]\[0\] po_0.regf_0.rf\[9\]\[0\] po_0.regf_0.rf\[10\]\[0\]
+ po_0.regf_0.rf\[11\]\[0\] _0405_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux4_1
XFILLER_1_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1769_ _0345_ _1466_ _1468_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__a21bo_1
X_3508_ net142 _0292_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3439_ net167 _0227_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfxtp_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput52 net52 VGND VGND VPWR VPWR D_addr[1] sky130_fd_sc_hd__clkbuf_4
Xoutput41 net41 VGND VGND VPWR VPWR D_W_data[15] sky130_fd_sc_hd__buf_2
Xoutput63 net63 VGND VGND VPWR VPWR I_addr[11] sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 VGND VGND VPWR VPWR I_addr[7] sky130_fd_sc_hd__buf_2
XFILLER_0_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2810_ po_0.regf_0.rf\[8\]\[15\] _0879_ _1116_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__mux2_1
X_2741_ _1096_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2672_ po_0.regf_0.w_addr\[2\] _0715_ po_0.regf_0.w_wr _0717_ VGND VGND VPWR VPWR
+ _1059_ sky130_fd_sc_hd__and4b_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1623_ uc_0.bc_0._55_\[1\] uc_0.bc_0._55_\[2\] uc_0.bc_0._55_\[3\] uc_0.bc_0._55_\[0\]
+ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__and4bb_1
X_3224_ po_0.regf_0._5_\[0\] net94 VGND VGND VPWR VPWR po_0._1_\[0\] sky130_fd_sc_hd__dlxtp_1
.ends

