// This is the unpowered netlist.
module vahid6i (D_rd,
    D_wr,
    I_rd,
    clock,
    led_clock,
    reset,
    D_R_data,
    D_W_data,
    D_addr,
    I_addr,
    I_data,
    leds);
 output D_rd;
 output D_wr;
 output I_rd;
 input clock;
 output led_clock;
 input reset;
 input [15:0] D_R_data;
 output [15:0] D_W_data;
 output [7:0] D_addr;
 output [15:0] I_addr;
 input [15:0] I_data;
 output [3:0] leds;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \po_0._1_[0] ;
 wire \po_0._1_[10] ;
 wire \po_0._1_[11] ;
 wire \po_0._1_[12] ;
 wire \po_0._1_[13] ;
 wire \po_0._1_[14] ;
 wire \po_0._1_[15] ;
 wire \po_0._1_[1] ;
 wire \po_0._1_[2] ;
 wire \po_0._1_[3] ;
 wire \po_0._1_[4] ;
 wire \po_0._1_[5] ;
 wire \po_0._1_[6] ;
 wire \po_0._1_[7] ;
 wire \po_0._1_[8] ;
 wire \po_0._1_[9] ;
 wire \po_0.alu_0._10_[0] ;
 wire \po_0.alu_0._10_[10] ;
 wire \po_0.alu_0._10_[11] ;
 wire \po_0.alu_0._10_[12] ;
 wire \po_0.alu_0._10_[13] ;
 wire \po_0.alu_0._10_[14] ;
 wire \po_0.alu_0._10_[15] ;
 wire \po_0.alu_0._10_[1] ;
 wire \po_0.alu_0._10_[2] ;
 wire \po_0.alu_0._10_[3] ;
 wire \po_0.alu_0._10_[4] ;
 wire \po_0.alu_0._10_[5] ;
 wire \po_0.alu_0._10_[6] ;
 wire \po_0.alu_0._10_[7] ;
 wire \po_0.alu_0._10_[8] ;
 wire \po_0.alu_0._10_[9] ;
 wire \po_0.alu_0._11_[0] ;
 wire \po_0.alu_0._11_[10] ;
 wire \po_0.alu_0._11_[11] ;
 wire \po_0.alu_0._11_[12] ;
 wire \po_0.alu_0._11_[13] ;
 wire \po_0.alu_0._11_[14] ;
 wire \po_0.alu_0._11_[15] ;
 wire \po_0.alu_0._11_[1] ;
 wire \po_0.alu_0._11_[2] ;
 wire \po_0.alu_0._11_[3] ;
 wire \po_0.alu_0._11_[4] ;
 wire \po_0.alu_0._11_[5] ;
 wire \po_0.alu_0._11_[6] ;
 wire \po_0.alu_0._11_[7] ;
 wire \po_0.alu_0._11_[8] ;
 wire \po_0.alu_0._11_[9] ;
 wire \po_0.alu_0.s0 ;
 wire \po_0.alu_0.s1 ;
 wire \po_0.muxf_0.rf_w_data[0] ;
 wire \po_0.muxf_0.rf_w_data[1] ;
 wire \po_0.muxf_0.rf_w_data[2] ;
 wire \po_0.muxf_0.rf_w_data[3] ;
 wire \po_0.muxf_0.rf_w_data[4] ;
 wire \po_0.muxf_0.rf_w_data[5] ;
 wire \po_0.muxf_0.rf_w_data[6] ;
 wire \po_0.muxf_0.rf_w_data[7] ;
 wire \po_0.muxf_0.s0 ;
 wire \po_0.muxf_0.s1 ;
 wire \po_0.regf_0._3_[0] ;
 wire \po_0.regf_0._3_[10] ;
 wire \po_0.regf_0._3_[11] ;
 wire \po_0.regf_0._3_[12] ;
 wire \po_0.regf_0._3_[13] ;
 wire \po_0.regf_0._3_[14] ;
 wire \po_0.regf_0._3_[15] ;
 wire \po_0.regf_0._3_[1] ;
 wire \po_0.regf_0._3_[2] ;
 wire \po_0.regf_0._3_[3] ;
 wire \po_0.regf_0._3_[4] ;
 wire \po_0.regf_0._3_[5] ;
 wire \po_0.regf_0._3_[6] ;
 wire \po_0.regf_0._3_[7] ;
 wire \po_0.regf_0._3_[8] ;
 wire \po_0.regf_0._3_[9] ;
 wire \po_0.regf_0._5_[0] ;
 wire \po_0.regf_0._5_[10] ;
 wire \po_0.regf_0._5_[11] ;
 wire \po_0.regf_0._5_[12] ;
 wire \po_0.regf_0._5_[13] ;
 wire \po_0.regf_0._5_[14] ;
 wire \po_0.regf_0._5_[15] ;
 wire \po_0.regf_0._5_[1] ;
 wire \po_0.regf_0._5_[2] ;
 wire \po_0.regf_0._5_[3] ;
 wire \po_0.regf_0._5_[4] ;
 wire \po_0.regf_0._5_[5] ;
 wire \po_0.regf_0._5_[6] ;
 wire \po_0.regf_0._5_[7] ;
 wire \po_0.regf_0._5_[8] ;
 wire \po_0.regf_0._5_[9] ;
 wire \po_0.regf_0.rf[0][0] ;
 wire \po_0.regf_0.rf[0][10] ;
 wire \po_0.regf_0.rf[0][11] ;
 wire \po_0.regf_0.rf[0][12] ;
 wire \po_0.regf_0.rf[0][13] ;
 wire \po_0.regf_0.rf[0][14] ;
 wire \po_0.regf_0.rf[0][15] ;
 wire \po_0.regf_0.rf[0][1] ;
 wire \po_0.regf_0.rf[0][2] ;
 wire \po_0.regf_0.rf[0][3] ;
 wire \po_0.regf_0.rf[0][4] ;
 wire \po_0.regf_0.rf[0][5] ;
 wire \po_0.regf_0.rf[0][6] ;
 wire \po_0.regf_0.rf[0][7] ;
 wire \po_0.regf_0.rf[0][8] ;
 wire \po_0.regf_0.rf[0][9] ;
 wire \po_0.regf_0.rf[10][0] ;
 wire \po_0.regf_0.rf[10][10] ;
 wire \po_0.regf_0.rf[10][11] ;
 wire \po_0.regf_0.rf[10][12] ;
 wire \po_0.regf_0.rf[10][13] ;
 wire \po_0.regf_0.rf[10][14] ;
 wire \po_0.regf_0.rf[10][15] ;
 wire \po_0.regf_0.rf[10][1] ;
 wire \po_0.regf_0.rf[10][2] ;
 wire \po_0.regf_0.rf[10][3] ;
 wire \po_0.regf_0.rf[10][4] ;
 wire \po_0.regf_0.rf[10][5] ;
 wire \po_0.regf_0.rf[10][6] ;
 wire \po_0.regf_0.rf[10][7] ;
 wire \po_0.regf_0.rf[10][8] ;
 wire \po_0.regf_0.rf[10][9] ;
 wire \po_0.regf_0.rf[11][0] ;
 wire \po_0.regf_0.rf[11][10] ;
 wire \po_0.regf_0.rf[11][11] ;
 wire \po_0.regf_0.rf[11][12] ;
 wire \po_0.regf_0.rf[11][13] ;
 wire \po_0.regf_0.rf[11][14] ;
 wire \po_0.regf_0.rf[11][15] ;
 wire \po_0.regf_0.rf[11][1] ;
 wire \po_0.regf_0.rf[11][2] ;
 wire \po_0.regf_0.rf[11][3] ;
 wire \po_0.regf_0.rf[11][4] ;
 wire \po_0.regf_0.rf[11][5] ;
 wire \po_0.regf_0.rf[11][6] ;
 wire \po_0.regf_0.rf[11][7] ;
 wire \po_0.regf_0.rf[11][8] ;
 wire \po_0.regf_0.rf[11][9] ;
 wire \po_0.regf_0.rf[12][0] ;
 wire \po_0.regf_0.rf[12][10] ;
 wire \po_0.regf_0.rf[12][11] ;
 wire \po_0.regf_0.rf[12][12] ;
 wire \po_0.regf_0.rf[12][13] ;
 wire \po_0.regf_0.rf[12][14] ;
 wire \po_0.regf_0.rf[12][15] ;
 wire \po_0.regf_0.rf[12][1] ;
 wire \po_0.regf_0.rf[12][2] ;
 wire \po_0.regf_0.rf[12][3] ;
 wire \po_0.regf_0.rf[12][4] ;
 wire \po_0.regf_0.rf[12][5] ;
 wire \po_0.regf_0.rf[12][6] ;
 wire \po_0.regf_0.rf[12][7] ;
 wire \po_0.regf_0.rf[12][8] ;
 wire \po_0.regf_0.rf[12][9] ;
 wire \po_0.regf_0.rf[13][0] ;
 wire \po_0.regf_0.rf[13][10] ;
 wire \po_0.regf_0.rf[13][11] ;
 wire \po_0.regf_0.rf[13][12] ;
 wire \po_0.regf_0.rf[13][13] ;
 wire \po_0.regf_0.rf[13][14] ;
 wire \po_0.regf_0.rf[13][15] ;
 wire \po_0.regf_0.rf[13][1] ;
 wire \po_0.regf_0.rf[13][2] ;
 wire \po_0.regf_0.rf[13][3] ;
 wire \po_0.regf_0.rf[13][4] ;
 wire \po_0.regf_0.rf[13][5] ;
 wire \po_0.regf_0.rf[13][6] ;
 wire \po_0.regf_0.rf[13][7] ;
 wire \po_0.regf_0.rf[13][8] ;
 wire \po_0.regf_0.rf[13][9] ;
 wire \po_0.regf_0.rf[14][0] ;
 wire \po_0.regf_0.rf[14][10] ;
 wire \po_0.regf_0.rf[14][11] ;
 wire \po_0.regf_0.rf[14][12] ;
 wire \po_0.regf_0.rf[14][13] ;
 wire \po_0.regf_0.rf[14][14] ;
 wire \po_0.regf_0.rf[14][15] ;
 wire \po_0.regf_0.rf[14][1] ;
 wire \po_0.regf_0.rf[14][2] ;
 wire \po_0.regf_0.rf[14][3] ;
 wire \po_0.regf_0.rf[14][4] ;
 wire \po_0.regf_0.rf[14][5] ;
 wire \po_0.regf_0.rf[14][6] ;
 wire \po_0.regf_0.rf[14][7] ;
 wire \po_0.regf_0.rf[14][8] ;
 wire \po_0.regf_0.rf[14][9] ;
 wire \po_0.regf_0.rf[15][0] ;
 wire \po_0.regf_0.rf[15][10] ;
 wire \po_0.regf_0.rf[15][11] ;
 wire \po_0.regf_0.rf[15][12] ;
 wire \po_0.regf_0.rf[15][13] ;
 wire \po_0.regf_0.rf[15][14] ;
 wire \po_0.regf_0.rf[15][15] ;
 wire \po_0.regf_0.rf[15][1] ;
 wire \po_0.regf_0.rf[15][2] ;
 wire \po_0.regf_0.rf[15][3] ;
 wire \po_0.regf_0.rf[15][4] ;
 wire \po_0.regf_0.rf[15][5] ;
 wire \po_0.regf_0.rf[15][6] ;
 wire \po_0.regf_0.rf[15][7] ;
 wire \po_0.regf_0.rf[15][8] ;
 wire \po_0.regf_0.rf[15][9] ;
 wire \po_0.regf_0.rf[1][0] ;
 wire \po_0.regf_0.rf[1][10] ;
 wire \po_0.regf_0.rf[1][11] ;
 wire \po_0.regf_0.rf[1][12] ;
 wire \po_0.regf_0.rf[1][13] ;
 wire \po_0.regf_0.rf[1][14] ;
 wire \po_0.regf_0.rf[1][15] ;
 wire \po_0.regf_0.rf[1][1] ;
 wire \po_0.regf_0.rf[1][2] ;
 wire \po_0.regf_0.rf[1][3] ;
 wire \po_0.regf_0.rf[1][4] ;
 wire \po_0.regf_0.rf[1][5] ;
 wire \po_0.regf_0.rf[1][6] ;
 wire \po_0.regf_0.rf[1][7] ;
 wire \po_0.regf_0.rf[1][8] ;
 wire \po_0.regf_0.rf[1][9] ;
 wire \po_0.regf_0.rf[2][0] ;
 wire \po_0.regf_0.rf[2][10] ;
 wire \po_0.regf_0.rf[2][11] ;
 wire \po_0.regf_0.rf[2][12] ;
 wire \po_0.regf_0.rf[2][13] ;
 wire \po_0.regf_0.rf[2][14] ;
 wire \po_0.regf_0.rf[2][15] ;
 wire \po_0.regf_0.rf[2][1] ;
 wire \po_0.regf_0.rf[2][2] ;
 wire \po_0.regf_0.rf[2][3] ;
 wire \po_0.regf_0.rf[2][4] ;
 wire \po_0.regf_0.rf[2][5] ;
 wire \po_0.regf_0.rf[2][6] ;
 wire \po_0.regf_0.rf[2][7] ;
 wire \po_0.regf_0.rf[2][8] ;
 wire \po_0.regf_0.rf[2][9] ;
 wire \po_0.regf_0.rf[3][0] ;
 wire \po_0.regf_0.rf[3][10] ;
 wire \po_0.regf_0.rf[3][11] ;
 wire \po_0.regf_0.rf[3][12] ;
 wire \po_0.regf_0.rf[3][13] ;
 wire \po_0.regf_0.rf[3][14] ;
 wire \po_0.regf_0.rf[3][15] ;
 wire \po_0.regf_0.rf[3][1] ;
 wire \po_0.regf_0.rf[3][2] ;
 wire \po_0.regf_0.rf[3][3] ;
 wire \po_0.regf_0.rf[3][4] ;
 wire \po_0.regf_0.rf[3][5] ;
 wire \po_0.regf_0.rf[3][6] ;
 wire \po_0.regf_0.rf[3][7] ;
 wire \po_0.regf_0.rf[3][8] ;
 wire \po_0.regf_0.rf[3][9] ;
 wire \po_0.regf_0.rf[4][0] ;
 wire \po_0.regf_0.rf[4][10] ;
 wire \po_0.regf_0.rf[4][11] ;
 wire \po_0.regf_0.rf[4][12] ;
 wire \po_0.regf_0.rf[4][13] ;
 wire \po_0.regf_0.rf[4][14] ;
 wire \po_0.regf_0.rf[4][15] ;
 wire \po_0.regf_0.rf[4][1] ;
 wire \po_0.regf_0.rf[4][2] ;
 wire \po_0.regf_0.rf[4][3] ;
 wire \po_0.regf_0.rf[4][4] ;
 wire \po_0.regf_0.rf[4][5] ;
 wire \po_0.regf_0.rf[4][6] ;
 wire \po_0.regf_0.rf[4][7] ;
 wire \po_0.regf_0.rf[4][8] ;
 wire \po_0.regf_0.rf[4][9] ;
 wire \po_0.regf_0.rf[5][0] ;
 wire \po_0.regf_0.rf[5][10] ;
 wire \po_0.regf_0.rf[5][11] ;
 wire \po_0.regf_0.rf[5][12] ;
 wire \po_0.regf_0.rf[5][13] ;
 wire \po_0.regf_0.rf[5][14] ;
 wire \po_0.regf_0.rf[5][15] ;
 wire \po_0.regf_0.rf[5][1] ;
 wire \po_0.regf_0.rf[5][2] ;
 wire \po_0.regf_0.rf[5][3] ;
 wire \po_0.regf_0.rf[5][4] ;
 wire \po_0.regf_0.rf[5][5] ;
 wire \po_0.regf_0.rf[5][6] ;
 wire \po_0.regf_0.rf[5][7] ;
 wire \po_0.regf_0.rf[5][8] ;
 wire \po_0.regf_0.rf[5][9] ;
 wire \po_0.regf_0.rf[6][0] ;
 wire \po_0.regf_0.rf[6][10] ;
 wire \po_0.regf_0.rf[6][11] ;
 wire \po_0.regf_0.rf[6][12] ;
 wire \po_0.regf_0.rf[6][13] ;
 wire \po_0.regf_0.rf[6][14] ;
 wire \po_0.regf_0.rf[6][15] ;
 wire \po_0.regf_0.rf[6][1] ;
 wire \po_0.regf_0.rf[6][2] ;
 wire \po_0.regf_0.rf[6][3] ;
 wire \po_0.regf_0.rf[6][4] ;
 wire \po_0.regf_0.rf[6][5] ;
 wire \po_0.regf_0.rf[6][6] ;
 wire \po_0.regf_0.rf[6][7] ;
 wire \po_0.regf_0.rf[6][8] ;
 wire \po_0.regf_0.rf[6][9] ;
 wire \po_0.regf_0.rf[7][0] ;
 wire \po_0.regf_0.rf[7][10] ;
 wire \po_0.regf_0.rf[7][11] ;
 wire \po_0.regf_0.rf[7][12] ;
 wire \po_0.regf_0.rf[7][13] ;
 wire \po_0.regf_0.rf[7][14] ;
 wire \po_0.regf_0.rf[7][15] ;
 wire \po_0.regf_0.rf[7][1] ;
 wire \po_0.regf_0.rf[7][2] ;
 wire \po_0.regf_0.rf[7][3] ;
 wire \po_0.regf_0.rf[7][4] ;
 wire \po_0.regf_0.rf[7][5] ;
 wire \po_0.regf_0.rf[7][6] ;
 wire \po_0.regf_0.rf[7][7] ;
 wire \po_0.regf_0.rf[7][8] ;
 wire \po_0.regf_0.rf[7][9] ;
 wire \po_0.regf_0.rf[8][0] ;
 wire \po_0.regf_0.rf[8][10] ;
 wire \po_0.regf_0.rf[8][11] ;
 wire \po_0.regf_0.rf[8][12] ;
 wire \po_0.regf_0.rf[8][13] ;
 wire \po_0.regf_0.rf[8][14] ;
 wire \po_0.regf_0.rf[8][15] ;
 wire \po_0.regf_0.rf[8][1] ;
 wire \po_0.regf_0.rf[8][2] ;
 wire \po_0.regf_0.rf[8][3] ;
 wire \po_0.regf_0.rf[8][4] ;
 wire \po_0.regf_0.rf[8][5] ;
 wire \po_0.regf_0.rf[8][6] ;
 wire \po_0.regf_0.rf[8][7] ;
 wire \po_0.regf_0.rf[8][8] ;
 wire \po_0.regf_0.rf[8][9] ;
 wire \po_0.regf_0.rf[9][0] ;
 wire \po_0.regf_0.rf[9][10] ;
 wire \po_0.regf_0.rf[9][11] ;
 wire \po_0.regf_0.rf[9][12] ;
 wire \po_0.regf_0.rf[9][13] ;
 wire \po_0.regf_0.rf[9][14] ;
 wire \po_0.regf_0.rf[9][15] ;
 wire \po_0.regf_0.rf[9][1] ;
 wire \po_0.regf_0.rf[9][2] ;
 wire \po_0.regf_0.rf[9][3] ;
 wire \po_0.regf_0.rf[9][4] ;
 wire \po_0.regf_0.rf[9][5] ;
 wire \po_0.regf_0.rf[9][6] ;
 wire \po_0.regf_0.rf[9][7] ;
 wire \po_0.regf_0.rf[9][8] ;
 wire \po_0.regf_0.rf[9][9] ;
 wire \po_0.regf_0.rp_addr[0] ;
 wire \po_0.regf_0.rp_addr[1] ;
 wire \po_0.regf_0.rp_addr[2] ;
 wire \po_0.regf_0.rp_addr[3] ;
 wire \po_0.regf_0.rp_rd ;
 wire \po_0.regf_0.rq_addr[0] ;
 wire \po_0.regf_0.rq_addr[1] ;
 wire \po_0.regf_0.rq_addr[2] ;
 wire \po_0.regf_0.rq_addr[3] ;
 wire \po_0.regf_0.rq_rd ;
 wire \po_0.regf_0.w_addr[0] ;
 wire \po_0.regf_0.w_addr[1] ;
 wire \po_0.regf_0.w_addr[2] ;
 wire \po_0.regf_0.w_addr[3] ;
 wire \po_0.regf_0.w_wr ;
 wire \uc_0._00_ ;
 wire \uc_0._01_ ;
 wire \uc_0._02_ ;
 wire \uc_0._03_ ;
 wire \uc_0._20_[10] ;
 wire \uc_0._20_[11] ;
 wire \uc_0._20_[8] ;
 wire \uc_0._20_[9] ;
 wire \uc_0.bc_0._54_[0] ;
 wire \uc_0.bc_0._54_[1] ;
 wire \uc_0.bc_0._54_[2] ;
 wire \uc_0.bc_0._54_[3] ;
 wire \uc_0.bc_0._55_[0] ;
 wire \uc_0.bc_0._55_[1] ;
 wire \uc_0.bc_0._55_[2] ;
 wire \uc_0.bc_0._55_[3] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net83));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__clkbuf_2 _1484_ (.A(\po_0.alu_0.s0 ),
    .X(_1313_));
 sky130_fd_sc_hd__clkbuf_2 _1485_ (.A(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__clkbuf_2 _1486_ (.A(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1487_ (.A(\po_0.alu_0.s1 ),
    .X(_1316_));
 sky130_fd_sc_hd__clkbuf_2 _1488_ (.A(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__buf_2 _1489_ (.A(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1490_ (.A(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__or2b_1 _1491_ (.A(_1315_),
    .B_N(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__clkbuf_1 _1492_ (.A(_1320_),
    .X(_1475_));
 sky130_fd_sc_hd__or2b_1 _1493_ (.A(_1315_),
    .B_N(_1319_),
    .X(_1321_));
 sky130_fd_sc_hd__clkbuf_1 _1494_ (.A(_1321_),
    .X(_1474_));
 sky130_fd_sc_hd__or2b_1 _1495_ (.A(_1315_),
    .B_N(_1319_),
    .X(_1322_));
 sky130_fd_sc_hd__clkbuf_1 _1496_ (.A(_1322_),
    .X(_1473_));
 sky130_fd_sc_hd__or2b_1 _1497_ (.A(_1315_),
    .B_N(_1319_),
    .X(_1323_));
 sky130_fd_sc_hd__clkbuf_1 _1498_ (.A(_1323_),
    .X(_1472_));
 sky130_fd_sc_hd__or2b_1 _1499_ (.A(_1315_),
    .B_N(_1319_),
    .X(_1324_));
 sky130_fd_sc_hd__clkbuf_1 _1500_ (.A(_1324_),
    .X(_1471_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1501_ (.A(_1314_),
    .X(_1325_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1502_ (.A(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__clkbuf_1 _1503_ (.A(_1318_),
    .X(_1327_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1504_ (.A(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__or2b_1 _1505_ (.A(_1326_),
    .B_N(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__clkbuf_1 _1506_ (.A(_1329_),
    .X(_1470_));
 sky130_fd_sc_hd__or2b_1 _1507_ (.A(_1326_),
    .B_N(_1328_),
    .X(_1330_));
 sky130_fd_sc_hd__clkbuf_1 _1508_ (.A(_1330_),
    .X(_1469_));
 sky130_fd_sc_hd__or2b_1 _1509_ (.A(_1326_),
    .B_N(_1328_),
    .X(_1331_));
 sky130_fd_sc_hd__clkbuf_1 _1510_ (.A(_1331_),
    .X(_1468_));
 sky130_fd_sc_hd__or2b_1 _1511_ (.A(_1326_),
    .B_N(_1328_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_1 _1512_ (.A(_1332_),
    .X(_1476_));
 sky130_fd_sc_hd__or2b_1 _1513_ (.A(_1326_),
    .B_N(_1328_),
    .X(_1333_));
 sky130_fd_sc_hd__clkbuf_1 _1514_ (.A(_1333_),
    .X(_1477_));
 sky130_fd_sc_hd__or2b_1 _1515_ (.A(_1326_),
    .B_N(_1328_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_1 _1516_ (.A(_1334_),
    .X(_1478_));
 sky130_fd_sc_hd__or2b_1 _1517_ (.A(_1325_),
    .B_N(_1327_),
    .X(_1335_));
 sky130_fd_sc_hd__clkbuf_1 _1518_ (.A(_1335_),
    .X(_1479_));
 sky130_fd_sc_hd__or2b_1 _1519_ (.A(_1325_),
    .B_N(_1327_),
    .X(_1336_));
 sky130_fd_sc_hd__clkbuf_1 _1520_ (.A(_1336_),
    .X(_1480_));
 sky130_fd_sc_hd__or2b_1 _1521_ (.A(_1325_),
    .B_N(_1327_),
    .X(_1337_));
 sky130_fd_sc_hd__clkbuf_1 _1522_ (.A(_1337_),
    .X(_1481_));
 sky130_fd_sc_hd__or2b_1 _1523_ (.A(_1325_),
    .B_N(_1327_),
    .X(_1338_));
 sky130_fd_sc_hd__clkbuf_1 _1524_ (.A(_1338_),
    .X(_1482_));
 sky130_fd_sc_hd__or2b_1 _1525_ (.A(_1325_),
    .B_N(_1327_),
    .X(_1339_));
 sky130_fd_sc_hd__clkbuf_1 _1526_ (.A(_1339_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_2 _1527_ (.A(net35),
    .X(_1340_));
 sky130_fd_sc_hd__or2_1 _1528_ (.A(\po_0._1_[0] ),
    .B(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__nand2_1 _1529_ (.A(\po_0._1_[0] ),
    .B(_1340_),
    .Y(_1342_));
 sky130_fd_sc_hd__and2_1 _1530_ (.A(_1341_),
    .B(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__clkbuf_1 _1531_ (.A(_1343_),
    .X(\po_0.alu_0._10_[0] ));
 sky130_fd_sc_hd__nor2_1 _1532_ (.A(\uc_0.bc_0._55_[2] ),
    .B(\uc_0.bc_0._55_[3] ),
    .Y(_1344_));
 sky130_fd_sc_hd__and3_1 _1533_ (.A(\uc_0.bc_0._55_[0] ),
    .B(\uc_0.bc_0._55_[1] ),
    .C(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__and4bb_1 _1534_ (.A_N(net80),
    .B_N(net94),
    .C(_1345_),
    .D(net95),
    .X(_1346_));
 sky130_fd_sc_hd__buf_2 _1535_ (.A(net47),
    .X(_1347_));
 sky130_fd_sc_hd__and4bb_1 _1536_ (.A_N(\uc_0.bc_0._55_[1] ),
    .B_N(\uc_0.bc_0._55_[2] ),
    .C(\uc_0.bc_0._55_[3] ),
    .D(\uc_0.bc_0._55_[0] ),
    .X(_1348_));
 sky130_fd_sc_hd__nor4_1 _1537_ (.A(net39),
    .B(net38),
    .C(net41),
    .D(net40),
    .Y(_1349_));
 sky130_fd_sc_hd__nor4_1 _1538_ (.A(net50),
    .B(net83),
    .C(net37),
    .D(net36),
    .Y(_1350_));
 sky130_fd_sc_hd__nand3_1 _1539_ (.A(_1348_),
    .B(_1349_),
    .C(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__or4_2 _1540_ (.A(net35),
    .B(net42),
    .C(net44),
    .D(net43),
    .X(_1352_));
 sky130_fd_sc_hd__or3_1 _1541_ (.A(net46),
    .B(net84),
    .C(net48),
    .X(_1353_));
 sky130_fd_sc_hd__nor4_4 _1542_ (.A(_1347_),
    .B(_1351_),
    .C(_1352_),
    .D(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__nor2_1 _1543_ (.A(_1346_),
    .B(_1354_),
    .Y(_1355_));
 sky130_fd_sc_hd__or2_1 _1544_ (.A(net34),
    .B(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__inv_2 _1545_ (.A(_1356_),
    .Y(\uc_0.bc_0._54_[3] ));
 sky130_fd_sc_hd__clkbuf_2 _1546_ (.A(net34),
    .X(_1357_));
 sky130_fd_sc_hd__a21bo_1 _1547_ (.A1(net80),
    .A2(net95),
    .B1_N(\uc_0.bc_0._55_[0] ),
    .X(_1358_));
 sky130_fd_sc_hd__o311a_1 _1548_ (.A1(net79),
    .A2(net94),
    .A3(_1358_),
    .B1(_1344_),
    .C1(\uc_0.bc_0._55_[1] ),
    .X(_1359_));
 sky130_fd_sc_hd__o21ba_1 _1549_ (.A1(_1344_),
    .A2(_1354_),
    .B1_N(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__clkbuf_2 _1550_ (.A(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__nor2_1 _1551_ (.A(_1357_),
    .B(_1361_),
    .Y(\uc_0.bc_0._54_[0] ));
 sky130_fd_sc_hd__or3b_1 _1552_ (.A(net95),
    .B(net94),
    .C_N(net80),
    .X(_1362_));
 sky130_fd_sc_hd__a311oi_4 _1553_ (.A1(_1362_),
    .A2(\uc_0.bc_0._55_[1] ),
    .A3(\uc_0.bc_0._55_[0] ),
    .B1(\uc_0.bc_0._55_[2] ),
    .C1(\uc_0.bc_0._55_[3] ),
    .Y(_1363_));
 sky130_fd_sc_hd__nor2_1 _1554_ (.A(_1354_),
    .B(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__clkbuf_2 _1555_ (.A(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__nor2_2 _1556_ (.A(net34),
    .B(_1365_),
    .Y(\uc_0.bc_0._54_[1] ));
 sky130_fd_sc_hd__or3b_2 _1557_ (.A(net95),
    .B(net94),
    .C_N(_1345_),
    .X(_1366_));
 sky130_fd_sc_hd__nor2_1 _1558_ (.A(_1357_),
    .B(_1366_),
    .Y(\uc_0.bc_0._54_[2] ));
 sky130_fd_sc_hd__a21oi_2 _1559_ (.A1(_1355_),
    .A2(_1366_),
    .B1(_1357_),
    .Y(_1367_));
 sky130_fd_sc_hd__nor4_4 _1560_ (.A(_1357_),
    .B(_1354_),
    .C(_1361_),
    .D(_1363_),
    .Y(_1368_));
 sky130_fd_sc_hd__nor3b_2 _1561_ (.A(net81),
    .B(net94),
    .C_N(_1345_),
    .Y(_1369_));
 sky130_fd_sc_hd__and3_1 _1562_ (.A(\uc_0.bc_0._54_[3] ),
    .B(_1360_),
    .C(_1364_),
    .X(_1370_));
 sky130_fd_sc_hd__a31o_1 _1563_ (.A1(_1361_),
    .A2(\uc_0.bc_0._54_[1] ),
    .A3(_1369_),
    .B1(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__a21oi_4 _1564_ (.A1(_1367_),
    .A2(_1368_),
    .B1(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__clkbuf_2 _1565_ (.A(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__mux2_1 _1566_ (.A0(\uc_0._20_[8] ),
    .A1(\po_0.regf_0.rp_addr[0] ),
    .S(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_1 _1567_ (.A(_1374_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _1568_ (.A0(\uc_0._20_[9] ),
    .A1(\po_0.regf_0.rp_addr[1] ),
    .S(_1373_),
    .X(_1375_));
 sky130_fd_sc_hd__clkbuf_1 _1569_ (.A(_1375_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _1570_ (.A0(\uc_0._20_[10] ),
    .A1(\po_0.regf_0.rp_addr[2] ),
    .S(_1373_),
    .X(_1376_));
 sky130_fd_sc_hd__clkbuf_1 _1571_ (.A(_1376_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _1572_ (.A0(\uc_0._20_[11] ),
    .A1(\po_0.regf_0.rp_addr[3] ),
    .S(_1373_),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_1 _1573_ (.A(_1377_),
    .X(_0011_));
 sky130_fd_sc_hd__clkbuf_2 _1574_ (.A(_0006_),
    .X(_1378_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1575_ (.A(_0004_),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_4 _1576_ (.A(_1379_),
    .X(_1380_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1577_ (.A(_0005_),
    .X(_1381_));
 sky130_fd_sc_hd__clkbuf_4 _1578_ (.A(_1381_),
    .X(_1382_));
 sky130_fd_sc_hd__mux4_1 _1579_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(\po_0.regf_0.rf[9][0] ),
    .A2(\po_0.regf_0.rf[10][0] ),
    .A3(\po_0.regf_0.rf[11][0] ),
    .S0(_1380_),
    .S1(_1382_),
    .X(_1383_));
 sky130_fd_sc_hd__and2b_1 _1580_ (.A_N(_1378_),
    .B(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__buf_2 _1581_ (.A(_0004_),
    .X(_1385_));
 sky130_fd_sc_hd__clkbuf_4 _1582_ (.A(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__buf_2 _1583_ (.A(_0005_),
    .X(_1387_));
 sky130_fd_sc_hd__buf_2 _1584_ (.A(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__mux4_1 _1585_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(\po_0.regf_0.rf[13][0] ),
    .A2(\po_0.regf_0.rf[14][0] ),
    .A3(\po_0.regf_0.rf[15][0] ),
    .S0(_1386_),
    .S1(_1388_),
    .X(_1389_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1586_ (.A(_0006_),
    .X(_1390_));
 sky130_fd_sc_hd__clkbuf_2 _1587_ (.A(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__clkinv_2 _1588_ (.A(_0007_),
    .Y(_1392_));
 sky130_fd_sc_hd__clkbuf_2 _1589_ (.A(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__a21o_1 _1590_ (.A1(_1389_),
    .A2(_1391_),
    .B1(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__buf_2 _1591_ (.A(_1390_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_4 _1592_ (.A(_1379_),
    .X(_1396_));
 sky130_fd_sc_hd__clkbuf_4 _1593_ (.A(_1381_),
    .X(_1397_));
 sky130_fd_sc_hd__mux4_1 _1594_ (.A0(\po_0.regf_0.rf[0][0] ),
    .A1(\po_0.regf_0.rf[1][0] ),
    .A2(\po_0.regf_0.rf[2][0] ),
    .A3(\po_0.regf_0.rf[3][0] ),
    .S0(_1396_),
    .S1(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__and2b_1 _1595_ (.A_N(_1395_),
    .B(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_4 _1596_ (.A(_1385_),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_4 _1597_ (.A(_1387_),
    .X(_1401_));
 sky130_fd_sc_hd__mux4_1 _1598_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(\po_0.regf_0.rf[5][0] ),
    .A2(\po_0.regf_0.rf[6][0] ),
    .A3(\po_0.regf_0.rf[7][0] ),
    .S0(_1400_),
    .S1(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__buf_2 _1599_ (.A(_1390_),
    .X(_1403_));
 sky130_fd_sc_hd__buf_2 _1600_ (.A(_0007_),
    .X(_1404_));
 sky130_fd_sc_hd__a21o_1 _1601_ (.A1(_1402_),
    .A2(_1403_),
    .B1(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__o22a_1 _1602_ (.A1(_1384_),
    .A2(_1394_),
    .B1(_1399_),
    .B2(_1405_),
    .X(\po_0.regf_0._5_[0] ));
 sky130_fd_sc_hd__clkbuf_4 _1603_ (.A(_1379_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_4 _1604_ (.A(_1381_),
    .X(_1407_));
 sky130_fd_sc_hd__mux4_1 _1605_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(\po_0.regf_0.rf[5][1] ),
    .A2(\po_0.regf_0.rf[6][1] ),
    .A3(\po_0.regf_0.rf[7][1] ),
    .S0(_1406_),
    .S1(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_2 _1606_ (.A(_1390_),
    .X(_1409_));
 sky130_fd_sc_hd__a21o_1 _1607_ (.A1(_1408_),
    .A2(_1409_),
    .B1(_0007_),
    .X(_1410_));
 sky130_fd_sc_hd__clkbuf_2 _1608_ (.A(_1390_),
    .X(_1411_));
 sky130_fd_sc_hd__clkbuf_4 _1609_ (.A(_1379_),
    .X(_1412_));
 sky130_fd_sc_hd__buf_2 _1610_ (.A(_1381_),
    .X(_1413_));
 sky130_fd_sc_hd__mux4_1 _1611_ (.A0(\po_0.regf_0.rf[0][1] ),
    .A1(\po_0.regf_0.rf[1][1] ),
    .A2(\po_0.regf_0.rf[2][1] ),
    .A3(\po_0.regf_0.rf[3][1] ),
    .S0(_1412_),
    .S1(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__and2b_1 _1612_ (.A_N(_1411_),
    .B(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__mux4_1 _1613_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(\po_0.regf_0.rf[13][1] ),
    .A2(\po_0.regf_0.rf[14][1] ),
    .A3(\po_0.regf_0.rf[15][1] ),
    .S0(_1386_),
    .S1(_1388_),
    .X(_1416_));
 sky130_fd_sc_hd__a21o_1 _1614_ (.A1(_1416_),
    .A2(_1391_),
    .B1(_1393_),
    .X(_1417_));
 sky130_fd_sc_hd__clkbuf_2 _1615_ (.A(_1390_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_4 _1616_ (.A(_1379_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_4 _1617_ (.A(_1381_),
    .X(_1420_));
 sky130_fd_sc_hd__mux4_1 _1618_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(\po_0.regf_0.rf[9][1] ),
    .A2(\po_0.regf_0.rf[10][1] ),
    .A3(\po_0.regf_0.rf[11][1] ),
    .S0(_1419_),
    .S1(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__and2b_1 _1619_ (.A_N(_1418_),
    .B(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__o22a_1 _1620_ (.A1(_1410_),
    .A2(_1415_),
    .B1(_1417_),
    .B2(_1422_),
    .X(\po_0.regf_0._5_[1] ));
 sky130_fd_sc_hd__mux4_1 _1621_ (.A0(\po_0.regf_0.rf[0][2] ),
    .A1(\po_0.regf_0.rf[1][2] ),
    .A2(\po_0.regf_0.rf[2][2] ),
    .A3(\po_0.regf_0.rf[3][2] ),
    .S0(_1380_),
    .S1(_1382_),
    .X(_1423_));
 sky130_fd_sc_hd__and2b_1 _1622_ (.A_N(_1378_),
    .B(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__mux4_1 _1623_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(\po_0.regf_0.rf[5][2] ),
    .A2(\po_0.regf_0.rf[6][2] ),
    .A3(\po_0.regf_0.rf[7][2] ),
    .S0(_1386_),
    .S1(_1388_),
    .X(_1425_));
 sky130_fd_sc_hd__a21o_1 _1624_ (.A1(_1425_),
    .A2(_1391_),
    .B1(_0007_),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_4 _1625_ (.A(_1379_),
    .X(_1427_));
 sky130_fd_sc_hd__buf_2 _1626_ (.A(_1381_),
    .X(_1428_));
 sky130_fd_sc_hd__mux4_1 _1627_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(\po_0.regf_0.rf[9][2] ),
    .A2(\po_0.regf_0.rf[10][2] ),
    .A3(\po_0.regf_0.rf[11][2] ),
    .S0(_1427_),
    .S1(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__buf_4 _1628_ (.A(_0004_),
    .X(_1430_));
 sky130_fd_sc_hd__clkbuf_4 _1629_ (.A(_0005_),
    .X(_1431_));
 sky130_fd_sc_hd__mux4_1 _1630_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(\po_0.regf_0.rf[13][2] ),
    .A2(\po_0.regf_0.rf[14][2] ),
    .A3(\po_0.regf_0.rf[15][2] ),
    .S0(_1430_),
    .S1(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__buf_2 _1631_ (.A(_0006_),
    .X(_1433_));
 sky130_fd_sc_hd__mux2_1 _1632_ (.A0(_1429_),
    .A1(_1432_),
    .S(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__o22a_1 _1633_ (.A1(_1424_),
    .A2(_1426_),
    .B1(_1393_),
    .B2(_1434_),
    .X(\po_0.regf_0._5_[2] ));
 sky130_fd_sc_hd__mux4_1 _1634_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(\po_0.regf_0.rf[13][3] ),
    .A2(\po_0.regf_0.rf[14][3] ),
    .A3(\po_0.regf_0.rf[15][3] ),
    .S0(_1406_),
    .S1(_1407_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_2 _1635_ (.A(_1392_),
    .X(_1436_));
 sky130_fd_sc_hd__a21o_1 _1636_ (.A1(_1435_),
    .A2(_1409_),
    .B1(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__mux4_1 _1637_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(\po_0.regf_0.rf[9][3] ),
    .A2(\po_0.regf_0.rf[10][3] ),
    .A3(\po_0.regf_0.rf[11][3] ),
    .S0(_1412_),
    .S1(_1413_),
    .X(_1438_));
 sky130_fd_sc_hd__and2b_1 _1638_ (.A_N(_1411_),
    .B(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__buf_2 _1639_ (.A(_0007_),
    .X(_1440_));
 sky130_fd_sc_hd__mux4_1 _1640_ (.A0(\po_0.regf_0.rf[0][3] ),
    .A1(\po_0.regf_0.rf[1][3] ),
    .A2(\po_0.regf_0.rf[2][3] ),
    .A3(\po_0.regf_0.rf[3][3] ),
    .S0(_1427_),
    .S1(_1428_),
    .X(_1441_));
 sky130_fd_sc_hd__buf_4 _1641_ (.A(_0004_),
    .X(_1442_));
 sky130_fd_sc_hd__clkbuf_4 _1642_ (.A(_0005_),
    .X(_1443_));
 sky130_fd_sc_hd__mux4_1 _1643_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(\po_0.regf_0.rf[5][3] ),
    .A2(\po_0.regf_0.rf[6][3] ),
    .A3(\po_0.regf_0.rf[7][3] ),
    .S0(_1442_),
    .S1(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_4 _1644_ (.A(_0006_),
    .X(_1445_));
 sky130_fd_sc_hd__mux2_1 _1645_ (.A0(_1441_),
    .A1(_1444_),
    .S(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__o22a_1 _1646_ (.A1(_1437_),
    .A2(_1439_),
    .B1(_1440_),
    .B2(_1446_),
    .X(\po_0.regf_0._5_[3] ));
 sky130_fd_sc_hd__mux4_1 _1647_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(\po_0.regf_0.rf[9][4] ),
    .A2(\po_0.regf_0.rf[10][4] ),
    .A3(\po_0.regf_0.rf[11][4] ),
    .S0(_1380_),
    .S1(_1382_),
    .X(_1447_));
 sky130_fd_sc_hd__and2b_1 _1648_ (.A_N(_1433_),
    .B(_1447_),
    .X(_1448_));
 sky130_fd_sc_hd__mux4_1 _1649_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(\po_0.regf_0.rf[13][4] ),
    .A2(\po_0.regf_0.rf[14][4] ),
    .A3(\po_0.regf_0.rf[15][4] ),
    .S0(_1386_),
    .S1(_1388_),
    .X(_1449_));
 sky130_fd_sc_hd__a21o_1 _1650_ (.A1(_1449_),
    .A2(_1391_),
    .B1(_1393_),
    .X(_1450_));
 sky130_fd_sc_hd__mux4_1 _1651_ (.A0(\po_0.regf_0.rf[0][4] ),
    .A1(\po_0.regf_0.rf[1][4] ),
    .A2(\po_0.regf_0.rf[2][4] ),
    .A3(\po_0.regf_0.rf[3][4] ),
    .S0(_1396_),
    .S1(_1397_),
    .X(_1451_));
 sky130_fd_sc_hd__and2b_1 _1652_ (.A_N(_1395_),
    .B(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__mux4_1 _1653_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(\po_0.regf_0.rf[5][4] ),
    .A2(\po_0.regf_0.rf[6][4] ),
    .A3(\po_0.regf_0.rf[7][4] ),
    .S0(_1400_),
    .S1(_1401_),
    .X(_1453_));
 sky130_fd_sc_hd__a21o_1 _1654_ (.A1(_1453_),
    .A2(_1403_),
    .B1(_1404_),
    .X(_1454_));
 sky130_fd_sc_hd__o22a_1 _1655_ (.A1(_1448_),
    .A2(_1450_),
    .B1(_1452_),
    .B2(_1454_),
    .X(\po_0.regf_0._5_[4] ));
 sky130_fd_sc_hd__mux4_1 _1656_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(\po_0.regf_0.rf[13][5] ),
    .A2(\po_0.regf_0.rf[14][5] ),
    .A3(\po_0.regf_0.rf[15][5] ),
    .S0(_1406_),
    .S1(_1407_),
    .X(_1455_));
 sky130_fd_sc_hd__a21o_1 _1657_ (.A1(_1455_),
    .A2(_1409_),
    .B1(_1436_),
    .X(_1456_));
 sky130_fd_sc_hd__mux4_1 _1658_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(\po_0.regf_0.rf[9][5] ),
    .A2(\po_0.regf_0.rf[10][5] ),
    .A3(\po_0.regf_0.rf[11][5] ),
    .S0(_1412_),
    .S1(_1413_),
    .X(_1457_));
 sky130_fd_sc_hd__and2b_1 _1659_ (.A_N(_1411_),
    .B(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__mux4_1 _1660_ (.A0(\po_0.regf_0.rf[0][5] ),
    .A1(\po_0.regf_0.rf[1][5] ),
    .A2(\po_0.regf_0.rf[2][5] ),
    .A3(\po_0.regf_0.rf[3][5] ),
    .S0(_1430_),
    .S1(_1431_),
    .X(_1459_));
 sky130_fd_sc_hd__mux4_1 _1661_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(\po_0.regf_0.rf[5][5] ),
    .A2(\po_0.regf_0.rf[6][5] ),
    .A3(\po_0.regf_0.rf[7][5] ),
    .S0(_1442_),
    .S1(_1443_),
    .X(_1460_));
 sky130_fd_sc_hd__mux2_1 _1662_ (.A0(_1459_),
    .A1(_1460_),
    .S(_1445_),
    .X(_1461_));
 sky130_fd_sc_hd__o22a_1 _1663_ (.A1(_1456_),
    .A2(_1458_),
    .B1(_1440_),
    .B2(_1461_),
    .X(\po_0.regf_0._5_[5] ));
 sky130_fd_sc_hd__mux4_1 _1664_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(\po_0.regf_0.rf[9][6] ),
    .A2(\po_0.regf_0.rf[10][6] ),
    .A3(\po_0.regf_0.rf[11][6] ),
    .S0(_1427_),
    .S1(_1428_),
    .X(_1462_));
 sky130_fd_sc_hd__and2b_1 _1665_ (.A_N(_1433_),
    .B(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__mux4_1 _1666_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(\po_0.regf_0.rf[13][6] ),
    .A2(\po_0.regf_0.rf[14][6] ),
    .A3(\po_0.regf_0.rf[15][6] ),
    .S0(_1386_),
    .S1(_1388_),
    .X(_1464_));
 sky130_fd_sc_hd__a21o_1 _1667_ (.A1(_1464_),
    .A2(_1391_),
    .B1(_1393_),
    .X(_1465_));
 sky130_fd_sc_hd__mux4_1 _1668_ (.A0(\po_0.regf_0.rf[0][6] ),
    .A1(\po_0.regf_0.rf[1][6] ),
    .A2(\po_0.regf_0.rf[2][6] ),
    .A3(\po_0.regf_0.rf[3][6] ),
    .S0(_1396_),
    .S1(_1397_),
    .X(_1466_));
 sky130_fd_sc_hd__and2b_1 _1669_ (.A_N(_1395_),
    .B(_1466_),
    .X(_1467_));
 sky130_fd_sc_hd__mux4_1 _1670_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(\po_0.regf_0.rf[5][6] ),
    .A2(\po_0.regf_0.rf[6][6] ),
    .A3(\po_0.regf_0.rf[7][6] ),
    .S0(_1400_),
    .S1(_1401_),
    .X(_0338_));
 sky130_fd_sc_hd__a21o_1 _1671_ (.A1(_0338_),
    .A2(_1403_),
    .B1(_1404_),
    .X(_0339_));
 sky130_fd_sc_hd__o22a_1 _1672_ (.A1(_1463_),
    .A2(_1465_),
    .B1(_1467_),
    .B2(_0339_),
    .X(\po_0.regf_0._5_[6] ));
 sky130_fd_sc_hd__mux4_1 _1673_ (.A0(\po_0.regf_0.rf[8][7] ),
    .A1(\po_0.regf_0.rf[9][7] ),
    .A2(\po_0.regf_0.rf[10][7] ),
    .A3(\po_0.regf_0.rf[11][7] ),
    .S0(_1427_),
    .S1(_1428_),
    .X(_0340_));
 sky130_fd_sc_hd__and2b_1 _1674_ (.A_N(_1433_),
    .B(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__mux4_1 _1675_ (.A0(\po_0.regf_0.rf[12][7] ),
    .A1(\po_0.regf_0.rf[13][7] ),
    .A2(\po_0.regf_0.rf[14][7] ),
    .A3(\po_0.regf_0.rf[15][7] ),
    .S0(_1406_),
    .S1(_1407_),
    .X(_0342_));
 sky130_fd_sc_hd__a21o_1 _1676_ (.A1(_0342_),
    .A2(_1418_),
    .B1(_1436_),
    .X(_0343_));
 sky130_fd_sc_hd__mux4_1 _1677_ (.A0(\po_0.regf_0.rf[0][7] ),
    .A1(\po_0.regf_0.rf[1][7] ),
    .A2(\po_0.regf_0.rf[2][7] ),
    .A3(\po_0.regf_0.rf[3][7] ),
    .S0(_1396_),
    .S1(_1397_),
    .X(_0344_));
 sky130_fd_sc_hd__and2b_1 _1678_ (.A_N(_1395_),
    .B(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__mux4_1 _1679_ (.A0(\po_0.regf_0.rf[4][7] ),
    .A1(\po_0.regf_0.rf[5][7] ),
    .A2(\po_0.regf_0.rf[6][7] ),
    .A3(\po_0.regf_0.rf[7][7] ),
    .S0(_1400_),
    .S1(_1401_),
    .X(_0346_));
 sky130_fd_sc_hd__a21o_1 _1680_ (.A1(_0346_),
    .A2(_1403_),
    .B1(_1404_),
    .X(_0347_));
 sky130_fd_sc_hd__o22a_1 _1681_ (.A1(_0341_),
    .A2(_0343_),
    .B1(_0345_),
    .B2(_0347_),
    .X(\po_0.regf_0._5_[7] ));
 sky130_fd_sc_hd__mux4_1 _1682_ (.A0(\po_0.regf_0.rf[8][8] ),
    .A1(\po_0.regf_0.rf[9][8] ),
    .A2(\po_0.regf_0.rf[10][8] ),
    .A3(\po_0.regf_0.rf[11][8] ),
    .S0(_1385_),
    .S1(_1387_),
    .X(_0348_));
 sky130_fd_sc_hd__mux4_1 _1683_ (.A0(\po_0.regf_0.rf[0][8] ),
    .A1(\po_0.regf_0.rf[1][8] ),
    .A2(\po_0.regf_0.rf[2][8] ),
    .A3(\po_0.regf_0.rf[3][8] ),
    .S0(_1385_),
    .S1(_1387_),
    .X(_0349_));
 sky130_fd_sc_hd__mux4_1 _1684_ (.A0(\po_0.regf_0.rf[12][8] ),
    .A1(\po_0.regf_0.rf[13][8] ),
    .A2(\po_0.regf_0.rf[14][8] ),
    .A3(\po_0.regf_0.rf[15][8] ),
    .S0(_1385_),
    .S1(_1387_),
    .X(_0350_));
 sky130_fd_sc_hd__mux4_1 _1685_ (.A0(\po_0.regf_0.rf[4][8] ),
    .A1(\po_0.regf_0.rf[5][8] ),
    .A2(\po_0.regf_0.rf[6][8] ),
    .A3(\po_0.regf_0.rf[7][8] ),
    .S0(_1385_),
    .S1(_1387_),
    .X(_0351_));
 sky130_fd_sc_hd__mux4_1 _1686_ (.A0(_0348_),
    .A1(_0349_),
    .A2(_0350_),
    .A3(_0351_),
    .S0(_1392_),
    .S1(_1418_),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_1 _1687_ (.A(_0352_),
    .X(\po_0.regf_0._5_[8] ));
 sky130_fd_sc_hd__mux4_1 _1688_ (.A0(\po_0.regf_0.rf[12][9] ),
    .A1(\po_0.regf_0.rf[13][9] ),
    .A2(\po_0.regf_0.rf[14][9] ),
    .A3(\po_0.regf_0.rf[15][9] ),
    .S0(_1419_),
    .S1(_1420_),
    .X(_0353_));
 sky130_fd_sc_hd__a21o_1 _1689_ (.A1(_0353_),
    .A2(_1409_),
    .B1(_1436_),
    .X(_0354_));
 sky130_fd_sc_hd__mux4_1 _1690_ (.A0(\po_0.regf_0.rf[8][9] ),
    .A1(\po_0.regf_0.rf[9][9] ),
    .A2(\po_0.regf_0.rf[10][9] ),
    .A3(\po_0.regf_0.rf[11][9] ),
    .S0(_1412_),
    .S1(_1413_),
    .X(_0355_));
 sky130_fd_sc_hd__and2b_1 _1691_ (.A_N(_1411_),
    .B(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__mux4_1 _1692_ (.A0(\po_0.regf_0.rf[0][9] ),
    .A1(\po_0.regf_0.rf[1][9] ),
    .A2(\po_0.regf_0.rf[2][9] ),
    .A3(\po_0.regf_0.rf[3][9] ),
    .S0(_1430_),
    .S1(_1431_),
    .X(_0357_));
 sky130_fd_sc_hd__mux4_1 _1693_ (.A0(\po_0.regf_0.rf[4][9] ),
    .A1(\po_0.regf_0.rf[5][9] ),
    .A2(\po_0.regf_0.rf[6][9] ),
    .A3(\po_0.regf_0.rf[7][9] ),
    .S0(_1442_),
    .S1(_1443_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _1694_ (.A0(_0357_),
    .A1(_0358_),
    .S(_1445_),
    .X(_0359_));
 sky130_fd_sc_hd__o22a_1 _1695_ (.A1(_0354_),
    .A2(_0356_),
    .B1(_1440_),
    .B2(_0359_),
    .X(\po_0.regf_0._5_[9] ));
 sky130_fd_sc_hd__mux4_1 _1696_ (.A0(\po_0.regf_0.rf[12][10] ),
    .A1(\po_0.regf_0.rf[13][10] ),
    .A2(\po_0.regf_0.rf[14][10] ),
    .A3(\po_0.regf_0.rf[15][10] ),
    .S0(_1419_),
    .S1(_1420_),
    .X(_0360_));
 sky130_fd_sc_hd__a21o_1 _1697_ (.A1(_0360_),
    .A2(_1409_),
    .B1(_1392_),
    .X(_0361_));
 sky130_fd_sc_hd__mux4_1 _1698_ (.A0(\po_0.regf_0.rf[8][10] ),
    .A1(\po_0.regf_0.rf[9][10] ),
    .A2(\po_0.regf_0.rf[10][10] ),
    .A3(\po_0.regf_0.rf[11][10] ),
    .S0(_1412_),
    .S1(_1413_),
    .X(_0362_));
 sky130_fd_sc_hd__and2b_1 _1699_ (.A_N(_1378_),
    .B(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__mux4_1 _1700_ (.A0(\po_0.regf_0.rf[0][10] ),
    .A1(\po_0.regf_0.rf[1][10] ),
    .A2(\po_0.regf_0.rf[2][10] ),
    .A3(\po_0.regf_0.rf[3][10] ),
    .S0(_1430_),
    .S1(_1431_),
    .X(_0364_));
 sky130_fd_sc_hd__mux4_1 _1701_ (.A0(\po_0.regf_0.rf[4][10] ),
    .A1(\po_0.regf_0.rf[5][10] ),
    .A2(\po_0.regf_0.rf[6][10] ),
    .A3(\po_0.regf_0.rf[7][10] ),
    .S0(_1442_),
    .S1(_1443_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _1702_ (.A0(_0364_),
    .A1(_0365_),
    .S(_1445_),
    .X(_0366_));
 sky130_fd_sc_hd__o22a_1 _1703_ (.A1(_0361_),
    .A2(_0363_),
    .B1(_1440_),
    .B2(_0366_),
    .X(\po_0.regf_0._5_[10] ));
 sky130_fd_sc_hd__mux4_1 _1704_ (.A0(\po_0.regf_0.rf[4][11] ),
    .A1(\po_0.regf_0.rf[5][11] ),
    .A2(\po_0.regf_0.rf[6][11] ),
    .A3(\po_0.regf_0.rf[7][11] ),
    .S0(_1419_),
    .S1(_1420_),
    .X(_0367_));
 sky130_fd_sc_hd__a21o_1 _1705_ (.A1(_0367_),
    .A2(_1409_),
    .B1(_0007_),
    .X(_0368_));
 sky130_fd_sc_hd__mux4_1 _1706_ (.A0(\po_0.regf_0.rf[0][11] ),
    .A1(\po_0.regf_0.rf[1][11] ),
    .A2(\po_0.regf_0.rf[2][11] ),
    .A3(\po_0.regf_0.rf[3][11] ),
    .S0(_1380_),
    .S1(_1382_),
    .X(_0369_));
 sky130_fd_sc_hd__and2b_1 _1707_ (.A_N(_1378_),
    .B(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__mux4_1 _1708_ (.A0(\po_0.regf_0.rf[12][11] ),
    .A1(\po_0.regf_0.rf[13][11] ),
    .A2(\po_0.regf_0.rf[14][11] ),
    .A3(\po_0.regf_0.rf[15][11] ),
    .S0(_1386_),
    .S1(_1388_),
    .X(_0371_));
 sky130_fd_sc_hd__a21o_1 _1709_ (.A1(_0371_),
    .A2(_1391_),
    .B1(_1393_),
    .X(_0372_));
 sky130_fd_sc_hd__mux4_1 _1710_ (.A0(\po_0.regf_0.rf[8][11] ),
    .A1(\po_0.regf_0.rf[9][11] ),
    .A2(\po_0.regf_0.rf[10][11] ),
    .A3(\po_0.regf_0.rf[11][11] ),
    .S0(_1396_),
    .S1(_1397_),
    .X(_0373_));
 sky130_fd_sc_hd__and2b_1 _1711_ (.A_N(_1418_),
    .B(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__o22a_1 _1712_ (.A1(_0368_),
    .A2(_0370_),
    .B1(_0372_),
    .B2(_0374_),
    .X(\po_0.regf_0._5_[11] ));
 sky130_fd_sc_hd__mux4_1 _1713_ (.A0(\po_0.regf_0.rf[8][12] ),
    .A1(\po_0.regf_0.rf[9][12] ),
    .A2(\po_0.regf_0.rf[10][12] ),
    .A3(\po_0.regf_0.rf[11][12] ),
    .S0(_1427_),
    .S1(_1428_),
    .X(_0375_));
 sky130_fd_sc_hd__and2b_1 _1714_ (.A_N(_1433_),
    .B(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__mux4_1 _1715_ (.A0(\po_0.regf_0.rf[12][12] ),
    .A1(\po_0.regf_0.rf[13][12] ),
    .A2(\po_0.regf_0.rf[14][12] ),
    .A3(\po_0.regf_0.rf[15][12] ),
    .S0(_1406_),
    .S1(_1407_),
    .X(_0377_));
 sky130_fd_sc_hd__a21o_1 _1716_ (.A1(_0377_),
    .A2(_1418_),
    .B1(_1436_),
    .X(_0378_));
 sky130_fd_sc_hd__mux4_1 _1717_ (.A0(\po_0.regf_0.rf[0][12] ),
    .A1(\po_0.regf_0.rf[1][12] ),
    .A2(\po_0.regf_0.rf[2][12] ),
    .A3(\po_0.regf_0.rf[3][12] ),
    .S0(_1396_),
    .S1(_1397_),
    .X(_0379_));
 sky130_fd_sc_hd__and2b_1 _1718_ (.A_N(_1411_),
    .B(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__mux4_1 _1719_ (.A0(\po_0.regf_0.rf[4][12] ),
    .A1(\po_0.regf_0.rf[5][12] ),
    .A2(\po_0.regf_0.rf[6][12] ),
    .A3(\po_0.regf_0.rf[7][12] ),
    .S0(_1400_),
    .S1(_1401_),
    .X(_0381_));
 sky130_fd_sc_hd__a21o_1 _1720_ (.A1(_0381_),
    .A2(_1403_),
    .B1(_1404_),
    .X(_0382_));
 sky130_fd_sc_hd__o22a_1 _1721_ (.A1(_0376_),
    .A2(_0378_),
    .B1(_0380_),
    .B2(_0382_),
    .X(\po_0.regf_0._5_[12] ));
 sky130_fd_sc_hd__mux4_1 _1722_ (.A0(\po_0.regf_0.rf[12][13] ),
    .A1(\po_0.regf_0.rf[13][13] ),
    .A2(\po_0.regf_0.rf[14][13] ),
    .A3(\po_0.regf_0.rf[15][13] ),
    .S0(_1419_),
    .S1(_1420_),
    .X(_0383_));
 sky130_fd_sc_hd__a21o_1 _1723_ (.A1(_0383_),
    .A2(_1395_),
    .B1(_1392_),
    .X(_0384_));
 sky130_fd_sc_hd__mux4_1 _1724_ (.A0(\po_0.regf_0.rf[8][13] ),
    .A1(\po_0.regf_0.rf[9][13] ),
    .A2(\po_0.regf_0.rf[10][13] ),
    .A3(\po_0.regf_0.rf[11][13] ),
    .S0(_1380_),
    .S1(_1382_),
    .X(_0385_));
 sky130_fd_sc_hd__and2b_1 _1725_ (.A_N(_1378_),
    .B(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__mux4_1 _1726_ (.A0(\po_0.regf_0.rf[0][13] ),
    .A1(\po_0.regf_0.rf[1][13] ),
    .A2(\po_0.regf_0.rf[2][13] ),
    .A3(\po_0.regf_0.rf[3][13] ),
    .S0(_1430_),
    .S1(_1431_),
    .X(_0387_));
 sky130_fd_sc_hd__mux4_1 _1727_ (.A0(\po_0.regf_0.rf[4][13] ),
    .A1(\po_0.regf_0.rf[5][13] ),
    .A2(\po_0.regf_0.rf[6][13] ),
    .A3(\po_0.regf_0.rf[7][13] ),
    .S0(_1442_),
    .S1(_1443_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _1728_ (.A0(_0387_),
    .A1(_0388_),
    .S(_1445_),
    .X(_0389_));
 sky130_fd_sc_hd__o22a_1 _1729_ (.A1(_0384_),
    .A2(_0386_),
    .B1(_1440_),
    .B2(_0389_),
    .X(\po_0.regf_0._5_[13] ));
 sky130_fd_sc_hd__mux4_1 _1730_ (.A0(\po_0.regf_0.rf[12][14] ),
    .A1(\po_0.regf_0.rf[13][14] ),
    .A2(\po_0.regf_0.rf[14][14] ),
    .A3(\po_0.regf_0.rf[15][14] ),
    .S0(_1419_),
    .S1(_1420_),
    .X(_0390_));
 sky130_fd_sc_hd__a21o_1 _1731_ (.A1(_0390_),
    .A2(_1395_),
    .B1(_1392_),
    .X(_0391_));
 sky130_fd_sc_hd__mux4_1 _1732_ (.A0(\po_0.regf_0.rf[8][14] ),
    .A1(\po_0.regf_0.rf[9][14] ),
    .A2(\po_0.regf_0.rf[10][14] ),
    .A3(\po_0.regf_0.rf[11][14] ),
    .S0(_1380_),
    .S1(_1382_),
    .X(_0392_));
 sky130_fd_sc_hd__and2b_1 _1733_ (.A_N(_1378_),
    .B(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__mux4_1 _1734_ (.A0(\po_0.regf_0.rf[0][14] ),
    .A1(\po_0.regf_0.rf[1][14] ),
    .A2(\po_0.regf_0.rf[2][14] ),
    .A3(\po_0.regf_0.rf[3][14] ),
    .S0(_1430_),
    .S1(_1431_),
    .X(_0394_));
 sky130_fd_sc_hd__mux4_1 _1735_ (.A0(\po_0.regf_0.rf[4][14] ),
    .A1(\po_0.regf_0.rf[5][14] ),
    .A2(\po_0.regf_0.rf[6][14] ),
    .A3(\po_0.regf_0.rf[7][14] ),
    .S0(_1442_),
    .S1(_1443_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _1736_ (.A0(_0394_),
    .A1(_0395_),
    .S(_1445_),
    .X(_0396_));
 sky130_fd_sc_hd__o22a_1 _1737_ (.A1(_0391_),
    .A2(_0393_),
    .B1(_1440_),
    .B2(_0396_),
    .X(\po_0.regf_0._5_[14] ));
 sky130_fd_sc_hd__mux4_1 _1738_ (.A0(\po_0.regf_0.rf[8][15] ),
    .A1(\po_0.regf_0.rf[9][15] ),
    .A2(\po_0.regf_0.rf[10][15] ),
    .A3(\po_0.regf_0.rf[11][15] ),
    .S0(_1427_),
    .S1(_1428_),
    .X(_0397_));
 sky130_fd_sc_hd__and2b_1 _1739_ (.A_N(_1433_),
    .B(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__mux4_1 _1740_ (.A0(\po_0.regf_0.rf[12][15] ),
    .A1(\po_0.regf_0.rf[13][15] ),
    .A2(\po_0.regf_0.rf[14][15] ),
    .A3(\po_0.regf_0.rf[15][15] ),
    .S0(_1406_),
    .S1(_1407_),
    .X(_0399_));
 sky130_fd_sc_hd__a21o_1 _1741_ (.A1(_0399_),
    .A2(_1418_),
    .B1(_1436_),
    .X(_0400_));
 sky130_fd_sc_hd__mux4_1 _1742_ (.A0(\po_0.regf_0.rf[0][15] ),
    .A1(\po_0.regf_0.rf[1][15] ),
    .A2(\po_0.regf_0.rf[2][15] ),
    .A3(\po_0.regf_0.rf[3][15] ),
    .S0(_1412_),
    .S1(_1413_),
    .X(_0401_));
 sky130_fd_sc_hd__and2b_1 _1743_ (.A_N(_1411_),
    .B(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__mux4_1 _1744_ (.A0(\po_0.regf_0.rf[4][15] ),
    .A1(\po_0.regf_0.rf[5][15] ),
    .A2(\po_0.regf_0.rf[6][15] ),
    .A3(\po_0.regf_0.rf[7][15] ),
    .S0(_1400_),
    .S1(_1401_),
    .X(_0403_));
 sky130_fd_sc_hd__a21o_1 _1745_ (.A1(_0403_),
    .A2(_1403_),
    .B1(_1404_),
    .X(_0404_));
 sky130_fd_sc_hd__o22a_1 _1746_ (.A1(_0398_),
    .A2(_0400_),
    .B1(_0402_),
    .B2(_0404_),
    .X(\po_0.regf_0._5_[15] ));
 sky130_fd_sc_hd__clkbuf_2 _1747_ (.A(_0000_),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_4 _1748_ (.A(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_2 _1749_ (.A(_0001_),
    .X(_0407_));
 sky130_fd_sc_hd__buf_2 _1750_ (.A(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__mux4_1 _1751_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(\po_0.regf_0.rf[13][0] ),
    .A2(\po_0.regf_0.rf[14][0] ),
    .A3(\po_0.regf_0.rf[15][0] ),
    .S0(_0406_),
    .S1(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__buf_2 _1752_ (.A(_0002_),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_2 _1753_ (.A(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_2 _1754_ (.A(_0003_),
    .X(_0412_));
 sky130_fd_sc_hd__a21bo_1 _1755_ (.A1(_0409_),
    .A2(_0411_),
    .B1_N(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__buf_2 _1756_ (.A(_0002_),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_2 _1757_ (.A(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_4 _1758_ (.A(_0405_),
    .X(_0416_));
 sky130_fd_sc_hd__buf_2 _1759_ (.A(_0407_),
    .X(_0417_));
 sky130_fd_sc_hd__mux4_1 _1760_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(\po_0.regf_0.rf[9][0] ),
    .A2(\po_0.regf_0.rf[10][0] ),
    .A3(\po_0.regf_0.rf[11][0] ),
    .S0(_0416_),
    .S1(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__and2b_1 _1761_ (.A_N(_0415_),
    .B(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__buf_2 _1762_ (.A(_0003_),
    .X(_0420_));
 sky130_fd_sc_hd__buf_2 _1763_ (.A(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__buf_2 _1764_ (.A(_0000_),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_4 _1765_ (.A(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__buf_2 _1766_ (.A(_0001_),
    .X(_0424_));
 sky130_fd_sc_hd__buf_2 _1767_ (.A(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__mux4_1 _1768_ (.A0(\po_0.regf_0.rf[0][0] ),
    .A1(\po_0.regf_0.rf[1][0] ),
    .A2(\po_0.regf_0.rf[2][0] ),
    .A3(\po_0.regf_0.rf[3][0] ),
    .S0(_0423_),
    .S1(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__buf_4 _1769_ (.A(_0422_),
    .X(_0427_));
 sky130_fd_sc_hd__buf_4 _1770_ (.A(_0424_),
    .X(_0428_));
 sky130_fd_sc_hd__mux4_1 _1771_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(\po_0.regf_0.rf[5][0] ),
    .A2(\po_0.regf_0.rf[6][0] ),
    .A3(\po_0.regf_0.rf[7][0] ),
    .S0(_0427_),
    .S1(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_2 _1772_ (.A(_0414_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _1773_ (.A0(_0426_),
    .A1(_0429_),
    .S(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__o22a_1 _1774_ (.A1(_0413_),
    .A2(_0419_),
    .B1(_0421_),
    .B2(_0431_),
    .X(\po_0.regf_0._3_[0] ));
 sky130_fd_sc_hd__mux4_1 _1775_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(\po_0.regf_0.rf[13][1] ),
    .A2(\po_0.regf_0.rf[14][1] ),
    .A3(\po_0.regf_0.rf[15][1] ),
    .S0(_0406_),
    .S1(_0408_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_2 _1776_ (.A(_0410_),
    .X(_0433_));
 sky130_fd_sc_hd__a21bo_1 _1777_ (.A1(_0432_),
    .A2(_0433_),
    .B1_N(_0412_),
    .X(_0434_));
 sky130_fd_sc_hd__mux4_1 _1778_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(\po_0.regf_0.rf[9][1] ),
    .A2(\po_0.regf_0.rf[10][1] ),
    .A3(\po_0.regf_0.rf[11][1] ),
    .S0(_0416_),
    .S1(_0417_),
    .X(_0435_));
 sky130_fd_sc_hd__and2b_1 _1779_ (.A_N(_0415_),
    .B(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__mux4_1 _1780_ (.A0(\po_0.regf_0.rf[0][1] ),
    .A1(\po_0.regf_0.rf[1][1] ),
    .A2(\po_0.regf_0.rf[2][1] ),
    .A3(\po_0.regf_0.rf[3][1] ),
    .S0(_0423_),
    .S1(_0425_),
    .X(_0437_));
 sky130_fd_sc_hd__mux4_1 _1781_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(\po_0.regf_0.rf[5][1] ),
    .A2(\po_0.regf_0.rf[6][1] ),
    .A3(\po_0.regf_0.rf[7][1] ),
    .S0(_0427_),
    .S1(_0428_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _1782_ (.A0(_0437_),
    .A1(_0438_),
    .S(_0430_),
    .X(_0439_));
 sky130_fd_sc_hd__o22a_1 _1783_ (.A1(_0434_),
    .A2(_0436_),
    .B1(_0421_),
    .B2(_0439_),
    .X(\po_0.regf_0._3_[1] ));
 sky130_fd_sc_hd__mux4_1 _1784_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(\po_0.regf_0.rf[5][2] ),
    .A2(\po_0.regf_0.rf[6][2] ),
    .A3(\po_0.regf_0.rf[7][2] ),
    .S0(_0406_),
    .S1(_0408_),
    .X(_0440_));
 sky130_fd_sc_hd__a21o_1 _1785_ (.A1(_0440_),
    .A2(_0411_),
    .B1(_0420_),
    .X(_0441_));
 sky130_fd_sc_hd__mux4_1 _1786_ (.A0(\po_0.regf_0.rf[0][2] ),
    .A1(\po_0.regf_0.rf[1][2] ),
    .A2(\po_0.regf_0.rf[2][2] ),
    .A3(\po_0.regf_0.rf[3][2] ),
    .S0(_0416_),
    .S1(_0417_),
    .X(_0442_));
 sky130_fd_sc_hd__and2b_1 _1787_ (.A_N(_0415_),
    .B(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__buf_4 _1788_ (.A(_0405_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_4 _1789_ (.A(_0407_),
    .X(_0445_));
 sky130_fd_sc_hd__mux4_1 _1790_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(\po_0.regf_0.rf[13][2] ),
    .A2(\po_0.regf_0.rf[14][2] ),
    .A3(\po_0.regf_0.rf[15][2] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__buf_2 _1791_ (.A(_0410_),
    .X(_0447_));
 sky130_fd_sc_hd__a21bo_1 _1792_ (.A1(_0446_),
    .A2(_0447_),
    .B1_N(_0420_),
    .X(_0448_));
 sky130_fd_sc_hd__buf_4 _1793_ (.A(_0405_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_4 _1794_ (.A(_0407_),
    .X(_0450_));
 sky130_fd_sc_hd__mux4_1 _1795_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(\po_0.regf_0.rf[9][2] ),
    .A2(\po_0.regf_0.rf[10][2] ),
    .A3(\po_0.regf_0.rf[11][2] ),
    .S0(_0449_),
    .S1(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__and2b_1 _1796_ (.A_N(_0411_),
    .B(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__o22a_1 _1797_ (.A1(_0441_),
    .A2(_0443_),
    .B1(_0448_),
    .B2(_0452_),
    .X(\po_0.regf_0._3_[2] ));
 sky130_fd_sc_hd__mux4_1 _1798_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(\po_0.regf_0.rf[9][3] ),
    .A2(\po_0.regf_0.rf[10][3] ),
    .A3(\po_0.regf_0.rf[11][3] ),
    .S0(_0423_),
    .S1(_0425_),
    .X(_0453_));
 sky130_fd_sc_hd__and2b_1 _1799_ (.A_N(_0430_),
    .B(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__mux4_1 _1800_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(\po_0.regf_0.rf[13][3] ),
    .A2(\po_0.regf_0.rf[14][3] ),
    .A3(\po_0.regf_0.rf[15][3] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0455_));
 sky130_fd_sc_hd__a21bo_1 _1801_ (.A1(_0455_),
    .A2(_0447_),
    .B1_N(_0412_),
    .X(_0456_));
 sky130_fd_sc_hd__buf_2 _1802_ (.A(_0410_),
    .X(_0457_));
 sky130_fd_sc_hd__mux4_1 _1803_ (.A0(\po_0.regf_0.rf[0][3] ),
    .A1(\po_0.regf_0.rf[1][3] ),
    .A2(\po_0.regf_0.rf[2][3] ),
    .A3(\po_0.regf_0.rf[3][3] ),
    .S0(_0449_),
    .S1(_0450_),
    .X(_0458_));
 sky130_fd_sc_hd__and2b_1 _1804_ (.A_N(_0457_),
    .B(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__mux4_1 _1805_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(\po_0.regf_0.rf[5][3] ),
    .A2(\po_0.regf_0.rf[6][3] ),
    .A3(\po_0.regf_0.rf[7][3] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0460_));
 sky130_fd_sc_hd__buf_2 _1806_ (.A(_0003_),
    .X(_0461_));
 sky130_fd_sc_hd__a21o_1 _1807_ (.A1(_0460_),
    .A2(_0447_),
    .B1(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__o22a_1 _1808_ (.A1(_0454_),
    .A2(_0456_),
    .B1(_0459_),
    .B2(_0462_),
    .X(\po_0.regf_0._3_[3] ));
 sky130_fd_sc_hd__mux4_1 _1809_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(\po_0.regf_0.rf[9][4] ),
    .A2(\po_0.regf_0.rf[10][4] ),
    .A3(\po_0.regf_0.rf[11][4] ),
    .S0(_0423_),
    .S1(_0425_),
    .X(_0463_));
 sky130_fd_sc_hd__and2b_1 _1810_ (.A_N(_0430_),
    .B(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__mux4_1 _1811_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(\po_0.regf_0.rf[13][4] ),
    .A2(\po_0.regf_0.rf[14][4] ),
    .A3(\po_0.regf_0.rf[15][4] ),
    .S0(_0406_),
    .S1(_0408_),
    .X(_0465_));
 sky130_fd_sc_hd__a21bo_1 _1812_ (.A1(_0465_),
    .A2(_0411_),
    .B1_N(_0412_),
    .X(_0466_));
 sky130_fd_sc_hd__mux4_1 _1813_ (.A0(\po_0.regf_0.rf[0][4] ),
    .A1(\po_0.regf_0.rf[1][4] ),
    .A2(\po_0.regf_0.rf[2][4] ),
    .A3(\po_0.regf_0.rf[3][4] ),
    .S0(_0449_),
    .S1(_0450_),
    .X(_0467_));
 sky130_fd_sc_hd__and2b_1 _1814_ (.A_N(_0457_),
    .B(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__mux4_1 _1815_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(\po_0.regf_0.rf[5][4] ),
    .A2(\po_0.regf_0.rf[6][4] ),
    .A3(\po_0.regf_0.rf[7][4] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0469_));
 sky130_fd_sc_hd__a21o_1 _1816_ (.A1(_0469_),
    .A2(_0447_),
    .B1(_0461_),
    .X(_0470_));
 sky130_fd_sc_hd__o22a_1 _1817_ (.A1(_0464_),
    .A2(_0466_),
    .B1(_0468_),
    .B2(_0470_),
    .X(\po_0.regf_0._3_[4] ));
 sky130_fd_sc_hd__clkbuf_4 _1818_ (.A(_0405_),
    .X(_0471_));
 sky130_fd_sc_hd__buf_2 _1819_ (.A(_0407_),
    .X(_0472_));
 sky130_fd_sc_hd__mux4_1 _1820_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(\po_0.regf_0.rf[13][5] ),
    .A2(\po_0.regf_0.rf[14][5] ),
    .A3(\po_0.regf_0.rf[15][5] ),
    .S0(_0471_),
    .S1(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_2 _1821_ (.A(_0003_),
    .X(_0474_));
 sky130_fd_sc_hd__a21bo_1 _1822_ (.A1(_0473_),
    .A2(_0433_),
    .B1_N(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__mux4_1 _1823_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(\po_0.regf_0.rf[9][5] ),
    .A2(\po_0.regf_0.rf[10][5] ),
    .A3(\po_0.regf_0.rf[11][5] ),
    .S0(_0416_),
    .S1(_0417_),
    .X(_0476_));
 sky130_fd_sc_hd__and2b_1 _1824_ (.A_N(_0415_),
    .B(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_4 _1825_ (.A(_0422_),
    .X(_0478_));
 sky130_fd_sc_hd__buf_2 _1826_ (.A(_0424_),
    .X(_0479_));
 sky130_fd_sc_hd__mux4_1 _1827_ (.A0(\po_0.regf_0.rf[0][5] ),
    .A1(\po_0.regf_0.rf[1][5] ),
    .A2(\po_0.regf_0.rf[2][5] ),
    .A3(\po_0.regf_0.rf[3][5] ),
    .S0(_0478_),
    .S1(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__mux4_1 _1828_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(\po_0.regf_0.rf[5][5] ),
    .A2(\po_0.regf_0.rf[6][5] ),
    .A3(\po_0.regf_0.rf[7][5] ),
    .S0(_0427_),
    .S1(_0428_),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_4 _1829_ (.A(_0414_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _1830_ (.A0(_0480_),
    .A1(_0481_),
    .S(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__o22a_1 _1831_ (.A1(_0475_),
    .A2(_0477_),
    .B1(_0421_),
    .B2(_0483_),
    .X(\po_0.regf_0._3_[5] ));
 sky130_fd_sc_hd__mux4_1 _1832_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(\po_0.regf_0.rf[13][6] ),
    .A2(\po_0.regf_0.rf[14][6] ),
    .A3(\po_0.regf_0.rf[15][6] ),
    .S0(_0471_),
    .S1(_0472_),
    .X(_0484_));
 sky130_fd_sc_hd__a21bo_1 _1833_ (.A1(_0484_),
    .A2(_0433_),
    .B1_N(_0474_),
    .X(_0485_));
 sky130_fd_sc_hd__mux4_1 _1834_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(\po_0.regf_0.rf[9][6] ),
    .A2(\po_0.regf_0.rf[10][6] ),
    .A3(\po_0.regf_0.rf[11][6] ),
    .S0(_0416_),
    .S1(_0417_),
    .X(_0486_));
 sky130_fd_sc_hd__and2b_1 _1835_ (.A_N(_0415_),
    .B(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__mux4_1 _1836_ (.A0(\po_0.regf_0.rf[0][6] ),
    .A1(\po_0.regf_0.rf[1][6] ),
    .A2(\po_0.regf_0.rf[2][6] ),
    .A3(\po_0.regf_0.rf[3][6] ),
    .S0(_0478_),
    .S1(_0479_),
    .X(_0488_));
 sky130_fd_sc_hd__mux4_1 _1837_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(\po_0.regf_0.rf[5][6] ),
    .A2(\po_0.regf_0.rf[6][6] ),
    .A3(\po_0.regf_0.rf[7][6] ),
    .S0(_0427_),
    .S1(_0428_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _1838_ (.A0(_0488_),
    .A1(_0489_),
    .S(_0482_),
    .X(_0490_));
 sky130_fd_sc_hd__o22a_1 _1839_ (.A1(_0485_),
    .A2(_0487_),
    .B1(_0421_),
    .B2(_0490_),
    .X(\po_0.regf_0._3_[6] ));
 sky130_fd_sc_hd__mux4_1 _1840_ (.A0(\po_0.regf_0.rf[8][7] ),
    .A1(\po_0.regf_0.rf[9][7] ),
    .A2(\po_0.regf_0.rf[10][7] ),
    .A3(\po_0.regf_0.rf[11][7] ),
    .S0(_0423_),
    .S1(_0425_),
    .X(_0491_));
 sky130_fd_sc_hd__and2b_1 _1841_ (.A_N(_0430_),
    .B(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__mux4_1 _1842_ (.A0(\po_0.regf_0.rf[12][7] ),
    .A1(\po_0.regf_0.rf[13][7] ),
    .A2(\po_0.regf_0.rf[14][7] ),
    .A3(\po_0.regf_0.rf[15][7] ),
    .S0(_0406_),
    .S1(_0408_),
    .X(_0493_));
 sky130_fd_sc_hd__a21bo_1 _1843_ (.A1(_0493_),
    .A2(_0411_),
    .B1_N(_0412_),
    .X(_0494_));
 sky130_fd_sc_hd__mux4_1 _1844_ (.A0(\po_0.regf_0.rf[0][7] ),
    .A1(\po_0.regf_0.rf[1][7] ),
    .A2(\po_0.regf_0.rf[2][7] ),
    .A3(\po_0.regf_0.rf[3][7] ),
    .S0(_0449_),
    .S1(_0450_),
    .X(_0495_));
 sky130_fd_sc_hd__and2b_1 _1845_ (.A_N(_0457_),
    .B(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__mux4_1 _1846_ (.A0(\po_0.regf_0.rf[4][7] ),
    .A1(\po_0.regf_0.rf[5][7] ),
    .A2(\po_0.regf_0.rf[6][7] ),
    .A3(\po_0.regf_0.rf[7][7] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0497_));
 sky130_fd_sc_hd__a21o_1 _1847_ (.A1(_0497_),
    .A2(_0447_),
    .B1(_0420_),
    .X(_0498_));
 sky130_fd_sc_hd__o22a_1 _1848_ (.A1(_0492_),
    .A2(_0494_),
    .B1(_0496_),
    .B2(_0498_),
    .X(\po_0.regf_0._3_[7] ));
 sky130_fd_sc_hd__mux4_1 _1849_ (.A0(\po_0.regf_0.rf[0][8] ),
    .A1(\po_0.regf_0.rf[1][8] ),
    .A2(\po_0.regf_0.rf[2][8] ),
    .A3(\po_0.regf_0.rf[3][8] ),
    .S0(_0422_),
    .S1(_0424_),
    .X(_0499_));
 sky130_fd_sc_hd__mux4_1 _1850_ (.A0(\po_0.regf_0.rf[4][8] ),
    .A1(\po_0.regf_0.rf[5][8] ),
    .A2(\po_0.regf_0.rf[6][8] ),
    .A3(\po_0.regf_0.rf[7][8] ),
    .S0(_0422_),
    .S1(_0424_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _1851_ (.A0(_0499_),
    .A1(_0500_),
    .S(_0414_),
    .X(_0501_));
 sky130_fd_sc_hd__mux4_1 _1852_ (.A0(\po_0.regf_0.rf[8][8] ),
    .A1(\po_0.regf_0.rf[9][8] ),
    .A2(\po_0.regf_0.rf[10][8] ),
    .A3(\po_0.regf_0.rf[11][8] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_0502_));
 sky130_fd_sc_hd__mux4_1 _1853_ (.A0(\po_0.regf_0.rf[12][8] ),
    .A1(\po_0.regf_0.rf[13][8] ),
    .A2(\po_0.regf_0.rf[14][8] ),
    .A3(\po_0.regf_0.rf[15][8] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _1854_ (.A0(_0502_),
    .A1(_0503_),
    .S(_0414_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _1855_ (.A0(_0501_),
    .A1(_0504_),
    .S(_0420_),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_1 _1856_ (.A(_0505_),
    .X(\po_0.regf_0._3_[8] ));
 sky130_fd_sc_hd__mux4_1 _1857_ (.A0(\po_0.regf_0.rf[12][9] ),
    .A1(\po_0.regf_0.rf[13][9] ),
    .A2(\po_0.regf_0.rf[14][9] ),
    .A3(\po_0.regf_0.rf[15][9] ),
    .S0(_0471_),
    .S1(_0472_),
    .X(_0506_));
 sky130_fd_sc_hd__a21bo_1 _1858_ (.A1(_0506_),
    .A2(_0433_),
    .B1_N(_0474_),
    .X(_0507_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1859_ (.A(_0414_),
    .X(_0508_));
 sky130_fd_sc_hd__buf_2 _1860_ (.A(_0405_),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_2 _1861_ (.A(_0407_),
    .X(_0510_));
 sky130_fd_sc_hd__mux4_1 _1862_ (.A0(\po_0.regf_0.rf[8][9] ),
    .A1(\po_0.regf_0.rf[9][9] ),
    .A2(\po_0.regf_0.rf[10][9] ),
    .A3(\po_0.regf_0.rf[11][9] ),
    .S0(_0509_),
    .S1(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__and2b_1 _1863_ (.A_N(_0508_),
    .B(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__mux4_1 _1864_ (.A0(\po_0.regf_0.rf[0][9] ),
    .A1(\po_0.regf_0.rf[1][9] ),
    .A2(\po_0.regf_0.rf[2][9] ),
    .A3(\po_0.regf_0.rf[3][9] ),
    .S0(_0478_),
    .S1(_0479_),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_4 _1865_ (.A(_0422_),
    .X(_0514_));
 sky130_fd_sc_hd__buf_2 _1866_ (.A(_0424_),
    .X(_0515_));
 sky130_fd_sc_hd__mux4_1 _1867_ (.A0(\po_0.regf_0.rf[4][9] ),
    .A1(\po_0.regf_0.rf[5][9] ),
    .A2(\po_0.regf_0.rf[6][9] ),
    .A3(\po_0.regf_0.rf[7][9] ),
    .S0(_0514_),
    .S1(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _1868_ (.A0(_0513_),
    .A1(_0516_),
    .S(_0482_),
    .X(_0517_));
 sky130_fd_sc_hd__o22a_1 _1869_ (.A1(_0507_),
    .A2(_0512_),
    .B1(_0421_),
    .B2(_0517_),
    .X(\po_0.regf_0._3_[9] ));
 sky130_fd_sc_hd__mux4_1 _1870_ (.A0(\po_0.regf_0.rf[8][10] ),
    .A1(\po_0.regf_0.rf[9][10] ),
    .A2(\po_0.regf_0.rf[10][10] ),
    .A3(\po_0.regf_0.rf[11][10] ),
    .S0(_0423_),
    .S1(_0425_),
    .X(_0518_));
 sky130_fd_sc_hd__and2b_1 _1871_ (.A_N(_0430_),
    .B(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__mux4_1 _1872_ (.A0(\po_0.regf_0.rf[12][10] ),
    .A1(\po_0.regf_0.rf[13][10] ),
    .A2(\po_0.regf_0.rf[14][10] ),
    .A3(\po_0.regf_0.rf[15][10] ),
    .S0(_0406_),
    .S1(_0408_),
    .X(_0520_));
 sky130_fd_sc_hd__a21bo_1 _1873_ (.A1(_0520_),
    .A2(_0411_),
    .B1_N(_0412_),
    .X(_0521_));
 sky130_fd_sc_hd__mux4_1 _1874_ (.A0(\po_0.regf_0.rf[0][10] ),
    .A1(\po_0.regf_0.rf[1][10] ),
    .A2(\po_0.regf_0.rf[2][10] ),
    .A3(\po_0.regf_0.rf[3][10] ),
    .S0(_0416_),
    .S1(_0417_),
    .X(_0522_));
 sky130_fd_sc_hd__and2b_1 _1875_ (.A_N(_0415_),
    .B(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__mux4_1 _1876_ (.A0(\po_0.regf_0.rf[4][10] ),
    .A1(\po_0.regf_0.rf[5][10] ),
    .A2(\po_0.regf_0.rf[6][10] ),
    .A3(\po_0.regf_0.rf[7][10] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0524_));
 sky130_fd_sc_hd__a21o_1 _1877_ (.A1(_0524_),
    .A2(_0447_),
    .B1(_0420_),
    .X(_0525_));
 sky130_fd_sc_hd__o22a_1 _1878_ (.A1(_0519_),
    .A2(_0521_),
    .B1(_0523_),
    .B2(_0525_),
    .X(\po_0.regf_0._3_[10] ));
 sky130_fd_sc_hd__mux4_1 _1879_ (.A0(\po_0.regf_0.rf[12][11] ),
    .A1(\po_0.regf_0.rf[13][11] ),
    .A2(\po_0.regf_0.rf[14][11] ),
    .A3(\po_0.regf_0.rf[15][11] ),
    .S0(_0471_),
    .S1(_0472_),
    .X(_0526_));
 sky130_fd_sc_hd__a21bo_1 _1880_ (.A1(_0526_),
    .A2(_0433_),
    .B1_N(_0474_),
    .X(_0527_));
 sky130_fd_sc_hd__mux4_1 _1881_ (.A0(\po_0.regf_0.rf[8][11] ),
    .A1(\po_0.regf_0.rf[9][11] ),
    .A2(\po_0.regf_0.rf[10][11] ),
    .A3(\po_0.regf_0.rf[11][11] ),
    .S0(_0509_),
    .S1(_0510_),
    .X(_0528_));
 sky130_fd_sc_hd__and2b_1 _1882_ (.A_N(_0508_),
    .B(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__mux4_1 _1883_ (.A0(\po_0.regf_0.rf[0][11] ),
    .A1(\po_0.regf_0.rf[1][11] ),
    .A2(\po_0.regf_0.rf[2][11] ),
    .A3(\po_0.regf_0.rf[3][11] ),
    .S0(_0478_),
    .S1(_0479_),
    .X(_0530_));
 sky130_fd_sc_hd__mux4_1 _1884_ (.A0(\po_0.regf_0.rf[4][11] ),
    .A1(\po_0.regf_0.rf[5][11] ),
    .A2(\po_0.regf_0.rf[6][11] ),
    .A3(\po_0.regf_0.rf[7][11] ),
    .S0(_0514_),
    .S1(_0515_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _1885_ (.A0(_0530_),
    .A1(_0531_),
    .S(_0482_),
    .X(_0532_));
 sky130_fd_sc_hd__o22a_1 _1886_ (.A1(_0527_),
    .A2(_0529_),
    .B1(_0421_),
    .B2(_0532_),
    .X(\po_0.regf_0._3_[11] ));
 sky130_fd_sc_hd__mux4_1 _1887_ (.A0(\po_0.regf_0.rf[12][12] ),
    .A1(\po_0.regf_0.rf[13][12] ),
    .A2(\po_0.regf_0.rf[14][12] ),
    .A3(\po_0.regf_0.rf[15][12] ),
    .S0(_0471_),
    .S1(_0472_),
    .X(_0533_));
 sky130_fd_sc_hd__a21bo_1 _1888_ (.A1(_0533_),
    .A2(_0433_),
    .B1_N(_0474_),
    .X(_0534_));
 sky130_fd_sc_hd__mux4_1 _1889_ (.A0(\po_0.regf_0.rf[8][12] ),
    .A1(\po_0.regf_0.rf[9][12] ),
    .A2(\po_0.regf_0.rf[10][12] ),
    .A3(\po_0.regf_0.rf[11][12] ),
    .S0(_0509_),
    .S1(_0510_),
    .X(_0535_));
 sky130_fd_sc_hd__and2b_1 _1890_ (.A_N(_0508_),
    .B(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__mux4_1 _1891_ (.A0(\po_0.regf_0.rf[0][12] ),
    .A1(\po_0.regf_0.rf[1][12] ),
    .A2(\po_0.regf_0.rf[2][12] ),
    .A3(\po_0.regf_0.rf[3][12] ),
    .S0(_0478_),
    .S1(_0479_),
    .X(_0537_));
 sky130_fd_sc_hd__mux4_1 _1892_ (.A0(\po_0.regf_0.rf[4][12] ),
    .A1(\po_0.regf_0.rf[5][12] ),
    .A2(\po_0.regf_0.rf[6][12] ),
    .A3(\po_0.regf_0.rf[7][12] ),
    .S0(_0514_),
    .S1(_0515_),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _1893_ (.A0(_0537_),
    .A1(_0538_),
    .S(_0482_),
    .X(_0539_));
 sky130_fd_sc_hd__o22a_1 _1894_ (.A1(_0534_),
    .A2(_0536_),
    .B1(_0461_),
    .B2(_0539_),
    .X(\po_0.regf_0._3_[12] ));
 sky130_fd_sc_hd__mux4_1 _1895_ (.A0(\po_0.regf_0.rf[12][13] ),
    .A1(\po_0.regf_0.rf[13][13] ),
    .A2(\po_0.regf_0.rf[14][13] ),
    .A3(\po_0.regf_0.rf[15][13] ),
    .S0(_0471_),
    .S1(_0472_),
    .X(_0540_));
 sky130_fd_sc_hd__a21bo_1 _1896_ (.A1(_0540_),
    .A2(_0457_),
    .B1_N(_0474_),
    .X(_0541_));
 sky130_fd_sc_hd__mux4_1 _1897_ (.A0(\po_0.regf_0.rf[8][13] ),
    .A1(\po_0.regf_0.rf[9][13] ),
    .A2(\po_0.regf_0.rf[10][13] ),
    .A3(\po_0.regf_0.rf[11][13] ),
    .S0(_0509_),
    .S1(_0510_),
    .X(_0542_));
 sky130_fd_sc_hd__and2b_1 _1898_ (.A_N(_0508_),
    .B(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__mux4_1 _1899_ (.A0(\po_0.regf_0.rf[0][13] ),
    .A1(\po_0.regf_0.rf[1][13] ),
    .A2(\po_0.regf_0.rf[2][13] ),
    .A3(\po_0.regf_0.rf[3][13] ),
    .S0(_0478_),
    .S1(_0479_),
    .X(_0544_));
 sky130_fd_sc_hd__mux4_1 _1900_ (.A0(\po_0.regf_0.rf[4][13] ),
    .A1(\po_0.regf_0.rf[5][13] ),
    .A2(\po_0.regf_0.rf[6][13] ),
    .A3(\po_0.regf_0.rf[7][13] ),
    .S0(_0514_),
    .S1(_0515_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _1901_ (.A0(_0544_),
    .A1(_0545_),
    .S(_0482_),
    .X(_0546_));
 sky130_fd_sc_hd__o22a_1 _1902_ (.A1(_0541_),
    .A2(_0543_),
    .B1(_0461_),
    .B2(_0546_),
    .X(\po_0.regf_0._3_[13] ));
 sky130_fd_sc_hd__mux4_1 _1903_ (.A0(\po_0.regf_0.rf[12][14] ),
    .A1(\po_0.regf_0.rf[13][14] ),
    .A2(\po_0.regf_0.rf[14][14] ),
    .A3(\po_0.regf_0.rf[15][14] ),
    .S0(_0449_),
    .S1(_0450_),
    .X(_0547_));
 sky130_fd_sc_hd__a21bo_1 _1904_ (.A1(_0547_),
    .A2(_0457_),
    .B1_N(_0003_),
    .X(_0548_));
 sky130_fd_sc_hd__mux4_1 _1905_ (.A0(\po_0.regf_0.rf[8][14] ),
    .A1(\po_0.regf_0.rf[9][14] ),
    .A2(\po_0.regf_0.rf[10][14] ),
    .A3(\po_0.regf_0.rf[11][14] ),
    .S0(_0509_),
    .S1(_0510_),
    .X(_0549_));
 sky130_fd_sc_hd__and2b_1 _1906_ (.A_N(_0508_),
    .B(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__mux4_1 _1907_ (.A0(\po_0.regf_0.rf[0][14] ),
    .A1(\po_0.regf_0.rf[1][14] ),
    .A2(\po_0.regf_0.rf[2][14] ),
    .A3(\po_0.regf_0.rf[3][14] ),
    .S0(_0427_),
    .S1(_0428_),
    .X(_0551_));
 sky130_fd_sc_hd__mux4_1 _1908_ (.A0(\po_0.regf_0.rf[4][14] ),
    .A1(\po_0.regf_0.rf[5][14] ),
    .A2(\po_0.regf_0.rf[6][14] ),
    .A3(\po_0.regf_0.rf[7][14] ),
    .S0(_0514_),
    .S1(_0515_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _1909_ (.A0(_0551_),
    .A1(_0552_),
    .S(_0410_),
    .X(_0553_));
 sky130_fd_sc_hd__o22a_1 _1910_ (.A1(_0548_),
    .A2(_0550_),
    .B1(_0461_),
    .B2(_0553_),
    .X(\po_0.regf_0._3_[14] ));
 sky130_fd_sc_hd__mux4_1 _1911_ (.A0(\po_0.regf_0.rf[12][15] ),
    .A1(\po_0.regf_0.rf[13][15] ),
    .A2(\po_0.regf_0.rf[14][15] ),
    .A3(\po_0.regf_0.rf[15][15] ),
    .S0(_0449_),
    .S1(_0450_),
    .X(_0554_));
 sky130_fd_sc_hd__a21bo_1 _1912_ (.A1(_0554_),
    .A2(_0457_),
    .B1_N(_0003_),
    .X(_0555_));
 sky130_fd_sc_hd__mux4_1 _1913_ (.A0(\po_0.regf_0.rf[8][15] ),
    .A1(\po_0.regf_0.rf[9][15] ),
    .A2(\po_0.regf_0.rf[10][15] ),
    .A3(\po_0.regf_0.rf[11][15] ),
    .S0(_0509_),
    .S1(_0510_),
    .X(_0556_));
 sky130_fd_sc_hd__and2b_1 _1914_ (.A_N(_0508_),
    .B(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__mux4_1 _1915_ (.A0(\po_0.regf_0.rf[0][15] ),
    .A1(\po_0.regf_0.rf[1][15] ),
    .A2(\po_0.regf_0.rf[2][15] ),
    .A3(\po_0.regf_0.rf[3][15] ),
    .S0(_0427_),
    .S1(_0428_),
    .X(_0558_));
 sky130_fd_sc_hd__mux4_1 _1916_ (.A0(\po_0.regf_0.rf[4][15] ),
    .A1(\po_0.regf_0.rf[5][15] ),
    .A2(\po_0.regf_0.rf[6][15] ),
    .A3(\po_0.regf_0.rf[7][15] ),
    .S0(_0514_),
    .S1(_0515_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _1917_ (.A0(_0558_),
    .A1(_0559_),
    .S(_0410_),
    .X(_0560_));
 sky130_fd_sc_hd__o22a_1 _1918_ (.A1(_0555_),
    .A2(_0557_),
    .B1(_0461_),
    .B2(_0560_),
    .X(\po_0.regf_0._3_[15] ));
 sky130_fd_sc_hd__buf_2 _1919_ (.A(\po_0.muxf_0.rf_w_data[4] ),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_4 _1920_ (.A(_1371_),
    .X(_0562_));
 sky130_fd_sc_hd__buf_2 _1921_ (.A(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _1922_ (.A0(\po_0.regf_0.rq_addr[0] ),
    .A1(_0561_),
    .S(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__clkbuf_1 _1923_ (.A(_0564_),
    .X(_0012_));
 sky130_fd_sc_hd__buf_2 _1924_ (.A(\po_0.muxf_0.rf_w_data[5] ),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _1925_ (.A0(\po_0.regf_0.rq_addr[1] ),
    .A1(_0565_),
    .S(_0563_),
    .X(_0566_));
 sky130_fd_sc_hd__clkbuf_1 _1926_ (.A(_0566_),
    .X(_0013_));
 sky130_fd_sc_hd__buf_2 _1927_ (.A(\po_0.muxf_0.rf_w_data[6] ),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_2 _1928_ (.A(_0562_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _1929_ (.A0(\po_0.regf_0.rq_addr[2] ),
    .A1(_0567_),
    .S(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__clkbuf_1 _1930_ (.A(_0569_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_4 _1931_ (.A(\po_0.muxf_0.rf_w_data[7] ),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _1932_ (.A0(\po_0.regf_0.rq_addr[3] ),
    .A1(_0570_),
    .S(_0568_),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_1 _1933_ (.A(_0571_),
    .X(_0015_));
 sky130_fd_sc_hd__and2b_1 _1934_ (.A_N(_1340_),
    .B(\po_0._1_[0] ),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_2 _1935_ (.A(\po_0._1_[1] ),
    .X(_0573_));
 sky130_fd_sc_hd__clkbuf_2 _1936_ (.A(net42),
    .X(_0574_));
 sky130_fd_sc_hd__or2b_1 _1937_ (.A(_0573_),
    .B_N(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__or2b_1 _1938_ (.A(net42),
    .B_N(\po_0._1_[1] ),
    .X(_0576_));
 sky130_fd_sc_hd__nand2_1 _1939_ (.A(_0575_),
    .B(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__xor2_1 _1940_ (.A(_0572_),
    .B(_0577_),
    .X(\po_0.alu_0._10_[1] ));
 sky130_fd_sc_hd__inv_2 _1941_ (.A(_0573_),
    .Y(_0578_));
 sky130_fd_sc_hd__clkbuf_2 _1942_ (.A(net43),
    .X(_0579_));
 sky130_fd_sc_hd__nand2b_2 _1943_ (.A_N(\po_0._1_[2] ),
    .B(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__or2b_1 _1944_ (.A(_0579_),
    .B_N(\po_0._1_[2] ),
    .X(_0581_));
 sky130_fd_sc_hd__inv_2 _1945_ (.A(_0574_),
    .Y(_0582_));
 sky130_fd_sc_hd__o21ai_1 _1946_ (.A1(_0573_),
    .A2(_0582_),
    .B1(_0572_),
    .Y(_0583_));
 sky130_fd_sc_hd__o2111ai_2 _1947_ (.A1(_0574_),
    .A2(_0578_),
    .B1(_0580_),
    .C1(_0581_),
    .D1(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__or2b_1 _1948_ (.A(_1340_),
    .B_N(\po_0._1_[0] ),
    .X(_0585_));
 sky130_fd_sc_hd__and2b_1 _1949_ (.A_N(_0573_),
    .B(net42),
    .X(_0586_));
 sky130_fd_sc_hd__a221o_1 _1950_ (.A1(_0585_),
    .A2(_0576_),
    .B1(_0580_),
    .B2(_0581_),
    .C1(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__and2_1 _1951_ (.A(_0584_),
    .B(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__clkbuf_1 _1952_ (.A(_0588_),
    .X(\po_0.alu_0._10_[2] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1953_ (.A(net44),
    .X(_0589_));
 sky130_fd_sc_hd__and2_1 _1954_ (.A(_0589_),
    .B(\po_0._1_[3] ),
    .X(_0590_));
 sky130_fd_sc_hd__nor2_1 _1955_ (.A(_0589_),
    .B(\po_0._1_[3] ),
    .Y(_0591_));
 sky130_fd_sc_hd__o2bb2ai_1 _1956_ (.A1_N(_0580_),
    .A2_N(_0584_),
    .B1(_0590_),
    .B2(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand2_1 _1957_ (.A(_0580_),
    .B(_0581_),
    .Y(_0593_));
 sky130_fd_sc_hd__a21oi_1 _1958_ (.A1(_0585_),
    .A2(_0576_),
    .B1(_0586_),
    .Y(_0594_));
 sky130_fd_sc_hd__nand2_1 _1959_ (.A(_0589_),
    .B(\po_0._1_[3] ),
    .Y(_0595_));
 sky130_fd_sc_hd__or2_1 _1960_ (.A(_0589_),
    .B(\po_0._1_[3] ),
    .X(_0596_));
 sky130_fd_sc_hd__o2111ai_1 _1961_ (.A1(_0593_),
    .A2(_0594_),
    .B1(_0595_),
    .C1(_0596_),
    .D1(_0580_),
    .Y(_0597_));
 sky130_fd_sc_hd__and2_1 _1962_ (.A(_0592_),
    .B(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__clkbuf_1 _1963_ (.A(_0598_),
    .X(\po_0.alu_0._10_[3] ));
 sky130_fd_sc_hd__and2_1 _1964_ (.A(net84),
    .B(\po_0._1_[4] ),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_1 _1965_ (.A(net84),
    .B(\po_0._1_[4] ),
    .Y(_0600_));
 sky130_fd_sc_hd__or2b_1 _1966_ (.A(\po_0._1_[3] ),
    .B_N(_0589_),
    .X(_0601_));
 sky130_fd_sc_hd__a2bb2oi_2 _1967_ (.A1_N(_0599_),
    .A2_N(_0600_),
    .B1(_0601_),
    .B2(_0592_),
    .Y(_0602_));
 sky130_fd_sc_hd__nor2_2 _1968_ (.A(_0599_),
    .B(_0600_),
    .Y(_0603_));
 sky130_fd_sc_hd__and3_1 _1969_ (.A(_0592_),
    .B(_0603_),
    .C(_0601_),
    .X(_0604_));
 sky130_fd_sc_hd__nor2_1 _1970_ (.A(_0602_),
    .B(_0604_),
    .Y(\po_0.alu_0._10_[4] ));
 sky130_fd_sc_hd__and2b_1 _1971_ (.A_N(\po_0._1_[4] ),
    .B(net84),
    .X(_0605_));
 sky130_fd_sc_hd__clkbuf_2 _1972_ (.A(net46),
    .X(_0606_));
 sky130_fd_sc_hd__nor2_2 _1973_ (.A(_0606_),
    .B(\po_0._1_[5] ),
    .Y(_0607_));
 sky130_fd_sc_hd__and2_1 _1974_ (.A(_0606_),
    .B(\po_0._1_[5] ),
    .X(_0608_));
 sky130_fd_sc_hd__nor2_2 _1975_ (.A(_0607_),
    .B(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__o21a_1 _1976_ (.A1(_0602_),
    .A2(_0605_),
    .B1(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__nor3_1 _1977_ (.A(_0602_),
    .B(_0609_),
    .C(_0605_),
    .Y(_0611_));
 sky130_fd_sc_hd__or2_1 _1978_ (.A(_0610_),
    .B(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__clkbuf_1 _1979_ (.A(_0612_),
    .X(\po_0.alu_0._10_[5] ));
 sky130_fd_sc_hd__and2_1 _1980_ (.A(net47),
    .B(\po_0._1_[6] ),
    .X(_0613_));
 sky130_fd_sc_hd__nor2_2 _1981_ (.A(_1347_),
    .B(\po_0._1_[6] ),
    .Y(_0614_));
 sky130_fd_sc_hd__or2b_1 _1982_ (.A(\po_0._1_[5] ),
    .B_N(_0606_),
    .X(_0615_));
 sky130_fd_sc_hd__o22ai_2 _1983_ (.A1(_0607_),
    .A2(_0608_),
    .B1(_0605_),
    .B2(_0602_),
    .Y(_0616_));
 sky130_fd_sc_hd__a2bb2oi_2 _1984_ (.A1_N(_0613_),
    .A2_N(_0614_),
    .B1(_0615_),
    .B2(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__nor2_1 _1985_ (.A(_0613_),
    .B(_0614_),
    .Y(_0618_));
 sky130_fd_sc_hd__nand3_1 _1986_ (.A(_0616_),
    .B(_0618_),
    .C(_0615_),
    .Y(_0619_));
 sky130_fd_sc_hd__and2b_1 _1987_ (.A_N(_0617_),
    .B(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__clkbuf_1 _1988_ (.A(_0620_),
    .X(\po_0.alu_0._10_[6] ));
 sky130_fd_sc_hd__clkbuf_2 _1989_ (.A(net48),
    .X(_0621_));
 sky130_fd_sc_hd__nor2_2 _1990_ (.A(_0621_),
    .B(\po_0._1_[7] ),
    .Y(_0622_));
 sky130_fd_sc_hd__and2_1 _1991_ (.A(_0621_),
    .B(\po_0._1_[7] ),
    .X(_0623_));
 sky130_fd_sc_hd__and2b_1 _1992_ (.A_N(\po_0._1_[6] ),
    .B(_1347_),
    .X(_0624_));
 sky130_fd_sc_hd__o22ai_4 _1993_ (.A1(_0622_),
    .A2(_0623_),
    .B1(_0624_),
    .B2(_0617_),
    .Y(_0625_));
 sky130_fd_sc_hd__inv_2 _1994_ (.A(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__nor4_1 _1995_ (.A(_0617_),
    .B(_0622_),
    .C(_0623_),
    .D(_0624_),
    .Y(_0627_));
 sky130_fd_sc_hd__nor2_1 _1996_ (.A(_0626_),
    .B(_0627_),
    .Y(\po_0.alu_0._10_[7] ));
 sky130_fd_sc_hd__nand2_1 _1997_ (.A(net83),
    .B(\po_0._1_[8] ),
    .Y(_0628_));
 sky130_fd_sc_hd__or2_1 _1998_ (.A(net83),
    .B(\po_0._1_[8] ),
    .X(_0629_));
 sky130_fd_sc_hd__nand2_1 _1999_ (.A(_0628_),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__inv_2 _2000_ (.A(_0621_),
    .Y(_0631_));
 sky130_fd_sc_hd__o21ai_4 _2001_ (.A1(_0631_),
    .A2(\po_0._1_[7] ),
    .B1(_0625_),
    .Y(_0632_));
 sky130_fd_sc_hd__xor2_1 _2002_ (.A(_0630_),
    .B(_0632_),
    .X(\po_0.alu_0._10_[8] ));
 sky130_fd_sc_hd__buf_2 _2003_ (.A(net50),
    .X(_0633_));
 sky130_fd_sc_hd__xnor2_2 _2004_ (.A(_0633_),
    .B(\po_0._1_[9] ),
    .Y(_0634_));
 sky130_fd_sc_hd__or2b_1 _2005_ (.A(\po_0._1_[8] ),
    .B_N(net83),
    .X(_0635_));
 sky130_fd_sc_hd__a21bo_1 _2006_ (.A1(_0630_),
    .A2(_0632_),
    .B1_N(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__xor2_1 _2007_ (.A(_0634_),
    .B(_0636_),
    .X(\po_0.alu_0._10_[9] ));
 sky130_fd_sc_hd__and2b_1 _2008_ (.A_N(net36),
    .B(\po_0._1_[10] ),
    .X(_0637_));
 sky130_fd_sc_hd__or2b_1 _2009_ (.A(\po_0._1_[10] ),
    .B_N(net36),
    .X(_0638_));
 sky130_fd_sc_hd__nand2b_2 _2010_ (.A_N(_0637_),
    .B(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__xor2_2 _2011_ (.A(net50),
    .B(\po_0._1_[9] ),
    .X(_0640_));
 sky130_fd_sc_hd__or2b_1 _2012_ (.A(\po_0._1_[9] ),
    .B_N(_0633_),
    .X(_0641_));
 sky130_fd_sc_hd__o21ai_1 _2013_ (.A1(_0635_),
    .A2(_0640_),
    .B1(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__a31oi_2 _2014_ (.A1(_0630_),
    .A2(_0632_),
    .A3(_0634_),
    .B1(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__xor2_1 _2015_ (.A(_0639_),
    .B(_0643_),
    .X(\po_0.alu_0._10_[10] ));
 sky130_fd_sc_hd__nor2_1 _2016_ (.A(net37),
    .B(\po_0._1_[11] ),
    .Y(_0644_));
 sky130_fd_sc_hd__and2_1 _2017_ (.A(net37),
    .B(\po_0._1_[11] ),
    .X(_0645_));
 sky130_fd_sc_hd__nor2_2 _2018_ (.A(_0644_),
    .B(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__o21ai_1 _2019_ (.A1(_0637_),
    .A2(_0643_),
    .B1(_0638_),
    .Y(_0647_));
 sky130_fd_sc_hd__xnor2_1 _2020_ (.A(_0646_),
    .B(_0647_),
    .Y(\po_0.alu_0._10_[11] ));
 sky130_fd_sc_hd__and2_1 _2021_ (.A(_0628_),
    .B(_0629_),
    .X(_0648_));
 sky130_fd_sc_hd__nor4_1 _2022_ (.A(_0648_),
    .B(_0640_),
    .C(_0639_),
    .D(_0646_),
    .Y(_0649_));
 sky130_fd_sc_hd__inv_2 _2023_ (.A(net37),
    .Y(_0650_));
 sky130_fd_sc_hd__o211a_1 _2024_ (.A1(_0635_),
    .A2(_0640_),
    .B1(_0641_),
    .C1(_0638_),
    .X(_0651_));
 sky130_fd_sc_hd__or3_1 _2025_ (.A(_0637_),
    .B(_0646_),
    .C(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__o21ai_1 _2026_ (.A1(_0650_),
    .A2(\po_0._1_[11] ),
    .B1(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__a21oi_2 _2027_ (.A1(_0632_),
    .A2(_0649_),
    .B1(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2028_ (.A(net38),
    .X(_0655_));
 sky130_fd_sc_hd__nand2_1 _2029_ (.A(_0655_),
    .B(\po_0._1_[12] ),
    .Y(_0656_));
 sky130_fd_sc_hd__or2_1 _2030_ (.A(_0655_),
    .B(\po_0._1_[12] ),
    .X(_0657_));
 sky130_fd_sc_hd__and2_1 _2031_ (.A(_0656_),
    .B(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__xor2_1 _2032_ (.A(_0654_),
    .B(_0658_),
    .X(\po_0.alu_0._10_[12] ));
 sky130_fd_sc_hd__buf_2 _2033_ (.A(net39),
    .X(_0659_));
 sky130_fd_sc_hd__xor2_2 _2034_ (.A(_0659_),
    .B(\po_0._1_[13] ),
    .X(_0660_));
 sky130_fd_sc_hd__or2b_1 _2035_ (.A(\po_0._1_[12] ),
    .B_N(_0655_),
    .X(_0661_));
 sky130_fd_sc_hd__o211a_1 _2036_ (.A1(_0654_),
    .A2(_0658_),
    .B1(_0660_),
    .C1(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__nand2_1 _2037_ (.A(_0632_),
    .B(_0649_),
    .Y(_0663_));
 sky130_fd_sc_hd__inv_2 _2038_ (.A(_0653_),
    .Y(_0664_));
 sky130_fd_sc_hd__a21o_1 _2039_ (.A1(_0656_),
    .A2(_0657_),
    .B1(_0660_),
    .X(_0665_));
 sky130_fd_sc_hd__a21oi_1 _2040_ (.A1(_0663_),
    .A2(_0664_),
    .B1(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__or3b_2 _2041_ (.A(\po_0._1_[12] ),
    .B(_0660_),
    .C_N(_0655_),
    .X(_0667_));
 sky130_fd_sc_hd__nor3b_1 _2042_ (.A(_0662_),
    .B(_0666_),
    .C_N(_0667_),
    .Y(\po_0.alu_0._10_[13] ));
 sky130_fd_sc_hd__and2_1 _2043_ (.A(net40),
    .B(\po_0._1_[14] ),
    .X(_0668_));
 sky130_fd_sc_hd__nor2_1 _2044_ (.A(net40),
    .B(\po_0._1_[14] ),
    .Y(_0669_));
 sky130_fd_sc_hd__or2_1 _2045_ (.A(_0668_),
    .B(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__inv_2 _2046_ (.A(_0659_),
    .Y(_0671_));
 sky130_fd_sc_hd__o221ai_4 _2047_ (.A1(_0671_),
    .A2(\po_0._1_[13] ),
    .B1(_0665_),
    .B2(_0654_),
    .C1(_0667_),
    .Y(_0672_));
 sky130_fd_sc_hd__xor2_1 _2048_ (.A(_0670_),
    .B(_0672_),
    .X(\po_0.alu_0._10_[14] ));
 sky130_fd_sc_hd__and2_1 _2049_ (.A(net41),
    .B(\po_0._1_[15] ),
    .X(_0673_));
 sky130_fd_sc_hd__nor2_1 _2050_ (.A(net41),
    .B(\po_0._1_[15] ),
    .Y(_0674_));
 sky130_fd_sc_hd__or2b_1 _2051_ (.A(\po_0._1_[14] ),
    .B_N(net40),
    .X(_0675_));
 sky130_fd_sc_hd__or3b_1 _2052_ (.A(_0673_),
    .B(_0674_),
    .C_N(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__a21oi_1 _2053_ (.A1(_0670_),
    .A2(_0672_),
    .B1(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__o21ai_1 _2054_ (.A1(_0671_),
    .A2(\po_0._1_[13] ),
    .B1(_0667_),
    .Y(_0678_));
 sky130_fd_sc_hd__o22ai_1 _2055_ (.A1(_0668_),
    .A2(_0669_),
    .B1(_0678_),
    .B2(_0666_),
    .Y(_0679_));
 sky130_fd_sc_hd__a2bb2oi_1 _2056_ (.A1_N(_0673_),
    .A2_N(_0674_),
    .B1(_0675_),
    .B2(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__nor2_1 _2057_ (.A(_0677_),
    .B(_0680_),
    .Y(\po_0.alu_0._10_[15] ));
 sky130_fd_sc_hd__clkbuf_4 _2058_ (.A(\po_0.muxf_0.rf_w_data[0] ),
    .X(_0681_));
 sky130_fd_sc_hd__and2b_1 _2059_ (.A_N(\po_0.muxf_0.s0 ),
    .B(\po_0.muxf_0.s1 ),
    .X(_0682_));
 sky130_fd_sc_hd__clkbuf_2 _2060_ (.A(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__and2b_1 _2061_ (.A_N(\po_0.muxf_0.s1 ),
    .B(\po_0.muxf_0.s0 ),
    .X(_0684_));
 sky130_fd_sc_hd__buf_2 _2062_ (.A(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__clkbuf_2 _2063_ (.A(_1316_),
    .X(_0686_));
 sky130_fd_sc_hd__nor2_2 _2064_ (.A(_0682_),
    .B(_0684_),
    .Y(_0687_));
 sky130_fd_sc_hd__nor2_2 _2065_ (.A(_1316_),
    .B(_1313_),
    .Y(_0688_));
 sky130_fd_sc_hd__and2b_1 _2066_ (.A_N(_1316_),
    .B(\po_0.alu_0.s0 ),
    .X(_0689_));
 sky130_fd_sc_hd__and3_1 _2067_ (.A(_1341_),
    .B(_1342_),
    .C(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__a211o_1 _2068_ (.A1(_1317_),
    .A2(\po_0.alu_0._11_[0] ),
    .B1(_0688_),
    .C1(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__o311a_1 _2069_ (.A1(_1340_),
    .A2(_0686_),
    .A3(_1314_),
    .B1(_0687_),
    .C1(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__a221o_2 _2070_ (.A1(_0681_),
    .A2(_0683_),
    .B1(_0685_),
    .B2(net1),
    .C1(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__clkbuf_2 _2071_ (.A(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2072_ (.A(\po_0.regf_0.w_addr[3] ),
    .X(_0695_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2073_ (.A(\po_0.regf_0.w_addr[1] ),
    .X(_0696_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2074_ (.A(\po_0.regf_0.w_addr[0] ),
    .X(_0697_));
 sky130_fd_sc_hd__and3_1 _2075_ (.A(_0696_),
    .B(_0697_),
    .C(\po_0.regf_0.w_wr ),
    .X(_0698_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2076_ (.A(\po_0.regf_0.w_addr[2] ),
    .X(_0699_));
 sky130_fd_sc_hd__and3b_4 _2077_ (.A_N(_0695_),
    .B(_0698_),
    .C(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__clkbuf_4 _2078_ (.A(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _2079_ (.A0(\po_0.regf_0.rf[7][0] ),
    .A1(_0694_),
    .S(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__clkbuf_1 _2080_ (.A(_0702_),
    .X(_0016_));
 sky130_fd_sc_hd__and2_1 _2081_ (.A(\po_0._1_[0] ),
    .B(_1340_),
    .X(_0703_));
 sky130_fd_sc_hd__and2b_1 _2082_ (.A_N(_0574_),
    .B(_0573_),
    .X(_0704_));
 sky130_fd_sc_hd__or3_1 _2083_ (.A(_0703_),
    .B(_0586_),
    .C(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__buf_2 _2084_ (.A(_0689_),
    .X(_0706_));
 sky130_fd_sc_hd__o21ai_2 _2085_ (.A1(_0586_),
    .A2(_0704_),
    .B1(_0703_),
    .Y(_0707_));
 sky130_fd_sc_hd__buf_2 _2086_ (.A(_1316_),
    .X(_0708_));
 sky130_fd_sc_hd__buf_2 _2087_ (.A(_0688_),
    .X(_0709_));
 sky130_fd_sc_hd__a22o_1 _2088_ (.A1(_0708_),
    .A2(\po_0.alu_0._11_[1] ),
    .B1(_0709_),
    .B2(_0574_),
    .X(_0710_));
 sky130_fd_sc_hd__a31o_1 _2089_ (.A1(_0705_),
    .A2(_0706_),
    .A3(_0707_),
    .B1(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__clkbuf_2 _2090_ (.A(_0687_),
    .X(_0712_));
 sky130_fd_sc_hd__clkbuf_2 _2091_ (.A(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__clkbuf_4 _2092_ (.A(\po_0.muxf_0.rf_w_data[1] ),
    .X(_0714_));
 sky130_fd_sc_hd__clkbuf_2 _2093_ (.A(_0684_),
    .X(_0715_));
 sky130_fd_sc_hd__a22o_1 _2094_ (.A1(_0714_),
    .A2(_0683_),
    .B1(_0715_),
    .B2(net8),
    .X(_0716_));
 sky130_fd_sc_hd__a21o_2 _2095_ (.A1(_0711_),
    .A2(_0713_),
    .B1(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__clkbuf_2 _2096_ (.A(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _2097_ (.A0(\po_0.regf_0.rf[7][1] ),
    .A1(_0718_),
    .S(_0701_),
    .X(_0719_));
 sky130_fd_sc_hd__clkbuf_1 _2098_ (.A(_0719_),
    .X(_0017_));
 sky130_fd_sc_hd__buf_2 _2099_ (.A(_0688_),
    .X(_0720_));
 sky130_fd_sc_hd__and2b_1 _2100_ (.A_N(\po_0._1_[2] ),
    .B(net43),
    .X(_0721_));
 sky130_fd_sc_hd__and2b_1 _2101_ (.A_N(_0579_),
    .B(\po_0._1_[2] ),
    .X(_0722_));
 sky130_fd_sc_hd__o21ai_2 _2102_ (.A1(_0582_),
    .A2(_0578_),
    .B1(_0707_),
    .Y(_0723_));
 sky130_fd_sc_hd__or2b_1 _2103_ (.A(\po_0.alu_0.s1 ),
    .B_N(_1313_),
    .X(_0724_));
 sky130_fd_sc_hd__buf_2 _2104_ (.A(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__a21oi_1 _2105_ (.A1(_0593_),
    .A2(_0723_),
    .B1(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__o31a_1 _2106_ (.A1(_0721_),
    .A2(_0722_),
    .A3(_0723_),
    .B1(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__a221o_1 _2107_ (.A1(_1318_),
    .A2(\po_0.alu_0._11_[2] ),
    .B1(_0720_),
    .B2(_0579_),
    .C1(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__clkbuf_4 _2108_ (.A(\po_0.muxf_0.rf_w_data[2] ),
    .X(_0729_));
 sky130_fd_sc_hd__a22o_1 _2109_ (.A1(_0729_),
    .A2(_0682_),
    .B1(_0715_),
    .B2(net9),
    .X(_0730_));
 sky130_fd_sc_hd__a21o_2 _2110_ (.A1(_0728_),
    .A2(_0713_),
    .B1(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__clkbuf_2 _2111_ (.A(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _2112_ (.A0(\po_0.regf_0.rf[7][2] ),
    .A1(_0732_),
    .S(_0701_),
    .X(_0733_));
 sky130_fd_sc_hd__clkbuf_1 _2113_ (.A(_0733_),
    .X(_0018_));
 sky130_fd_sc_hd__nor2_1 _2114_ (.A(_0590_),
    .B(_0591_),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_1 _2115_ (.A(_0579_),
    .B(\po_0._1_[2] ),
    .Y(_0735_));
 sky130_fd_sc_hd__a21bo_1 _2116_ (.A1(_0593_),
    .A2(_0723_),
    .B1_N(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__o21ai_1 _2117_ (.A1(_0734_),
    .A2(_0736_),
    .B1(_0689_),
    .Y(_0737_));
 sky130_fd_sc_hd__a21oi_1 _2118_ (.A1(_0734_),
    .A2(_0736_),
    .B1(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__a211o_1 _2119_ (.A1(_1317_),
    .A2(\po_0.alu_0._11_[3] ),
    .B1(_0688_),
    .C1(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__o311a_1 _2120_ (.A1(_0589_),
    .A2(_0686_),
    .A3(_1314_),
    .B1(_0687_),
    .C1(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__a221o_2 _2121_ (.A1(\po_0.muxf_0.rf_w_data[3] ),
    .A2(_0683_),
    .B1(_0685_),
    .B2(net10),
    .C1(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2122_ (.A(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _2123_ (.A0(\po_0.regf_0.rf[7][3] ),
    .A1(_0742_),
    .S(_0701_),
    .X(_0743_));
 sky130_fd_sc_hd__clkbuf_1 _2124_ (.A(_0743_),
    .X(_0019_));
 sky130_fd_sc_hd__a22o_1 _2125_ (.A1(_1317_),
    .A2(\po_0.alu_0._11_[4] ),
    .B1(_0688_),
    .B2(net84),
    .X(_0744_));
 sky130_fd_sc_hd__o211a_1 _2126_ (.A1(_0721_),
    .A2(_0722_),
    .B1(_0595_),
    .C1(_0596_),
    .X(_0745_));
 sky130_fd_sc_hd__a31o_1 _2127_ (.A1(_0596_),
    .A2(\po_0._1_[2] ),
    .A3(_0579_),
    .B1(_0590_),
    .X(_0746_));
 sky130_fd_sc_hd__a21oi_1 _2128_ (.A1(_0723_),
    .A2(_0745_),
    .B1(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__nand2_1 _2129_ (.A(_0574_),
    .B(_0573_),
    .Y(_0748_));
 sky130_fd_sc_hd__o21ai_1 _2130_ (.A1(_0721_),
    .A2(_0722_),
    .B1(_0734_),
    .Y(_0749_));
 sky130_fd_sc_hd__a21oi_1 _2131_ (.A1(_0707_),
    .A2(_0748_),
    .B1(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__o31a_1 _2132_ (.A1(_0603_),
    .A2(_0746_),
    .A3(_0750_),
    .B1(_0689_),
    .X(_0751_));
 sky130_fd_sc_hd__o31a_1 _2133_ (.A1(_0599_),
    .A2(_0600_),
    .A3(_0747_),
    .B1(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__o21a_1 _2134_ (.A1(_0744_),
    .A2(_0752_),
    .B1(_0712_),
    .X(_0753_));
 sky130_fd_sc_hd__a221o_2 _2135_ (.A1(_0561_),
    .A2(_0683_),
    .B1(_0685_),
    .B2(net11),
    .C1(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__clkbuf_2 _2136_ (.A(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _2137_ (.A0(\po_0.regf_0.rf[7][4] ),
    .A1(_0755_),
    .S(_0701_),
    .X(_0756_));
 sky130_fd_sc_hd__clkbuf_1 _2138_ (.A(_0756_),
    .X(_0020_));
 sky130_fd_sc_hd__o21a_1 _2139_ (.A1(_0746_),
    .A2(_0750_),
    .B1(_0603_),
    .X(_0757_));
 sky130_fd_sc_hd__or3_1 _2140_ (.A(_0599_),
    .B(_0609_),
    .C(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__o21ai_1 _2141_ (.A1(_0599_),
    .A2(_0757_),
    .B1(_0609_),
    .Y(_0759_));
 sky130_fd_sc_hd__and3_1 _2142_ (.A(_0758_),
    .B(_0689_),
    .C(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__a211o_1 _2143_ (.A1(_1318_),
    .A2(\po_0.alu_0._11_[5] ),
    .B1(_0720_),
    .C1(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__or3_1 _2144_ (.A(_0606_),
    .B(_0708_),
    .C(_1313_),
    .X(_0762_));
 sky130_fd_sc_hd__a22o_1 _2145_ (.A1(_0565_),
    .A2(_0682_),
    .B1(_0715_),
    .B2(net12),
    .X(_0763_));
 sky130_fd_sc_hd__a31o_2 _2146_ (.A1(_0761_),
    .A2(_0712_),
    .A3(_0762_),
    .B1(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2147_ (.A(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _2148_ (.A0(\po_0.regf_0.rf[7][5] ),
    .A1(_0765_),
    .S(_0701_),
    .X(_0766_));
 sky130_fd_sc_hd__clkbuf_1 _2149_ (.A(_0766_),
    .X(_0021_));
 sky130_fd_sc_hd__a21boi_1 _2150_ (.A1(_0577_),
    .A2(_0703_),
    .B1_N(_0748_),
    .Y(_0767_));
 sky130_fd_sc_hd__o21bai_2 _2151_ (.A1(_0749_),
    .A2(_0767_),
    .B1_N(_0746_),
    .Y(_0768_));
 sky130_fd_sc_hd__a22o_1 _2152_ (.A1(net45),
    .A2(\po_0._1_[4] ),
    .B1(\po_0._1_[5] ),
    .B2(_0606_),
    .X(_0769_));
 sky130_fd_sc_hd__a21oi_1 _2153_ (.A1(_0768_),
    .A2(_0603_),
    .B1(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__o22ai_1 _2154_ (.A1(_0613_),
    .A2(_0614_),
    .B1(_0770_),
    .B2(_0607_),
    .Y(_0771_));
 sky130_fd_sc_hd__o221ai_2 _2155_ (.A1(_0606_),
    .A2(\po_0._1_[5] ),
    .B1(_0769_),
    .B2(_0757_),
    .C1(_0618_),
    .Y(_0772_));
 sky130_fd_sc_hd__a22o_1 _2156_ (.A1(_0708_),
    .A2(\po_0.alu_0._11_[6] ),
    .B1(_0709_),
    .B2(_1347_),
    .X(_0773_));
 sky130_fd_sc_hd__a31o_1 _2157_ (.A1(_0771_),
    .A2(_0772_),
    .A3(_0706_),
    .B1(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_1 _2158_ (.A1(_0567_),
    .A2(_0682_),
    .B1(_0715_),
    .B2(net13),
    .X(_0775_));
 sky130_fd_sc_hd__a21o_2 _2159_ (.A1(_0774_),
    .A2(_0713_),
    .B1(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2160_ (.A(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__buf_2 _2161_ (.A(_0700_),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_1 _2162_ (.A0(\po_0.regf_0.rf[7][6] ),
    .A1(_0777_),
    .S(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__clkbuf_1 _2163_ (.A(_0779_),
    .X(_0022_));
 sky130_fd_sc_hd__nand2_1 _2164_ (.A(_1347_),
    .B(\po_0._1_[6] ),
    .Y(_0780_));
 sky130_fd_sc_hd__nor2_1 _2165_ (.A(_0622_),
    .B(_0623_),
    .Y(_0781_));
 sky130_fd_sc_hd__a21oi_1 _2166_ (.A1(_0780_),
    .A2(_0772_),
    .B1(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__o311a_1 _2167_ (.A1(_0607_),
    .A2(_0614_),
    .A3(_0770_),
    .B1(_0781_),
    .C1(_0780_),
    .X(_0783_));
 sky130_fd_sc_hd__or2b_1 _2168_ (.A(\po_0.alu_0._11_[7] ),
    .B_N(_1316_),
    .X(_0784_));
 sky130_fd_sc_hd__o311a_1 _2169_ (.A1(_0621_),
    .A2(_1317_),
    .A3(_1313_),
    .B1(_0784_),
    .C1(_0687_),
    .X(_0785_));
 sky130_fd_sc_hd__o31a_1 _2170_ (.A1(_0725_),
    .A2(_0782_),
    .A3(_0783_),
    .B1(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__a221o_2 _2171_ (.A1(\po_0.muxf_0.rf_w_data[7] ),
    .A2(_0683_),
    .B1(_0685_),
    .B2(net14),
    .C1(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2172_ (.A(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__mux2_1 _2173_ (.A0(\po_0.regf_0.rf[7][7] ),
    .A1(_0788_),
    .S(_0778_),
    .X(_0789_));
 sky130_fd_sc_hd__clkbuf_1 _2174_ (.A(_0789_),
    .X(_0023_));
 sky130_fd_sc_hd__buf_2 _2175_ (.A(_0715_),
    .X(_0790_));
 sky130_fd_sc_hd__nand4_1 _2176_ (.A(_0603_),
    .B(_0609_),
    .C(_0618_),
    .D(_0781_),
    .Y(_0791_));
 sky130_fd_sc_hd__a22o_1 _2177_ (.A1(_1347_),
    .A2(\po_0._1_[6] ),
    .B1(\po_0._1_[7] ),
    .B2(_0621_),
    .X(_0792_));
 sky130_fd_sc_hd__nor4b_1 _2178_ (.A(_0607_),
    .B(_0613_),
    .C(_0614_),
    .D_N(_0769_),
    .Y(_0793_));
 sky130_fd_sc_hd__o22a_1 _2179_ (.A1(_0621_),
    .A2(\po_0._1_[7] ),
    .B1(_0792_),
    .B2(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__o21bai_1 _2180_ (.A1(_0791_),
    .A2(_0747_),
    .B1_N(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__nand2_2 _2181_ (.A(_0795_),
    .B(_0648_),
    .Y(_0796_));
 sky130_fd_sc_hd__and4_1 _2182_ (.A(_0603_),
    .B(_0609_),
    .C(_0618_),
    .D(_0781_),
    .X(_0797_));
 sky130_fd_sc_hd__a211o_1 _2183_ (.A1(_0768_),
    .A2(_0797_),
    .B1(_0794_),
    .C1(_0648_),
    .X(_0798_));
 sky130_fd_sc_hd__a22o_1 _2184_ (.A1(_0708_),
    .A2(\po_0.alu_0._11_[8] ),
    .B1(_0709_),
    .B2(net83),
    .X(_0799_));
 sky130_fd_sc_hd__a31o_1 _2185_ (.A1(_0796_),
    .A2(_0706_),
    .A3(_0798_),
    .B1(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__a22o_2 _2186_ (.A1(net15),
    .A2(_0790_),
    .B1(_0800_),
    .B2(_0713_),
    .X(_0801_));
 sky130_fd_sc_hd__clkbuf_2 _2187_ (.A(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _2188_ (.A0(\po_0.regf_0.rf[7][8] ),
    .A1(_0802_),
    .S(_0778_),
    .X(_0803_));
 sky130_fd_sc_hd__clkbuf_1 _2189_ (.A(_0803_),
    .X(_0024_));
 sky130_fd_sc_hd__a21oi_1 _2190_ (.A1(_0628_),
    .A2(_0796_),
    .B1(_0634_),
    .Y(_0804_));
 sky130_fd_sc_hd__a31o_1 _2191_ (.A1(_0628_),
    .A2(_0634_),
    .A3(_0796_),
    .B1(_0724_),
    .X(_0805_));
 sky130_fd_sc_hd__nor2_1 _2192_ (.A(_0804_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__a211o_1 _2193_ (.A1(\po_0.alu_0._11_[9] ),
    .A2(_0725_),
    .B1(_0720_),
    .C1(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__o31a_1 _2194_ (.A1(_0633_),
    .A2(_0686_),
    .A3(_1314_),
    .B1(_0712_),
    .X(_0808_));
 sky130_fd_sc_hd__a22o_2 _2195_ (.A1(net16),
    .A2(_0790_),
    .B1(_0807_),
    .B2(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2196_ (.A(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _2197_ (.A0(\po_0.regf_0.rf[7][9] ),
    .A1(_0810_),
    .S(_0778_),
    .X(_0811_));
 sky130_fd_sc_hd__clkbuf_1 _2198_ (.A(_0811_),
    .X(_0025_));
 sky130_fd_sc_hd__a22oi_2 _2199_ (.A1(net49),
    .A2(\po_0._1_[8] ),
    .B1(\po_0._1_[9] ),
    .B2(_0633_),
    .Y(_0812_));
 sky130_fd_sc_hd__o21ai_1 _2200_ (.A1(_0633_),
    .A2(\po_0._1_[9] ),
    .B1(_0639_),
    .Y(_0813_));
 sky130_fd_sc_hd__a21oi_2 _2201_ (.A1(_0796_),
    .A2(_0812_),
    .B1(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__o2bb2a_1 _2202_ (.A1_N(_0812_),
    .A2_N(_0796_),
    .B1(\po_0._1_[9] ),
    .B2(_0633_),
    .X(_0815_));
 sky130_fd_sc_hd__nor2_1 _2203_ (.A(_0639_),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__a22oi_1 _2204_ (.A1(_0686_),
    .A2(\po_0.alu_0._11_[10] ),
    .B1(_0709_),
    .B2(net36),
    .Y(_0817_));
 sky130_fd_sc_hd__o31ai_1 _2205_ (.A1(_0814_),
    .A2(_0725_),
    .A3(_0816_),
    .B1(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__a22o_2 _2206_ (.A1(net2),
    .A2(_0790_),
    .B1(_0818_),
    .B2(_0713_),
    .X(_0819_));
 sky130_fd_sc_hd__clkbuf_2 _2207_ (.A(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _2208_ (.A0(\po_0.regf_0.rf[7][10] ),
    .A1(_0820_),
    .S(_0778_),
    .X(_0821_));
 sky130_fd_sc_hd__clkbuf_1 _2209_ (.A(_0821_),
    .X(_0026_));
 sky130_fd_sc_hd__a211o_1 _2210_ (.A1(_0650_),
    .A2(_0720_),
    .B1(_0683_),
    .C1(_0715_),
    .X(_0822_));
 sky130_fd_sc_hd__and2_1 _2211_ (.A(net36),
    .B(\po_0._1_[10] ),
    .X(_0823_));
 sky130_fd_sc_hd__o31a_1 _2212_ (.A1(_0823_),
    .A2(_0646_),
    .A3(_0814_),
    .B1(_0706_),
    .X(_0824_));
 sky130_fd_sc_hd__o21ai_2 _2213_ (.A1(_0823_),
    .A2(_0814_),
    .B1(_0646_),
    .Y(_0825_));
 sky130_fd_sc_hd__a221oi_4 _2214_ (.A1(_1318_),
    .A2(\po_0.alu_0._11_[11] ),
    .B1(_0824_),
    .B2(_0825_),
    .C1(_0720_),
    .Y(_0826_));
 sky130_fd_sc_hd__o2bb2ai_4 _2215_ (.A1_N(net3),
    .A2_N(_0790_),
    .B1(_0822_),
    .B2(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__clkbuf_2 _2216_ (.A(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_1 _2217_ (.A0(\po_0.regf_0.rf[7][11] ),
    .A1(_0828_),
    .S(_0778_),
    .X(_0829_));
 sky130_fd_sc_hd__clkbuf_1 _2218_ (.A(_0829_),
    .X(_0027_));
 sky130_fd_sc_hd__a21oi_1 _2219_ (.A1(net37),
    .A2(\po_0._1_[11] ),
    .B1(_0823_),
    .Y(_0830_));
 sky130_fd_sc_hd__o21a_1 _2220_ (.A1(_0812_),
    .A2(_0813_),
    .B1(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__nand4_1 _2221_ (.A(_0648_),
    .B(_0640_),
    .C(_0639_),
    .D(_0646_),
    .Y(_0832_));
 sky130_fd_sc_hd__a21oi_1 _2222_ (.A1(_0768_),
    .A2(_0797_),
    .B1(_0794_),
    .Y(_0833_));
 sky130_fd_sc_hd__o22ai_2 _2223_ (.A1(_0644_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__a21o_1 _2224_ (.A1(_0656_),
    .A2(_0657_),
    .B1(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__nand2_1 _2225_ (.A(_0834_),
    .B(_0658_),
    .Y(_0836_));
 sky130_fd_sc_hd__a22o_1 _2226_ (.A1(_0708_),
    .A2(\po_0.alu_0._11_[12] ),
    .B1(_0709_),
    .B2(_0655_),
    .X(_0837_));
 sky130_fd_sc_hd__a31o_1 _2227_ (.A1(_0835_),
    .A2(_0836_),
    .A3(_0706_),
    .B1(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__a22o_2 _2228_ (.A1(net4),
    .A2(_0685_),
    .B1(_0838_),
    .B2(_0713_),
    .X(_0839_));
 sky130_fd_sc_hd__clkbuf_2 _2229_ (.A(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _2230_ (.A0(\po_0.regf_0.rf[7][12] ),
    .A1(_0840_),
    .S(_0700_),
    .X(_0841_));
 sky130_fd_sc_hd__clkbuf_1 _2231_ (.A(_0841_),
    .X(_0028_));
 sky130_fd_sc_hd__xnor2_1 _2232_ (.A(_0659_),
    .B(\po_0._1_[13] ),
    .Y(_0842_));
 sky130_fd_sc_hd__a21oi_1 _2233_ (.A1(_0656_),
    .A2(_0836_),
    .B1(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__a31o_1 _2234_ (.A1(_0656_),
    .A2(_0842_),
    .A3(_0836_),
    .B1(_0725_),
    .X(_0844_));
 sky130_fd_sc_hd__a21oi_1 _2235_ (.A1(_1318_),
    .A2(\po_0.alu_0._11_[13] ),
    .B1(_0709_),
    .Y(_0845_));
 sky130_fd_sc_hd__o21ai_1 _2236_ (.A1(_0843_),
    .A2(_0844_),
    .B1(_0845_),
    .Y(_0846_));
 sky130_fd_sc_hd__or3_1 _2237_ (.A(_0659_),
    .B(_0708_),
    .C(_1313_),
    .X(_0847_));
 sky130_fd_sc_hd__a32o_2 _2238_ (.A1(_0846_),
    .A2(_0847_),
    .A3(_0712_),
    .B1(_0790_),
    .B2(net5),
    .X(_0848_));
 sky130_fd_sc_hd__clkbuf_2 _2239_ (.A(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _2240_ (.A0(\po_0.regf_0.rf[7][13] ),
    .A1(_0849_),
    .S(_0700_),
    .X(_0850_));
 sky130_fd_sc_hd__clkbuf_1 _2241_ (.A(_0850_),
    .X(_0029_));
 sky130_fd_sc_hd__and3_1 _2242_ (.A(_0660_),
    .B(_0657_),
    .C(_0656_),
    .X(_0851_));
 sky130_fd_sc_hd__nand2_1 _2243_ (.A(_0834_),
    .B(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__o211a_1 _2244_ (.A1(_0659_),
    .A2(\po_0._1_[13] ),
    .B1(\po_0._1_[12] ),
    .C1(_0655_),
    .X(_0853_));
 sky130_fd_sc_hd__a21oi_1 _2245_ (.A1(_0659_),
    .A2(\po_0._1_[13] ),
    .B1(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__a21oi_1 _2246_ (.A1(_0852_),
    .A2(_0854_),
    .B1(_0670_),
    .Y(_0855_));
 sky130_fd_sc_hd__a31o_1 _2247_ (.A1(_0670_),
    .A2(_0852_),
    .A3(_0854_),
    .B1(_0725_),
    .X(_0856_));
 sky130_fd_sc_hd__a22oi_1 _2248_ (.A1(_0686_),
    .A2(\po_0.alu_0._11_[14] ),
    .B1(_0720_),
    .B2(net40),
    .Y(_0857_));
 sky130_fd_sc_hd__o21ai_1 _2249_ (.A1(_0855_),
    .A2(_0856_),
    .B1(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__a22o_2 _2250_ (.A1(net6),
    .A2(_0685_),
    .B1(_0858_),
    .B2(_0712_),
    .X(_0859_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2251_ (.A(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _2252_ (.A0(\po_0.regf_0.rf[7][14] ),
    .A1(_0860_),
    .S(_0700_),
    .X(_0861_));
 sky130_fd_sc_hd__clkbuf_1 _2253_ (.A(_0861_),
    .X(_0030_));
 sky130_fd_sc_hd__nand2_1 _2254_ (.A(net7),
    .B(_0790_),
    .Y(_0862_));
 sky130_fd_sc_hd__o22a_1 _2255_ (.A1(_0673_),
    .A2(_0674_),
    .B1(_0855_),
    .B2(_0668_),
    .X(_0863_));
 sky130_fd_sc_hd__or2_1 _2256_ (.A(_0673_),
    .B(_0674_),
    .X(_0864_));
 sky130_fd_sc_hd__o31ai_1 _2257_ (.A1(_0668_),
    .A2(_0864_),
    .A3(_0855_),
    .B1(_0706_),
    .Y(_0865_));
 sky130_fd_sc_hd__or2b_1 _2258_ (.A(\po_0.alu_0._11_[15] ),
    .B_N(_1317_),
    .X(_0866_));
 sky130_fd_sc_hd__o311a_1 _2259_ (.A1(net41),
    .A2(_0686_),
    .A3(_1314_),
    .B1(_0866_),
    .C1(_0687_),
    .X(_0867_));
 sky130_fd_sc_hd__o21ai_1 _2260_ (.A1(_0863_),
    .A2(_0865_),
    .B1(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__nand2_2 _2261_ (.A(_0862_),
    .B(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__clkbuf_2 _2262_ (.A(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_1 _2263_ (.A0(\po_0.regf_0.rf[7][15] ),
    .A1(_0870_),
    .S(_0700_),
    .X(_0871_));
 sky130_fd_sc_hd__clkbuf_1 _2264_ (.A(_0871_),
    .X(_0031_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2265_ (.A(\po_0.regf_0.w_wr ),
    .X(_0872_));
 sky130_fd_sc_hd__clkbuf_2 _2266_ (.A(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__and2b_1 _2267_ (.A_N(\po_0.regf_0.w_addr[1] ),
    .B(\po_0.regf_0.w_addr[0] ),
    .X(_0874_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2268_ (.A(\po_0.regf_0.w_addr[2] ),
    .X(_0875_));
 sky130_fd_sc_hd__and4b_4 _2269_ (.A_N(_0695_),
    .B(_0873_),
    .C(_0874_),
    .D(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__clkbuf_4 _2270_ (.A(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _2271_ (.A0(\po_0.regf_0.rf[5][0] ),
    .A1(_0694_),
    .S(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__clkbuf_1 _2272_ (.A(_0878_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2273_ (.A0(\po_0.regf_0.rf[5][1] ),
    .A1(_0718_),
    .S(_0877_),
    .X(_0879_));
 sky130_fd_sc_hd__clkbuf_1 _2274_ (.A(_0879_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _2275_ (.A0(\po_0.regf_0.rf[5][2] ),
    .A1(_0732_),
    .S(_0877_),
    .X(_0880_));
 sky130_fd_sc_hd__clkbuf_1 _2276_ (.A(_0880_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2277_ (.A0(\po_0.regf_0.rf[5][3] ),
    .A1(_0742_),
    .S(_0877_),
    .X(_0881_));
 sky130_fd_sc_hd__clkbuf_1 _2278_ (.A(_0881_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2279_ (.A0(\po_0.regf_0.rf[5][4] ),
    .A1(_0755_),
    .S(_0877_),
    .X(_0882_));
 sky130_fd_sc_hd__clkbuf_1 _2280_ (.A(_0882_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2281_ (.A0(\po_0.regf_0.rf[5][5] ),
    .A1(_0765_),
    .S(_0877_),
    .X(_0883_));
 sky130_fd_sc_hd__clkbuf_1 _2282_ (.A(_0883_),
    .X(_0037_));
 sky130_fd_sc_hd__buf_2 _2283_ (.A(_0876_),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _2284_ (.A0(\po_0.regf_0.rf[5][6] ),
    .A1(_0777_),
    .S(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__clkbuf_1 _2285_ (.A(_0885_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2286_ (.A0(\po_0.regf_0.rf[5][7] ),
    .A1(_0788_),
    .S(_0884_),
    .X(_0886_));
 sky130_fd_sc_hd__clkbuf_1 _2287_ (.A(_0886_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2288_ (.A0(\po_0.regf_0.rf[5][8] ),
    .A1(_0802_),
    .S(_0884_),
    .X(_0887_));
 sky130_fd_sc_hd__clkbuf_1 _2289_ (.A(_0887_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2290_ (.A0(\po_0.regf_0.rf[5][9] ),
    .A1(_0810_),
    .S(_0884_),
    .X(_0888_));
 sky130_fd_sc_hd__clkbuf_1 _2291_ (.A(_0888_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _2292_ (.A0(\po_0.regf_0.rf[5][10] ),
    .A1(_0820_),
    .S(_0884_),
    .X(_0889_));
 sky130_fd_sc_hd__clkbuf_1 _2293_ (.A(_0889_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _2294_ (.A0(\po_0.regf_0.rf[5][11] ),
    .A1(_0828_),
    .S(_0884_),
    .X(_0890_));
 sky130_fd_sc_hd__clkbuf_1 _2295_ (.A(_0890_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _2296_ (.A0(\po_0.regf_0.rf[5][12] ),
    .A1(_0840_),
    .S(_0876_),
    .X(_0891_));
 sky130_fd_sc_hd__clkbuf_1 _2297_ (.A(_0891_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _2298_ (.A0(\po_0.regf_0.rf[5][13] ),
    .A1(_0849_),
    .S(_0876_),
    .X(_0892_));
 sky130_fd_sc_hd__clkbuf_1 _2299_ (.A(_0892_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2300_ (.A0(\po_0.regf_0.rf[5][14] ),
    .A1(_0860_),
    .S(_0876_),
    .X(_0893_));
 sky130_fd_sc_hd__clkbuf_1 _2301_ (.A(_0893_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2302_ (.A0(\po_0.regf_0.rf[5][15] ),
    .A1(_0870_),
    .S(_0876_),
    .X(_0894_));
 sky130_fd_sc_hd__clkbuf_1 _2303_ (.A(_0894_),
    .X(_0047_));
 sky130_fd_sc_hd__and2b_1 _2304_ (.A_N(\po_0.regf_0.w_addr[0] ),
    .B(\po_0.regf_0.w_addr[1] ),
    .X(_0895_));
 sky130_fd_sc_hd__and4b_4 _2305_ (.A_N(_0695_),
    .B(_0873_),
    .C(_0895_),
    .D(_0875_),
    .X(_0896_));
 sky130_fd_sc_hd__clkbuf_4 _2306_ (.A(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _2307_ (.A0(\po_0.regf_0.rf[6][0] ),
    .A1(_0694_),
    .S(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__clkbuf_1 _2308_ (.A(_0898_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _2309_ (.A0(\po_0.regf_0.rf[6][1] ),
    .A1(_0718_),
    .S(_0897_),
    .X(_0899_));
 sky130_fd_sc_hd__clkbuf_1 _2310_ (.A(_0899_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _2311_ (.A0(\po_0.regf_0.rf[6][2] ),
    .A1(_0732_),
    .S(_0897_),
    .X(_0900_));
 sky130_fd_sc_hd__clkbuf_1 _2312_ (.A(_0900_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _2313_ (.A0(\po_0.regf_0.rf[6][3] ),
    .A1(_0742_),
    .S(_0897_),
    .X(_0901_));
 sky130_fd_sc_hd__clkbuf_1 _2314_ (.A(_0901_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _2315_ (.A0(\po_0.regf_0.rf[6][4] ),
    .A1(_0755_),
    .S(_0897_),
    .X(_0902_));
 sky130_fd_sc_hd__clkbuf_1 _2316_ (.A(_0902_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _2317_ (.A0(\po_0.regf_0.rf[6][5] ),
    .A1(_0765_),
    .S(_0897_),
    .X(_0903_));
 sky130_fd_sc_hd__clkbuf_1 _2318_ (.A(_0903_),
    .X(_0053_));
 sky130_fd_sc_hd__clkbuf_4 _2319_ (.A(_0896_),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _2320_ (.A0(\po_0.regf_0.rf[6][6] ),
    .A1(_0777_),
    .S(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__clkbuf_1 _2321_ (.A(_0905_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2322_ (.A0(\po_0.regf_0.rf[6][7] ),
    .A1(_0788_),
    .S(_0904_),
    .X(_0906_));
 sky130_fd_sc_hd__clkbuf_1 _2323_ (.A(_0906_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2324_ (.A0(\po_0.regf_0.rf[6][8] ),
    .A1(_0802_),
    .S(_0904_),
    .X(_0907_));
 sky130_fd_sc_hd__clkbuf_1 _2325_ (.A(_0907_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2326_ (.A0(\po_0.regf_0.rf[6][9] ),
    .A1(_0810_),
    .S(_0904_),
    .X(_0908_));
 sky130_fd_sc_hd__clkbuf_1 _2327_ (.A(_0908_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2328_ (.A0(\po_0.regf_0.rf[6][10] ),
    .A1(_0820_),
    .S(_0904_),
    .X(_0909_));
 sky130_fd_sc_hd__clkbuf_1 _2329_ (.A(_0909_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _2330_ (.A0(\po_0.regf_0.rf[6][11] ),
    .A1(_0828_),
    .S(_0904_),
    .X(_0910_));
 sky130_fd_sc_hd__clkbuf_1 _2331_ (.A(_0910_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _2332_ (.A0(\po_0.regf_0.rf[6][12] ),
    .A1(_0840_),
    .S(_0896_),
    .X(_0911_));
 sky130_fd_sc_hd__clkbuf_1 _2333_ (.A(_0911_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _2334_ (.A0(\po_0.regf_0.rf[6][13] ),
    .A1(_0849_),
    .S(_0896_),
    .X(_0912_));
 sky130_fd_sc_hd__clkbuf_1 _2335_ (.A(_0912_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2336_ (.A0(\po_0.regf_0.rf[6][14] ),
    .A1(_0860_),
    .S(_0896_),
    .X(_0913_));
 sky130_fd_sc_hd__clkbuf_1 _2337_ (.A(_0913_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2338_ (.A0(\po_0.regf_0.rf[6][15] ),
    .A1(_0870_),
    .S(_0896_),
    .X(_0914_));
 sky130_fd_sc_hd__clkbuf_1 _2339_ (.A(_0914_),
    .X(_0063_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2340_ (.A(\po_0.regf_0.w_addr[3] ),
    .X(_0915_));
 sky130_fd_sc_hd__and4b_4 _2341_ (.A_N(_0875_),
    .B(_0915_),
    .C(_0873_),
    .D(_0874_),
    .X(_0916_));
 sky130_fd_sc_hd__clkbuf_4 _2342_ (.A(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _2343_ (.A0(\po_0.regf_0.rf[9][0] ),
    .A1(_0694_),
    .S(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__clkbuf_1 _2344_ (.A(_0918_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _2345_ (.A0(\po_0.regf_0.rf[9][1] ),
    .A1(_0718_),
    .S(_0917_),
    .X(_0919_));
 sky130_fd_sc_hd__clkbuf_1 _2346_ (.A(_0919_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _2347_ (.A0(\po_0.regf_0.rf[9][2] ),
    .A1(_0732_),
    .S(_0917_),
    .X(_0920_));
 sky130_fd_sc_hd__clkbuf_1 _2348_ (.A(_0920_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _2349_ (.A0(\po_0.regf_0.rf[9][3] ),
    .A1(_0742_),
    .S(_0917_),
    .X(_0921_));
 sky130_fd_sc_hd__clkbuf_1 _2350_ (.A(_0921_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _2351_ (.A0(\po_0.regf_0.rf[9][4] ),
    .A1(_0755_),
    .S(_0917_),
    .X(_0922_));
 sky130_fd_sc_hd__clkbuf_1 _2352_ (.A(_0922_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2353_ (.A0(\po_0.regf_0.rf[9][5] ),
    .A1(_0765_),
    .S(_0917_),
    .X(_0923_));
 sky130_fd_sc_hd__clkbuf_1 _2354_ (.A(_0923_),
    .X(_0069_));
 sky130_fd_sc_hd__clkbuf_4 _2355_ (.A(_0916_),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_1 _2356_ (.A0(\po_0.regf_0.rf[9][6] ),
    .A1(_0777_),
    .S(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_1 _2357_ (.A(_0925_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _2358_ (.A0(\po_0.regf_0.rf[9][7] ),
    .A1(_0788_),
    .S(_0924_),
    .X(_0926_));
 sky130_fd_sc_hd__clkbuf_1 _2359_ (.A(_0926_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _2360_ (.A0(\po_0.regf_0.rf[9][8] ),
    .A1(_0802_),
    .S(_0924_),
    .X(_0927_));
 sky130_fd_sc_hd__clkbuf_1 _2361_ (.A(_0927_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _2362_ (.A0(\po_0.regf_0.rf[9][9] ),
    .A1(_0810_),
    .S(_0924_),
    .X(_0928_));
 sky130_fd_sc_hd__clkbuf_1 _2363_ (.A(_0928_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2364_ (.A0(\po_0.regf_0.rf[9][10] ),
    .A1(_0820_),
    .S(_0924_),
    .X(_0929_));
 sky130_fd_sc_hd__clkbuf_1 _2365_ (.A(_0929_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _2366_ (.A0(\po_0.regf_0.rf[9][11] ),
    .A1(_0828_),
    .S(_0924_),
    .X(_0930_));
 sky130_fd_sc_hd__clkbuf_1 _2367_ (.A(_0930_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _2368_ (.A0(\po_0.regf_0.rf[9][12] ),
    .A1(_0840_),
    .S(_0916_),
    .X(_0931_));
 sky130_fd_sc_hd__clkbuf_1 _2369_ (.A(_0931_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2370_ (.A0(\po_0.regf_0.rf[9][13] ),
    .A1(_0849_),
    .S(_0916_),
    .X(_0932_));
 sky130_fd_sc_hd__clkbuf_1 _2371_ (.A(_0932_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2372_ (.A0(\po_0.regf_0.rf[9][14] ),
    .A1(_0860_),
    .S(_0916_),
    .X(_0933_));
 sky130_fd_sc_hd__clkbuf_1 _2373_ (.A(_0933_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _2374_ (.A0(\po_0.regf_0.rf[9][15] ),
    .A1(_0870_),
    .S(_0916_),
    .X(_0934_));
 sky130_fd_sc_hd__clkbuf_1 _2375_ (.A(_0934_),
    .X(_0079_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2376_ (.A(_0872_),
    .X(_0935_));
 sky130_fd_sc_hd__nor2_1 _2377_ (.A(\po_0.regf_0.w_addr[2] ),
    .B(\po_0.regf_0.w_addr[3] ),
    .Y(_0936_));
 sky130_fd_sc_hd__and3_4 _2378_ (.A(_0935_),
    .B(_0874_),
    .C(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__clkbuf_4 _2379_ (.A(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_1 _2380_ (.A0(\po_0.regf_0.rf[1][0] ),
    .A1(_0694_),
    .S(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__clkbuf_1 _2381_ (.A(_0939_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2382_ (.A0(\po_0.regf_0.rf[1][1] ),
    .A1(_0718_),
    .S(_0938_),
    .X(_0940_));
 sky130_fd_sc_hd__clkbuf_1 _2383_ (.A(_0940_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2384_ (.A0(\po_0.regf_0.rf[1][2] ),
    .A1(_0732_),
    .S(_0938_),
    .X(_0941_));
 sky130_fd_sc_hd__clkbuf_1 _2385_ (.A(_0941_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2386_ (.A0(\po_0.regf_0.rf[1][3] ),
    .A1(_0742_),
    .S(_0938_),
    .X(_0942_));
 sky130_fd_sc_hd__clkbuf_1 _2387_ (.A(_0942_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2388_ (.A0(\po_0.regf_0.rf[1][4] ),
    .A1(_0755_),
    .S(_0938_),
    .X(_0943_));
 sky130_fd_sc_hd__clkbuf_1 _2389_ (.A(_0943_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2390_ (.A0(\po_0.regf_0.rf[1][5] ),
    .A1(_0765_),
    .S(_0938_),
    .X(_0944_));
 sky130_fd_sc_hd__clkbuf_1 _2391_ (.A(_0944_),
    .X(_0085_));
 sky130_fd_sc_hd__buf_2 _2392_ (.A(_0937_),
    .X(_0945_));
 sky130_fd_sc_hd__mux2_1 _2393_ (.A0(\po_0.regf_0.rf[1][6] ),
    .A1(_0777_),
    .S(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__clkbuf_1 _2394_ (.A(_0946_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2395_ (.A0(\po_0.regf_0.rf[1][7] ),
    .A1(_0788_),
    .S(_0945_),
    .X(_0947_));
 sky130_fd_sc_hd__clkbuf_1 _2396_ (.A(_0947_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2397_ (.A0(\po_0.regf_0.rf[1][8] ),
    .A1(_0802_),
    .S(_0945_),
    .X(_0948_));
 sky130_fd_sc_hd__clkbuf_1 _2398_ (.A(_0948_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2399_ (.A0(\po_0.regf_0.rf[1][9] ),
    .A1(_0810_),
    .S(_0945_),
    .X(_0949_));
 sky130_fd_sc_hd__clkbuf_1 _2400_ (.A(_0949_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2401_ (.A0(\po_0.regf_0.rf[1][10] ),
    .A1(_0820_),
    .S(_0945_),
    .X(_0950_));
 sky130_fd_sc_hd__clkbuf_1 _2402_ (.A(_0950_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(\po_0.regf_0.rf[1][11] ),
    .A1(_0828_),
    .S(_0945_),
    .X(_0951_));
 sky130_fd_sc_hd__clkbuf_1 _2404_ (.A(_0951_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _2405_ (.A0(\po_0.regf_0.rf[1][12] ),
    .A1(_0840_),
    .S(_0937_),
    .X(_0952_));
 sky130_fd_sc_hd__clkbuf_1 _2406_ (.A(_0952_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2407_ (.A0(\po_0.regf_0.rf[1][13] ),
    .A1(_0849_),
    .S(_0937_),
    .X(_0953_));
 sky130_fd_sc_hd__clkbuf_1 _2408_ (.A(_0953_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2409_ (.A0(\po_0.regf_0.rf[1][14] ),
    .A1(_0860_),
    .S(_0937_),
    .X(_0954_));
 sky130_fd_sc_hd__clkbuf_1 _2410_ (.A(_0954_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(\po_0.regf_0.rf[1][15] ),
    .A1(_0870_),
    .S(_0937_),
    .X(_0955_));
 sky130_fd_sc_hd__clkbuf_1 _2412_ (.A(_0955_),
    .X(_0095_));
 sky130_fd_sc_hd__clkbuf_2 _2413_ (.A(_0693_),
    .X(_0956_));
 sky130_fd_sc_hd__and3_1 _2414_ (.A(\po_0.regf_0.w_addr[2] ),
    .B(\po_0.regf_0.w_addr[3] ),
    .C(_0872_),
    .X(_0957_));
 sky130_fd_sc_hd__and3_2 _2415_ (.A(_0696_),
    .B(_0697_),
    .C(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__buf_2 _2416_ (.A(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _2417_ (.A0(\po_0.regf_0.rf[15][0] ),
    .A1(_0956_),
    .S(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__clkbuf_1 _2418_ (.A(_0960_),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_2 _2419_ (.A(_0717_),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _2420_ (.A0(\po_0.regf_0.rf[15][1] ),
    .A1(_0961_),
    .S(_0959_),
    .X(_0962_));
 sky130_fd_sc_hd__clkbuf_1 _2421_ (.A(_0962_),
    .X(_0097_));
 sky130_fd_sc_hd__clkbuf_2 _2422_ (.A(_0731_),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_1 _2423_ (.A0(\po_0.regf_0.rf[15][2] ),
    .A1(_0963_),
    .S(_0959_),
    .X(_0964_));
 sky130_fd_sc_hd__clkbuf_1 _2424_ (.A(_0964_),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_2 _2425_ (.A(_0741_),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_1 _2426_ (.A0(\po_0.regf_0.rf[15][3] ),
    .A1(_0965_),
    .S(_0959_),
    .X(_0966_));
 sky130_fd_sc_hd__clkbuf_1 _2427_ (.A(_0966_),
    .X(_0099_));
 sky130_fd_sc_hd__clkbuf_2 _2428_ (.A(_0754_),
    .X(_0967_));
 sky130_fd_sc_hd__mux2_1 _2429_ (.A0(\po_0.regf_0.rf[15][4] ),
    .A1(_0967_),
    .S(_0959_),
    .X(_0968_));
 sky130_fd_sc_hd__clkbuf_1 _2430_ (.A(_0968_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_2 _2431_ (.A(_0764_),
    .X(_0969_));
 sky130_fd_sc_hd__mux2_1 _2432_ (.A0(\po_0.regf_0.rf[15][5] ),
    .A1(_0969_),
    .S(_0959_),
    .X(_0970_));
 sky130_fd_sc_hd__clkbuf_1 _2433_ (.A(_0970_),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_2 _2434_ (.A(_0776_),
    .X(_0971_));
 sky130_fd_sc_hd__buf_2 _2435_ (.A(_0958_),
    .X(_0972_));
 sky130_fd_sc_hd__mux2_1 _2436_ (.A0(\po_0.regf_0.rf[15][6] ),
    .A1(_0971_),
    .S(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__clkbuf_1 _2437_ (.A(_0973_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_2 _2438_ (.A(_0787_),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_1 _2439_ (.A0(\po_0.regf_0.rf[15][7] ),
    .A1(_0974_),
    .S(_0972_),
    .X(_0975_));
 sky130_fd_sc_hd__clkbuf_1 _2440_ (.A(_0975_),
    .X(_0103_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2441_ (.A(_0801_),
    .X(_0976_));
 sky130_fd_sc_hd__mux2_1 _2442_ (.A0(\po_0.regf_0.rf[15][8] ),
    .A1(_0976_),
    .S(_0972_),
    .X(_0977_));
 sky130_fd_sc_hd__clkbuf_1 _2443_ (.A(_0977_),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_2 _2444_ (.A(_0809_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _2445_ (.A0(\po_0.regf_0.rf[15][9] ),
    .A1(_0978_),
    .S(_0972_),
    .X(_0979_));
 sky130_fd_sc_hd__clkbuf_1 _2446_ (.A(_0979_),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_2 _2447_ (.A(_0819_),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_1 _2448_ (.A0(\po_0.regf_0.rf[15][10] ),
    .A1(_0980_),
    .S(_0972_),
    .X(_0981_));
 sky130_fd_sc_hd__clkbuf_1 _2449_ (.A(_0981_),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_2 _2450_ (.A(_0827_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _2451_ (.A0(\po_0.regf_0.rf[15][11] ),
    .A1(_0982_),
    .S(_0972_),
    .X(_0983_));
 sky130_fd_sc_hd__clkbuf_1 _2452_ (.A(_0983_),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_2 _2453_ (.A(_0839_),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _2454_ (.A0(\po_0.regf_0.rf[15][12] ),
    .A1(_0984_),
    .S(_0958_),
    .X(_0985_));
 sky130_fd_sc_hd__clkbuf_1 _2455_ (.A(_0985_),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_2 _2456_ (.A(_0848_),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_1 _2457_ (.A0(\po_0.regf_0.rf[15][13] ),
    .A1(_0986_),
    .S(_0958_),
    .X(_0987_));
 sky130_fd_sc_hd__clkbuf_1 _2458_ (.A(_0987_),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_2 _2459_ (.A(_0859_),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_1 _2460_ (.A0(\po_0.regf_0.rf[15][14] ),
    .A1(_0988_),
    .S(_0958_),
    .X(_0989_));
 sky130_fd_sc_hd__clkbuf_1 _2461_ (.A(_0989_),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_2 _2462_ (.A(_0869_),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_1 _2463_ (.A0(\po_0.regf_0.rf[15][15] ),
    .A1(_0990_),
    .S(_0958_),
    .X(_0991_));
 sky130_fd_sc_hd__clkbuf_1 _2464_ (.A(_0991_),
    .X(_0111_));
 sky130_fd_sc_hd__and4_2 _2465_ (.A(_0699_),
    .B(_0915_),
    .C(_0935_),
    .D(_0895_),
    .X(_0992_));
 sky130_fd_sc_hd__buf_2 _2466_ (.A(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__mux2_1 _2467_ (.A0(\po_0.regf_0.rf[14][0] ),
    .A1(_0956_),
    .S(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__clkbuf_1 _2468_ (.A(_0994_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _2469_ (.A0(\po_0.regf_0.rf[14][1] ),
    .A1(_0961_),
    .S(_0993_),
    .X(_0995_));
 sky130_fd_sc_hd__clkbuf_1 _2470_ (.A(_0995_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _2471_ (.A0(\po_0.regf_0.rf[14][2] ),
    .A1(_0963_),
    .S(_0993_),
    .X(_0996_));
 sky130_fd_sc_hd__clkbuf_1 _2472_ (.A(_0996_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _2473_ (.A0(\po_0.regf_0.rf[14][3] ),
    .A1(_0965_),
    .S(_0993_),
    .X(_0997_));
 sky130_fd_sc_hd__clkbuf_1 _2474_ (.A(_0997_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _2475_ (.A0(\po_0.regf_0.rf[14][4] ),
    .A1(_0967_),
    .S(_0993_),
    .X(_0998_));
 sky130_fd_sc_hd__clkbuf_1 _2476_ (.A(_0998_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _2477_ (.A0(\po_0.regf_0.rf[14][5] ),
    .A1(_0969_),
    .S(_0993_),
    .X(_0999_));
 sky130_fd_sc_hd__clkbuf_1 _2478_ (.A(_0999_),
    .X(_0117_));
 sky130_fd_sc_hd__buf_2 _2479_ (.A(_0992_),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_1 _2480_ (.A0(\po_0.regf_0.rf[14][6] ),
    .A1(_0971_),
    .S(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__clkbuf_1 _2481_ (.A(_1001_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _2482_ (.A0(\po_0.regf_0.rf[14][7] ),
    .A1(_0974_),
    .S(_1000_),
    .X(_1002_));
 sky130_fd_sc_hd__clkbuf_1 _2483_ (.A(_1002_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _2484_ (.A0(\po_0.regf_0.rf[14][8] ),
    .A1(_0976_),
    .S(_1000_),
    .X(_1003_));
 sky130_fd_sc_hd__clkbuf_1 _2485_ (.A(_1003_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _2486_ (.A0(\po_0.regf_0.rf[14][9] ),
    .A1(_0978_),
    .S(_1000_),
    .X(_1004_));
 sky130_fd_sc_hd__clkbuf_1 _2487_ (.A(_1004_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2488_ (.A0(\po_0.regf_0.rf[14][10] ),
    .A1(_0980_),
    .S(_1000_),
    .X(_1005_));
 sky130_fd_sc_hd__clkbuf_1 _2489_ (.A(_1005_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _2490_ (.A0(\po_0.regf_0.rf[14][11] ),
    .A1(_0982_),
    .S(_1000_),
    .X(_1006_));
 sky130_fd_sc_hd__clkbuf_1 _2491_ (.A(_1006_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _2492_ (.A0(\po_0.regf_0.rf[14][12] ),
    .A1(_0984_),
    .S(_0992_),
    .X(_1007_));
 sky130_fd_sc_hd__clkbuf_1 _2493_ (.A(_1007_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _2494_ (.A0(\po_0.regf_0.rf[14][13] ),
    .A1(_0986_),
    .S(_0992_),
    .X(_1008_));
 sky130_fd_sc_hd__clkbuf_1 _2495_ (.A(_1008_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2496_ (.A0(\po_0.regf_0.rf[14][14] ),
    .A1(_0988_),
    .S(_0992_),
    .X(_1009_));
 sky130_fd_sc_hd__clkbuf_1 _2497_ (.A(_1009_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _2498_ (.A0(\po_0.regf_0.rf[14][15] ),
    .A1(_0990_),
    .S(_0992_),
    .X(_1010_));
 sky130_fd_sc_hd__clkbuf_1 _2499_ (.A(_1010_),
    .X(_0127_));
 sky130_fd_sc_hd__and4_2 _2500_ (.A(_0699_),
    .B(_0915_),
    .C(_0935_),
    .D(_0874_),
    .X(_1011_));
 sky130_fd_sc_hd__buf_2 _2501_ (.A(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_1 _2502_ (.A0(\po_0.regf_0.rf[13][0] ),
    .A1(_0956_),
    .S(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__clkbuf_1 _2503_ (.A(_1013_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(\po_0.regf_0.rf[13][1] ),
    .A1(_0961_),
    .S(_1012_),
    .X(_1014_));
 sky130_fd_sc_hd__clkbuf_1 _2505_ (.A(_1014_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(\po_0.regf_0.rf[13][2] ),
    .A1(_0963_),
    .S(_1012_),
    .X(_1015_));
 sky130_fd_sc_hd__clkbuf_1 _2507_ (.A(_1015_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _2508_ (.A0(\po_0.regf_0.rf[13][3] ),
    .A1(_0965_),
    .S(_1012_),
    .X(_1016_));
 sky130_fd_sc_hd__clkbuf_1 _2509_ (.A(_1016_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(\po_0.regf_0.rf[13][4] ),
    .A1(_0967_),
    .S(_1012_),
    .X(_1017_));
 sky130_fd_sc_hd__clkbuf_1 _2511_ (.A(_1017_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(\po_0.regf_0.rf[13][5] ),
    .A1(_0969_),
    .S(_1012_),
    .X(_1018_));
 sky130_fd_sc_hd__clkbuf_1 _2513_ (.A(_1018_),
    .X(_0133_));
 sky130_fd_sc_hd__buf_2 _2514_ (.A(_1011_),
    .X(_1019_));
 sky130_fd_sc_hd__mux2_1 _2515_ (.A0(\po_0.regf_0.rf[13][6] ),
    .A1(_0971_),
    .S(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__clkbuf_1 _2516_ (.A(_1020_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(\po_0.regf_0.rf[13][7] ),
    .A1(_0974_),
    .S(_1019_),
    .X(_1021_));
 sky130_fd_sc_hd__clkbuf_1 _2518_ (.A(_1021_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _2519_ (.A0(\po_0.regf_0.rf[13][8] ),
    .A1(_0976_),
    .S(_1019_),
    .X(_1022_));
 sky130_fd_sc_hd__clkbuf_1 _2520_ (.A(_1022_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _2521_ (.A0(\po_0.regf_0.rf[13][9] ),
    .A1(_0978_),
    .S(_1019_),
    .X(_1023_));
 sky130_fd_sc_hd__clkbuf_1 _2522_ (.A(_1023_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(\po_0.regf_0.rf[13][10] ),
    .A1(_0980_),
    .S(_1019_),
    .X(_1024_));
 sky130_fd_sc_hd__clkbuf_1 _2524_ (.A(_1024_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(\po_0.regf_0.rf[13][11] ),
    .A1(_0982_),
    .S(_1019_),
    .X(_1025_));
 sky130_fd_sc_hd__clkbuf_1 _2526_ (.A(_1025_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _2527_ (.A0(\po_0.regf_0.rf[13][12] ),
    .A1(_0984_),
    .S(_1011_),
    .X(_1026_));
 sky130_fd_sc_hd__clkbuf_1 _2528_ (.A(_1026_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _2529_ (.A0(\po_0.regf_0.rf[13][13] ),
    .A1(_0986_),
    .S(_1011_),
    .X(_1027_));
 sky130_fd_sc_hd__clkbuf_1 _2530_ (.A(_1027_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(\po_0.regf_0.rf[13][14] ),
    .A1(_0988_),
    .S(_1011_),
    .X(_1028_));
 sky130_fd_sc_hd__clkbuf_1 _2532_ (.A(_1028_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _2533_ (.A0(\po_0.regf_0.rf[13][15] ),
    .A1(_0990_),
    .S(_1011_),
    .X(_1029_));
 sky130_fd_sc_hd__clkbuf_1 _2534_ (.A(_1029_),
    .X(_0143_));
 sky130_fd_sc_hd__nor2_1 _2535_ (.A(_0696_),
    .B(_0697_),
    .Y(_1030_));
 sky130_fd_sc_hd__and4_2 _2536_ (.A(_0699_),
    .B(_0915_),
    .C(_0873_),
    .D(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__buf_2 _2537_ (.A(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(_0956_),
    .S(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__clkbuf_1 _2539_ (.A(_1033_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2540_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(_0961_),
    .S(_1032_),
    .X(_1034_));
 sky130_fd_sc_hd__clkbuf_1 _2541_ (.A(_1034_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(_0963_),
    .S(_1032_),
    .X(_1035_));
 sky130_fd_sc_hd__clkbuf_1 _2543_ (.A(_1035_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2544_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(_0965_),
    .S(_1032_),
    .X(_1036_));
 sky130_fd_sc_hd__clkbuf_1 _2545_ (.A(_1036_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(_0967_),
    .S(_1032_),
    .X(_1037_));
 sky130_fd_sc_hd__clkbuf_1 _2547_ (.A(_1037_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(_0969_),
    .S(_1032_),
    .X(_1038_));
 sky130_fd_sc_hd__clkbuf_1 _2549_ (.A(_1038_),
    .X(_0149_));
 sky130_fd_sc_hd__buf_2 _2550_ (.A(_1031_),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(_0971_),
    .S(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__clkbuf_1 _2552_ (.A(_1040_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2553_ (.A0(\po_0.regf_0.rf[12][7] ),
    .A1(_0974_),
    .S(_1039_),
    .X(_1041_));
 sky130_fd_sc_hd__clkbuf_1 _2554_ (.A(_1041_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(\po_0.regf_0.rf[12][8] ),
    .A1(_0976_),
    .S(_1039_),
    .X(_1042_));
 sky130_fd_sc_hd__clkbuf_1 _2556_ (.A(_1042_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(\po_0.regf_0.rf[12][9] ),
    .A1(_0978_),
    .S(_1039_),
    .X(_1043_));
 sky130_fd_sc_hd__clkbuf_1 _2558_ (.A(_1043_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2559_ (.A0(\po_0.regf_0.rf[12][10] ),
    .A1(_0980_),
    .S(_1039_),
    .X(_1044_));
 sky130_fd_sc_hd__clkbuf_1 _2560_ (.A(_1044_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(\po_0.regf_0.rf[12][11] ),
    .A1(_0982_),
    .S(_1039_),
    .X(_1045_));
 sky130_fd_sc_hd__clkbuf_1 _2562_ (.A(_1045_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2563_ (.A0(\po_0.regf_0.rf[12][12] ),
    .A1(_0984_),
    .S(_1031_),
    .X(_1046_));
 sky130_fd_sc_hd__clkbuf_1 _2564_ (.A(_1046_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(\po_0.regf_0.rf[12][13] ),
    .A1(_0986_),
    .S(_1031_),
    .X(_1047_));
 sky130_fd_sc_hd__clkbuf_1 _2566_ (.A(_1047_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(\po_0.regf_0.rf[12][14] ),
    .A1(_0988_),
    .S(_1031_),
    .X(_1048_));
 sky130_fd_sc_hd__clkbuf_1 _2568_ (.A(_1048_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(\po_0.regf_0.rf[12][15] ),
    .A1(_0990_),
    .S(_1031_),
    .X(_1049_));
 sky130_fd_sc_hd__clkbuf_1 _2570_ (.A(_1049_),
    .X(_0159_));
 sky130_fd_sc_hd__and3b_1 _2571_ (.A_N(\po_0.regf_0.w_addr[2] ),
    .B(\po_0.regf_0.w_addr[3] ),
    .C(_0872_),
    .X(_1050_));
 sky130_fd_sc_hd__and3_2 _2572_ (.A(_0696_),
    .B(_0697_),
    .C(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__clkbuf_4 _2573_ (.A(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(\po_0.regf_0.rf[11][0] ),
    .A1(_0956_),
    .S(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__clkbuf_1 _2575_ (.A(_1053_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(\po_0.regf_0.rf[11][1] ),
    .A1(_0961_),
    .S(_1052_),
    .X(_1054_));
 sky130_fd_sc_hd__clkbuf_1 _2577_ (.A(_1054_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(\po_0.regf_0.rf[11][2] ),
    .A1(_0963_),
    .S(_1052_),
    .X(_1055_));
 sky130_fd_sc_hd__clkbuf_1 _2579_ (.A(_1055_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(\po_0.regf_0.rf[11][3] ),
    .A1(_0965_),
    .S(_1052_),
    .X(_1056_));
 sky130_fd_sc_hd__clkbuf_1 _2581_ (.A(_1056_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(\po_0.regf_0.rf[11][4] ),
    .A1(_0967_),
    .S(_1052_),
    .X(_1057_));
 sky130_fd_sc_hd__clkbuf_1 _2583_ (.A(_1057_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2584_ (.A0(\po_0.regf_0.rf[11][5] ),
    .A1(_0969_),
    .S(_1052_),
    .X(_1058_));
 sky130_fd_sc_hd__clkbuf_1 _2585_ (.A(_1058_),
    .X(_0165_));
 sky130_fd_sc_hd__buf_2 _2586_ (.A(_1051_),
    .X(_1059_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(\po_0.regf_0.rf[11][6] ),
    .A1(_0971_),
    .S(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__clkbuf_1 _2588_ (.A(_1060_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2589_ (.A0(\po_0.regf_0.rf[11][7] ),
    .A1(_0974_),
    .S(_1059_),
    .X(_1061_));
 sky130_fd_sc_hd__clkbuf_1 _2590_ (.A(_1061_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2591_ (.A0(\po_0.regf_0.rf[11][8] ),
    .A1(_0976_),
    .S(_1059_),
    .X(_1062_));
 sky130_fd_sc_hd__clkbuf_1 _2592_ (.A(_1062_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2593_ (.A0(\po_0.regf_0.rf[11][9] ),
    .A1(_0978_),
    .S(_1059_),
    .X(_1063_));
 sky130_fd_sc_hd__clkbuf_1 _2594_ (.A(_1063_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _2595_ (.A0(\po_0.regf_0.rf[11][10] ),
    .A1(_0980_),
    .S(_1059_),
    .X(_1064_));
 sky130_fd_sc_hd__clkbuf_1 _2596_ (.A(_1064_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2597_ (.A0(\po_0.regf_0.rf[11][11] ),
    .A1(_0982_),
    .S(_1059_),
    .X(_1065_));
 sky130_fd_sc_hd__clkbuf_1 _2598_ (.A(_1065_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _2599_ (.A0(\po_0.regf_0.rf[11][12] ),
    .A1(_0984_),
    .S(_1051_),
    .X(_1066_));
 sky130_fd_sc_hd__clkbuf_1 _2600_ (.A(_1066_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2601_ (.A0(\po_0.regf_0.rf[11][13] ),
    .A1(_0986_),
    .S(_1051_),
    .X(_1067_));
 sky130_fd_sc_hd__clkbuf_1 _2602_ (.A(_1067_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2603_ (.A0(\po_0.regf_0.rf[11][14] ),
    .A1(_0988_),
    .S(_1051_),
    .X(_1068_));
 sky130_fd_sc_hd__clkbuf_1 _2604_ (.A(_1068_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _2605_ (.A0(\po_0.regf_0.rf[11][15] ),
    .A1(_0990_),
    .S(_1051_),
    .X(_1069_));
 sky130_fd_sc_hd__clkbuf_1 _2606_ (.A(_1069_),
    .X(_0175_));
 sky130_fd_sc_hd__and4b_2 _2607_ (.A_N(_0875_),
    .B(_0915_),
    .C(_0872_),
    .D(_0895_),
    .X(_1070_));
 sky130_fd_sc_hd__clkbuf_4 _2608_ (.A(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(\po_0.regf_0.rf[10][0] ),
    .A1(_0956_),
    .S(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__clkbuf_1 _2610_ (.A(_1072_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(\po_0.regf_0.rf[10][1] ),
    .A1(_0961_),
    .S(_1071_),
    .X(_1073_));
 sky130_fd_sc_hd__clkbuf_1 _2612_ (.A(_1073_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2613_ (.A0(\po_0.regf_0.rf[10][2] ),
    .A1(_0963_),
    .S(_1071_),
    .X(_1074_));
 sky130_fd_sc_hd__clkbuf_1 _2614_ (.A(_1074_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2615_ (.A0(\po_0.regf_0.rf[10][3] ),
    .A1(_0965_),
    .S(_1071_),
    .X(_1075_));
 sky130_fd_sc_hd__clkbuf_1 _2616_ (.A(_1075_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _2617_ (.A0(\po_0.regf_0.rf[10][4] ),
    .A1(_0967_),
    .S(_1071_),
    .X(_1076_));
 sky130_fd_sc_hd__clkbuf_1 _2618_ (.A(_1076_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2619_ (.A0(\po_0.regf_0.rf[10][5] ),
    .A1(_0969_),
    .S(_1071_),
    .X(_1077_));
 sky130_fd_sc_hd__clkbuf_1 _2620_ (.A(_1077_),
    .X(_0181_));
 sky130_fd_sc_hd__buf_2 _2621_ (.A(_1070_),
    .X(_1078_));
 sky130_fd_sc_hd__mux2_1 _2622_ (.A0(\po_0.regf_0.rf[10][6] ),
    .A1(_0971_),
    .S(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__clkbuf_1 _2623_ (.A(_1079_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2624_ (.A0(\po_0.regf_0.rf[10][7] ),
    .A1(_0974_),
    .S(_1078_),
    .X(_1080_));
 sky130_fd_sc_hd__clkbuf_1 _2625_ (.A(_1080_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2626_ (.A0(\po_0.regf_0.rf[10][8] ),
    .A1(_0976_),
    .S(_1078_),
    .X(_1081_));
 sky130_fd_sc_hd__clkbuf_1 _2627_ (.A(_1081_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _2628_ (.A0(\po_0.regf_0.rf[10][9] ),
    .A1(_0978_),
    .S(_1078_),
    .X(_1082_));
 sky130_fd_sc_hd__clkbuf_1 _2629_ (.A(_1082_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _2630_ (.A0(\po_0.regf_0.rf[10][10] ),
    .A1(_0980_),
    .S(_1078_),
    .X(_1083_));
 sky130_fd_sc_hd__clkbuf_1 _2631_ (.A(_1083_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(\po_0.regf_0.rf[10][11] ),
    .A1(_0982_),
    .S(_1078_),
    .X(_1084_));
 sky130_fd_sc_hd__clkbuf_1 _2633_ (.A(_1084_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(\po_0.regf_0.rf[10][12] ),
    .A1(_0984_),
    .S(_1070_),
    .X(_1085_));
 sky130_fd_sc_hd__clkbuf_1 _2635_ (.A(_1085_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(\po_0.regf_0.rf[10][13] ),
    .A1(_0986_),
    .S(_1070_),
    .X(_1086_));
 sky130_fd_sc_hd__clkbuf_1 _2637_ (.A(_1086_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _2638_ (.A0(\po_0.regf_0.rf[10][14] ),
    .A1(_0988_),
    .S(_1070_),
    .X(_1087_));
 sky130_fd_sc_hd__clkbuf_1 _2639_ (.A(_1087_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _2640_ (.A0(\po_0.regf_0.rf[10][15] ),
    .A1(_0990_),
    .S(_1070_),
    .X(_1088_));
 sky130_fd_sc_hd__clkbuf_1 _2641_ (.A(_1088_),
    .X(_0191_));
 sky130_fd_sc_hd__or4bb_4 _2642_ (.A(_0699_),
    .B(_0695_),
    .C_N(_0935_),
    .D_N(_1030_),
    .X(_1089_));
 sky130_fd_sc_hd__clkbuf_4 _2643_ (.A(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__mux2_1 _2644_ (.A0(_0694_),
    .A1(\po_0.regf_0.rf[0][0] ),
    .S(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__clkbuf_1 _2645_ (.A(_1091_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _2646_ (.A0(_0718_),
    .A1(\po_0.regf_0.rf[0][1] ),
    .S(_1090_),
    .X(_1092_));
 sky130_fd_sc_hd__clkbuf_1 _2647_ (.A(_1092_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _2648_ (.A0(_0732_),
    .A1(\po_0.regf_0.rf[0][2] ),
    .S(_1090_),
    .X(_1093_));
 sky130_fd_sc_hd__clkbuf_1 _2649_ (.A(_1093_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _2650_ (.A0(_0742_),
    .A1(\po_0.regf_0.rf[0][3] ),
    .S(_1090_),
    .X(_1094_));
 sky130_fd_sc_hd__clkbuf_1 _2651_ (.A(_1094_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _2652_ (.A0(_0755_),
    .A1(\po_0.regf_0.rf[0][4] ),
    .S(_1090_),
    .X(_1095_));
 sky130_fd_sc_hd__clkbuf_1 _2653_ (.A(_1095_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _2654_ (.A0(_0765_),
    .A1(\po_0.regf_0.rf[0][5] ),
    .S(_1090_),
    .X(_1096_));
 sky130_fd_sc_hd__clkbuf_1 _2655_ (.A(_1096_),
    .X(_0197_));
 sky130_fd_sc_hd__buf_2 _2656_ (.A(_1089_),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_1 _2657_ (.A0(_0777_),
    .A1(\po_0.regf_0.rf[0][6] ),
    .S(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__clkbuf_1 _2658_ (.A(_1098_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2659_ (.A0(_0788_),
    .A1(\po_0.regf_0.rf[0][7] ),
    .S(_1097_),
    .X(_1099_));
 sky130_fd_sc_hd__clkbuf_1 _2660_ (.A(_1099_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _2661_ (.A0(_0802_),
    .A1(\po_0.regf_0.rf[0][8] ),
    .S(_1097_),
    .X(_1100_));
 sky130_fd_sc_hd__clkbuf_1 _2662_ (.A(_1100_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2663_ (.A0(_0810_),
    .A1(\po_0.regf_0.rf[0][9] ),
    .S(_1097_),
    .X(_1101_));
 sky130_fd_sc_hd__clkbuf_1 _2664_ (.A(_1101_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2665_ (.A0(_0820_),
    .A1(\po_0.regf_0.rf[0][10] ),
    .S(_1097_),
    .X(_1102_));
 sky130_fd_sc_hd__clkbuf_1 _2666_ (.A(_1102_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _2667_ (.A0(_0828_),
    .A1(\po_0.regf_0.rf[0][11] ),
    .S(_1097_),
    .X(_1103_));
 sky130_fd_sc_hd__clkbuf_1 _2668_ (.A(_1103_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _2669_ (.A0(_0840_),
    .A1(\po_0.regf_0.rf[0][12] ),
    .S(_1089_),
    .X(_1104_));
 sky130_fd_sc_hd__clkbuf_1 _2670_ (.A(_1104_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _2671_ (.A0(_0849_),
    .A1(\po_0.regf_0.rf[0][13] ),
    .S(_1089_),
    .X(_1105_));
 sky130_fd_sc_hd__clkbuf_1 _2672_ (.A(_1105_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _2673_ (.A0(_0860_),
    .A1(\po_0.regf_0.rf[0][14] ),
    .S(_1089_),
    .X(_1106_));
 sky130_fd_sc_hd__clkbuf_1 _2674_ (.A(_1106_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _2675_ (.A0(_0870_),
    .A1(\po_0.regf_0.rf[0][15] ),
    .S(_1089_),
    .X(_1107_));
 sky130_fd_sc_hd__clkbuf_1 _2676_ (.A(_1107_),
    .X(_0207_));
 sky130_fd_sc_hd__and4b_4 _2677_ (.A_N(_0875_),
    .B(_0695_),
    .C(_0872_),
    .D(_1030_),
    .X(_1108_));
 sky130_fd_sc_hd__buf_2 _2678_ (.A(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__mux2_1 _2679_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(_0693_),
    .S(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__clkbuf_1 _2680_ (.A(_1110_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _2681_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(_0717_),
    .S(_1109_),
    .X(_1111_));
 sky130_fd_sc_hd__clkbuf_1 _2682_ (.A(_1111_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _2683_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(_0731_),
    .S(_1109_),
    .X(_1112_));
 sky130_fd_sc_hd__clkbuf_1 _2684_ (.A(_1112_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _2685_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(_0741_),
    .S(_1109_),
    .X(_1113_));
 sky130_fd_sc_hd__clkbuf_1 _2686_ (.A(_1113_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _2687_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(_0754_),
    .S(_1109_),
    .X(_1114_));
 sky130_fd_sc_hd__clkbuf_1 _2688_ (.A(_1114_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _2689_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(_0764_),
    .S(_1109_),
    .X(_1115_));
 sky130_fd_sc_hd__clkbuf_1 _2690_ (.A(_1115_),
    .X(_0213_));
 sky130_fd_sc_hd__buf_2 _2691_ (.A(_1108_),
    .X(_1116_));
 sky130_fd_sc_hd__mux2_1 _2692_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(_0776_),
    .S(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__clkbuf_1 _2693_ (.A(_1117_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(\po_0.regf_0.rf[8][7] ),
    .A1(_0787_),
    .S(_1116_),
    .X(_1118_));
 sky130_fd_sc_hd__clkbuf_1 _2695_ (.A(_1118_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _2696_ (.A0(\po_0.regf_0.rf[8][8] ),
    .A1(_0801_),
    .S(_1116_),
    .X(_1119_));
 sky130_fd_sc_hd__clkbuf_1 _2697_ (.A(_1119_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _2698_ (.A0(\po_0.regf_0.rf[8][9] ),
    .A1(_0809_),
    .S(_1116_),
    .X(_1120_));
 sky130_fd_sc_hd__clkbuf_1 _2699_ (.A(_1120_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2700_ (.A0(\po_0.regf_0.rf[8][10] ),
    .A1(_0819_),
    .S(_1116_),
    .X(_1121_));
 sky130_fd_sc_hd__clkbuf_1 _2701_ (.A(_1121_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _2702_ (.A0(\po_0.regf_0.rf[8][11] ),
    .A1(_0827_),
    .S(_1116_),
    .X(_1122_));
 sky130_fd_sc_hd__clkbuf_1 _2703_ (.A(_1122_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _2704_ (.A0(\po_0.regf_0.rf[8][12] ),
    .A1(_0839_),
    .S(_1108_),
    .X(_1123_));
 sky130_fd_sc_hd__clkbuf_1 _2705_ (.A(_1123_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _2706_ (.A0(\po_0.regf_0.rf[8][13] ),
    .A1(_0848_),
    .S(_1108_),
    .X(_1124_));
 sky130_fd_sc_hd__clkbuf_1 _2707_ (.A(_1124_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _2708_ (.A0(\po_0.regf_0.rf[8][14] ),
    .A1(_0859_),
    .S(_1108_),
    .X(_1125_));
 sky130_fd_sc_hd__clkbuf_1 _2709_ (.A(_1125_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _2710_ (.A0(\po_0.regf_0.rf[8][15] ),
    .A1(_0869_),
    .S(_1108_),
    .X(_1126_));
 sky130_fd_sc_hd__clkbuf_1 _2711_ (.A(_1126_),
    .X(_0223_));
 sky130_fd_sc_hd__buf_2 _2712_ (.A(\uc_0._03_ ),
    .X(_1127_));
 sky130_fd_sc_hd__mux2_1 _2713_ (.A0(_0681_),
    .A1(net17),
    .S(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__clkbuf_1 _2714_ (.A(_1128_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _2715_ (.A0(_0714_),
    .A1(net24),
    .S(_1127_),
    .X(_1129_));
 sky130_fd_sc_hd__clkbuf_1 _2716_ (.A(_1129_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _2717_ (.A0(_0729_),
    .A1(net25),
    .S(_1127_),
    .X(_1130_));
 sky130_fd_sc_hd__clkbuf_1 _2718_ (.A(_1130_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _2719_ (.A0(\po_0.muxf_0.rf_w_data[3] ),
    .A1(net26),
    .S(_1127_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_1 _2720_ (.A(_1131_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _2721_ (.A0(_0561_),
    .A1(net27),
    .S(_1127_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _2722_ (.A(_1132_),
    .X(_0228_));
 sky130_fd_sc_hd__buf_4 _2723_ (.A(\uc_0._03_ ),
    .X(_1133_));
 sky130_fd_sc_hd__buf_2 _2724_ (.A(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__mux2_1 _2725_ (.A0(_0565_),
    .A1(net28),
    .S(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_1 _2726_ (.A(_1135_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _2727_ (.A0(_0567_),
    .A1(net29),
    .S(_1134_),
    .X(_1136_));
 sky130_fd_sc_hd__clkbuf_1 _2728_ (.A(_1136_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _2729_ (.A0(_0570_),
    .A1(net30),
    .S(_1134_),
    .X(_1137_));
 sky130_fd_sc_hd__clkbuf_1 _2730_ (.A(_1137_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _2731_ (.A0(\uc_0._20_[8] ),
    .A1(net31),
    .S(_1134_),
    .X(_1138_));
 sky130_fd_sc_hd__clkbuf_1 _2732_ (.A(_1138_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _2733_ (.A0(\uc_0._20_[9] ),
    .A1(net32),
    .S(_1134_),
    .X(_1139_));
 sky130_fd_sc_hd__clkbuf_1 _2734_ (.A(_1139_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _2735_ (.A0(\uc_0._20_[10] ),
    .A1(net18),
    .S(_1134_),
    .X(_1140_));
 sky130_fd_sc_hd__clkbuf_1 _2736_ (.A(_1140_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _2737_ (.A0(\uc_0._20_[11] ),
    .A1(net19),
    .S(_1133_),
    .X(_1141_));
 sky130_fd_sc_hd__clkbuf_1 _2738_ (.A(_1141_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _2739_ (.A0(net79),
    .A1(net20),
    .S(_1133_),
    .X(_1142_));
 sky130_fd_sc_hd__clkbuf_1 _2740_ (.A(_1142_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _2741_ (.A0(net80),
    .A1(net21),
    .S(_1133_),
    .X(_1143_));
 sky130_fd_sc_hd__clkbuf_1 _2742_ (.A(_1143_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _2743_ (.A0(net95),
    .A1(net22),
    .S(_1133_),
    .X(_1144_));
 sky130_fd_sc_hd__clkbuf_1 _2744_ (.A(_1144_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _2745_ (.A0(net82),
    .A1(net23),
    .S(_1133_),
    .X(_1145_));
 sky130_fd_sc_hd__clkbuf_1 _2746_ (.A(_1145_),
    .X(_0239_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2747_ (.A(\uc_0._02_ ),
    .X(_1146_));
 sky130_fd_sc_hd__or2_2 _2748_ (.A(\uc_0._00_ ),
    .B(\uc_0._02_ ),
    .X(_1147_));
 sky130_fd_sc_hd__nor2_1 _2749_ (.A(\uc_0._01_ ),
    .B(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__clkbuf_2 _2750_ (.A(net93),
    .X(_1149_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(_1146_),
    .A1(_1148_),
    .S(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__or2_1 _2752_ (.A(_1149_),
    .B(_0681_),
    .X(_1151_));
 sky130_fd_sc_hd__nand2_1 _2753_ (.A(_1149_),
    .B(_0681_),
    .Y(_1152_));
 sky130_fd_sc_hd__clkbuf_2 _2754_ (.A(\uc_0._01_ ),
    .X(_1153_));
 sky130_fd_sc_hd__nor2_1 _2755_ (.A(\uc_0._00_ ),
    .B(\uc_0._02_ ),
    .Y(_1154_));
 sky130_fd_sc_hd__and4_1 _2756_ (.A(_1151_),
    .B(_1152_),
    .C(_1153_),
    .D(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__or4_1 _2757_ (.A(net74),
    .B(net73),
    .C(net72),
    .D(net71),
    .X(_1156_));
 sky130_fd_sc_hd__or4_1 _2758_ (.A(net63),
    .B(net62),
    .C(net76),
    .D(net75),
    .X(_1157_));
 sky130_fd_sc_hd__or4_1 _2759_ (.A(net67),
    .B(net64),
    .C(_1156_),
    .D(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__clkbuf_2 _2760_ (.A(net69),
    .X(_1159_));
 sky130_fd_sc_hd__nand4_1 _2761_ (.A(net70),
    .B(_1159_),
    .C(net92),
    .D(net93),
    .Y(_1160_));
 sky130_fd_sc_hd__nor4b_1 _2762_ (.A(net66),
    .B(net65),
    .C(_1158_),
    .D_N(_1160_),
    .Y(_1161_));
 sky130_fd_sc_hd__clkbuf_2 _2763_ (.A(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__o21a_1 _2764_ (.A1(_1150_),
    .A2(_1155_),
    .B1(_1162_),
    .X(_0240_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2765_ (.A(net92),
    .X(_1163_));
 sky130_fd_sc_hd__o21ba_1 _2766_ (.A1(\uc_0._01_ ),
    .A2(\uc_0._00_ ),
    .B1_N(_1146_),
    .X(_1164_));
 sky130_fd_sc_hd__and3_1 _2767_ (.A(_1163_),
    .B(_1149_),
    .C(_1146_),
    .X(_1165_));
 sky130_fd_sc_hd__nor2_1 _2768_ (.A(_1163_),
    .B(_1149_),
    .Y(_1166_));
 sky130_fd_sc_hd__or2_1 _2769_ (.A(net92),
    .B(\po_0.muxf_0.rf_w_data[1] ),
    .X(_1167_));
 sky130_fd_sc_hd__nand2_1 _2770_ (.A(net92),
    .B(\po_0.muxf_0.rf_w_data[1] ),
    .Y(_1168_));
 sky130_fd_sc_hd__and4_1 _2771_ (.A(_1167_),
    .B(\po_0.muxf_0.rf_w_data[0] ),
    .C(net93),
    .D(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__a22o_1 _2772_ (.A1(net93),
    .A2(\po_0.muxf_0.rf_w_data[0] ),
    .B1(_1168_),
    .B2(_1167_),
    .X(_1170_));
 sky130_fd_sc_hd__or4b_1 _2773_ (.A(\uc_0._00_ ),
    .B(\uc_0._02_ ),
    .C(_1169_),
    .D_N(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__o31ai_1 _2774_ (.A1(_1164_),
    .A2(_1165_),
    .A3(_1166_),
    .B1(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__o311a_1 _2775_ (.A1(_1163_),
    .A2(_1153_),
    .A3(_1147_),
    .B1(_1172_),
    .C1(_1162_),
    .X(_0241_));
 sky130_fd_sc_hd__a21oi_1 _2776_ (.A1(net92),
    .A2(_0714_),
    .B1(_1169_),
    .Y(_1173_));
 sky130_fd_sc_hd__nor2_1 _2777_ (.A(net69),
    .B(\po_0.muxf_0.rf_w_data[2] ),
    .Y(_1174_));
 sky130_fd_sc_hd__nand2_1 _2778_ (.A(net69),
    .B(_0729_),
    .Y(_1175_));
 sky130_fd_sc_hd__or3b_1 _2779_ (.A(_1173_),
    .B(_1174_),
    .C_N(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__or2_1 _2780_ (.A(_1159_),
    .B(_0729_),
    .X(_1177_));
 sky130_fd_sc_hd__a221o_1 _2781_ (.A1(_1163_),
    .A2(_0714_),
    .B1(_1177_),
    .B2(_1175_),
    .C1(_1169_),
    .X(_1178_));
 sky130_fd_sc_hd__nand3_1 _2782_ (.A(_1159_),
    .B(_1163_),
    .C(net93),
    .Y(_1179_));
 sky130_fd_sc_hd__a21o_1 _2783_ (.A1(net68),
    .A2(net61),
    .B1(_1159_),
    .X(_1180_));
 sky130_fd_sc_hd__a31o_1 _2784_ (.A1(_1146_),
    .A2(_1179_),
    .A3(_1180_),
    .B1(_1148_),
    .X(_1181_));
 sky130_fd_sc_hd__a31o_1 _2785_ (.A1(_1176_),
    .A2(_1178_),
    .A3(_1154_),
    .B1(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__o311a_1 _2786_ (.A1(_1159_),
    .A2(_1153_),
    .A3(_1147_),
    .B1(_1162_),
    .C1(_1182_),
    .X(_0242_));
 sky130_fd_sc_hd__a31o_1 _2787_ (.A1(_1159_),
    .A2(_1163_),
    .A3(_1149_),
    .B1(net70),
    .X(_1183_));
 sky130_fd_sc_hd__or2_1 _2788_ (.A(net70),
    .B(\po_0.muxf_0.rf_w_data[3] ),
    .X(_1184_));
 sky130_fd_sc_hd__nand2_1 _2789_ (.A(net70),
    .B(\po_0.muxf_0.rf_w_data[3] ),
    .Y(_1185_));
 sky130_fd_sc_hd__o21ai_1 _2790_ (.A1(_1173_),
    .A2(_1174_),
    .B1(_1175_),
    .Y(_1186_));
 sky130_fd_sc_hd__a21oi_1 _2791_ (.A1(_1184_),
    .A2(_1185_),
    .B1(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__a31o_1 _2792_ (.A1(_1186_),
    .A2(_1185_),
    .A3(_1184_),
    .B1(_1147_),
    .X(_1188_));
 sky130_fd_sc_hd__nor2_1 _2793_ (.A(_1187_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__a311o_1 _2794_ (.A1(_1146_),
    .A2(_1160_),
    .A3(_1183_),
    .B1(_1189_),
    .C1(_1148_),
    .X(_1190_));
 sky130_fd_sc_hd__o311a_1 _2795_ (.A1(net70),
    .A2(_1153_),
    .A3(_1147_),
    .B1(_1162_),
    .C1(_1190_),
    .X(_0243_));
 sky130_fd_sc_hd__and2_1 _2796_ (.A(net71),
    .B(\po_0.muxf_0.rf_w_data[4] ),
    .X(_1191_));
 sky130_fd_sc_hd__nor2_1 _2797_ (.A(net71),
    .B(\po_0.muxf_0.rf_w_data[4] ),
    .Y(_1192_));
 sky130_fd_sc_hd__a21boi_1 _2798_ (.A1(_1186_),
    .A2(_1184_),
    .B1_N(_1185_),
    .Y(_1193_));
 sky130_fd_sc_hd__o21ai_1 _2799_ (.A1(_1191_),
    .A2(_1192_),
    .B1(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__and3_1 _2800_ (.A(\uc_0._01_ ),
    .B(_1154_),
    .C(_1162_),
    .X(_1195_));
 sky130_fd_sc_hd__o311a_1 _2801_ (.A1(_1191_),
    .A2(_1192_),
    .A3(_1193_),
    .B1(_1194_),
    .C1(_1195_),
    .X(_0244_));
 sky130_fd_sc_hd__nand2_1 _2802_ (.A(net72),
    .B(_0565_),
    .Y(_1196_));
 sky130_fd_sc_hd__or2_1 _2803_ (.A(net72),
    .B(\po_0.muxf_0.rf_w_data[5] ),
    .X(_1197_));
 sky130_fd_sc_hd__or2_1 _2804_ (.A(_1191_),
    .B(_1192_),
    .X(_1198_));
 sky130_fd_sc_hd__nor2_1 _2805_ (.A(_1198_),
    .B(_1193_),
    .Y(_1199_));
 sky130_fd_sc_hd__a221o_1 _2806_ (.A1(net71),
    .A2(_0561_),
    .B1(_1196_),
    .B2(_1197_),
    .C1(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__o211ai_2 _2807_ (.A1(_1191_),
    .A2(_1199_),
    .B1(_1196_),
    .C1(_1197_),
    .Y(_1201_));
 sky130_fd_sc_hd__and3_1 _2808_ (.A(_1200_),
    .B(_1195_),
    .C(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__clkbuf_1 _2809_ (.A(_1202_),
    .X(_0245_));
 sky130_fd_sc_hd__and2_1 _2810_ (.A(net73),
    .B(\po_0.muxf_0.rf_w_data[6] ),
    .X(_1203_));
 sky130_fd_sc_hd__nor2_1 _2811_ (.A(net73),
    .B(\po_0.muxf_0.rf_w_data[6] ),
    .Y(_1204_));
 sky130_fd_sc_hd__or2_1 _2812_ (.A(_1203_),
    .B(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__a21oi_1 _2813_ (.A1(_1196_),
    .A2(_1201_),
    .B1(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__or4bb_1 _2814_ (.A(\uc_0._00_ ),
    .B(\uc_0._02_ ),
    .C_N(_1161_),
    .D_N(\uc_0._01_ ),
    .X(_1207_));
 sky130_fd_sc_hd__a31o_1 _2815_ (.A1(_1196_),
    .A2(_1201_),
    .A3(_1205_),
    .B1(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__nor2_1 _2816_ (.A(_1206_),
    .B(_1208_),
    .Y(_0246_));
 sky130_fd_sc_hd__nand2_1 _2817_ (.A(net74),
    .B(_0570_),
    .Y(_1209_));
 sky130_fd_sc_hd__or2_1 _2818_ (.A(net74),
    .B(\po_0.muxf_0.rf_w_data[7] ),
    .X(_1210_));
 sky130_fd_sc_hd__o211a_1 _2819_ (.A1(_1203_),
    .A2(_1206_),
    .B1(_1209_),
    .C1(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__a221o_1 _2820_ (.A1(net73),
    .A2(_0567_),
    .B1(_1209_),
    .B2(_1210_),
    .C1(_1206_),
    .X(_1212_));
 sky130_fd_sc_hd__and3b_1 _2821_ (.A_N(_1211_),
    .B(_1212_),
    .C(_1195_),
    .X(_1213_));
 sky130_fd_sc_hd__clkbuf_1 _2822_ (.A(_1213_),
    .X(_0247_));
 sky130_fd_sc_hd__a21o_1 _2823_ (.A1(net74),
    .A2(_0570_),
    .B1(net75),
    .X(_1214_));
 sky130_fd_sc_hd__o2111a_1 _2824_ (.A1(_1214_),
    .A2(_1211_),
    .B1(_1154_),
    .C1(_1153_),
    .D1(_1162_),
    .X(_0248_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2825_ (.A(_1357_),
    .X(_1215_));
 sky130_fd_sc_hd__o211a_1 _2826_ (.A1(_1215_),
    .A2(_1366_),
    .B1(_1368_),
    .C1(_1356_),
    .X(_1216_));
 sky130_fd_sc_hd__o2111a_1 _2827_ (.A1(_1215_),
    .A2(_1366_),
    .B1(\uc_0.bc_0._54_[1] ),
    .C1(_1361_),
    .D1(_1356_),
    .X(_1217_));
 sky130_fd_sc_hd__nor2_1 _2828_ (.A(_1216_),
    .B(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__buf_2 _2829_ (.A(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__o21a_1 _2830_ (.A1(_1215_),
    .A2(\uc_0._00_ ),
    .B1(_1219_),
    .X(_0256_));
 sky130_fd_sc_hd__and4b_4 _2831_ (.A_N(_0695_),
    .B(_0873_),
    .C(_1030_),
    .D(_0875_),
    .X(_1220_));
 sky130_fd_sc_hd__clkbuf_4 _2832_ (.A(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__mux2_1 _2833_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(_0693_),
    .S(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__clkbuf_1 _2834_ (.A(_1222_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _2835_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(_0717_),
    .S(_1221_),
    .X(_1223_));
 sky130_fd_sc_hd__clkbuf_1 _2836_ (.A(_1223_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _2837_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(_0731_),
    .S(_1221_),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_1 _2838_ (.A(_1224_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _2839_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(_0741_),
    .S(_1221_),
    .X(_1225_));
 sky130_fd_sc_hd__clkbuf_1 _2840_ (.A(_1225_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _2841_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(_0754_),
    .S(_1221_),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_1 _2842_ (.A(_1226_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _2843_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(_0764_),
    .S(_1221_),
    .X(_1227_));
 sky130_fd_sc_hd__clkbuf_1 _2844_ (.A(_1227_),
    .X(_0262_));
 sky130_fd_sc_hd__buf_2 _2845_ (.A(_1220_),
    .X(_1228_));
 sky130_fd_sc_hd__mux2_1 _2846_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(_0776_),
    .S(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _2847_ (.A(_1229_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _2848_ (.A0(\po_0.regf_0.rf[4][7] ),
    .A1(_0787_),
    .S(_1228_),
    .X(_1230_));
 sky130_fd_sc_hd__clkbuf_1 _2849_ (.A(_1230_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _2850_ (.A0(\po_0.regf_0.rf[4][8] ),
    .A1(_0801_),
    .S(_1228_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _2851_ (.A(_1231_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _2852_ (.A0(\po_0.regf_0.rf[4][9] ),
    .A1(_0809_),
    .S(_1228_),
    .X(_1232_));
 sky130_fd_sc_hd__clkbuf_1 _2853_ (.A(_1232_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _2854_ (.A0(\po_0.regf_0.rf[4][10] ),
    .A1(_0819_),
    .S(_1228_),
    .X(_1233_));
 sky130_fd_sc_hd__clkbuf_1 _2855_ (.A(_1233_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _2856_ (.A0(\po_0.regf_0.rf[4][11] ),
    .A1(_0827_),
    .S(_1228_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _2857_ (.A(_1234_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _2858_ (.A0(\po_0.regf_0.rf[4][12] ),
    .A1(_0839_),
    .S(_1220_),
    .X(_1235_));
 sky130_fd_sc_hd__clkbuf_1 _2859_ (.A(_1235_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _2860_ (.A0(\po_0.regf_0.rf[4][13] ),
    .A1(_0848_),
    .S(_1220_),
    .X(_1236_));
 sky130_fd_sc_hd__clkbuf_1 _2861_ (.A(_1236_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _2862_ (.A0(\po_0.regf_0.rf[4][14] ),
    .A1(_0859_),
    .S(_1220_),
    .X(_1237_));
 sky130_fd_sc_hd__clkbuf_1 _2863_ (.A(_1237_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _2864_ (.A0(\po_0.regf_0.rf[4][15] ),
    .A1(_0869_),
    .S(_1220_),
    .X(_1238_));
 sky130_fd_sc_hd__clkbuf_1 _2865_ (.A(_1238_),
    .X(_0272_));
 sky130_fd_sc_hd__and4_4 _2866_ (.A(_0696_),
    .B(_0697_),
    .C(_0873_),
    .D(_0936_),
    .X(_1239_));
 sky130_fd_sc_hd__clkbuf_4 _2867_ (.A(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(\po_0.regf_0.rf[3][0] ),
    .A1(_0693_),
    .S(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__clkbuf_1 _2869_ (.A(_1241_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _2870_ (.A0(\po_0.regf_0.rf[3][1] ),
    .A1(_0717_),
    .S(_1240_),
    .X(_1242_));
 sky130_fd_sc_hd__clkbuf_1 _2871_ (.A(_1242_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _2872_ (.A0(\po_0.regf_0.rf[3][2] ),
    .A1(_0731_),
    .S(_1240_),
    .X(_1243_));
 sky130_fd_sc_hd__clkbuf_1 _2873_ (.A(_1243_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(\po_0.regf_0.rf[3][3] ),
    .A1(_0741_),
    .S(_1240_),
    .X(_1244_));
 sky130_fd_sc_hd__clkbuf_1 _2875_ (.A(_1244_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(\po_0.regf_0.rf[3][4] ),
    .A1(_0754_),
    .S(_1240_),
    .X(_1245_));
 sky130_fd_sc_hd__clkbuf_1 _2877_ (.A(_1245_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _2878_ (.A0(\po_0.regf_0.rf[3][5] ),
    .A1(_0764_),
    .S(_1240_),
    .X(_1246_));
 sky130_fd_sc_hd__clkbuf_1 _2879_ (.A(_1246_),
    .X(_0278_));
 sky130_fd_sc_hd__buf_2 _2880_ (.A(_1239_),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _2881_ (.A0(\po_0.regf_0.rf[3][6] ),
    .A1(_0776_),
    .S(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__clkbuf_1 _2882_ (.A(_1248_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _2883_ (.A0(\po_0.regf_0.rf[3][7] ),
    .A1(_0787_),
    .S(_1247_),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_1 _2884_ (.A(_1249_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _2885_ (.A0(\po_0.regf_0.rf[3][8] ),
    .A1(_0801_),
    .S(_1247_),
    .X(_1250_));
 sky130_fd_sc_hd__clkbuf_1 _2886_ (.A(_1250_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _2887_ (.A0(\po_0.regf_0.rf[3][9] ),
    .A1(_0809_),
    .S(_1247_),
    .X(_1251_));
 sky130_fd_sc_hd__clkbuf_1 _2888_ (.A(_1251_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _2889_ (.A0(\po_0.regf_0.rf[3][10] ),
    .A1(_0819_),
    .S(_1247_),
    .X(_1252_));
 sky130_fd_sc_hd__clkbuf_1 _2890_ (.A(_1252_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _2891_ (.A0(\po_0.regf_0.rf[3][11] ),
    .A1(_0827_),
    .S(_1247_),
    .X(_1253_));
 sky130_fd_sc_hd__clkbuf_1 _2892_ (.A(_1253_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _2893_ (.A0(\po_0.regf_0.rf[3][12] ),
    .A1(_0839_),
    .S(_1239_),
    .X(_1254_));
 sky130_fd_sc_hd__clkbuf_1 _2894_ (.A(_1254_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _2895_ (.A0(\po_0.regf_0.rf[3][13] ),
    .A1(_0848_),
    .S(_1239_),
    .X(_1255_));
 sky130_fd_sc_hd__clkbuf_1 _2896_ (.A(_1255_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _2897_ (.A0(\po_0.regf_0.rf[3][14] ),
    .A1(_0859_),
    .S(_1239_),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_1 _2898_ (.A(_1256_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _2899_ (.A0(\po_0.regf_0.rf[3][15] ),
    .A1(_0869_),
    .S(_1239_),
    .X(_1257_));
 sky130_fd_sc_hd__clkbuf_1 _2900_ (.A(_1257_),
    .X(_0288_));
 sky130_fd_sc_hd__and3_4 _2901_ (.A(_0935_),
    .B(_0895_),
    .C(_0936_),
    .X(_1258_));
 sky130_fd_sc_hd__clkbuf_4 _2902_ (.A(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__mux2_1 _2903_ (.A0(\po_0.regf_0.rf[2][0] ),
    .A1(_0693_),
    .S(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__clkbuf_1 _2904_ (.A(_1260_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _2905_ (.A0(\po_0.regf_0.rf[2][1] ),
    .A1(_0717_),
    .S(_1259_),
    .X(_1261_));
 sky130_fd_sc_hd__clkbuf_1 _2906_ (.A(_1261_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _2907_ (.A0(\po_0.regf_0.rf[2][2] ),
    .A1(_0731_),
    .S(_1259_),
    .X(_1262_));
 sky130_fd_sc_hd__clkbuf_1 _2908_ (.A(_1262_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _2909_ (.A0(\po_0.regf_0.rf[2][3] ),
    .A1(_0741_),
    .S(_1259_),
    .X(_1263_));
 sky130_fd_sc_hd__clkbuf_1 _2910_ (.A(_1263_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _2911_ (.A0(\po_0.regf_0.rf[2][4] ),
    .A1(_0754_),
    .S(_1259_),
    .X(_1264_));
 sky130_fd_sc_hd__clkbuf_1 _2912_ (.A(_1264_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _2913_ (.A0(\po_0.regf_0.rf[2][5] ),
    .A1(_0764_),
    .S(_1259_),
    .X(_1265_));
 sky130_fd_sc_hd__clkbuf_1 _2914_ (.A(_1265_),
    .X(_0294_));
 sky130_fd_sc_hd__buf_2 _2915_ (.A(_1258_),
    .X(_1266_));
 sky130_fd_sc_hd__mux2_1 _2916_ (.A0(\po_0.regf_0.rf[2][6] ),
    .A1(_0776_),
    .S(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__clkbuf_1 _2917_ (.A(_1267_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _2918_ (.A0(\po_0.regf_0.rf[2][7] ),
    .A1(_0787_),
    .S(_1266_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_1 _2919_ (.A(_1268_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _2920_ (.A0(\po_0.regf_0.rf[2][8] ),
    .A1(_0801_),
    .S(_1266_),
    .X(_1269_));
 sky130_fd_sc_hd__clkbuf_1 _2921_ (.A(_1269_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _2922_ (.A0(\po_0.regf_0.rf[2][9] ),
    .A1(_0809_),
    .S(_1266_),
    .X(_1270_));
 sky130_fd_sc_hd__clkbuf_1 _2923_ (.A(_1270_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _2924_ (.A0(\po_0.regf_0.rf[2][10] ),
    .A1(_0819_),
    .S(_1266_),
    .X(_1271_));
 sky130_fd_sc_hd__clkbuf_1 _2925_ (.A(_1271_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _2926_ (.A0(\po_0.regf_0.rf[2][11] ),
    .A1(_0827_),
    .S(_1266_),
    .X(_1272_));
 sky130_fd_sc_hd__clkbuf_1 _2927_ (.A(_1272_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _2928_ (.A0(\po_0.regf_0.rf[2][12] ),
    .A1(_0839_),
    .S(_1258_),
    .X(_1273_));
 sky130_fd_sc_hd__clkbuf_1 _2929_ (.A(_1273_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _2930_ (.A0(\po_0.regf_0.rf[2][13] ),
    .A1(_0848_),
    .S(_1258_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _2931_ (.A(_1274_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _2932_ (.A0(\po_0.regf_0.rf[2][14] ),
    .A1(_0859_),
    .S(_1258_),
    .X(_1275_));
 sky130_fd_sc_hd__clkbuf_1 _2933_ (.A(_1275_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _2934_ (.A0(\po_0.regf_0.rf[2][15] ),
    .A1(_0869_),
    .S(_1258_),
    .X(_1276_));
 sky130_fd_sc_hd__clkbuf_1 _2935_ (.A(_1276_),
    .X(_0304_));
 sky130_fd_sc_hd__or4_1 _2936_ (.A(_1215_),
    .B(_1359_),
    .C(_1365_),
    .D(_1366_),
    .X(_1277_));
 sky130_fd_sc_hd__a21o_1 _2937_ (.A1(_1277_),
    .A2(_1319_),
    .B1(_1370_),
    .X(_0305_));
 sky130_fd_sc_hd__o21ba_1 _2938_ (.A1(_1315_),
    .A2(_0563_),
    .B1_N(_1370_),
    .X(_0306_));
 sky130_fd_sc_hd__a21o_1 _2939_ (.A1(net91),
    .A2(_1219_),
    .B1(_0563_),
    .X(_0307_));
 sky130_fd_sc_hd__a221o_1 _2940_ (.A1(_1367_),
    .A2(_1368_),
    .B1(_1218_),
    .B2(\po_0.regf_0.rp_rd ),
    .C1(_0563_),
    .X(_0308_));
 sky130_fd_sc_hd__o211a_1 _2941_ (.A1(_1354_),
    .A2(_1363_),
    .B1(_1369_),
    .C1(\uc_0.bc_0._54_[0] ),
    .X(_1278_));
 sky130_fd_sc_hd__and3_1 _2942_ (.A(_1361_),
    .B(_1365_),
    .C(\uc_0.bc_0._54_[2] ),
    .X(_1279_));
 sky130_fd_sc_hd__or3_4 _2943_ (.A(_1278_),
    .B(_1279_),
    .C(_1371_),
    .X(_1280_));
 sky130_fd_sc_hd__a21o_1 _2944_ (.A1(_0935_),
    .A2(_1219_),
    .B1(_1280_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _2945_ (.A0(\po_0.regf_0.rq_addr[0] ),
    .A1(_0561_),
    .S(_0568_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_1 _2946_ (.A(_1281_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _2947_ (.A0(\po_0.regf_0.rq_addr[1] ),
    .A1(_0565_),
    .S(_0568_),
    .X(_1282_));
 sky130_fd_sc_hd__clkbuf_1 _2948_ (.A(_1282_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _2949_ (.A0(\po_0.regf_0.rq_addr[2] ),
    .A1(_0567_),
    .S(_0568_),
    .X(_1283_));
 sky130_fd_sc_hd__clkbuf_1 _2950_ (.A(_1283_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2951_ (.A0(\po_0.regf_0.rq_addr[3] ),
    .A1(_0570_),
    .S(_0568_),
    .X(_1284_));
 sky130_fd_sc_hd__clkbuf_1 _2952_ (.A(_1284_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2953_ (.A0(\uc_0._20_[8] ),
    .A1(\po_0.regf_0.rp_addr[0] ),
    .S(_1373_),
    .X(_1285_));
 sky130_fd_sc_hd__clkbuf_1 _2954_ (.A(_1285_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _2955_ (.A0(\uc_0._20_[9] ),
    .A1(\po_0.regf_0.rp_addr[1] ),
    .S(_1373_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_1 _2956_ (.A(_1286_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _2957_ (.A0(\uc_0._20_[10] ),
    .A1(\po_0.regf_0.rp_addr[2] ),
    .S(_1372_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_1 _2958_ (.A(_1287_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _2959_ (.A0(\uc_0._20_[11] ),
    .A1(\po_0.regf_0.rp_addr[3] ),
    .S(_1372_),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_1 _2960_ (.A(_1288_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _2961_ (.A0(\uc_0._20_[8] ),
    .A1(_0681_),
    .S(_0562_),
    .X(_1289_));
 sky130_fd_sc_hd__mux2_1 _2962_ (.A0(_0697_),
    .A1(_1289_),
    .S(_1280_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _2963_ (.A(_1290_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _2964_ (.A0(\uc_0._20_[9] ),
    .A1(_0714_),
    .S(_0562_),
    .X(_1291_));
 sky130_fd_sc_hd__mux2_1 _2965_ (.A0(_0696_),
    .A1(_1291_),
    .S(_1280_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _2966_ (.A(_1292_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(\uc_0._20_[10] ),
    .A1(_0729_),
    .S(_0562_),
    .X(_1293_));
 sky130_fd_sc_hd__mux2_1 _2968_ (.A0(_0699_),
    .A1(_1293_),
    .S(_1280_),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _2969_ (.A(_1294_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _2970_ (.A0(\uc_0._20_[11] ),
    .A1(\po_0.muxf_0.rf_w_data[3] ),
    .S(_0562_),
    .X(_1295_));
 sky130_fd_sc_hd__mux2_1 _2971_ (.A0(_0915_),
    .A1(_1295_),
    .S(_1280_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _2972_ (.A(_1296_),
    .X(_0321_));
 sky130_fd_sc_hd__a21oi_1 _2973_ (.A1(\uc_0.bc_0._54_[1] ),
    .A2(_1369_),
    .B1(_1370_),
    .Y(_1297_));
 sky130_fd_sc_hd__o21a_1 _2974_ (.A1(\po_0.muxf_0.s0 ),
    .A2(_1279_),
    .B1(_1297_),
    .X(_0322_));
 sky130_fd_sc_hd__nor2_1 _2975_ (.A(_1279_),
    .B(_0563_),
    .Y(_1298_));
 sky130_fd_sc_hd__o21a_1 _2976_ (.A1(\po_0.muxf_0.s1 ),
    .A2(_1278_),
    .B1(_1298_),
    .X(_0323_));
 sky130_fd_sc_hd__a32o_1 _2977_ (.A1(\uc_0.bc_0._54_[0] ),
    .A2(_1365_),
    .A3(_1369_),
    .B1(_1219_),
    .B2(net60),
    .X(_0324_));
 sky130_fd_sc_hd__or3_1 _2978_ (.A(_1357_),
    .B(_1363_),
    .C(_1366_),
    .X(_1299_));
 sky130_fd_sc_hd__clkbuf_4 _2979_ (.A(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__a2bb2o_1 _2980_ (.A1_N(_1300_),
    .A2_N(\uc_0.bc_0._54_[0] ),
    .B1(net59),
    .B2(_1219_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _2981_ (.A0(_0681_),
    .A1(net51),
    .S(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_1 _2982_ (.A(_1301_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _2983_ (.A0(_0714_),
    .A1(net52),
    .S(_1300_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _2984_ (.A(_1302_),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_8 _2985_ (.A(_1299_),
    .X(_1303_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(_0729_),
    .A1(net53),
    .S(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_1 _2987_ (.A(_1304_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(\po_0.muxf_0.rf_w_data[3] ),
    .A1(net54),
    .S(_1303_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_1 _2989_ (.A(_1305_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _2990_ (.A0(_0561_),
    .A1(net55),
    .S(_1303_),
    .X(_1306_));
 sky130_fd_sc_hd__clkbuf_1 _2991_ (.A(_1306_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _2992_ (.A0(_0565_),
    .A1(net56),
    .S(_1303_),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_1 _2993_ (.A(_1307_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _2994_ (.A0(_0567_),
    .A1(net57),
    .S(_1303_),
    .X(_1308_));
 sky130_fd_sc_hd__clkbuf_1 _2995_ (.A(_1308_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _2996_ (.A0(_0570_),
    .A1(net58),
    .S(_1303_),
    .X(_1309_));
 sky130_fd_sc_hd__clkbuf_1 _2997_ (.A(_1309_),
    .X(_0333_));
 sky130_fd_sc_hd__or4_1 _2998_ (.A(_1215_),
    .B(_1361_),
    .C(_1365_),
    .D(_1367_),
    .X(_1310_));
 sky130_fd_sc_hd__o311a_1 _2999_ (.A1(net77),
    .A2(_1216_),
    .A3(_1217_),
    .B1(_1300_),
    .C1(_1310_),
    .X(_0334_));
 sky130_fd_sc_hd__o211a_1 _3000_ (.A1(_1127_),
    .A2(_1217_),
    .B1(_1300_),
    .C1(_1310_),
    .X(_0335_));
 sky130_fd_sc_hd__inv_2 _3001_ (.A(\uc_0.bc_0._54_[1] ),
    .Y(_1311_));
 sky130_fd_sc_hd__o221a_1 _3002_ (.A1(_1311_),
    .A2(_1367_),
    .B1(_1216_),
    .B2(_1146_),
    .C1(_1300_),
    .X(_0336_));
 sky130_fd_sc_hd__or3_1 _3003_ (.A(_1215_),
    .B(_1359_),
    .C(_1365_),
    .X(_1312_));
 sky130_fd_sc_hd__a2bb2o_1 _3004_ (.A1_N(_1312_),
    .A2_N(_1355_),
    .B1(_1153_),
    .B2(_1219_),
    .X(_0337_));
 sky130_fd_sc_hd__dfxtp_1 _3005_ (.CLK(net169),
    .D(_0016_),
    .Q(\po_0.regf_0.rf[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3006_ (.CLK(net143),
    .D(_0017_),
    .Q(\po_0.regf_0.rf[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3007_ (.CLK(net147),
    .D(_0018_),
    .Q(\po_0.regf_0.rf[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3008_ (.CLK(net161),
    .D(_0019_),
    .Q(\po_0.regf_0.rf[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3009_ (.CLK(net165),
    .D(_0020_),
    .Q(\po_0.regf_0.rf[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3010_ (.CLK(net163),
    .D(_0021_),
    .Q(\po_0.regf_0.rf[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3011_ (.CLK(net132),
    .D(_0022_),
    .Q(\po_0.regf_0.rf[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3012_ (.CLK(net133),
    .D(_0023_),
    .Q(\po_0.regf_0.rf[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3013_ (.CLK(net129),
    .D(_0024_),
    .Q(\po_0.regf_0.rf[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3014_ (.CLK(net126),
    .D(_0025_),
    .Q(\po_0.regf_0.rf[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3015_ (.CLK(net133),
    .D(_0026_),
    .Q(\po_0.regf_0.rf[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3016_ (.CLK(net121),
    .D(_0027_),
    .Q(\po_0.regf_0.rf[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3017_ (.CLK(net124),
    .D(_0028_),
    .Q(\po_0.regf_0.rf[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3018_ (.CLK(net124),
    .D(_0029_),
    .Q(\po_0.regf_0.rf[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3019_ (.CLK(net118),
    .D(_0030_),
    .Q(\po_0.regf_0.rf[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3020_ (.CLK(net118),
    .D(_0031_),
    .Q(\po_0.regf_0.rf[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3021_ (.CLK(net169),
    .D(_0032_),
    .Q(\po_0.regf_0.rf[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3022_ (.CLK(net143),
    .D(_0033_),
    .Q(\po_0.regf_0.rf[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3023_ (.CLK(net150),
    .D(_0034_),
    .Q(\po_0.regf_0.rf[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3024_ (.CLK(net161),
    .D(_0035_),
    .Q(\po_0.regf_0.rf[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3025_ (.CLK(net169),
    .D(_0036_),
    .Q(\po_0.regf_0.rf[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3026_ (.CLK(net163),
    .D(_0037_),
    .Q(\po_0.regf_0.rf[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3027_ (.CLK(net132),
    .D(_0038_),
    .Q(\po_0.regf_0.rf[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3028_ (.CLK(net134),
    .D(_0039_),
    .Q(\po_0.regf_0.rf[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3029_ (.CLK(net130),
    .D(_0040_),
    .Q(\po_0.regf_0.rf[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3030_ (.CLK(net126),
    .D(_0041_),
    .Q(\po_0.regf_0.rf[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3031_ (.CLK(net134),
    .D(_0042_),
    .Q(\po_0.regf_0.rf[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3032_ (.CLK(net121),
    .D(_0043_),
    .Q(\po_0.regf_0.rf[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3033_ (.CLK(net124),
    .D(_0044_),
    .Q(\po_0.regf_0.rf[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3034_ (.CLK(net125),
    .D(_0045_),
    .Q(\po_0.regf_0.rf[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3035_ (.CLK(net118),
    .D(_0046_),
    .Q(\po_0.regf_0.rf[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3036_ (.CLK(net119),
    .D(_0047_),
    .Q(\po_0.regf_0.rf[5][15] ));
 sky130_fd_sc_hd__dlxtp_1 _3037_ (.D(\po_0.regf_0._5_[0] ),
    .GATE(net90),
    .Q(\po_0._1_[0] ));
 sky130_fd_sc_hd__dlxtp_1 _3038_ (.D(\po_0.regf_0._5_[1] ),
    .GATE(net91),
    .Q(\po_0._1_[1] ));
 sky130_fd_sc_hd__dlxtp_1 _3039_ (.D(\po_0.regf_0._5_[2] ),
    .GATE(net90),
    .Q(\po_0._1_[2] ));
 sky130_fd_sc_hd__dlxtp_1 _3040_ (.D(\po_0.regf_0._5_[3] ),
    .GATE(net90),
    .Q(\po_0._1_[3] ));
 sky130_fd_sc_hd__dlxtp_1 _3041_ (.D(\po_0.regf_0._5_[4] ),
    .GATE(net90),
    .Q(\po_0._1_[4] ));
 sky130_fd_sc_hd__dlxtp_1 _3042_ (.D(\po_0.regf_0._5_[5] ),
    .GATE(net90),
    .Q(\po_0._1_[5] ));
 sky130_fd_sc_hd__dlxtp_1 _3043_ (.D(\po_0.regf_0._5_[6] ),
    .GATE(net89),
    .Q(\po_0._1_[6] ));
 sky130_fd_sc_hd__dlxtp_1 _3044_ (.D(\po_0.regf_0._5_[7] ),
    .GATE(net90),
    .Q(\po_0._1_[7] ));
 sky130_fd_sc_hd__dlxtp_1 _3045_ (.D(\po_0.regf_0._5_[8] ),
    .GATE(net88),
    .Q(\po_0._1_[8] ));
 sky130_fd_sc_hd__dlxtp_1 _3046_ (.D(\po_0.regf_0._5_[9] ),
    .GATE(net89),
    .Q(\po_0._1_[9] ));
 sky130_fd_sc_hd__dlxtp_1 _3047_ (.D(\po_0.regf_0._5_[10] ),
    .GATE(net89),
    .Q(\po_0._1_[10] ));
 sky130_fd_sc_hd__dlxtp_1 _3048_ (.D(\po_0.regf_0._5_[11] ),
    .GATE(net88),
    .Q(\po_0._1_[11] ));
 sky130_fd_sc_hd__dlxtp_1 _3049_ (.D(\po_0.regf_0._5_[12] ),
    .GATE(net88),
    .Q(\po_0._1_[12] ));
 sky130_fd_sc_hd__dlxtp_1 _3050_ (.D(\po_0.regf_0._5_[13] ),
    .GATE(net88),
    .Q(\po_0._1_[13] ));
 sky130_fd_sc_hd__dlxtp_1 _3051_ (.D(\po_0.regf_0._5_[14] ),
    .GATE(net88),
    .Q(\po_0._1_[14] ));
 sky130_fd_sc_hd__dlxtp_1 _3052_ (.D(\po_0.regf_0._5_[15] ),
    .GATE(net88),
    .Q(\po_0._1_[15] ));
 sky130_fd_sc_hd__dlxtp_1 _3053_ (.D(\po_0.regf_0._3_[0] ),
    .GATE(\po_0.regf_0.rp_rd ),
    .Q(net35));
 sky130_fd_sc_hd__dlxtp_1 _3054_ (.D(\po_0.regf_0._3_[1] ),
    .GATE(net87),
    .Q(net42));
 sky130_fd_sc_hd__dlxtp_1 _3055_ (.D(\po_0.regf_0._3_[2] ),
    .GATE(net87),
    .Q(net43));
 sky130_fd_sc_hd__dlxtp_1 _3056_ (.D(\po_0.regf_0._3_[3] ),
    .GATE(net87),
    .Q(net44));
 sky130_fd_sc_hd__dlxtp_1 _3057_ (.D(\po_0.regf_0._3_[4] ),
    .GATE(net87),
    .Q(net45));
 sky130_fd_sc_hd__dlxtp_1 _3058_ (.D(\po_0.regf_0._3_[5] ),
    .GATE(net85),
    .Q(net46));
 sky130_fd_sc_hd__dlxtp_1 _3059_ (.D(\po_0.regf_0._3_[6] ),
    .GATE(net86),
    .Q(net47));
 sky130_fd_sc_hd__dlxtp_1 _3060_ (.D(\po_0.regf_0._3_[7] ),
    .GATE(net85),
    .Q(net48));
 sky130_fd_sc_hd__dlxtp_1 _3061_ (.D(\po_0.regf_0._3_[8] ),
    .GATE(net85),
    .Q(net49));
 sky130_fd_sc_hd__dlxtp_1 _3062_ (.D(\po_0.regf_0._3_[9] ),
    .GATE(net85),
    .Q(net50));
 sky130_fd_sc_hd__dlxtp_1 _3063_ (.D(\po_0.regf_0._3_[10] ),
    .GATE(net86),
    .Q(net36));
 sky130_fd_sc_hd__dlxtp_1 _3064_ (.D(\po_0.regf_0._3_[11] ),
    .GATE(net86),
    .Q(net37));
 sky130_fd_sc_hd__dlxtp_1 _3065_ (.D(\po_0.regf_0._3_[12] ),
    .GATE(net85),
    .Q(net38));
 sky130_fd_sc_hd__dlxtp_1 _3066_ (.D(\po_0.regf_0._3_[13] ),
    .GATE(net86),
    .Q(net39));
 sky130_fd_sc_hd__dlxtp_1 _3067_ (.D(\po_0.regf_0._3_[14] ),
    .GATE(net86),
    .Q(net40));
 sky130_fd_sc_hd__dlxtp_1 _3068_ (.D(\po_0.regf_0._3_[15] ),
    .GATE(net85),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _3069_ (.CLK(net169),
    .D(_0048_),
    .Q(\po_0.regf_0.rf[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3070_ (.CLK(net143),
    .D(_0049_),
    .Q(\po_0.regf_0.rf[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3071_ (.CLK(net148),
    .D(_0050_),
    .Q(\po_0.regf_0.rf[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3072_ (.CLK(net161),
    .D(_0051_),
    .Q(\po_0.regf_0.rf[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3073_ (.CLK(net159),
    .D(_0052_),
    .Q(\po_0.regf_0.rf[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3074_ (.CLK(net163),
    .D(_0053_),
    .Q(\po_0.regf_0.rf[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3075_ (.CLK(net132),
    .D(_0054_),
    .Q(\po_0.regf_0.rf[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3076_ (.CLK(net133),
    .D(_0055_),
    .Q(\po_0.regf_0.rf[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3077_ (.CLK(net129),
    .D(_0056_),
    .Q(\po_0.regf_0.rf[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3078_ (.CLK(net126),
    .D(_0057_),
    .Q(\po_0.regf_0.rf[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3079_ (.CLK(net133),
    .D(_0058_),
    .Q(\po_0.regf_0.rf[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3080_ (.CLK(net121),
    .D(_0059_),
    .Q(\po_0.regf_0.rf[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3081_ (.CLK(net124),
    .D(_0060_),
    .Q(\po_0.regf_0.rf[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3082_ (.CLK(net124),
    .D(_0061_),
    .Q(\po_0.regf_0.rf[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3083_ (.CLK(net100),
    .D(_0062_),
    .Q(\po_0.regf_0.rf[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3084_ (.CLK(net118),
    .D(_0063_),
    .Q(\po_0.regf_0.rf[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3085_ (.CLK(net109),
    .D(_0008_),
    .Q(_0000_));
 sky130_fd_sc_hd__dfxtp_1 _3086_ (.CLK(net109),
    .D(_0009_),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_1 _3087_ (.CLK(net109),
    .D(_0010_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_2 _3088_ (.CLK(net138),
    .D(_0011_),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_1 _3089_ (.CLK(net164),
    .D(_0064_),
    .Q(\po_0.regf_0.rf[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3090_ (.CLK(net143),
    .D(_0065_),
    .Q(\po_0.regf_0.rf[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3091_ (.CLK(net150),
    .D(_0066_),
    .Q(\po_0.regf_0.rf[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3092_ (.CLK(net156),
    .D(_0067_),
    .Q(\po_0.regf_0.rf[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3093_ (.CLK(net165),
    .D(_0068_),
    .Q(\po_0.regf_0.rf[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3094_ (.CLK(net156),
    .D(_0069_),
    .Q(\po_0.regf_0.rf[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3095_ (.CLK(net133),
    .D(_0070_),
    .Q(\po_0.regf_0.rf[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3096_ (.CLK(net134),
    .D(_0071_),
    .Q(\po_0.regf_0.rf[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3097_ (.CLK(net113),
    .D(_0072_),
    .Q(\po_0.regf_0.rf[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3098_ (.CLK(net132),
    .D(_0073_),
    .Q(\po_0.regf_0.rf[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3099_ (.CLK(net130),
    .D(_0074_),
    .Q(\po_0.regf_0.rf[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3100_ (.CLK(net103),
    .D(_0075_),
    .Q(\po_0.regf_0.rf[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3101_ (.CLK(net100),
    .D(_0076_),
    .Q(\po_0.regf_0.rf[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3102_ (.CLK(net100),
    .D(_0077_),
    .Q(\po_0.regf_0.rf[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3103_ (.CLK(net100),
    .D(_0078_),
    .Q(\po_0.regf_0.rf[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3104_ (.CLK(net100),
    .D(_0079_),
    .Q(\po_0.regf_0.rf[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3105_ (.CLK(net164),
    .D(_0080_),
    .Q(\po_0.regf_0.rf[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3106_ (.CLK(net143),
    .D(_0081_),
    .Q(\po_0.regf_0.rf[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3107_ (.CLK(net151),
    .D(_0082_),
    .Q(\po_0.regf_0.rf[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3108_ (.CLK(net159),
    .D(_0083_),
    .Q(\po_0.regf_0.rf[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3109_ (.CLK(net165),
    .D(_0084_),
    .Q(\po_0.regf_0.rf[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3110_ (.CLK(net156),
    .D(_0085_),
    .Q(\po_0.regf_0.rf[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3111_ (.CLK(net132),
    .D(_0086_),
    .Q(\po_0.regf_0.rf[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3112_ (.CLK(net133),
    .D(_0087_),
    .Q(\po_0.regf_0.rf[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3113_ (.CLK(net128),
    .D(_0088_),
    .Q(\po_0.regf_0.rf[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3114_ (.CLK(net126),
    .D(_0089_),
    .Q(\po_0.regf_0.rf[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3115_ (.CLK(net130),
    .D(_0090_),
    .Q(\po_0.regf_0.rf[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3116_ (.CLK(net121),
    .D(_0091_),
    .Q(\po_0.regf_0.rf[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3117_ (.CLK(net119),
    .D(_0092_),
    .Q(\po_0.regf_0.rf[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3118_ (.CLK(net125),
    .D(_0093_),
    .Q(\po_0.regf_0.rf[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3119_ (.CLK(net99),
    .D(_0094_),
    .Q(\po_0.regf_0.rf[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3120_ (.CLK(net118),
    .D(_0095_),
    .Q(\po_0.regf_0.rf[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3121_ (.CLK(net147),
    .D(_0096_),
    .Q(\po_0.regf_0.rf[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3122_ (.CLK(net140),
    .D(_0097_),
    .Q(\po_0.regf_0.rf[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3123_ (.CLK(net141),
    .D(_0098_),
    .Q(\po_0.regf_0.rf[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3124_ (.CLK(net141),
    .D(_0099_),
    .Q(\po_0.regf_0.rf[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3125_ (.CLK(net140),
    .D(_0100_),
    .Q(\po_0.regf_0.rf[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3126_ (.CLK(net137),
    .D(_0101_),
    .Q(\po_0.regf_0.rf[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3127_ (.CLK(net108),
    .D(_0102_),
    .Q(\po_0.regf_0.rf[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3128_ (.CLK(net108),
    .D(_0103_),
    .Q(\po_0.regf_0.rf[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3129_ (.CLK(net107),
    .D(_0104_),
    .Q(\po_0.regf_0.rf[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3130_ (.CLK(net106),
    .D(_0105_),
    .Q(\po_0.regf_0.rf[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3131_ (.CLK(net109),
    .D(_0106_),
    .Q(\po_0.regf_0.rf[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3132_ (.CLK(net106),
    .D(_0107_),
    .Q(\po_0.regf_0.rf[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3133_ (.CLK(net96),
    .D(_0108_),
    .Q(\po_0.regf_0.rf[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3134_ (.CLK(net96),
    .D(_0109_),
    .Q(\po_0.regf_0.rf[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3135_ (.CLK(net96),
    .D(_0110_),
    .Q(\po_0.regf_0.rf[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3136_ (.CLK(net97),
    .D(_0111_),
    .Q(\po_0.regf_0.rf[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3137_ (.CLK(net147),
    .D(_0112_),
    .Q(\po_0.regf_0.rf[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3138_ (.CLK(net140),
    .D(_0113_),
    .Q(\po_0.regf_0.rf[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3139_ (.CLK(net141),
    .D(_0114_),
    .Q(\po_0.regf_0.rf[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3140_ (.CLK(net141),
    .D(_0115_),
    .Q(\po_0.regf_0.rf[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3141_ (.CLK(net140),
    .D(_0116_),
    .Q(\po_0.regf_0.rf[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3142_ (.CLK(net137),
    .D(_0117_),
    .Q(\po_0.regf_0.rf[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3143_ (.CLK(net108),
    .D(_0118_),
    .Q(\po_0.regf_0.rf[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3144_ (.CLK(net108),
    .D(_0119_),
    .Q(\po_0.regf_0.rf[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3145_ (.CLK(net107),
    .D(_0120_),
    .Q(\po_0.regf_0.rf[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3146_ (.CLK(net106),
    .D(_0121_),
    .Q(\po_0.regf_0.rf[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3147_ (.CLK(net109),
    .D(_0122_),
    .Q(\po_0.regf_0.rf[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3148_ (.CLK(net106),
    .D(_0123_),
    .Q(\po_0.regf_0.rf[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3149_ (.CLK(net96),
    .D(_0124_),
    .Q(\po_0.regf_0.rf[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3150_ (.CLK(net96),
    .D(_0125_),
    .Q(\po_0.regf_0.rf[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3151_ (.CLK(net97),
    .D(_0126_),
    .Q(\po_0.regf_0.rf[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3152_ (.CLK(net97),
    .D(_0127_),
    .Q(\po_0.regf_0.rf[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3153_ (.CLK(net148),
    .D(_0128_),
    .Q(\po_0.regf_0.rf[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3154_ (.CLK(net142),
    .D(_0129_),
    .Q(\po_0.regf_0.rf[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3155_ (.CLK(net142),
    .D(_0130_),
    .Q(\po_0.regf_0.rf[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3156_ (.CLK(net141),
    .D(_0131_),
    .Q(\po_0.regf_0.rf[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3157_ (.CLK(net147),
    .D(_0132_),
    .Q(\po_0.regf_0.rf[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3158_ (.CLK(net137),
    .D(_0133_),
    .Q(\po_0.regf_0.rf[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3159_ (.CLK(net108),
    .D(_0134_),
    .Q(\po_0.regf_0.rf[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3160_ (.CLK(net110),
    .D(_0135_),
    .Q(\po_0.regf_0.rf[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3161_ (.CLK(net107),
    .D(_0136_),
    .Q(\po_0.regf_0.rf[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3162_ (.CLK(net107),
    .D(_0137_),
    .Q(\po_0.regf_0.rf[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3163_ (.CLK(net110),
    .D(_0138_),
    .Q(\po_0.regf_0.rf[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3164_ (.CLK(net106),
    .D(_0139_),
    .Q(\po_0.regf_0.rf[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3165_ (.CLK(net96),
    .D(_0140_),
    .Q(\po_0.regf_0.rf[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3166_ (.CLK(net98),
    .D(_0141_),
    .Q(\po_0.regf_0.rf[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3167_ (.CLK(net98),
    .D(_0142_),
    .Q(\po_0.regf_0.rf[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3168_ (.CLK(net97),
    .D(_0143_),
    .Q(\po_0.regf_0.rf[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3169_ (.CLK(net148),
    .D(_0144_),
    .Q(\po_0.regf_0.rf[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3170_ (.CLK(net140),
    .D(_0145_),
    .Q(\po_0.regf_0.rf[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3171_ (.CLK(net142),
    .D(_0146_),
    .Q(\po_0.regf_0.rf[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3172_ (.CLK(net141),
    .D(_0147_),
    .Q(\po_0.regf_0.rf[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3173_ (.CLK(net147),
    .D(_0148_),
    .Q(\po_0.regf_0.rf[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3174_ (.CLK(net137),
    .D(_0149_),
    .Q(\po_0.regf_0.rf[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3175_ (.CLK(net108),
    .D(_0150_),
    .Q(\po_0.regf_0.rf[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3176_ (.CLK(net110),
    .D(_0151_),
    .Q(\po_0.regf_0.rf[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3177_ (.CLK(net111),
    .D(_0152_),
    .Q(\po_0.regf_0.rf[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3178_ (.CLK(net111),
    .D(_0153_),
    .Q(\po_0.regf_0.rf[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3179_ (.CLK(net109),
    .D(_0154_),
    .Q(\po_0.regf_0.rf[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3180_ (.CLK(net106),
    .D(_0155_),
    .Q(\po_0.regf_0.rf[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3181_ (.CLK(net97),
    .D(_0156_),
    .Q(\po_0.regf_0.rf[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3182_ (.CLK(net98),
    .D(_0157_),
    .Q(\po_0.regf_0.rf[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3183_ (.CLK(net98),
    .D(_0158_),
    .Q(\po_0.regf_0.rf[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3184_ (.CLK(net103),
    .D(_0159_),
    .Q(\po_0.regf_0.rf[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3185_ (.CLK(net151),
    .D(_0160_),
    .Q(\po_0.regf_0.rf[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3186_ (.CLK(net145),
    .D(_0161_),
    .Q(\po_0.regf_0.rf[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3187_ (.CLK(net150),
    .D(_0162_),
    .Q(\po_0.regf_0.rf[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3188_ (.CLK(net158),
    .D(_0163_),
    .Q(\po_0.regf_0.rf[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3189_ (.CLK(net158),
    .D(_0164_),
    .Q(\po_0.regf_0.rf[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3190_ (.CLK(net156),
    .D(_0165_),
    .Q(\po_0.regf_0.rf[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3191_ (.CLK(net114),
    .D(_0166_),
    .Q(\po_0.regf_0.rf[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3192_ (.CLK(net114),
    .D(_0167_),
    .Q(\po_0.regf_0.rf[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3193_ (.CLK(net112),
    .D(_0168_),
    .Q(\po_0.regf_0.rf[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3194_ (.CLK(net112),
    .D(_0169_),
    .Q(\po_0.regf_0.rf[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3195_ (.CLK(net114),
    .D(_0170_),
    .Q(\po_0.regf_0.rf[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3196_ (.CLK(net112),
    .D(_0171_),
    .Q(\po_0.regf_0.rf[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3197_ (.CLK(net103),
    .D(_0172_),
    .Q(\po_0.regf_0.rf[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3198_ (.CLK(net99),
    .D(_0173_),
    .Q(\po_0.regf_0.rf[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3199_ (.CLK(net99),
    .D(_0174_),
    .Q(\po_0.regf_0.rf[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3200_ (.CLK(net103),
    .D(_0175_),
    .Q(\po_0.regf_0.rf[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3201_ (.CLK(net151),
    .D(_0176_),
    .Q(\po_0.regf_0.rf[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3202_ (.CLK(net145),
    .D(_0177_),
    .Q(\po_0.regf_0.rf[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3203_ (.CLK(net150),
    .D(_0178_),
    .Q(\po_0.regf_0.rf[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3204_ (.CLK(net158),
    .D(_0179_),
    .Q(\po_0.regf_0.rf[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3205_ (.CLK(net158),
    .D(_0180_),
    .Q(\po_0.regf_0.rf[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3206_ (.CLK(net156),
    .D(_0181_),
    .Q(\po_0.regf_0.rf[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3207_ (.CLK(net114),
    .D(_0182_),
    .Q(\po_0.regf_0.rf[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3208_ (.CLK(net114),
    .D(_0183_),
    .Q(\po_0.regf_0.rf[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3209_ (.CLK(net112),
    .D(_0184_),
    .Q(\po_0.regf_0.rf[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3210_ (.CLK(net112),
    .D(_0185_),
    .Q(\po_0.regf_0.rf[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3211_ (.CLK(net115),
    .D(_0186_),
    .Q(\po_0.regf_0.rf[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3212_ (.CLK(net112),
    .D(_0187_),
    .Q(\po_0.regf_0.rf[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3213_ (.CLK(net103),
    .D(_0188_),
    .Q(\po_0.regf_0.rf[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3214_ (.CLK(net101),
    .D(_0189_),
    .Q(\po_0.regf_0.rf[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3215_ (.CLK(net102),
    .D(_0190_),
    .Q(\po_0.regf_0.rf[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3216_ (.CLK(net103),
    .D(_0191_),
    .Q(\po_0.regf_0.rf[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3217_ (.CLK(net164),
    .D(_0192_),
    .Q(\po_0.regf_0.rf[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3218_ (.CLK(net144),
    .D(_0193_),
    .Q(\po_0.regf_0.rf[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3219_ (.CLK(net151),
    .D(_0194_),
    .Q(\po_0.regf_0.rf[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3220_ (.CLK(net159),
    .D(_0195_),
    .Q(\po_0.regf_0.rf[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3221_ (.CLK(net165),
    .D(_0196_),
    .Q(\po_0.regf_0.rf[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3222_ (.CLK(net157),
    .D(_0197_),
    .Q(\po_0.regf_0.rf[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3223_ (.CLK(net132),
    .D(_0198_),
    .Q(\po_0.regf_0.rf[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3224_ (.CLK(net134),
    .D(_0199_),
    .Q(\po_0.regf_0.rf[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3225_ (.CLK(net128),
    .D(_0200_),
    .Q(\po_0.regf_0.rf[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3226_ (.CLK(net126),
    .D(_0201_),
    .Q(\po_0.regf_0.rf[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3227_ (.CLK(net130),
    .D(_0202_),
    .Q(\po_0.regf_0.rf[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3228_ (.CLK(net121),
    .D(_0203_),
    .Q(\po_0.regf_0.rf[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3229_ (.CLK(net119),
    .D(_0204_),
    .Q(\po_0.regf_0.rf[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3230_ (.CLK(net119),
    .D(_0205_),
    .Q(\po_0.regf_0.rf[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3231_ (.CLK(net99),
    .D(_0206_),
    .Q(\po_0.regf_0.rf[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3232_ (.CLK(net120),
    .D(_0207_),
    .Q(\po_0.regf_0.rf[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3233_ (.CLK(net164),
    .D(_0208_),
    .Q(\po_0.regf_0.rf[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3234_ (.CLK(net145),
    .D(_0209_),
    .Q(\po_0.regf_0.rf[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3235_ (.CLK(net154),
    .D(_0210_),
    .Q(\po_0.regf_0.rf[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3236_ (.CLK(net158),
    .D(_0211_),
    .Q(\po_0.regf_0.rf[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3237_ (.CLK(net159),
    .D(_0212_),
    .Q(\po_0.regf_0.rf[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3238_ (.CLK(net156),
    .D(_0213_),
    .Q(\po_0.regf_0.rf[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3239_ (.CLK(net115),
    .D(_0214_),
    .Q(\po_0.regf_0.rf[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3240_ (.CLK(net115),
    .D(_0215_),
    .Q(\po_0.regf_0.rf[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3241_ (.CLK(net113),
    .D(_0216_),
    .Q(\po_0.regf_0.rf[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3242_ (.CLK(net113),
    .D(_0217_),
    .Q(\po_0.regf_0.rf[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3243_ (.CLK(net115),
    .D(_0218_),
    .Q(\po_0.regf_0.rf[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3244_ (.CLK(net113),
    .D(_0219_),
    .Q(\po_0.regf_0.rf[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3245_ (.CLK(net104),
    .D(_0220_),
    .Q(\po_0.regf_0.rf[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3246_ (.CLK(net101),
    .D(_0221_),
    .Q(\po_0.regf_0.rf[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3247_ (.CLK(net101),
    .D(_0222_),
    .Q(\po_0.regf_0.rf[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3248_ (.CLK(net104),
    .D(_0223_),
    .Q(\po_0.regf_0.rf[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3249_ (.CLK(net171),
    .D(_0224_),
    .Q(\po_0.muxf_0.rf_w_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3250_ (.CLK(net172),
    .D(_0225_),
    .Q(\po_0.muxf_0.rf_w_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3251_ (.CLK(net171),
    .D(_0226_),
    .Q(\po_0.muxf_0.rf_w_data[2] ));
 sky130_fd_sc_hd__dfxtp_4 _3252_ (.CLK(net171),
    .D(_0227_),
    .Q(\po_0.muxf_0.rf_w_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3253_ (.CLK(net166),
    .D(_0228_),
    .Q(\po_0.muxf_0.rf_w_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3254_ (.CLK(net153),
    .D(_0229_),
    .Q(\po_0.muxf_0.rf_w_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3255_ (.CLK(net153),
    .D(_0230_),
    .Q(\po_0.muxf_0.rf_w_data[6] ));
 sky130_fd_sc_hd__dfxtp_2 _3256_ (.CLK(net137),
    .D(_0231_),
    .Q(\po_0.muxf_0.rf_w_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3257_ (.CLK(net138),
    .D(_0232_),
    .Q(\uc_0._20_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3258_ (.CLK(net114),
    .D(_0233_),
    .Q(\uc_0._20_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3259_ (.CLK(net140),
    .D(_0234_),
    .Q(\uc_0._20_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3260_ (.CLK(net137),
    .D(_0235_),
    .Q(\uc_0._20_[11] ));
 sky130_fd_sc_hd__dfxtp_2 _3261_ (.CLK(net147),
    .D(_0236_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_2 _3262_ (.CLK(net172),
    .D(_0237_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_2 _3263_ (.CLK(net107),
    .D(_0238_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _3264_ (.CLK(net164),
    .D(_0239_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _3265_ (.CLK(net152),
    .D(_0012_),
    .Q(_0004_));
 sky130_fd_sc_hd__dfxtp_1 _3266_ (.CLK(net154),
    .D(_0013_),
    .Q(_0005_));
 sky130_fd_sc_hd__dfxtp_1 _3267_ (.CLK(net152),
    .D(_0014_),
    .Q(_0006_));
 sky130_fd_sc_hd__dfxtp_2 _3268_ (.CLK(net152),
    .D(_0015_),
    .Q(_0007_));
 sky130_fd_sc_hd__dfxtp_1 _3269_ (.CLK(net166),
    .D(_0240_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _3270_ (.CLK(net172),
    .D(_0241_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_2 _3271_ (.CLK(net167),
    .D(_0242_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_2 _3272_ (.CLK(net167),
    .D(_0243_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _3273_ (.CLK(net166),
    .D(_0244_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_2 _3274_ (.CLK(net166),
    .D(_0245_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_2 _3275_ (.CLK(net152),
    .D(_0246_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_2 _3276_ (.CLK(net166),
    .D(_0247_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _3277_ (.CLK(net166),
    .D(_0248_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _3278_ (.CLK(net167),
    .D(net182),
    .Q(net76));
 sky130_fd_sc_hd__conb_1 _3278__182 (.LO(net182));
 sky130_fd_sc_hd__dfxtp_1 _3279_ (.CLK(net119),
    .D(net181),
    .Q(net62));
 sky130_fd_sc_hd__conb_1 _3279__181 (.LO(net181));
 sky130_fd_sc_hd__dfxtp_1 _3280_ (.CLK(net149),
    .D(net180),
    .Q(net63));
 sky130_fd_sc_hd__conb_1 _3280__180 (.LO(net180));
 sky130_fd_sc_hd__dfxtp_2 _3281_ (.CLK(net125),
    .D(net179),
    .Q(net64));
 sky130_fd_sc_hd__conb_1 _3281__179 (.LO(net179));
 sky130_fd_sc_hd__dfxtp_1 _3282_ (.CLK(net154),
    .D(net178),
    .Q(net65));
 sky130_fd_sc_hd__conb_1 _3282__178 (.LO(net178));
 sky130_fd_sc_hd__dfxtp_2 _3283_ (.CLK(net126),
    .D(net177),
    .Q(net66));
 sky130_fd_sc_hd__conb_1 _3283__177 (.LO(net177));
 sky130_fd_sc_hd__dfxtp_1 _3284_ (.CLK(net172),
    .D(net176),
    .Q(net67));
 sky130_fd_sc_hd__conb_1 _3284__176 (.LO(net176));
 sky130_fd_sc_hd__dfxtp_1 _3285_ (.CLK(net171),
    .D(_0256_),
    .Q(\uc_0._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _3286_ (.CLK(net169),
    .D(_0257_),
    .Q(\po_0.regf_0.rf[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3287_ (.CLK(net143),
    .D(_0258_),
    .Q(\po_0.regf_0.rf[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3288_ (.CLK(net150),
    .D(_0259_),
    .Q(\po_0.regf_0.rf[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3289_ (.CLK(net161),
    .D(_0260_),
    .Q(\po_0.regf_0.rf[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3290_ (.CLK(net161),
    .D(_0261_),
    .Q(\po_0.regf_0.rf[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3291_ (.CLK(net163),
    .D(_0262_),
    .Q(\po_0.regf_0.rf[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3292_ (.CLK(net135),
    .D(_0263_),
    .Q(\po_0.regf_0.rf[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3293_ (.CLK(net134),
    .D(_0264_),
    .Q(\po_0.regf_0.rf[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3294_ (.CLK(net135),
    .D(_0265_),
    .Q(\po_0.regf_0.rf[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3295_ (.CLK(net127),
    .D(_0266_),
    .Q(\po_0.regf_0.rf[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3296_ (.CLK(net135),
    .D(_0267_),
    .Q(\po_0.regf_0.rf[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3297_ (.CLK(net127),
    .D(_0268_),
    .Q(\po_0.regf_0.rf[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3298_ (.CLK(net125),
    .D(_0269_),
    .Q(\po_0.regf_0.rf[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3299_ (.CLK(net125),
    .D(_0270_),
    .Q(\po_0.regf_0.rf[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3300_ (.CLK(net118),
    .D(_0271_),
    .Q(\po_0.regf_0.rf[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3301_ (.CLK(net119),
    .D(_0272_),
    .Q(\po_0.regf_0.rf[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3302_ (.CLK(net164),
    .D(_0273_),
    .Q(\po_0.regf_0.rf[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3303_ (.CLK(net144),
    .D(_0274_),
    .Q(\po_0.regf_0.rf[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3304_ (.CLK(net150),
    .D(_0275_),
    .Q(\po_0.regf_0.rf[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3305_ (.CLK(net159),
    .D(_0276_),
    .Q(\po_0.regf_0.rf[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3306_ (.CLK(net168),
    .D(_0277_),
    .Q(\po_0.regf_0.rf[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3307_ (.CLK(net157),
    .D(_0278_),
    .Q(\po_0.regf_0.rf[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3308_ (.CLK(net128),
    .D(_0279_),
    .Q(\po_0.regf_0.rf[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3309_ (.CLK(net131),
    .D(_0280_),
    .Q(\po_0.regf_0.rf[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3310_ (.CLK(net128),
    .D(_0281_),
    .Q(\po_0.regf_0.rf[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3311_ (.CLK(net128),
    .D(_0282_),
    .Q(\po_0.regf_0.rf[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3312_ (.CLK(net130),
    .D(_0283_),
    .Q(\po_0.regf_0.rf[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3313_ (.CLK(net128),
    .D(_0284_),
    .Q(\po_0.regf_0.rf[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3314_ (.CLK(net122),
    .D(_0285_),
    .Q(\po_0.regf_0.rf[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3315_ (.CLK(net120),
    .D(_0286_),
    .Q(\po_0.regf_0.rf[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3316_ (.CLK(net99),
    .D(_0287_),
    .Q(\po_0.regf_0.rf[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3317_ (.CLK(net121),
    .D(_0288_),
    .Q(\po_0.regf_0.rf[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3318_ (.CLK(net165),
    .D(_0289_),
    .Q(\po_0.regf_0.rf[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3319_ (.CLK(net144),
    .D(_0290_),
    .Q(\po_0.regf_0.rf[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3320_ (.CLK(net151),
    .D(_0291_),
    .Q(\po_0.regf_0.rf[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3321_ (.CLK(net158),
    .D(_0292_),
    .Q(\po_0.regf_0.rf[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3322_ (.CLK(net168),
    .D(_0293_),
    .Q(\po_0.regf_0.rf[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3323_ (.CLK(net157),
    .D(_0294_),
    .Q(\po_0.regf_0.rf[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3324_ (.CLK(net129),
    .D(_0295_),
    .Q(\po_0.regf_0.rf[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3325_ (.CLK(net131),
    .D(_0296_),
    .Q(\po_0.regf_0.rf[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3326_ (.CLK(net129),
    .D(_0297_),
    .Q(\po_0.regf_0.rf[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3327_ (.CLK(net122),
    .D(_0298_),
    .Q(\po_0.regf_0.rf[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3328_ (.CLK(net130),
    .D(_0299_),
    .Q(\po_0.regf_0.rf[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3329_ (.CLK(net122),
    .D(_0300_),
    .Q(\po_0.regf_0.rf[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3330_ (.CLK(net122),
    .D(_0301_),
    .Q(\po_0.regf_0.rf[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3331_ (.CLK(net120),
    .D(_0302_),
    .Q(\po_0.regf_0.rf[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3332_ (.CLK(net99),
    .D(_0303_),
    .Q(\po_0.regf_0.rf[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3333_ (.CLK(net120),
    .D(_0304_),
    .Q(\po_0.regf_0.rf[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3334_ (.CLK(net161),
    .D(_0305_),
    .Q(\po_0.alu_0.s1 ));
 sky130_fd_sc_hd__dfxtp_1 _3335_ (.CLK(net162),
    .D(_0306_),
    .Q(\po_0.alu_0.s0 ));
 sky130_fd_sc_hd__dfxtp_1 _3336_ (.CLK(net162),
    .D(_0307_),
    .Q(\po_0.regf_0.rq_rd ));
 sky130_fd_sc_hd__dfxtp_1 _3337_ (.CLK(net170),
    .D(_0308_),
    .Q(\po_0.regf_0.rp_rd ));
 sky130_fd_sc_hd__dfxtp_1 _3338_ (.CLK(net145),
    .D(_0309_),
    .Q(\po_0.regf_0.w_wr ));
 sky130_fd_sc_hd__dfxtp_1 _3339_ (.CLK(net152),
    .D(_0310_),
    .Q(\po_0.regf_0.rq_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3340_ (.CLK(net152),
    .D(_0311_),
    .Q(\po_0.regf_0.rq_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3341_ (.CLK(net153),
    .D(_0312_),
    .Q(\po_0.regf_0.rq_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3342_ (.CLK(net153),
    .D(_0313_),
    .Q(\po_0.regf_0.rq_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3343_ (.CLK(net138),
    .D(_0314_),
    .Q(\po_0.regf_0.rp_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3344_ (.CLK(net110),
    .D(_0315_),
    .Q(\po_0.regf_0.rp_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3345_ (.CLK(net139),
    .D(_0316_),
    .Q(\po_0.regf_0.rp_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3346_ (.CLK(net139),
    .D(_0317_),
    .Q(\po_0.regf_0.rp_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3347_ (.CLK(net138),
    .D(_0318_),
    .Q(\po_0.regf_0.w_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3348_ (.CLK(net145),
    .D(_0319_),
    .Q(\po_0.regf_0.w_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3349_ (.CLK(net138),
    .D(_0320_),
    .Q(\po_0.regf_0.w_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3350_ (.CLK(net138),
    .D(_0321_),
    .Q(\po_0.regf_0.w_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3351_ (.CLK(net162),
    .D(_0322_),
    .Q(\po_0.muxf_0.s0 ));
 sky130_fd_sc_hd__dfxtp_1 _3352_ (.CLK(net162),
    .D(_0323_),
    .Q(\po_0.muxf_0.s1 ));
 sky130_fd_sc_hd__dfxtp_1 _3353_ (.CLK(net170),
    .D(_0324_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _3354_ (.CLK(net169),
    .D(_0325_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _3355_ (.CLK(net148),
    .D(_0326_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _3356_ (.CLK(net167),
    .D(_0327_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _3357_ (.CLK(net100),
    .D(_0328_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _3358_ (.CLK(net124),
    .D(_0329_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _3359_ (.CLK(net170),
    .D(_0330_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _3360_ (.CLK(net153),
    .D(_0331_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _3361_ (.CLK(net139),
    .D(_0332_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _3362_ (.CLK(net98),
    .D(_0333_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _3363_ (.CLK(net172),
    .D(_0334_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _3364_ (.CLK(net173),
    .D(_0335_),
    .Q(\uc_0._03_ ));
 sky130_fd_sc_hd__dfxtp_1 _3365_ (.CLK(net171),
    .D(_0336_),
    .Q(\uc_0._02_ ));
 sky130_fd_sc_hd__dfxtp_1 _3366_ (.CLK(net171),
    .D(_0337_),
    .Q(\uc_0._01_ ));
 sky130_fd_sc_hd__dfxtp_1 _3367_ (.CLK(net170),
    .D(\uc_0.bc_0._54_[0] ),
    .Q(\uc_0.bc_0._55_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3368_ (.CLK(net173),
    .D(\uc_0.bc_0._54_[1] ),
    .Q(\uc_0.bc_0._55_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3369_ (.CLK(net170),
    .D(\uc_0.bc_0._54_[2] ),
    .Q(\uc_0.bc_0._55_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3370_ (.CLK(net173),
    .D(\uc_0.bc_0._54_[3] ),
    .Q(\uc_0.bc_0._55_[3] ));
 sky130_fd_sc_hd__clkbuf_1 _3378_ (.A(net149),
    .X(net78));
 sky130_fd_sc_hd__ebufn_1 _3379_ (.A(\po_0.alu_0._10_[0] ),
    .TE_B(_1468_),
    .Z(\po_0.alu_0._11_[0] ));
 sky130_fd_sc_hd__ebufn_1 _3380_ (.A(\po_0.alu_0._10_[1] ),
    .TE_B(_1469_),
    .Z(\po_0.alu_0._11_[1] ));
 sky130_fd_sc_hd__ebufn_1 _3381_ (.A(\po_0.alu_0._10_[2] ),
    .TE_B(_1470_),
    .Z(\po_0.alu_0._11_[2] ));
 sky130_fd_sc_hd__ebufn_1 _3382_ (.A(\po_0.alu_0._10_[3] ),
    .TE_B(_1471_),
    .Z(\po_0.alu_0._11_[3] ));
 sky130_fd_sc_hd__ebufn_1 _3383_ (.A(\po_0.alu_0._10_[4] ),
    .TE_B(_1472_),
    .Z(\po_0.alu_0._11_[4] ));
 sky130_fd_sc_hd__ebufn_1 _3384_ (.A(\po_0.alu_0._10_[5] ),
    .TE_B(_1473_),
    .Z(\po_0.alu_0._11_[5] ));
 sky130_fd_sc_hd__ebufn_1 _3385_ (.A(\po_0.alu_0._10_[6] ),
    .TE_B(_1474_),
    .Z(\po_0.alu_0._11_[6] ));
 sky130_fd_sc_hd__ebufn_1 _3386_ (.A(\po_0.alu_0._10_[7] ),
    .TE_B(_1475_),
    .Z(\po_0.alu_0._11_[7] ));
 sky130_fd_sc_hd__ebufn_1 _3387_ (.A(\po_0.alu_0._10_[8] ),
    .TE_B(_1476_),
    .Z(\po_0.alu_0._11_[8] ));
 sky130_fd_sc_hd__ebufn_1 _3388_ (.A(\po_0.alu_0._10_[9] ),
    .TE_B(_1477_),
    .Z(\po_0.alu_0._11_[9] ));
 sky130_fd_sc_hd__ebufn_1 _3389_ (.A(\po_0.alu_0._10_[10] ),
    .TE_B(_1478_),
    .Z(\po_0.alu_0._11_[10] ));
 sky130_fd_sc_hd__ebufn_2 _3390_ (.A(\po_0.alu_0._10_[11] ),
    .TE_B(_1479_),
    .Z(\po_0.alu_0._11_[11] ));
 sky130_fd_sc_hd__ebufn_1 _3391_ (.A(\po_0.alu_0._10_[12] ),
    .TE_B(_1480_),
    .Z(\po_0.alu_0._11_[12] ));
 sky130_fd_sc_hd__ebufn_1 _3392_ (.A(\po_0.alu_0._10_[13] ),
    .TE_B(_1481_),
    .Z(\po_0.alu_0._11_[13] ));
 sky130_fd_sc_hd__ebufn_1 _3393_ (.A(\po_0.alu_0._10_[14] ),
    .TE_B(_1482_),
    .Z(\po_0.alu_0._11_[14] ));
 sky130_fd_sc_hd__ebufn_1 _3394_ (.A(\po_0.alu_0._10_[15] ),
    .TE_B(_1483_),
    .Z(\po_0.alu_0._11_[15] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout100 (.A(net102),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 fanout101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout102 (.A(net104),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout105 (.A(net117),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout107 (.A(net111),
    .X(net107));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout108 (.A(net110),
    .X(net108));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout111 (.A(net117),
    .X(net111));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout112 (.A(net116),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 fanout113 (.A(net116),
    .X(net113));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout114 (.A(net116),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout117 (.A(net175),
    .X(net117));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout118 (.A(net120),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout120 (.A(net123),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 fanout121 (.A(net123),
    .X(net121));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 fanout123 (.A(net136),
    .X(net123));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(net127),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout127 (.A(net136),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout129 (.A(net131),
    .X(net129));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 fanout131 (.A(net136),
    .X(net131));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout132 (.A(net135),
    .X(net132));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 fanout136 (.A(net175),
    .X(net136));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout137 (.A(net139),
    .X(net137));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout139 (.A(net146),
    .X(net139));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout140 (.A(net142),
    .X(net140));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout142 (.A(net146),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 fanout143 (.A(net146),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout146 (.A(net155),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 fanout147 (.A(net149),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout149 (.A(net155),
    .X(net149));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout151 (.A(net154),
    .X(net151));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout155 (.A(net175),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 fanout156 (.A(net160),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 fanout157 (.A(net160),
    .X(net157));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 fanout160 (.A(net174),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 fanout161 (.A(net163),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 fanout163 (.A(net174),
    .X(net163));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout165 (.A(net168),
    .X(net165));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout168 (.A(net174),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 fanout170 (.A(net173),
    .X(net170));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__buf_2 fanout175 (.A(net33),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(net49),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 fanout84 (.A(net45),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 fanout85 (.A(net87),
    .X(net85));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_2 fanout87 (.A(\po_0.regf_0.rp_rd ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 fanout88 (.A(net91),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 fanout89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(\po_0.regf_0.rq_rd ),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(net68),
    .X(net92));
 sky130_fd_sc_hd__buf_2 fanout93 (.A(net61),
    .X(net93));
 sky130_fd_sc_hd__buf_2 fanout94 (.A(net82),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 fanout95 (.A(net81),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 fanout96 (.A(net105),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 fanout97 (.A(net98),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 fanout98 (.A(net105),
    .X(net98));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout99 (.A(net102),
    .X(net99));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(D_R_data[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(D_R_data[3]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(D_R_data[4]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(D_R_data[5]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(D_R_data[6]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(D_R_data[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(D_R_data[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(D_R_data[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(I_data[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(I_data[10]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(I_data[11]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(D_R_data[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(I_data[12]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(I_data[13]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(I_data[14]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(I_data[15]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(I_data[1]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(I_data[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(I_data[3]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(I_data[4]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(I_data[5]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(I_data[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input3 (.A(D_R_data[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(I_data[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(I_data[8]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(I_data[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(clock),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(reset),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(D_R_data[12]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(D_R_data[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(D_R_data[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(D_R_data[15]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(D_R_data[1]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(D_R_data[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(D_W_data[0]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(D_W_data[10]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(D_W_data[11]));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net38),
    .X(D_W_data[12]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(D_W_data[13]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(D_W_data[14]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(D_W_data[15]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(D_W_data[1]));
 sky130_fd_sc_hd__clkbuf_4 output43 (.A(net43),
    .X(D_W_data[2]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(D_W_data[3]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net84),
    .X(D_W_data[4]));
 sky130_fd_sc_hd__clkbuf_4 output46 (.A(net46),
    .X(D_W_data[5]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(D_W_data[6]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(D_W_data[7]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net83),
    .X(D_W_data[8]));
 sky130_fd_sc_hd__clkbuf_4 output50 (.A(net50),
    .X(D_W_data[9]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(D_addr[0]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(D_addr[1]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(D_addr[2]));
 sky130_fd_sc_hd__clkbuf_4 output54 (.A(net54),
    .X(D_addr[3]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(D_addr[4]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(D_addr[5]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(D_addr[6]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(D_addr[7]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(D_rd));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(D_wr));
 sky130_fd_sc_hd__buf_2 output61 (.A(net93),
    .X(I_addr[0]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(I_addr[10]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(I_addr[11]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(I_addr[12]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(I_addr[13]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(I_addr[14]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(I_addr[15]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net92),
    .X(I_addr[1]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(I_addr[2]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(I_addr[3]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(I_addr[4]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(I_addr[5]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(I_addr[6]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(I_addr[7]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(I_addr[8]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(I_addr[9]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(I_rd));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(led_clock));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(leds[0]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(leds[1]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net95),
    .X(leds[2]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net94),
    .X(leds[3]));
endmodule

