magic
tech sky130A
magscale 1 2
timestamp 1680041752
<< checkpaint >>
rect -3932 -3932 52212 54356
<< viali >>
rect 1777 47753 1811 47787
rect 3525 47753 3559 47787
rect 6101 47753 6135 47787
rect 10609 47753 10643 47787
rect 13185 47753 13219 47787
rect 15761 47753 15795 47787
rect 17509 47753 17543 47787
rect 17969 47753 18003 47787
rect 20361 47753 20395 47787
rect 22845 47753 22879 47787
rect 29285 47753 29319 47787
rect 32321 47753 32355 47787
rect 34437 47753 34471 47787
rect 36369 47753 36403 47787
rect 41521 47753 41555 47787
rect 6009 47685 6043 47719
rect 27261 47685 27295 47719
rect 1685 47617 1719 47651
rect 3341 47617 3375 47651
rect 8677 47617 8711 47651
rect 10425 47617 10459 47651
rect 13001 47617 13035 47651
rect 15577 47617 15611 47651
rect 17325 47617 17359 47651
rect 18245 47617 18279 47651
rect 19349 47617 19383 47651
rect 20177 47617 20211 47651
rect 22661 47617 22695 47651
rect 24593 47617 24627 47651
rect 29101 47617 29135 47651
rect 32229 47617 32263 47651
rect 34253 47617 34287 47651
rect 36185 47617 36219 47651
rect 38945 47617 38979 47651
rect 41429 47617 41463 47651
rect 43269 47617 43303 47651
rect 45845 47617 45879 47651
rect 45937 47617 45971 47651
rect 24869 47549 24903 47583
rect 43545 47549 43579 47583
rect 46213 47549 46247 47583
rect 8493 47481 8527 47515
rect 27445 47481 27479 47515
rect 18475 47413 18509 47447
rect 19441 47413 19475 47447
rect 38761 47413 38795 47447
rect 45661 47413 45695 47447
rect 3065 47209 3099 47243
rect 20637 47209 20671 47243
rect 25789 47209 25823 47243
rect 27261 47209 27295 47243
rect 29929 47209 29963 47243
rect 2145 47141 2179 47175
rect 30021 47141 30055 47175
rect 31125 47141 31159 47175
rect 17785 47073 17819 47107
rect 21741 47073 21775 47107
rect 27353 47073 27387 47107
rect 28273 47073 28307 47107
rect 31585 47073 31619 47107
rect 31769 47073 31803 47107
rect 1685 47005 1719 47039
rect 1961 47005 1995 47039
rect 3249 47005 3283 47039
rect 4629 47005 4663 47039
rect 18153 47005 18187 47039
rect 18245 47005 18279 47039
rect 18521 47005 18555 47039
rect 19257 47005 19291 47039
rect 21097 47005 21131 47039
rect 24225 47005 24259 47039
rect 24409 47005 24443 47039
rect 25881 47005 25915 47039
rect 27629 47005 27663 47039
rect 28549 47005 28583 47039
rect 29193 47005 29227 47039
rect 29377 47005 29411 47039
rect 29561 47005 29595 47039
rect 30205 47005 30239 47039
rect 30297 47005 30331 47039
rect 31493 47005 31527 47039
rect 31953 47005 31987 47039
rect 32229 47005 32263 47039
rect 34989 47005 35023 47039
rect 46765 47005 46799 47039
rect 4896 46937 4930 46971
rect 19502 46937 19536 46971
rect 22008 46937 22042 46971
rect 24654 46937 24688 46971
rect 26148 46937 26182 46971
rect 29745 46937 29779 46971
rect 30021 46937 30055 46971
rect 33609 46937 33643 46971
rect 6009 46869 6043 46903
rect 17141 46869 17175 46903
rect 17509 46869 17543 46903
rect 17601 46869 17635 46903
rect 20913 46869 20947 46903
rect 23121 46869 23155 46903
rect 29285 46869 29319 46903
rect 34805 46869 34839 46903
rect 46581 46869 46615 46903
rect 1593 46665 1627 46699
rect 18061 46665 18095 46699
rect 19625 46665 19659 46699
rect 21557 46665 21591 46699
rect 22385 46665 22419 46699
rect 25145 46665 25179 46699
rect 26525 46665 26559 46699
rect 32137 46665 32171 46699
rect 35449 46665 35483 46699
rect 1501 46597 1535 46631
rect 20444 46597 20478 46631
rect 23397 46597 23431 46631
rect 26433 46597 26467 46631
rect 34244 46597 34278 46631
rect 5089 46529 5123 46563
rect 16948 46529 16982 46563
rect 18501 46529 18535 46563
rect 22569 46529 22603 46563
rect 22845 46529 22879 46563
rect 23029 46529 23063 46563
rect 23121 46529 23155 46563
rect 23489 46529 23523 46563
rect 23756 46529 23790 46563
rect 25513 46529 25547 46563
rect 25697 46529 25731 46563
rect 25789 46529 25823 46563
rect 26985 46529 27019 46563
rect 27252 46529 27286 46563
rect 29653 46529 29687 46563
rect 29837 46529 29871 46563
rect 30205 46529 30239 46563
rect 30461 46529 30495 46563
rect 32321 46529 32355 46563
rect 35817 46529 35851 46563
rect 35909 46529 35943 46563
rect 36737 46529 36771 46563
rect 16681 46461 16715 46495
rect 18245 46461 18279 46495
rect 20177 46461 20211 46495
rect 22661 46461 22695 46495
rect 23213 46461 23247 46495
rect 23397 46461 23431 46495
rect 26709 46461 26743 46495
rect 29009 46461 29043 46495
rect 29193 46461 29227 46495
rect 29285 46461 29319 46495
rect 29377 46461 29411 46495
rect 29469 46461 29503 46495
rect 33057 46461 33091 46495
rect 33333 46461 33367 46495
rect 33977 46461 34011 46495
rect 36001 46461 36035 46495
rect 22753 46393 22787 46427
rect 25973 46393 26007 46427
rect 24869 46325 24903 46359
rect 25789 46325 25823 46359
rect 26065 46325 26099 46359
rect 28365 46325 28399 46359
rect 29653 46325 29687 46359
rect 31585 46325 31619 46359
rect 35357 46325 35391 46359
rect 36553 46325 36587 46359
rect 16957 46121 16991 46155
rect 21189 46121 21223 46155
rect 21373 46121 21407 46155
rect 23029 46121 23063 46155
rect 25329 46121 25363 46155
rect 26157 46121 26191 46155
rect 27353 46121 27387 46155
rect 30113 46121 30147 46155
rect 17417 46053 17451 46087
rect 28641 46053 28675 46087
rect 30481 46053 30515 46087
rect 17969 45985 18003 46019
rect 18245 45985 18279 46019
rect 20177 45985 20211 46019
rect 22937 45985 22971 46019
rect 24685 45985 24719 46019
rect 27721 45985 27755 46019
rect 28457 45985 28491 46019
rect 30389 45985 30423 46019
rect 36093 45985 36127 46019
rect 17141 45917 17175 45951
rect 17785 45917 17819 45951
rect 18521 45917 18555 45951
rect 20361 45917 20395 45951
rect 20637 45917 20671 45951
rect 20821 45917 20855 45951
rect 22569 45917 22603 45951
rect 22753 45917 22787 45951
rect 23029 45917 23063 45951
rect 23213 45917 23247 45951
rect 23305 45917 23339 45951
rect 23489 45917 23523 45951
rect 24409 45917 24443 45951
rect 25605 45917 25639 45951
rect 25789 45917 25823 45951
rect 25973 45917 26007 45951
rect 26065 45917 26099 45951
rect 26341 45917 26375 45951
rect 27537 45917 27571 45951
rect 27629 45917 27663 45951
rect 27813 45917 27847 45951
rect 27997 45917 28031 45951
rect 28917 45917 28951 45951
rect 30297 45917 30331 45951
rect 30573 45917 30607 45951
rect 30757 45917 30791 45951
rect 30849 45917 30883 45951
rect 33057 45917 33091 45951
rect 33517 45917 33551 45951
rect 33701 45917 33735 45951
rect 34805 45917 34839 45951
rect 36360 45917 36394 45951
rect 21189 45849 21223 45883
rect 33241 45849 33275 45883
rect 17877 45781 17911 45815
rect 20545 45781 20579 45815
rect 23397 45781 23431 45815
rect 25697 45781 25731 45815
rect 28825 45781 28859 45815
rect 31033 45781 31067 45815
rect 33425 45781 33459 45815
rect 33701 45781 33735 45815
rect 34897 45781 34931 45815
rect 37473 45781 37507 45815
rect 28457 45577 28491 45611
rect 31677 45577 31711 45611
rect 33793 45577 33827 45611
rect 37657 45577 37691 45611
rect 33425 45509 33459 45543
rect 33609 45509 33643 45543
rect 36737 45509 36771 45543
rect 17049 45441 17083 45475
rect 18061 45441 18095 45475
rect 19993 45441 20027 45475
rect 20177 45441 20211 45475
rect 28641 45441 28675 45475
rect 28733 45441 28767 45475
rect 28825 45441 28859 45475
rect 29009 45441 29043 45475
rect 29101 45441 29135 45475
rect 31309 45441 31343 45475
rect 31769 45441 31803 45475
rect 32781 45441 32815 45475
rect 32965 45441 32999 45475
rect 33057 45441 33091 45475
rect 33149 45441 33183 45475
rect 33701 45441 33735 45475
rect 46765 45441 46799 45475
rect 17141 45373 17175 45407
rect 17325 45373 17359 45407
rect 29193 45373 29227 45407
rect 29377 45373 29411 45407
rect 29469 45373 29503 45407
rect 29561 45373 29595 45407
rect 29653 45373 29687 45407
rect 30389 45373 30423 45407
rect 30665 45373 30699 45407
rect 37749 45373 37783 45407
rect 37841 45373 37875 45407
rect 17877 45305 17911 45339
rect 37289 45305 37323 45339
rect 46581 45305 46615 45339
rect 16681 45237 16715 45271
rect 20085 45237 20119 45271
rect 31447 45237 31481 45271
rect 31585 45237 31619 45271
rect 33333 45237 33367 45271
rect 33977 45237 34011 45271
rect 37013 45237 37047 45271
rect 20821 45033 20855 45067
rect 23305 45033 23339 45067
rect 25513 45033 25547 45067
rect 30849 45033 30883 45067
rect 31033 45033 31067 45067
rect 31125 45033 31159 45067
rect 32505 45033 32539 45067
rect 32965 45033 32999 45067
rect 16405 44965 16439 44999
rect 20913 44965 20947 44999
rect 25697 44965 25731 44999
rect 28641 44965 28675 44999
rect 30389 44965 30423 44999
rect 16957 44897 16991 44931
rect 17141 44897 17175 44931
rect 22017 44897 22051 44931
rect 22109 44897 22143 44931
rect 26709 44897 26743 44931
rect 26893 44897 26927 44931
rect 32689 44897 32723 44931
rect 15025 44829 15059 44863
rect 16865 44829 16899 44863
rect 20177 44829 20211 44863
rect 20270 44829 20304 44863
rect 20407 44829 20441 44863
rect 20642 44829 20676 44863
rect 21189 44829 21223 44863
rect 21281 44829 21315 44863
rect 21373 44829 21407 44863
rect 21557 44829 21591 44863
rect 22201 44829 22235 44863
rect 22293 44829 22327 44863
rect 22937 44829 22971 44863
rect 23121 44829 23155 44863
rect 25789 44829 25823 44863
rect 26617 44829 26651 44863
rect 26801 44829 26835 44863
rect 27629 44829 27663 44863
rect 27813 44829 27847 44863
rect 28181 44829 28215 44863
rect 28549 44829 28583 44863
rect 28917 44829 28951 44863
rect 29193 44829 29227 44863
rect 29377 44829 29411 44863
rect 30389 44829 30423 44863
rect 30573 44829 30607 44863
rect 31309 44829 31343 44863
rect 31585 44829 31619 44863
rect 31769 44829 31803 44863
rect 32321 44829 32355 44863
rect 32781 44829 32815 44863
rect 38853 44829 38887 44863
rect 25559 44795 25593 44829
rect 15292 44761 15326 44795
rect 20545 44761 20579 44795
rect 25329 44761 25363 44795
rect 26433 44761 26467 44795
rect 27997 44761 28031 44795
rect 28365 44761 28399 44795
rect 30665 44761 30699 44795
rect 16497 44693 16531 44727
rect 21833 44693 21867 44727
rect 25973 44693 26007 44727
rect 27721 44693 27755 44727
rect 28641 44693 28675 44727
rect 28733 44693 28767 44727
rect 29285 44693 29319 44727
rect 30875 44693 30909 44727
rect 39037 44693 39071 44727
rect 15393 44489 15427 44523
rect 16865 44489 16899 44523
rect 20085 44489 20119 44523
rect 27721 44489 27755 44523
rect 28641 44489 28675 44523
rect 33333 44489 33367 44523
rect 36369 44489 36403 44523
rect 37473 44489 37507 44523
rect 38393 44489 38427 44523
rect 17662 44421 17696 44455
rect 22937 44421 22971 44455
rect 23029 44421 23063 44455
rect 23229 44421 23263 44455
rect 29745 44421 29779 44455
rect 35256 44421 35290 44455
rect 38853 44421 38887 44455
rect 1409 44353 1443 44387
rect 15577 44353 15611 44387
rect 17049 44353 17083 44387
rect 19717 44353 19751 44387
rect 19901 44353 19935 44387
rect 20637 44353 20671 44387
rect 20821 44353 20855 44387
rect 22293 44353 22327 44387
rect 22661 44353 22695 44387
rect 25421 44353 25455 44387
rect 25605 44353 25639 44387
rect 25789 44353 25823 44387
rect 27077 44353 27111 44387
rect 27169 44353 27203 44387
rect 27537 44353 27571 44387
rect 28549 44353 28583 44387
rect 29561 44353 29595 44387
rect 29837 44353 29871 44387
rect 33241 44353 33275 44387
rect 33517 44353 33551 44387
rect 34989 44353 35023 44387
rect 37289 44353 37323 44387
rect 38301 44353 38335 44387
rect 38669 44353 38703 44387
rect 39773 44353 39807 44387
rect 17417 44285 17451 44319
rect 25973 44285 26007 44319
rect 28825 44285 28859 44319
rect 33793 44285 33827 44319
rect 39497 44285 39531 44319
rect 1593 44217 1627 44251
rect 22109 44217 22143 44251
rect 22661 44217 22695 44251
rect 25513 44217 25547 44251
rect 28181 44217 28215 44251
rect 18797 44149 18831 44183
rect 20637 44149 20671 44183
rect 23213 44149 23247 44183
rect 23397 44149 23431 44183
rect 27537 44149 27571 44183
rect 29837 44149 29871 44183
rect 20177 43945 20211 43979
rect 22569 43945 22603 43979
rect 24225 43945 24259 43979
rect 26157 43945 26191 43979
rect 33793 43945 33827 43979
rect 35081 43945 35115 43979
rect 37473 43945 37507 43979
rect 35449 43877 35483 43911
rect 20269 43809 20303 43843
rect 24777 43809 24811 43843
rect 28181 43809 28215 43843
rect 28273 43809 28307 43843
rect 28825 43809 28859 43843
rect 29285 43809 29319 43843
rect 29561 43809 29595 43843
rect 29837 43809 29871 43843
rect 29929 43809 29963 43843
rect 30021 43809 30055 43843
rect 38209 43809 38243 43843
rect 40417 43809 40451 43843
rect 15117 43741 15151 43775
rect 16865 43741 16899 43775
rect 16957 43741 16991 43775
rect 18889 43741 18923 43775
rect 19073 43741 19107 43775
rect 19349 43741 19383 43775
rect 19533 43741 19567 43775
rect 19717 43741 19751 43775
rect 20536 43741 20570 43775
rect 21925 43741 21959 43775
rect 22018 43741 22052 43775
rect 22201 43741 22235 43775
rect 22431 43741 22465 43775
rect 22845 43741 22879 43775
rect 24415 43741 24449 43775
rect 26433 43741 26467 43775
rect 26985 43741 27019 43775
rect 27169 43741 27203 43775
rect 28089 43735 28123 43769
rect 28365 43741 28399 43775
rect 28549 43741 28583 43775
rect 29009 43741 29043 43775
rect 29101 43741 29135 43775
rect 29193 43741 29227 43775
rect 29745 43741 29779 43775
rect 30205 43741 30239 43775
rect 30389 43741 30423 43775
rect 30665 43741 30699 43775
rect 32413 43741 32447 43775
rect 35265 43741 35299 43775
rect 35357 43741 35391 43775
rect 35541 43741 35575 43775
rect 35725 43741 35759 43775
rect 36093 43741 36127 43775
rect 37565 43741 37599 43775
rect 40325 43741 40359 43775
rect 3893 43673 3927 43707
rect 4261 43673 4295 43707
rect 17202 43673 17236 43707
rect 18981 43673 19015 43707
rect 19809 43673 19843 43707
rect 19993 43673 20027 43707
rect 22293 43673 22327 43707
rect 23112 43673 23146 43707
rect 25044 43673 25078 43707
rect 26249 43673 26283 43707
rect 26617 43673 26651 43707
rect 30573 43673 30607 43707
rect 32680 43673 32714 43707
rect 36338 43673 36372 43707
rect 37841 43673 37875 43707
rect 38476 43673 38510 43707
rect 40233 43673 40267 43707
rect 15301 43605 15335 43639
rect 16681 43605 16715 43639
rect 18337 43605 18371 43639
rect 21649 43605 21683 43639
rect 24593 43605 24627 43639
rect 26525 43605 26559 43639
rect 26801 43605 26835 43639
rect 27905 43605 27939 43639
rect 39589 43605 39623 43639
rect 39865 43605 39899 43639
rect 13461 43401 13495 43435
rect 15117 43401 15151 43435
rect 16313 43401 16347 43435
rect 18153 43401 18187 43435
rect 21281 43401 21315 43435
rect 21649 43401 21683 43435
rect 24133 43401 24167 43435
rect 25513 43401 25547 43435
rect 26433 43401 26467 43435
rect 27445 43401 27479 43435
rect 30389 43401 30423 43435
rect 30665 43401 30699 43435
rect 34805 43401 34839 43435
rect 35725 43401 35759 43435
rect 37657 43401 37691 43435
rect 38761 43401 38795 43435
rect 40417 43401 40451 43435
rect 13982 43333 14016 43367
rect 16926 43333 16960 43367
rect 18613 43333 18647 43367
rect 20545 43333 20579 43367
rect 20729 43333 20763 43367
rect 26985 43333 27019 43367
rect 29653 43333 29687 43367
rect 30481 43333 30515 43367
rect 33692 43333 33726 43367
rect 13645 43265 13679 43299
rect 16497 43265 16531 43299
rect 16681 43265 16715 43299
rect 18521 43265 18555 43299
rect 20361 43265 20395 43299
rect 21097 43265 21131 43299
rect 21373 43265 21407 43299
rect 21465 43265 21499 43299
rect 21649 43265 21683 43299
rect 21833 43265 21867 43299
rect 22109 43265 22143 43299
rect 23009 43265 23043 43299
rect 25697 43265 25731 43299
rect 25881 43265 25915 43299
rect 25973 43265 26007 43299
rect 26065 43265 26099 43299
rect 26249 43265 26283 43299
rect 27261 43265 27295 43299
rect 29377 43265 29411 43299
rect 29745 43265 29779 43299
rect 29838 43265 29872 43299
rect 30021 43265 30055 43299
rect 30113 43265 30147 43299
rect 30251 43265 30285 43299
rect 30757 43265 30791 43299
rect 33425 43265 33459 43299
rect 34897 43265 34931 43299
rect 35081 43265 35115 43299
rect 35449 43265 35483 43299
rect 36001 43265 36035 43299
rect 36093 43265 36127 43299
rect 36185 43265 36219 43299
rect 36369 43265 36403 43299
rect 36737 43265 36771 43299
rect 38945 43265 38979 43299
rect 39304 43265 39338 43299
rect 46489 43265 46523 43299
rect 13737 43197 13771 43231
rect 18705 43197 18739 43231
rect 21925 43197 21959 43231
rect 22661 43197 22695 43231
rect 22753 43197 22787 43231
rect 27077 43197 27111 43231
rect 29653 43197 29687 43231
rect 35173 43197 35207 43231
rect 35265 43197 35299 43231
rect 37749 43197 37783 43231
rect 37841 43197 37875 43231
rect 39037 43197 39071 43231
rect 21097 43129 21131 43163
rect 22293 43129 22327 43163
rect 29469 43129 29503 43163
rect 35633 43129 35667 43163
rect 37289 43129 37323 43163
rect 18061 43061 18095 43095
rect 21833 43061 21867 43095
rect 27077 43061 27111 43095
rect 30481 43061 30515 43095
rect 36553 43061 36587 43095
rect 46673 43061 46707 43095
rect 15485 42857 15519 42891
rect 16589 42857 16623 42891
rect 17601 42857 17635 42891
rect 22569 42857 22603 42891
rect 29929 42857 29963 42891
rect 35265 42857 35299 42891
rect 39589 42857 39623 42891
rect 30113 42789 30147 42823
rect 14105 42721 14139 42755
rect 16037 42721 16071 42755
rect 16221 42721 16255 42755
rect 17233 42721 17267 42755
rect 19717 42721 19751 42755
rect 19901 42721 19935 42755
rect 26985 42721 27019 42755
rect 29377 42721 29411 42755
rect 16957 42653 16991 42687
rect 19625 42653 19659 42687
rect 22753 42653 22787 42687
rect 27252 42653 27286 42687
rect 29561 42653 29595 42687
rect 29929 42653 29963 42687
rect 30389 42653 30423 42687
rect 31677 42653 31711 42687
rect 32781 42653 32815 42687
rect 32965 42653 32999 42687
rect 33057 42653 33091 42687
rect 35173 42653 35207 42687
rect 37473 42653 37507 42687
rect 14350 42585 14384 42619
rect 17509 42585 17543 42619
rect 29193 42585 29227 42619
rect 30205 42585 30239 42619
rect 37718 42585 37752 42619
rect 15577 42517 15611 42551
rect 15945 42517 15979 42551
rect 17049 42517 17083 42551
rect 19257 42517 19291 42551
rect 28365 42517 28399 42551
rect 30573 42517 30607 42551
rect 31493 42517 31527 42551
rect 32597 42517 32631 42551
rect 38853 42517 38887 42551
rect 13277 42313 13311 42347
rect 15853 42313 15887 42347
rect 18981 42313 19015 42347
rect 19073 42313 19107 42347
rect 31953 42313 31987 42347
rect 33517 42313 33551 42347
rect 33609 42313 33643 42347
rect 29469 42245 29503 42279
rect 30021 42245 30055 42279
rect 32404 42245 32438 42279
rect 34253 42245 34287 42279
rect 13461 42177 13495 42211
rect 13993 42177 14027 42211
rect 15669 42177 15703 42211
rect 19625 42177 19659 42211
rect 29377 42177 29411 42211
rect 29561 42177 29595 42211
rect 29929 42177 29963 42211
rect 30113 42177 30147 42211
rect 30573 42177 30607 42211
rect 30840 42177 30874 42211
rect 33885 42177 33919 42211
rect 35357 42177 35391 42211
rect 13737 42109 13771 42143
rect 19165 42109 19199 42143
rect 32137 42109 32171 42143
rect 33793 42109 33827 42143
rect 34161 42109 34195 42143
rect 35449 42109 35483 42143
rect 15117 42041 15151 42075
rect 35725 42041 35759 42075
rect 18613 41973 18647 42007
rect 19441 41973 19475 42007
rect 35541 41973 35575 42007
rect 13461 41769 13495 41803
rect 32137 41769 32171 41803
rect 34897 41769 34931 41803
rect 35173 41769 35207 41803
rect 37197 41769 37231 41803
rect 38761 41769 38795 41803
rect 20637 41701 20671 41735
rect 33149 41701 33183 41735
rect 36645 41701 36679 41735
rect 11345 41633 11379 41667
rect 17417 41633 17451 41667
rect 19257 41633 19291 41667
rect 32781 41633 32815 41667
rect 34897 41633 34931 41667
rect 35909 41633 35943 41667
rect 1409 41565 1443 41599
rect 1961 41565 1995 41599
rect 11069 41565 11103 41599
rect 13645 41565 13679 41599
rect 17141 41565 17175 41599
rect 19073 41565 19107 41599
rect 19524 41565 19558 41599
rect 20913 41565 20947 41599
rect 22109 41565 22143 41599
rect 24409 41565 24443 41599
rect 32965 41565 32999 41599
rect 34345 41565 34379 41599
rect 34529 41565 34563 41599
rect 34989 41565 35023 41599
rect 35541 41565 35575 41599
rect 35633 41565 35667 41599
rect 36001 41565 36035 41599
rect 37013 41565 37047 41599
rect 24654 41497 24688 41531
rect 31217 41497 31251 41531
rect 34713 41497 34747 41531
rect 35265 41497 35299 41531
rect 38577 41497 38611 41531
rect 1593 41429 1627 41463
rect 18889 41429 18923 41463
rect 20729 41429 20763 41463
rect 21925 41429 21959 41463
rect 25789 41429 25823 41463
rect 31493 41429 31527 41463
rect 32505 41429 32539 41463
rect 32597 41429 32631 41463
rect 34437 41429 34471 41463
rect 35725 41429 35759 41463
rect 38777 41429 38811 41463
rect 38945 41429 38979 41463
rect 23949 41225 23983 41259
rect 34989 41225 35023 41259
rect 37381 41225 37415 41259
rect 11621 41157 11655 41191
rect 19042 41157 19076 41191
rect 20536 41157 20570 41191
rect 22100 41157 22134 41191
rect 24746 41157 24780 41191
rect 36185 41157 36219 41191
rect 38945 41157 38979 41191
rect 11069 41089 11103 41123
rect 12817 41089 12851 41123
rect 12909 41089 12943 41123
rect 14464 41089 14498 41123
rect 16957 41089 16991 41123
rect 17316 41089 17350 41123
rect 18797 41089 18831 41123
rect 20269 41089 20303 41123
rect 24133 41089 24167 41123
rect 24409 41089 24443 41123
rect 33977 41089 34011 41123
rect 35265 41089 35299 41123
rect 35357 41089 35391 41123
rect 35449 41089 35483 41123
rect 35633 41089 35667 41123
rect 35725 41089 35759 41123
rect 35909 41089 35943 41123
rect 36921 41089 36955 41123
rect 37289 41089 37323 41123
rect 37657 41089 37691 41123
rect 38117 41089 38151 41123
rect 38393 41089 38427 41123
rect 38669 41089 38703 41123
rect 38853 41089 38887 41123
rect 13093 41021 13127 41055
rect 14197 41021 14231 41055
rect 17049 41021 17083 41055
rect 21833 41021 21867 41055
rect 24501 41021 24535 41055
rect 27905 41021 27939 41055
rect 28181 41021 28215 41055
rect 36645 41021 36679 41055
rect 36737 41021 36771 41055
rect 39313 41021 39347 41055
rect 39405 41021 39439 41055
rect 12449 40953 12483 40987
rect 21649 40953 21683 40987
rect 24225 40953 24259 40987
rect 36185 40953 36219 40987
rect 38485 40953 38519 40987
rect 38577 40953 38611 40987
rect 39589 40953 39623 40987
rect 10885 40885 10919 40919
rect 11713 40885 11747 40919
rect 15577 40885 15611 40919
rect 16773 40885 16807 40919
rect 18429 40885 18463 40919
rect 20177 40885 20211 40919
rect 23213 40885 23247 40919
rect 25881 40885 25915 40919
rect 34161 40885 34195 40919
rect 35725 40885 35759 40919
rect 38209 40885 38243 40919
rect 3525 40681 3559 40715
rect 12173 40681 12207 40715
rect 20177 40681 20211 40715
rect 21833 40681 21867 40715
rect 36921 40681 36955 40715
rect 39957 40681 39991 40715
rect 17785 40613 17819 40647
rect 38853 40613 38887 40647
rect 10793 40545 10827 40579
rect 14565 40545 14599 40579
rect 15853 40545 15887 40579
rect 18245 40545 18279 40579
rect 18429 40545 18463 40579
rect 20729 40545 20763 40579
rect 22477 40545 22511 40579
rect 24777 40545 24811 40579
rect 35127 40545 35161 40579
rect 36553 40545 36587 40579
rect 40141 40545 40175 40579
rect 2053 40477 2087 40511
rect 2145 40477 2179 40511
rect 8953 40477 8987 40511
rect 10701 40477 10735 40511
rect 12449 40477 12483 40511
rect 12541 40477 12575 40511
rect 14289 40477 14323 40511
rect 16313 40477 16347 40511
rect 16580 40477 16614 40511
rect 18797 40477 18831 40511
rect 20545 40477 20579 40511
rect 22201 40477 22235 40511
rect 22661 40477 22695 40511
rect 24501 40477 24535 40511
rect 25697 40477 25731 40511
rect 27353 40477 27387 40511
rect 27445 40477 27479 40511
rect 29101 40477 29135 40511
rect 30205 40477 30239 40511
rect 32965 40477 32999 40511
rect 34989 40477 35023 40511
rect 35357 40477 35391 40511
rect 35541 40477 35575 40511
rect 35817 40477 35851 40511
rect 36921 40477 36955 40511
rect 37657 40477 37691 40511
rect 37933 40477 37967 40511
rect 38117 40477 38151 40511
rect 39865 40477 39899 40511
rect 46489 40477 46523 40511
rect 2390 40409 2424 40443
rect 9198 40409 9232 40443
rect 11038 40409 11072 40443
rect 12786 40409 12820 40443
rect 15669 40409 15703 40443
rect 22928 40409 22962 40443
rect 25964 40409 25998 40443
rect 27690 40409 27724 40443
rect 30472 40409 30506 40443
rect 33232 40409 33266 40443
rect 38853 40409 38887 40443
rect 39313 40409 39347 40443
rect 1869 40341 1903 40375
rect 5825 40341 5859 40375
rect 6193 40341 6227 40375
rect 6561 40341 6595 40375
rect 6929 40341 6963 40375
rect 7205 40341 7239 40375
rect 7573 40341 7607 40375
rect 10333 40341 10367 40375
rect 10517 40341 10551 40375
rect 12265 40341 12299 40375
rect 13921 40341 13955 40375
rect 15209 40341 15243 40375
rect 15577 40341 15611 40375
rect 17693 40341 17727 40375
rect 18153 40341 18187 40375
rect 18613 40341 18647 40375
rect 20637 40341 20671 40375
rect 22293 40341 22327 40375
rect 24041 40341 24075 40375
rect 27077 40341 27111 40375
rect 27169 40341 27203 40375
rect 28825 40341 28859 40375
rect 28917 40341 28951 40375
rect 31585 40341 31619 40375
rect 34345 40341 34379 40375
rect 34989 40341 35023 40375
rect 36737 40341 36771 40375
rect 37473 40341 37507 40375
rect 39405 40341 39439 40375
rect 39589 40341 39623 40375
rect 40417 40341 40451 40375
rect 46673 40341 46707 40375
rect 2237 40137 2271 40171
rect 2605 40137 2639 40171
rect 8861 40137 8895 40171
rect 9689 40137 9723 40171
rect 11161 40137 11195 40171
rect 12909 40137 12943 40171
rect 13185 40137 13219 40171
rect 13553 40137 13587 40171
rect 14657 40137 14691 40171
rect 17325 40137 17359 40171
rect 17693 40137 17727 40171
rect 23029 40137 23063 40171
rect 24041 40137 24075 40171
rect 24869 40137 24903 40171
rect 25329 40137 25363 40171
rect 26249 40137 26283 40171
rect 26985 40137 27019 40171
rect 27353 40137 27387 40171
rect 29377 40137 29411 40171
rect 30573 40137 30607 40171
rect 30849 40137 30883 40171
rect 31217 40137 31251 40171
rect 34069 40137 34103 40171
rect 36921 40137 36955 40171
rect 38485 40137 38519 40171
rect 10057 40069 10091 40103
rect 11774 40069 11808 40103
rect 28172 40069 28206 40103
rect 33701 40069 33735 40103
rect 33793 40069 33827 40103
rect 35541 40069 35575 40103
rect 35725 40069 35759 40103
rect 37381 40069 37415 40103
rect 1409 40001 1443 40035
rect 9045 40001 9079 40035
rect 10149 40001 10183 40035
rect 11345 40001 11379 40035
rect 11529 40001 11563 40035
rect 14841 40001 14875 40035
rect 23213 40001 23247 40035
rect 24409 40001 24443 40035
rect 25237 40001 25271 40035
rect 26433 40001 26467 40035
rect 27905 40001 27939 40035
rect 29745 40001 29779 40035
rect 30757 40001 30791 40035
rect 33425 40001 33459 40035
rect 33573 40001 33607 40035
rect 33931 40001 33965 40035
rect 36185 40001 36219 40035
rect 36461 40001 36495 40035
rect 36737 40001 36771 40035
rect 38393 40001 38427 40035
rect 38577 40001 38611 40035
rect 38761 40001 38795 40035
rect 39037 40001 39071 40035
rect 39681 40001 39715 40035
rect 40233 40001 40267 40035
rect 2697 39933 2731 39967
rect 2881 39933 2915 39967
rect 10241 39933 10275 39967
rect 13645 39933 13679 39967
rect 13829 39933 13863 39967
rect 17785 39933 17819 39967
rect 17877 39933 17911 39967
rect 24501 39933 24535 39967
rect 24685 39933 24719 39967
rect 25513 39933 25547 39967
rect 27445 39933 27479 39967
rect 27537 39933 27571 39967
rect 29837 39933 29871 39967
rect 30021 39933 30055 39967
rect 31309 39933 31343 39967
rect 31401 39933 31435 39967
rect 35909 39933 35943 39967
rect 36553 39933 36587 39967
rect 39773 39933 39807 39967
rect 29285 39865 29319 39899
rect 36277 39865 36311 39899
rect 40141 39865 40175 39899
rect 1593 39797 1627 39831
rect 2053 39797 2087 39831
rect 6929 39797 6963 39831
rect 7297 39797 7331 39831
rect 7665 39797 7699 39831
rect 8033 39797 8067 39831
rect 8401 39797 8435 39831
rect 8769 39797 8803 39831
rect 9321 39797 9355 39831
rect 36737 39797 36771 39831
rect 37473 39797 37507 39831
rect 23213 39593 23247 39627
rect 27905 39593 27939 39627
rect 32413 39593 32447 39627
rect 36553 39593 36587 39627
rect 38025 39593 38059 39627
rect 39681 39593 39715 39627
rect 2053 39525 2087 39559
rect 2421 39525 2455 39559
rect 6929 39525 6963 39559
rect 11805 39525 11839 39559
rect 37105 39525 37139 39559
rect 2789 39457 2823 39491
rect 12357 39457 12391 39491
rect 23765 39457 23799 39491
rect 28365 39457 28399 39491
rect 28549 39457 28583 39491
rect 30941 39457 30975 39491
rect 32965 39457 32999 39491
rect 36185 39457 36219 39491
rect 38301 39457 38335 39491
rect 15393 39389 15427 39423
rect 23581 39389 23615 39423
rect 28273 39389 28307 39423
rect 30849 39389 30883 39423
rect 36369 39389 36403 39423
rect 36553 39389 36587 39423
rect 36829 39389 36863 39423
rect 37013 39389 37047 39423
rect 37749 39389 37783 39423
rect 14749 39321 14783 39355
rect 15660 39321 15694 39355
rect 31186 39321 31220 39355
rect 36001 39321 36035 39355
rect 37565 39321 37599 39355
rect 37841 39321 37875 39355
rect 38546 39321 38580 39355
rect 9321 39253 9355 39287
rect 12173 39253 12207 39287
rect 12265 39253 12299 39287
rect 14841 39253 14875 39287
rect 16773 39253 16807 39287
rect 23673 39253 23707 39287
rect 30665 39253 30699 39287
rect 32321 39253 32355 39287
rect 32781 39253 32815 39287
rect 32873 39253 32907 39287
rect 36737 39253 36771 39287
rect 38041 39253 38075 39287
rect 38209 39253 38243 39287
rect 34437 39049 34471 39083
rect 35541 39049 35575 39083
rect 37657 39049 37691 39083
rect 30297 38981 30331 39015
rect 31217 38981 31251 39015
rect 31401 38981 31435 39015
rect 38393 38981 38427 39015
rect 7573 38913 7607 38947
rect 9505 38913 9539 38947
rect 15117 38913 15151 38947
rect 15384 38913 15418 38947
rect 17049 38913 17083 38947
rect 17693 38913 17727 38947
rect 19533 38913 19567 38947
rect 20085 38913 20119 38947
rect 21833 38913 21867 38947
rect 22100 38913 22134 38947
rect 24501 38913 24535 38947
rect 30205 38913 30239 38947
rect 33324 38913 33358 38947
rect 34713 38913 34747 38947
rect 34805 38913 34839 38947
rect 34897 38913 34931 38947
rect 35015 38913 35049 38947
rect 35173 38913 35207 38947
rect 35725 38913 35759 38947
rect 36185 38913 36219 38947
rect 36461 38913 36495 38947
rect 36829 38913 36863 38947
rect 37289 38913 37323 38947
rect 37473 38913 37507 38947
rect 37565 38913 37599 38947
rect 37749 38913 37783 38947
rect 17141 38845 17175 38879
rect 17325 38845 17359 38879
rect 20177 38845 20211 38879
rect 20269 38845 20303 38879
rect 24593 38845 24627 38879
rect 24777 38845 24811 38879
rect 30481 38845 30515 38879
rect 33057 38845 33091 38879
rect 16497 38777 16531 38811
rect 17509 38777 17543 38811
rect 7389 38709 7423 38743
rect 9321 38709 9355 38743
rect 16681 38709 16715 38743
rect 19349 38709 19383 38743
rect 19717 38709 19751 38743
rect 23213 38709 23247 38743
rect 24133 38709 24167 38743
rect 29837 38709 29871 38743
rect 34529 38709 34563 38743
rect 37289 38709 37323 38743
rect 38485 38709 38519 38743
rect 16037 38505 16071 38539
rect 16405 38505 16439 38539
rect 20637 38505 20671 38539
rect 25789 38505 25823 38539
rect 30941 38505 30975 38539
rect 35541 38505 35575 38539
rect 39313 38505 39347 38539
rect 33517 38437 33551 38471
rect 14105 38369 14139 38403
rect 16957 38369 16991 38403
rect 17233 38369 17267 38403
rect 17877 38369 17911 38403
rect 18153 38369 18187 38403
rect 18270 38369 18304 38403
rect 21189 38369 21223 38403
rect 21833 38369 21867 38403
rect 22109 38369 22143 38403
rect 23581 38369 23615 38403
rect 23765 38369 23799 38403
rect 24409 38369 24443 38403
rect 28365 38369 28399 38403
rect 29561 38369 29595 38403
rect 31677 38369 31711 38403
rect 34437 38369 34471 38403
rect 35173 38369 35207 38403
rect 37105 38369 37139 38403
rect 37197 38369 37231 38403
rect 37289 38369 37323 38403
rect 37381 38369 37415 38403
rect 4353 38301 4387 38335
rect 5641 38301 5675 38335
rect 7113 38301 7147 38335
rect 7380 38301 7414 38335
rect 9045 38301 9079 38335
rect 9312 38301 9346 38335
rect 11161 38301 11195 38335
rect 12817 38301 12851 38335
rect 13645 38301 13679 38335
rect 13921 38301 13955 38335
rect 16221 38301 16255 38335
rect 16773 38301 16807 38335
rect 17417 38301 17451 38335
rect 18429 38301 18463 38335
rect 19257 38301 19291 38335
rect 20913 38301 20947 38335
rect 21373 38301 21407 38335
rect 22226 38301 22260 38335
rect 22385 38301 22419 38335
rect 23489 38301 23523 38335
rect 24133 38301 24167 38335
rect 26341 38301 26375 38335
rect 31585 38301 31619 38335
rect 33609 38301 33643 38335
rect 33977 38301 34011 38335
rect 35081 38301 35115 38335
rect 35265 38301 35299 38335
rect 35449 38301 35483 38335
rect 35909 38301 35943 38335
rect 37933 38301 37967 38335
rect 5908 38233 5942 38267
rect 11428 38233 11462 38267
rect 14350 38233 14384 38267
rect 19524 38233 19558 38267
rect 24654 38233 24688 38267
rect 26608 38233 26642 38267
rect 28273 38233 28307 38267
rect 29828 38233 29862 38267
rect 31922 38233 31956 38267
rect 36645 38233 36679 38267
rect 38178 38233 38212 38267
rect 4169 38165 4203 38199
rect 7021 38165 7055 38199
rect 8493 38165 8527 38199
rect 10425 38165 10459 38199
rect 12541 38165 12575 38199
rect 12633 38165 12667 38199
rect 13461 38165 13495 38199
rect 13737 38165 13771 38199
rect 15485 38165 15519 38199
rect 16865 38165 16899 38199
rect 19073 38165 19107 38199
rect 20729 38165 20763 38199
rect 23029 38165 23063 38199
rect 23121 38165 23155 38199
rect 23949 38165 23983 38199
rect 27721 38165 27755 38199
rect 27813 38165 27847 38199
rect 28181 38165 28215 38199
rect 31401 38165 31435 38199
rect 33057 38165 33091 38199
rect 36921 38165 36955 38199
rect 6009 37961 6043 37995
rect 10517 37961 10551 37995
rect 10885 37961 10919 37995
rect 10977 37961 11011 37995
rect 15025 37961 15059 37995
rect 15393 37961 15427 37995
rect 21005 37961 21039 37995
rect 26525 37961 26559 37995
rect 29745 37961 29779 37995
rect 30665 37961 30699 37995
rect 32137 37961 32171 37995
rect 32505 37961 32539 37995
rect 32597 37961 32631 37995
rect 33333 37961 33367 37995
rect 37489 37961 37523 37995
rect 39589 37961 39623 37995
rect 4068 37893 4102 37927
rect 19340 37893 19374 37927
rect 20913 37893 20947 37927
rect 33241 37893 33275 37927
rect 37289 37893 37323 37927
rect 38454 37893 38488 37927
rect 3709 37825 3743 37859
rect 3801 37825 3835 37859
rect 6193 37825 6227 37859
rect 6633 37825 6667 37859
rect 8585 37825 8619 37859
rect 8769 37825 8803 37859
rect 9622 37825 9656 37859
rect 11713 37825 11747 37859
rect 12449 37825 12483 37859
rect 13553 37825 13587 37859
rect 13820 37825 13854 37859
rect 16957 37825 16991 37859
rect 17141 37825 17175 37859
rect 17877 37825 17911 37859
rect 17994 37825 18028 37859
rect 19073 37825 19107 37859
rect 21649 37825 21683 37859
rect 21833 37825 21867 37859
rect 22753 37825 22787 37859
rect 24409 37825 24443 37859
rect 25329 37825 25363 37859
rect 26709 37825 26743 37859
rect 27261 37825 27295 37859
rect 27629 37825 27663 37859
rect 29929 37825 29963 37859
rect 30573 37825 30607 37859
rect 36461 37825 36495 37859
rect 36553 37825 36587 37859
rect 36645 37825 36679 37859
rect 36829 37825 36863 37859
rect 46489 37825 46523 37859
rect 6377 37757 6411 37791
rect 9505 37757 9539 37791
rect 9781 37757 9815 37791
rect 11069 37757 11103 37791
rect 11529 37757 11563 37791
rect 12566 37757 12600 37791
rect 12725 37757 12759 37791
rect 15485 37757 15519 37791
rect 15669 37757 15703 37791
rect 17601 37757 17635 37791
rect 18153 37757 18187 37791
rect 22017 37757 22051 37791
rect 22870 37757 22904 37791
rect 23029 37757 23063 37791
rect 24593 37757 24627 37791
rect 25446 37757 25480 37791
rect 25605 37757 25639 37791
rect 27813 37757 27847 37791
rect 28549 37757 28583 37791
rect 28687 37757 28721 37791
rect 28825 37757 28859 37791
rect 30849 37757 30883 37791
rect 32689 37757 32723 37791
rect 38209 37757 38243 37791
rect 7757 37689 7791 37723
rect 9229 37689 9263 37723
rect 12173 37689 12207 37723
rect 21465 37689 21499 37723
rect 22477 37689 22511 37723
rect 25053 37689 25087 37723
rect 28273 37689 28307 37723
rect 3525 37621 3559 37655
rect 5181 37621 5215 37655
rect 10425 37621 10459 37655
rect 13369 37621 13403 37655
rect 14933 37621 14967 37655
rect 18797 37621 18831 37655
rect 20453 37621 20487 37655
rect 23673 37621 23707 37655
rect 26249 37621 26283 37655
rect 27077 37621 27111 37655
rect 29469 37621 29503 37655
rect 30205 37621 30239 37655
rect 36185 37621 36219 37655
rect 37473 37621 37507 37655
rect 37657 37621 37691 37655
rect 46673 37621 46707 37655
rect 5273 37417 5307 37451
rect 10793 37417 10827 37451
rect 13185 37417 13219 37451
rect 14289 37417 14323 37451
rect 26525 37417 26559 37451
rect 31401 37417 31435 37451
rect 6285 37349 6319 37383
rect 6653 37349 6687 37383
rect 11897 37349 11931 37383
rect 3801 37281 3835 37315
rect 5917 37281 5951 37315
rect 7205 37281 7239 37315
rect 8217 37281 8251 37315
rect 8953 37281 8987 37315
rect 9597 37281 9631 37315
rect 9873 37281 9907 37315
rect 9990 37281 10024 37315
rect 11253 37281 11287 37315
rect 12173 37281 12207 37315
rect 12290 37281 12324 37315
rect 13093 37281 13127 37315
rect 13737 37281 13771 37315
rect 14841 37281 14875 37315
rect 20177 37281 20211 37315
rect 24409 37281 24443 37315
rect 24593 37281 24627 37315
rect 25053 37281 25087 37315
rect 25329 37281 25363 37315
rect 25446 37281 25480 37315
rect 26249 37281 26283 37315
rect 27077 37281 27111 37315
rect 27997 37281 28031 37315
rect 28273 37281 28307 37315
rect 28390 37281 28424 37315
rect 29193 37281 29227 37315
rect 33977 37281 34011 37315
rect 38945 37281 38979 37315
rect 1593 37213 1627 37247
rect 4068 37213 4102 37247
rect 5641 37213 5675 37247
rect 6469 37213 6503 37247
rect 7021 37213 7055 37247
rect 8033 37213 8067 37247
rect 9137 37213 9171 37247
rect 10149 37213 10183 37247
rect 11437 37213 11471 37247
rect 12449 37213 12483 37247
rect 14657 37213 14691 37247
rect 19901 37213 19935 37247
rect 25605 37213 25639 37247
rect 27353 37213 27387 37247
rect 27537 37213 27571 37247
rect 28549 37213 28583 37247
rect 29929 37213 29963 37247
rect 30021 37213 30055 37247
rect 33793 37213 33827 37247
rect 34713 37213 34747 37247
rect 36461 37213 36495 37247
rect 36737 37213 36771 37247
rect 39405 37213 39439 37247
rect 7113 37145 7147 37179
rect 19993 37145 20027 37179
rect 26893 37145 26927 37179
rect 30266 37145 30300 37179
rect 34958 37145 34992 37179
rect 36645 37145 36679 37179
rect 1409 37077 1443 37111
rect 5181 37077 5215 37111
rect 5733 37077 5767 37111
rect 7665 37077 7699 37111
rect 8125 37077 8159 37111
rect 13553 37077 13587 37111
rect 13645 37077 13679 37111
rect 14749 37077 14783 37111
rect 19533 37077 19567 37111
rect 26985 37077 27019 37111
rect 29745 37077 29779 37111
rect 36093 37077 36127 37111
rect 36559 37077 36593 37111
rect 38393 37077 38427 37111
rect 38761 37077 38795 37111
rect 38853 37077 38887 37111
rect 39221 37077 39255 37111
rect 4077 36873 4111 36907
rect 4445 36873 4479 36907
rect 4537 36873 4571 36907
rect 6653 36873 6687 36907
rect 7021 36873 7055 36907
rect 16681 36873 16715 36907
rect 17141 36873 17175 36907
rect 28365 36873 28399 36907
rect 34529 36873 34563 36907
rect 36553 36873 36587 36907
rect 40233 36873 40267 36907
rect 7113 36805 7147 36839
rect 27230 36805 27264 36839
rect 30113 36805 30147 36839
rect 30297 36805 30331 36839
rect 35173 36805 35207 36839
rect 39120 36805 39154 36839
rect 16505 36741 16539 36775
rect 17049 36737 17083 36771
rect 23121 36737 23155 36771
rect 26985 36737 27019 36771
rect 32597 36737 32631 36771
rect 32864 36737 32898 36771
rect 34805 36737 34839 36771
rect 36093 36737 36127 36771
rect 36369 36737 36403 36771
rect 38853 36737 38887 36771
rect 4721 36669 4755 36703
rect 7297 36669 7331 36703
rect 17325 36669 17359 36703
rect 19257 36669 19291 36703
rect 23305 36669 23339 36703
rect 34713 36669 34747 36703
rect 35081 36669 35115 36703
rect 19533 36601 19567 36635
rect 36185 36601 36219 36635
rect 16313 36533 16347 36567
rect 19717 36533 19751 36567
rect 33977 36533 34011 36567
rect 17509 36329 17543 36363
rect 29745 36329 29779 36363
rect 34713 36329 34747 36363
rect 36737 36329 36771 36363
rect 37289 36329 37323 36363
rect 18705 36261 18739 36295
rect 20269 36261 20303 36295
rect 21649 36261 21683 36295
rect 23029 36261 23063 36295
rect 23673 36261 23707 36295
rect 2513 36193 2547 36227
rect 4445 36193 4479 36227
rect 10057 36193 10091 36227
rect 11253 36193 11287 36227
rect 15761 36193 15795 36227
rect 16221 36193 16255 36227
rect 16614 36193 16648 36227
rect 16773 36193 16807 36227
rect 18153 36193 18187 36227
rect 19717 36193 19751 36227
rect 22569 36193 22603 36227
rect 22753 36193 22787 36227
rect 31953 36193 31987 36227
rect 32413 36193 32447 36227
rect 32689 36193 32723 36227
rect 32827 36193 32861 36227
rect 34253 36193 34287 36227
rect 2237 36125 2271 36159
rect 4261 36125 4295 36159
rect 9781 36125 9815 36159
rect 15577 36125 15611 36159
rect 16497 36125 16531 36159
rect 18337 36125 18371 36159
rect 19901 36125 19935 36159
rect 20177 36125 20211 36159
rect 20453 36125 20487 36159
rect 20729 36125 20763 36159
rect 21833 36125 21867 36159
rect 22385 36125 22419 36159
rect 29285 36125 29319 36159
rect 31769 36125 31803 36159
rect 32965 36125 32999 36159
rect 34897 36125 34931 36159
rect 35817 36125 35851 36159
rect 36001 36125 36035 36159
rect 36277 36125 36311 36159
rect 36553 36125 36587 36159
rect 36829 36125 36863 36159
rect 37105 36125 37139 36159
rect 37381 36125 37415 36159
rect 14197 36057 14231 36091
rect 17417 36057 17451 36091
rect 17877 36057 17911 36091
rect 20085 36057 20119 36091
rect 23305 36057 23339 36091
rect 29653 36057 29687 36091
rect 34069 36057 34103 36091
rect 35909 36057 35943 36091
rect 3801 35989 3835 36023
rect 4169 35989 4203 36023
rect 10701 35989 10735 36023
rect 11069 35989 11103 36023
rect 11161 35989 11195 36023
rect 14289 35989 14323 36023
rect 17969 35989 18003 36023
rect 18797 35989 18831 36023
rect 20637 35989 20671 36023
rect 21925 35989 21959 36023
rect 22293 35989 22327 36023
rect 23213 35989 23247 36023
rect 23765 35989 23799 36023
rect 29101 35989 29135 36023
rect 33609 35989 33643 36023
rect 33701 35989 33735 36023
rect 34161 35989 34195 36023
rect 36093 35989 36127 36023
rect 36369 35989 36403 36023
rect 36921 35989 36955 36023
rect 1869 35785 1903 35819
rect 3525 35785 3559 35819
rect 7113 35785 7147 35819
rect 13461 35785 13495 35819
rect 18061 35785 18095 35819
rect 20913 35785 20947 35819
rect 21373 35785 21407 35819
rect 23213 35785 23247 35819
rect 30389 35785 30423 35819
rect 30849 35785 30883 35819
rect 33977 35785 34011 35819
rect 37105 35785 37139 35819
rect 2390 35717 2424 35751
rect 7573 35717 7607 35751
rect 9934 35717 9968 35751
rect 22100 35717 22134 35751
rect 23765 35717 23799 35751
rect 35992 35717 36026 35751
rect 2053 35649 2087 35683
rect 3801 35649 3835 35683
rect 4261 35649 4295 35683
rect 5298 35649 5332 35683
rect 7021 35649 7055 35683
rect 7481 35649 7515 35683
rect 8401 35649 8435 35683
rect 9597 35649 9631 35683
rect 13277 35649 13311 35683
rect 13553 35649 13587 35683
rect 14657 35649 14691 35683
rect 15577 35649 15611 35683
rect 15694 35649 15728 35683
rect 16681 35649 16715 35683
rect 16937 35649 16971 35683
rect 18245 35649 18279 35683
rect 19349 35649 19383 35683
rect 19441 35649 19475 35683
rect 19717 35649 19751 35683
rect 19993 35649 20027 35683
rect 20177 35649 20211 35683
rect 20269 35649 20303 35683
rect 20821 35649 20855 35683
rect 21281 35649 21315 35683
rect 23673 35649 23707 35683
rect 25053 35649 25087 35683
rect 27169 35649 27203 35683
rect 27261 35649 27295 35683
rect 27537 35649 27571 35683
rect 28457 35649 28491 35683
rect 29009 35649 29043 35683
rect 29276 35649 29310 35683
rect 30941 35649 30975 35683
rect 32137 35649 32171 35683
rect 32321 35649 32355 35683
rect 33174 35649 33208 35683
rect 40049 35649 40083 35683
rect 46489 35649 46523 35683
rect 2145 35581 2179 35615
rect 4445 35581 4479 35615
rect 4905 35581 4939 35615
rect 5181 35581 5215 35615
rect 5457 35581 5491 35615
rect 7665 35581 7699 35615
rect 9689 35581 9723 35615
rect 13737 35581 13771 35615
rect 14841 35581 14875 35615
rect 15853 35581 15887 35615
rect 18521 35581 18555 35615
rect 19165 35581 19199 35615
rect 21465 35581 21499 35615
rect 21833 35581 21867 35615
rect 23857 35581 23891 35615
rect 24133 35581 24167 35615
rect 24317 35581 24351 35615
rect 25191 35581 25225 35615
rect 25329 35581 25363 35615
rect 26157 35581 26191 35615
rect 26617 35581 26651 35615
rect 26985 35581 27019 35615
rect 31125 35581 31159 35615
rect 33057 35581 33091 35615
rect 33333 35581 33367 35615
rect 35725 35581 35759 35615
rect 39773 35581 39807 35615
rect 14105 35513 14139 35547
rect 15301 35513 15335 35547
rect 19625 35513 19659 35547
rect 24777 35513 24811 35547
rect 26433 35513 26467 35547
rect 27445 35513 27479 35547
rect 28825 35513 28859 35547
rect 32781 35513 32815 35547
rect 3617 35445 3651 35479
rect 6101 35445 6135 35479
rect 6837 35445 6871 35479
rect 8217 35445 8251 35479
rect 9413 35445 9447 35479
rect 11069 35445 11103 35479
rect 13093 35445 13127 35479
rect 14197 35445 14231 35479
rect 16497 35445 16531 35479
rect 19809 35445 19843 35479
rect 20637 35445 20671 35479
rect 23305 35445 23339 35479
rect 25973 35445 26007 35479
rect 28917 35445 28951 35479
rect 30481 35445 30515 35479
rect 40785 35445 40819 35479
rect 46673 35445 46707 35479
rect 8953 35241 8987 35275
rect 11897 35241 11931 35275
rect 14565 35241 14599 35275
rect 23489 35241 23523 35275
rect 27537 35241 27571 35275
rect 29561 35241 29595 35275
rect 37381 35241 37415 35275
rect 3525 35173 3559 35207
rect 7941 35173 7975 35207
rect 10707 35173 10741 35207
rect 12633 35173 12667 35207
rect 19625 35173 19659 35207
rect 20361 35173 20395 35207
rect 22201 35173 22235 35207
rect 26249 35173 26283 35207
rect 26617 35173 26651 35207
rect 27169 35173 27203 35207
rect 27353 35173 27387 35207
rect 4261 35105 4295 35139
rect 4905 35105 4939 35139
rect 5181 35105 5215 35139
rect 5298 35105 5332 35139
rect 5457 35105 5491 35139
rect 6101 35105 6135 35139
rect 8585 35105 8619 35139
rect 9505 35105 9539 35139
rect 11094 35105 11128 35139
rect 12357 35105 12391 35139
rect 20821 35105 20855 35139
rect 24409 35105 24443 35139
rect 25053 35105 25087 35139
rect 29285 35105 29319 35139
rect 30573 35105 30607 35139
rect 30849 35105 30883 35139
rect 30966 35105 31000 35139
rect 2145 35037 2179 35071
rect 2412 35037 2446 35071
rect 4445 35037 4479 35071
rect 6469 35037 6503 35071
rect 6561 35037 6595 35071
rect 6828 35037 6862 35071
rect 9321 35037 9355 35071
rect 10057 35037 10091 35071
rect 10241 35037 10275 35071
rect 10977 35037 11011 35071
rect 11253 35037 11287 35071
rect 12449 35037 12483 35071
rect 13553 35037 13587 35071
rect 13645 35037 13679 35071
rect 13829 35037 13863 35071
rect 14289 35037 14323 35071
rect 14381 35037 14415 35071
rect 14657 35037 14691 35071
rect 17693 35037 17727 35071
rect 19441 35037 19475 35071
rect 21077 35037 21111 35071
rect 23213 35037 23247 35071
rect 23305 35037 23339 35071
rect 23581 35037 23615 35071
rect 24041 35037 24075 35071
rect 24593 35037 24627 35071
rect 25329 35037 25363 35071
rect 25446 35037 25480 35071
rect 25605 35037 25639 35071
rect 26893 35037 26927 35071
rect 27721 35037 27755 35071
rect 27905 35037 27939 35071
rect 27997 35037 28031 35071
rect 28825 35037 28859 35071
rect 29009 35037 29043 35071
rect 29101 35037 29135 35071
rect 29377 35037 29411 35071
rect 29745 35037 29779 35071
rect 29929 35037 29963 35071
rect 30113 35037 30147 35071
rect 31125 35037 31159 35071
rect 34253 35037 34287 35071
rect 34713 35037 34747 35071
rect 34989 35037 35023 35071
rect 36001 35037 36035 35071
rect 36268 35037 36302 35071
rect 39221 35037 39255 35071
rect 39865 35037 39899 35071
rect 40141 35037 40175 35071
rect 8401 34969 8435 35003
rect 14105 34969 14139 35003
rect 17960 34969 17994 35003
rect 20177 34969 20211 35003
rect 26341 34969 26375 35003
rect 38301 34969 38335 35003
rect 6285 34901 6319 34935
rect 8033 34901 8067 34935
rect 8493 34901 8527 34935
rect 9413 34901 9447 34935
rect 11989 34901 12023 34935
rect 13185 34901 13219 34935
rect 19073 34901 19107 34935
rect 23029 34901 23063 34935
rect 23857 34901 23891 34935
rect 26801 34901 26835 34935
rect 31769 34901 31803 34935
rect 34437 34901 34471 34935
rect 35725 34901 35759 34935
rect 38393 34901 38427 34935
rect 39313 34901 39347 34935
rect 40877 34901 40911 34935
rect 3065 34697 3099 34731
rect 7941 34697 7975 34731
rect 9413 34697 9447 34731
rect 11345 34697 11379 34731
rect 14473 34697 14507 34731
rect 14933 34697 14967 34731
rect 16129 34697 16163 34731
rect 25237 34697 25271 34731
rect 25605 34697 25639 34731
rect 28549 34697 28583 34731
rect 29377 34697 29411 34731
rect 29745 34697 29779 34731
rect 31769 34697 31803 34731
rect 35449 34697 35483 34731
rect 37749 34697 37783 34731
rect 39497 34697 39531 34731
rect 40601 34697 40635 34731
rect 1501 34629 1535 34663
rect 3433 34629 3467 34663
rect 3525 34629 3559 34663
rect 6806 34629 6840 34663
rect 12357 34629 12391 34663
rect 16926 34629 16960 34663
rect 18245 34629 18279 34663
rect 19441 34629 19475 34663
rect 29009 34629 29043 34663
rect 37381 34629 37415 34663
rect 38362 34629 38396 34663
rect 6561 34561 6595 34595
rect 8300 34561 8334 34595
rect 9505 34561 9539 34595
rect 9689 34561 9723 34595
rect 10425 34561 10459 34595
rect 12081 34561 12115 34595
rect 13360 34561 13394 34595
rect 15025 34561 15059 34595
rect 16313 34561 16347 34595
rect 18429 34561 18463 34595
rect 23940 34561 23974 34595
rect 25697 34561 25731 34595
rect 27629 34561 27663 34595
rect 27721 34561 27755 34595
rect 27997 34561 28031 34595
rect 28089 34561 28123 34595
rect 28825 34561 28859 34595
rect 29101 34561 29135 34595
rect 29561 34561 29595 34595
rect 29837 34561 29871 34595
rect 29929 34561 29963 34595
rect 30849 34561 30883 34595
rect 30966 34561 31000 34595
rect 34713 34561 34747 34595
rect 35633 34561 35667 34595
rect 37565 34561 37599 34595
rect 37841 34561 37875 34595
rect 39589 34561 39623 34595
rect 39865 34561 39899 34595
rect 41245 34561 41279 34595
rect 41797 34561 41831 34595
rect 42533 34561 42567 34595
rect 43361 34561 43395 34595
rect 3617 34493 3651 34527
rect 8033 34493 8067 34527
rect 10149 34493 10183 34527
rect 10542 34493 10576 34527
rect 10701 34493 10735 34527
rect 11713 34493 11747 34527
rect 12173 34493 12207 34527
rect 13093 34493 13127 34527
rect 15117 34493 15151 34527
rect 16681 34493 16715 34527
rect 19533 34493 19567 34527
rect 19717 34493 19751 34527
rect 23673 34493 23707 34527
rect 25789 34493 25823 34527
rect 27445 34493 27479 34527
rect 28641 34493 28675 34527
rect 30113 34493 30147 34527
rect 30573 34493 30607 34527
rect 31125 34493 31159 34527
rect 34437 34493 34471 34527
rect 35817 34493 35851 34527
rect 38117 34493 38151 34527
rect 41521 34493 41555 34527
rect 25053 34425 25087 34459
rect 28457 34425 28491 34459
rect 42165 34425 42199 34459
rect 42257 34425 42291 34459
rect 1593 34357 1627 34391
rect 14565 34357 14599 34391
rect 18061 34357 18095 34391
rect 19073 34357 19107 34391
rect 27905 34357 27939 34391
rect 41613 34357 41647 34391
rect 42625 34357 42659 34391
rect 43453 34357 43487 34391
rect 43821 34357 43855 34391
rect 13369 34153 13403 34187
rect 16313 34153 16347 34187
rect 18337 34153 18371 34187
rect 36093 34153 36127 34187
rect 21005 34085 21039 34119
rect 42257 34085 42291 34119
rect 45017 34085 45051 34119
rect 5089 34017 5123 34051
rect 16865 34017 16899 34051
rect 4905 33949 4939 33983
rect 13553 33949 13587 33983
rect 16681 33949 16715 33983
rect 18521 33949 18555 33983
rect 21281 33949 21315 33983
rect 21925 33949 21959 33983
rect 31677 33949 31711 33983
rect 31769 33949 31803 33983
rect 34253 33949 34287 33983
rect 34529 33949 34563 33983
rect 34713 33949 34747 33983
rect 37381 33949 37415 33983
rect 37657 33949 37691 33983
rect 37841 33949 37875 33983
rect 40969 33949 41003 33983
rect 41061 33949 41095 33983
rect 43177 33949 43211 33983
rect 43361 33949 43395 33983
rect 45293 33949 45327 33983
rect 4813 33881 4847 33915
rect 20821 33881 20855 33915
rect 21557 33881 21591 33915
rect 32014 33881 32048 33915
rect 34069 33881 34103 33915
rect 34958 33881 34992 33915
rect 41981 33881 42015 33915
rect 45017 33881 45051 33915
rect 4445 33813 4479 33847
rect 16773 33813 16807 33847
rect 22109 33813 22143 33847
rect 31493 33813 31527 33847
rect 33149 33813 33183 33847
rect 34437 33813 34471 33847
rect 37197 33813 37231 33847
rect 41245 33813 41279 33847
rect 42441 33813 42475 33847
rect 43269 33813 43303 33847
rect 45201 33813 45235 33847
rect 2605 33609 2639 33643
rect 3065 33609 3099 33643
rect 3709 33609 3743 33643
rect 5365 33609 5399 33643
rect 24317 33609 24351 33643
rect 32137 33609 32171 33643
rect 32505 33609 32539 33643
rect 41613 33609 41647 33643
rect 41797 33609 41831 33643
rect 46213 33609 46247 33643
rect 4230 33541 4264 33575
rect 13093 33541 13127 33575
rect 18981 33541 19015 33575
rect 37810 33541 37844 33575
rect 45385 33541 45419 33575
rect 2421 33473 2455 33507
rect 2973 33473 3007 33507
rect 3893 33473 3927 33507
rect 3985 33473 4019 33507
rect 9413 33473 9447 33507
rect 12449 33473 12483 33507
rect 13001 33473 13035 33507
rect 18797 33473 18831 33507
rect 22293 33473 22327 33507
rect 22560 33473 22594 33507
rect 24133 33473 24167 33507
rect 24501 33473 24535 33507
rect 25421 33473 25455 33507
rect 25688 33473 25722 33507
rect 34713 33473 34747 33507
rect 37565 33473 37599 33507
rect 39313 33473 39347 33507
rect 39405 33473 39439 33507
rect 40325 33473 40359 33507
rect 40785 33473 40819 33507
rect 40877 33473 40911 33507
rect 41337 33473 41371 33507
rect 41705 33473 41739 33507
rect 42073 33473 42107 33507
rect 42165 33473 42199 33507
rect 42717 33473 42751 33507
rect 42809 33473 42843 33507
rect 42901 33473 42935 33507
rect 43085 33473 43119 33507
rect 43913 33473 43947 33507
rect 44189 33473 44223 33507
rect 44465 33473 44499 33507
rect 44557 33473 44591 33507
rect 44925 33473 44959 33507
rect 45017 33473 45051 33507
rect 45110 33473 45144 33507
rect 45293 33473 45327 33507
rect 45482 33473 45516 33507
rect 45753 33473 45787 33507
rect 46489 33473 46523 33507
rect 3157 33405 3191 33439
rect 9689 33405 9723 33439
rect 13185 33405 13219 33439
rect 24777 33405 24811 33439
rect 32597 33405 32631 33439
rect 32781 33405 32815 33439
rect 34437 33405 34471 33439
rect 39589 33405 39623 33439
rect 41889 33405 41923 33439
rect 46305 33405 46339 33439
rect 12633 33337 12667 33371
rect 39129 33337 39163 33371
rect 40141 33337 40175 33371
rect 44005 33337 44039 33371
rect 45661 33337 45695 33371
rect 2237 33269 2271 33303
rect 12265 33269 12299 33303
rect 18613 33269 18647 33303
rect 19073 33269 19107 33303
rect 23673 33269 23707 33303
rect 26801 33269 26835 33303
rect 35449 33269 35483 33303
rect 38945 33269 38979 33303
rect 40049 33269 40083 33303
rect 41153 33269 41187 33303
rect 41245 33269 41279 33303
rect 42441 33269 42475 33303
rect 45845 33269 45879 33303
rect 46673 33269 46707 33303
rect 3157 33065 3191 33099
rect 13277 33065 13311 33099
rect 16037 33065 16071 33099
rect 23213 33065 23247 33099
rect 26065 33065 26099 33099
rect 38669 33065 38703 33099
rect 38945 33065 38979 33099
rect 41061 33065 41095 33099
rect 44373 33065 44407 33099
rect 45109 33065 45143 33099
rect 45477 33065 45511 33099
rect 46029 33065 46063 33099
rect 4721 32997 4755 33031
rect 7021 32997 7055 33031
rect 18061 32997 18095 33031
rect 26341 32997 26375 33031
rect 37197 32997 37231 33031
rect 41613 32997 41647 33031
rect 42533 32997 42567 33031
rect 45845 32997 45879 33031
rect 4077 32929 4111 32963
rect 5114 32929 5148 32963
rect 5273 32929 5307 32963
rect 7665 32929 7699 32963
rect 8401 32929 8435 32963
rect 14197 32929 14231 32963
rect 14841 32929 14875 32963
rect 15117 32929 15151 32963
rect 16957 32929 16991 32963
rect 17785 32929 17819 32963
rect 18889 32929 18923 32963
rect 21189 32929 21223 32963
rect 21373 32929 21407 32963
rect 22937 32929 22971 32963
rect 26801 32929 26835 32963
rect 26985 32929 27019 32963
rect 30021 32929 30055 32963
rect 30113 32929 30147 32963
rect 36829 32929 36863 32963
rect 40877 32929 40911 32963
rect 41981 32929 42015 32963
rect 1685 32861 1719 32895
rect 1777 32861 1811 32895
rect 2044 32861 2078 32895
rect 4261 32861 4295 32895
rect 4997 32861 5031 32895
rect 6929 32861 6963 32895
rect 9229 32861 9263 32895
rect 9321 32861 9355 32895
rect 11897 32861 11931 32895
rect 12164 32861 12198 32895
rect 14381 32861 14415 32895
rect 15234 32861 15268 32895
rect 15393 32861 15427 32895
rect 18245 32861 18279 32895
rect 19257 32861 19291 32895
rect 19513 32861 19547 32895
rect 23397 32861 23431 32895
rect 24501 32861 24535 32895
rect 26249 32861 26283 32895
rect 26709 32861 26743 32895
rect 29377 32861 29411 32895
rect 32137 32861 32171 32895
rect 32229 32861 32263 32895
rect 35725 32861 35759 32895
rect 36001 32861 36035 32895
rect 38485 32861 38519 32895
rect 40969 32861 41003 32895
rect 41153 32861 41187 32895
rect 41797 32861 41831 32895
rect 41890 32861 41924 32895
rect 42073 32861 42107 32895
rect 42257 32861 42291 32895
rect 42441 32861 42475 32895
rect 42717 32861 42751 32895
rect 42809 32861 42843 32895
rect 44281 32861 44315 32895
rect 45017 32861 45051 32895
rect 46489 32861 46523 32895
rect 5917 32793 5951 32827
rect 7481 32793 7515 32827
rect 9566 32793 9600 32827
rect 16773 32793 16807 32827
rect 17601 32793 17635 32827
rect 22845 32793 22879 32827
rect 24768 32793 24802 32827
rect 32485 32793 32519 32827
rect 38117 32793 38151 32827
rect 38301 32793 38335 32827
rect 40509 32793 40543 32827
rect 40693 32793 40727 32827
rect 42533 32793 42567 32827
rect 44649 32793 44683 32827
rect 45569 32793 45603 32827
rect 1501 32725 1535 32759
rect 6745 32725 6779 32759
rect 7389 32725 7423 32759
rect 7849 32725 7883 32759
rect 8217 32725 8251 32759
rect 8309 32725 8343 32759
rect 9045 32725 9079 32759
rect 10701 32725 10735 32759
rect 17233 32725 17267 32759
rect 17693 32725 17727 32759
rect 18337 32725 18371 32759
rect 18705 32725 18739 32759
rect 18797 32725 18831 32759
rect 20637 32725 20671 32759
rect 20729 32725 20763 32759
rect 21097 32725 21131 32759
rect 22385 32725 22419 32759
rect 22753 32725 22787 32759
rect 25881 32725 25915 32759
rect 29193 32725 29227 32759
rect 29561 32725 29595 32759
rect 29929 32725 29963 32759
rect 31953 32725 31987 32759
rect 33609 32725 33643 32759
rect 36737 32725 36771 32759
rect 37289 32725 37323 32759
rect 42441 32725 42475 32759
rect 44741 32725 44775 32759
rect 46673 32725 46707 32759
rect 3157 32521 3191 32555
rect 3525 32521 3559 32555
rect 5917 32521 5951 32555
rect 7757 32521 7791 32555
rect 11529 32521 11563 32555
rect 13185 32521 13219 32555
rect 15761 32521 15795 32555
rect 18061 32521 18095 32555
rect 18613 32521 18647 32555
rect 20821 32521 20855 32555
rect 24777 32521 24811 32555
rect 25421 32521 25455 32555
rect 30389 32521 30423 32555
rect 30757 32521 30791 32555
rect 32137 32521 32171 32555
rect 32505 32521 32539 32555
rect 42441 32521 42475 32555
rect 44833 32521 44867 32555
rect 1930 32453 1964 32487
rect 3617 32453 3651 32487
rect 6644 32453 6678 32487
rect 16926 32453 16960 32487
rect 25513 32453 25547 32487
rect 32597 32453 32631 32487
rect 36645 32453 36679 32487
rect 40785 32453 40819 32487
rect 43177 32453 43211 32487
rect 44465 32453 44499 32487
rect 1685 32385 1719 32419
rect 4077 32385 4111 32419
rect 4997 32385 5031 32419
rect 6193 32385 6227 32419
rect 8208 32385 8242 32419
rect 9689 32385 9723 32419
rect 10542 32385 10576 32419
rect 10701 32385 10735 32419
rect 11713 32385 11747 32419
rect 12072 32385 12106 32419
rect 13829 32385 13863 32419
rect 13921 32385 13955 32419
rect 14958 32385 14992 32419
rect 15117 32385 15151 32419
rect 16221 32385 16255 32419
rect 16497 32385 16531 32419
rect 18521 32385 18555 32419
rect 18981 32385 19015 32419
rect 19165 32385 19199 32419
rect 20913 32385 20947 32419
rect 21097 32385 21131 32419
rect 21189 32385 21223 32419
rect 21465 32385 21499 32419
rect 22201 32385 22235 32419
rect 23581 32385 23615 32419
rect 24961 32385 24995 32419
rect 28022 32385 28056 32419
rect 28917 32385 28951 32419
rect 29184 32385 29218 32419
rect 37381 32385 37415 32419
rect 37657 32385 37691 32419
rect 40417 32385 40451 32419
rect 40693 32385 40727 32419
rect 40877 32385 40911 32419
rect 41245 32385 41279 32419
rect 41441 32385 41475 32419
rect 41889 32385 41923 32419
rect 42165 32385 42199 32419
rect 42809 32385 42843 32419
rect 43361 32385 43395 32419
rect 43453 32385 43487 32419
rect 44097 32385 44131 32419
rect 44557 32385 44591 32419
rect 45017 32385 45051 32419
rect 45477 32385 45511 32419
rect 46029 32385 46063 32419
rect 46213 32385 46247 32419
rect 3709 32317 3743 32351
rect 4261 32317 4295 32351
rect 5114 32317 5148 32351
rect 5273 32317 5307 32351
rect 6377 32317 6411 32351
rect 7941 32317 7975 32351
rect 9505 32317 9539 32351
rect 10425 32317 10459 32351
rect 11805 32317 11839 32351
rect 14105 32317 14139 32351
rect 14841 32317 14875 32351
rect 16681 32317 16715 32351
rect 18797 32317 18831 32351
rect 19901 32317 19935 32351
rect 20018 32317 20052 32351
rect 20177 32317 20211 32351
rect 25697 32317 25731 32351
rect 26985 32317 27019 32351
rect 27169 32317 27203 32351
rect 27905 32317 27939 32351
rect 28181 32317 28215 32351
rect 30849 32317 30883 32351
rect 31033 32317 31067 32351
rect 32689 32317 32723 32351
rect 37565 32317 37599 32351
rect 40233 32317 40267 32351
rect 41981 32317 42015 32351
rect 42901 32317 42935 32351
rect 44281 32317 44315 32351
rect 44649 32317 44683 32351
rect 44833 32317 44867 32351
rect 45937 32317 45971 32351
rect 3065 32249 3099 32283
rect 4721 32249 4755 32283
rect 9321 32249 9355 32283
rect 10149 32249 10183 32283
rect 14565 32249 14599 32283
rect 16313 32249 16347 32283
rect 19625 32249 19659 32283
rect 25053 32249 25087 32283
rect 27629 32249 27663 32283
rect 36921 32249 36955 32283
rect 40601 32249 40635 32283
rect 42073 32249 42107 32283
rect 43177 32249 43211 32283
rect 44097 32249 44131 32283
rect 46121 32249 46155 32283
rect 6009 32181 6043 32215
rect 11345 32181 11379 32215
rect 13645 32181 13679 32215
rect 16037 32181 16071 32215
rect 18153 32181 18187 32215
rect 21373 32181 21407 32215
rect 22017 32181 22051 32215
rect 23673 32181 23707 32215
rect 28825 32181 28859 32215
rect 30297 32181 30331 32215
rect 37105 32181 37139 32215
rect 37657 32181 37691 32215
rect 37841 32181 37875 32215
rect 41245 32181 41279 32215
rect 41705 32181 41739 32215
rect 43085 32181 43119 32215
rect 45109 32181 45143 32215
rect 45569 32181 45603 32215
rect 7757 31977 7791 32011
rect 8953 31977 8987 32011
rect 17785 31977 17819 32011
rect 29193 31977 29227 32011
rect 30941 31977 30975 32011
rect 36829 31977 36863 32011
rect 42441 31977 42475 32011
rect 45109 31977 45143 32011
rect 8033 31909 8067 31943
rect 9873 31909 9907 31943
rect 11069 31909 11103 31943
rect 15577 31909 15611 31943
rect 27261 31909 27295 31943
rect 28457 31909 28491 31943
rect 28825 31909 28859 31943
rect 31263 31909 31297 31943
rect 35357 31909 35391 31943
rect 38669 31909 38703 31943
rect 1409 31841 1443 31875
rect 1685 31841 1719 31875
rect 6377 31841 6411 31875
rect 8677 31841 8711 31875
rect 9229 31841 9263 31875
rect 9413 31841 9447 31875
rect 10149 31841 10183 31875
rect 10287 31841 10321 31875
rect 12265 31841 12299 31875
rect 12357 31841 12391 31875
rect 12541 31841 12575 31875
rect 13093 31841 13127 31875
rect 13277 31841 13311 31875
rect 14197 31841 14231 31875
rect 16405 31841 16439 31875
rect 19257 31841 19291 31875
rect 19441 31841 19475 31875
rect 19901 31841 19935 31875
rect 20177 31841 20211 31875
rect 20294 31841 20328 31875
rect 21833 31841 21867 31875
rect 26617 31841 26651 31875
rect 26801 31841 26835 31875
rect 27537 31841 27571 31875
rect 27675 31841 27709 31875
rect 28549 31841 28583 31875
rect 37657 31841 37691 31875
rect 39865 31841 39899 31875
rect 42625 31841 42659 31875
rect 6644 31773 6678 31807
rect 9137 31773 9171 31807
rect 10425 31773 10459 31807
rect 13001 31773 13035 31807
rect 14453 31773 14487 31807
rect 15945 31773 15979 31807
rect 16661 31773 16695 31807
rect 20453 31773 20487 31807
rect 21373 31773 21407 31807
rect 21557 31773 21591 31807
rect 21649 31773 21683 31807
rect 22100 31773 22134 31807
rect 27813 31773 27847 31807
rect 29377 31773 29411 31807
rect 29561 31773 29595 31807
rect 29817 31773 29851 31807
rect 31033 31773 31067 31807
rect 34161 31773 34195 31807
rect 34713 31773 34747 31807
rect 34861 31773 34895 31807
rect 35081 31773 35115 31807
rect 35219 31773 35253 31807
rect 35817 31773 35851 31807
rect 36093 31773 36127 31807
rect 37933 31773 37967 31807
rect 40141 31773 40175 31807
rect 42349 31773 42383 31807
rect 45017 31773 45051 31807
rect 8401 31705 8435 31739
rect 11897 31705 11931 31739
rect 34989 31705 35023 31739
rect 42625 31705 42659 31739
rect 8493 31637 8527 31671
rect 12633 31637 12667 31671
rect 16037 31637 16071 31671
rect 21097 31637 21131 31671
rect 21189 31637 21223 31671
rect 23213 31637 23247 31671
rect 29009 31637 29043 31671
rect 33977 31637 34011 31671
rect 9689 31433 9723 31467
rect 10057 31433 10091 31467
rect 11805 31433 11839 31467
rect 14933 31433 14967 31467
rect 15301 31433 15335 31467
rect 15393 31433 15427 31467
rect 21465 31433 21499 31467
rect 22385 31433 22419 31467
rect 22477 31433 22511 31467
rect 31585 31433 31619 31467
rect 32597 31433 32631 31467
rect 35173 31433 35207 31467
rect 35633 31433 35667 31467
rect 41521 31433 41555 31467
rect 45201 31433 45235 31467
rect 20453 31365 20487 31399
rect 28549 31365 28583 31399
rect 33968 31365 34002 31399
rect 2237 31297 2271 31331
rect 12173 31297 12207 31331
rect 20637 31297 20671 31331
rect 20729 31297 20763 31331
rect 21005 31297 21039 31331
rect 21097 31297 21131 31331
rect 21281 31297 21315 31331
rect 21557 31297 21591 31331
rect 27721 31297 27755 31331
rect 27813 31297 27847 31331
rect 28089 31297 28123 31331
rect 28365 31297 28399 31331
rect 28641 31297 28675 31331
rect 31033 31297 31067 31331
rect 31493 31297 31527 31331
rect 32505 31297 32539 31331
rect 35541 31297 35575 31331
rect 36461 31297 36495 31331
rect 36737 31297 36771 31331
rect 37565 31297 37599 31331
rect 41337 31297 41371 31331
rect 41613 31297 41647 31331
rect 41705 31297 41739 31331
rect 41797 31297 41831 31331
rect 10149 31229 10183 31263
rect 10241 31229 10275 31263
rect 12265 31229 12299 31263
rect 15577 31229 15611 31263
rect 22569 31229 22603 31263
rect 23581 31229 23615 31263
rect 23765 31229 23799 31263
rect 24225 31229 24259 31263
rect 24501 31229 24535 31263
rect 24618 31229 24652 31263
rect 24777 31229 24811 31263
rect 25697 31229 25731 31263
rect 26157 31229 26191 31263
rect 28181 31229 28215 31263
rect 31677 31229 31711 31263
rect 32689 31229 32723 31263
rect 33701 31229 33735 31263
rect 35725 31229 35759 31263
rect 41981 31229 42015 31263
rect 44741 31229 44775 31263
rect 22017 31161 22051 31195
rect 25421 31161 25455 31195
rect 25973 31161 26007 31195
rect 31125 31161 31159 31195
rect 32137 31161 32171 31195
rect 35081 31161 35115 31195
rect 41889 31161 41923 31195
rect 45109 31161 45143 31195
rect 2053 31093 2087 31127
rect 12449 31093 12483 31127
rect 20913 31093 20947 31127
rect 27537 31093 27571 31127
rect 27997 31093 28031 31127
rect 30849 31093 30883 31127
rect 36553 31093 36587 31127
rect 36921 31093 36955 31127
rect 37657 31093 37691 31127
rect 41337 31093 41371 31127
rect 13093 30889 13127 30923
rect 21097 30889 21131 30923
rect 22201 30889 22235 30923
rect 24225 30889 24259 30923
rect 31953 30889 31987 30923
rect 33977 30889 34011 30923
rect 35357 30889 35391 30923
rect 38393 30889 38427 30923
rect 40601 30889 40635 30923
rect 4077 30821 4111 30855
rect 21005 30821 21039 30855
rect 24409 30821 24443 30855
rect 36093 30821 36127 30855
rect 4721 30753 4755 30787
rect 10977 30753 11011 30787
rect 13645 30753 13679 30787
rect 22845 30753 22879 30787
rect 24869 30753 24903 30787
rect 24961 30753 24995 30787
rect 27813 30753 27847 30787
rect 30573 30753 30607 30787
rect 32137 30753 32171 30787
rect 32781 30753 32815 30787
rect 45385 30753 45419 30787
rect 45845 30753 45879 30787
rect 1777 30685 1811 30719
rect 2044 30685 2078 30719
rect 3985 30685 4019 30719
rect 4997 30685 5031 30719
rect 20637 30685 20671 30719
rect 21925 30685 21959 30719
rect 24777 30685 24811 30719
rect 25421 30685 25455 30719
rect 27629 30685 27663 30719
rect 30481 30685 30515 30719
rect 30840 30685 30874 30719
rect 32321 30685 32355 30719
rect 33057 30685 33091 30719
rect 33174 30685 33208 30719
rect 33333 30685 33367 30719
rect 34713 30685 34747 30719
rect 34806 30685 34840 30719
rect 35081 30685 35115 30719
rect 35178 30685 35212 30719
rect 35541 30685 35575 30719
rect 35817 30685 35851 30719
rect 35909 30685 35943 30719
rect 36185 30685 36219 30719
rect 36461 30685 36495 30719
rect 36553 30685 36587 30719
rect 36921 30685 36955 30719
rect 37197 30685 37231 30719
rect 37381 30685 37415 30719
rect 37657 30685 37691 30719
rect 40049 30685 40083 30719
rect 40141 30685 40175 30719
rect 40325 30685 40359 30719
rect 40417 30685 40451 30719
rect 40509 30685 40543 30719
rect 45477 30685 45511 30719
rect 46121 30685 46155 30719
rect 4445 30617 4479 30651
rect 5264 30617 5298 30651
rect 10793 30617 10827 30651
rect 10885 30617 10919 30651
rect 13461 30617 13495 30651
rect 21741 30617 21775 30651
rect 22109 30617 22143 30651
rect 23112 30617 23146 30651
rect 34989 30617 35023 30651
rect 35725 30617 35759 30651
rect 36369 30617 36403 30651
rect 3157 30549 3191 30583
rect 3801 30549 3835 30583
rect 4537 30549 4571 30583
rect 6377 30549 6411 30583
rect 10425 30549 10459 30583
rect 13553 30549 13587 30583
rect 25237 30549 25271 30583
rect 27261 30549 27295 30583
rect 27721 30549 27755 30583
rect 30297 30549 30331 30583
rect 36737 30549 36771 30583
rect 37197 30549 37231 30583
rect 39865 30549 39899 30583
rect 40969 30549 41003 30583
rect 45937 30549 45971 30583
rect 1961 30345 1995 30379
rect 4721 30345 4755 30379
rect 5457 30345 5491 30379
rect 6837 30345 6871 30379
rect 18797 30345 18831 30379
rect 19809 30345 19843 30379
rect 31953 30345 31987 30379
rect 38761 30345 38795 30379
rect 40785 30345 40819 30379
rect 42257 30345 42291 30379
rect 44925 30345 44959 30379
rect 2421 30277 2455 30311
rect 3608 30277 3642 30311
rect 6745 30277 6779 30311
rect 16037 30277 16071 30311
rect 17141 30277 17175 30311
rect 18061 30277 18095 30311
rect 30840 30277 30874 30311
rect 37381 30277 37415 30311
rect 38209 30277 38243 30311
rect 43361 30277 43395 30311
rect 2329 30209 2363 30243
rect 2973 30209 3007 30243
rect 5641 30209 5675 30243
rect 8208 30209 8242 30243
rect 10333 30209 10367 30243
rect 11989 30209 12023 30243
rect 13645 30209 13679 30243
rect 15945 30209 15979 30243
rect 17049 30209 17083 30243
rect 18705 30209 18739 30243
rect 20913 30209 20947 30243
rect 21373 30209 21407 30243
rect 21557 30209 21591 30243
rect 21649 30209 21683 30243
rect 21833 30209 21867 30243
rect 23029 30209 23063 30243
rect 23489 30209 23523 30243
rect 24409 30209 24443 30243
rect 24547 30209 24581 30243
rect 25789 30209 25823 30243
rect 25881 30209 25915 30243
rect 26157 30209 26191 30243
rect 26801 30209 26835 30243
rect 26985 30209 27019 30243
rect 27252 30209 27286 30243
rect 32137 30209 32171 30243
rect 33174 30209 33208 30243
rect 36369 30209 36403 30243
rect 36553 30209 36587 30243
rect 36645 30209 36679 30243
rect 38393 30209 38427 30243
rect 38669 30209 38703 30243
rect 38945 30209 38979 30243
rect 39221 30209 39255 30243
rect 39405 30209 39439 30243
rect 40233 30209 40267 30243
rect 40417 30209 40451 30243
rect 40509 30209 40543 30243
rect 40601 30209 40635 30243
rect 41613 30209 41647 30243
rect 41761 30209 41795 30243
rect 41889 30209 41923 30243
rect 41981 30209 42015 30243
rect 42119 30209 42153 30243
rect 43085 30209 43119 30243
rect 43637 30209 43671 30243
rect 43729 30209 43763 30243
rect 43913 30209 43947 30243
rect 44097 30209 44131 30243
rect 44189 30209 44223 30243
rect 44281 30209 44315 30243
rect 44465 30209 44499 30243
rect 44741 30209 44775 30243
rect 45017 30209 45051 30243
rect 45661 30209 45695 30243
rect 2513 30141 2547 30175
rect 3341 30141 3375 30175
rect 7021 30141 7055 30175
rect 7941 30141 7975 30175
rect 10057 30141 10091 30175
rect 13737 30141 13771 30175
rect 13829 30141 13863 30175
rect 16221 30141 16255 30175
rect 17325 30141 17359 30175
rect 18981 30141 19015 30175
rect 19349 30141 19383 30175
rect 22109 30141 22143 30175
rect 23673 30141 23707 30175
rect 24685 30141 24719 30175
rect 30573 30141 30607 30175
rect 32321 30141 32355 30175
rect 33057 30141 33091 30175
rect 33333 30141 33367 30175
rect 39497 30141 39531 30175
rect 39681 30141 39715 30175
rect 40141 30141 40175 30175
rect 44373 30141 44407 30175
rect 44557 30141 44591 30175
rect 45109 30141 45143 30175
rect 45845 30141 45879 30175
rect 3157 30073 3191 30107
rect 6377 30073 6411 30107
rect 13277 30073 13311 30107
rect 19625 30073 19659 30107
rect 24133 30073 24167 30107
rect 25605 30073 25639 30107
rect 26617 30073 26651 30107
rect 32781 30073 32815 30107
rect 38577 30073 38611 30107
rect 39037 30073 39071 30107
rect 39129 30073 39163 30107
rect 45385 30073 45419 30107
rect 46029 30073 46063 30107
rect 9321 30005 9355 30039
rect 11805 30005 11839 30039
rect 15577 30005 15611 30039
rect 16681 30005 16715 30039
rect 18337 30005 18371 30039
rect 21005 30005 21039 30039
rect 21189 30005 21223 30039
rect 23213 30005 23247 30039
rect 25329 30005 25363 30039
rect 26065 30005 26099 30039
rect 28365 30005 28399 30039
rect 33977 30005 34011 30039
rect 36185 30005 36219 30039
rect 37473 30005 37507 30039
rect 43913 30005 43947 30039
rect 45569 30005 45603 30039
rect 8585 29801 8619 29835
rect 17141 29801 17175 29835
rect 20729 29801 20763 29835
rect 25697 29801 25731 29835
rect 27169 29801 27203 29835
rect 38577 29801 38611 29835
rect 39037 29801 39071 29835
rect 40785 29801 40819 29835
rect 42165 29801 42199 29835
rect 45661 29801 45695 29835
rect 17883 29733 17917 29767
rect 19073 29733 19107 29767
rect 20545 29733 20579 29767
rect 23765 29733 23799 29767
rect 25513 29733 25547 29767
rect 29377 29733 29411 29767
rect 39589 29733 39623 29767
rect 43085 29733 43119 29767
rect 46305 29733 46339 29767
rect 1685 29665 1719 29699
rect 7113 29665 7147 29699
rect 7297 29665 7331 29699
rect 7849 29665 7883 29699
rect 9873 29665 9907 29699
rect 10057 29665 10091 29699
rect 10425 29665 10459 29699
rect 10701 29665 10735 29699
rect 17233 29665 17267 29699
rect 18153 29665 18187 29699
rect 18429 29665 18463 29699
rect 22201 29665 22235 29699
rect 27721 29665 27755 29699
rect 29561 29665 29595 29699
rect 38761 29665 38795 29699
rect 41061 29665 41095 29699
rect 42441 29665 42475 29699
rect 42533 29665 42567 29699
rect 45017 29665 45051 29699
rect 1409 29597 1443 29631
rect 5641 29597 5675 29631
rect 7021 29597 7055 29631
rect 8769 29597 8803 29631
rect 9781 29597 9815 29631
rect 11345 29597 11379 29631
rect 11612 29597 11646 29631
rect 15393 29597 15427 29631
rect 15669 29597 15703 29631
rect 15761 29597 15795 29631
rect 17417 29597 17451 29631
rect 18291 29597 18325 29631
rect 20913 29597 20947 29631
rect 21189 29597 21223 29631
rect 21925 29597 21959 29631
rect 22477 29597 22511 29631
rect 23581 29597 23615 29631
rect 27629 29597 27663 29631
rect 29193 29597 29227 29631
rect 35449 29597 35483 29631
rect 35633 29597 35667 29631
rect 35725 29597 35759 29631
rect 35817 29597 35851 29631
rect 38301 29597 38335 29631
rect 39221 29597 39255 29631
rect 39865 29597 39899 29631
rect 41245 29597 41279 29631
rect 41797 29597 41831 29631
rect 42073 29597 42107 29631
rect 42349 29597 42383 29631
rect 42625 29597 42659 29631
rect 42809 29597 42843 29631
rect 42993 29597 43027 29631
rect 43177 29597 43211 29631
rect 43269 29597 43303 29631
rect 45201 29597 45235 29631
rect 45477 29597 45511 29631
rect 45661 29597 45695 29631
rect 46121 29597 46155 29631
rect 46305 29597 46339 29631
rect 46673 29597 46707 29631
rect 7665 29529 7699 29563
rect 16006 29529 16040 29563
rect 20269 29529 20303 29563
rect 21465 29529 21499 29563
rect 25237 29529 25271 29563
rect 29828 29529 29862 29563
rect 37749 29529 37783 29563
rect 39405 29529 39439 29563
rect 40601 29529 40635 29563
rect 40817 29529 40851 29563
rect 45385 29529 45419 29563
rect 5457 29461 5491 29495
rect 6653 29461 6687 29495
rect 9413 29461 9447 29495
rect 12725 29461 12759 29495
rect 15209 29461 15243 29495
rect 15485 29461 15519 29495
rect 21005 29461 21039 29495
rect 22661 29461 22695 29495
rect 27537 29461 27571 29495
rect 30941 29461 30975 29495
rect 36001 29461 36035 29495
rect 37841 29461 37875 29495
rect 40049 29461 40083 29495
rect 40969 29461 41003 29495
rect 41521 29461 41555 29495
rect 45845 29461 45879 29495
rect 6377 29257 6411 29291
rect 9597 29257 9631 29291
rect 11529 29257 11563 29291
rect 12449 29257 12483 29291
rect 13185 29257 13219 29291
rect 16497 29257 16531 29291
rect 19257 29257 19291 29291
rect 20729 29257 20763 29291
rect 29193 29257 29227 29291
rect 36737 29257 36771 29291
rect 38485 29257 38519 29291
rect 40969 29257 41003 29291
rect 46673 29257 46707 29291
rect 5080 29189 5114 29223
rect 10232 29189 10266 29223
rect 15362 29189 15396 29223
rect 37565 29189 37599 29223
rect 6745 29121 6779 29155
rect 7840 29121 7874 29155
rect 9505 29121 9539 29155
rect 11713 29121 11747 29155
rect 13093 29121 13127 29155
rect 13820 29121 13854 29155
rect 17417 29121 17451 29155
rect 17601 29121 17635 29155
rect 18475 29121 18509 29155
rect 19605 29121 19639 29155
rect 29561 29121 29595 29155
rect 29653 29121 29687 29155
rect 30205 29121 30239 29155
rect 33609 29121 33643 29155
rect 33876 29121 33910 29155
rect 36093 29121 36127 29155
rect 36186 29121 36220 29155
rect 36369 29121 36403 29155
rect 36461 29121 36495 29155
rect 36599 29121 36633 29155
rect 37289 29121 37323 29155
rect 37473 29121 37507 29155
rect 37657 29121 37691 29155
rect 38117 29121 38151 29155
rect 38669 29121 38703 29155
rect 38761 29121 38795 29155
rect 38945 29121 38979 29155
rect 39129 29121 39163 29155
rect 40877 29121 40911 29155
rect 41061 29121 41095 29155
rect 41521 29121 41555 29155
rect 41717 29121 41751 29155
rect 41889 29121 41923 29155
rect 42073 29121 42107 29155
rect 42625 29121 42659 29155
rect 42809 29121 42843 29155
rect 42901 29121 42935 29155
rect 46489 29121 46523 29155
rect 4813 29053 4847 29087
rect 6837 29053 6871 29087
rect 7021 29053 7055 29087
rect 7573 29053 7607 29087
rect 9781 29053 9815 29087
rect 9965 29053 9999 29087
rect 13369 29053 13403 29087
rect 13553 29053 13587 29087
rect 15117 29053 15151 29087
rect 18337 29053 18371 29087
rect 18613 29053 18647 29087
rect 19349 29053 19383 29087
rect 29745 29053 29779 29087
rect 41613 29053 41647 29087
rect 6193 28985 6227 29019
rect 9137 28985 9171 29019
rect 18061 28985 18095 29019
rect 30021 28985 30055 29019
rect 34989 28985 35023 29019
rect 38853 28985 38887 29019
rect 42073 28985 42107 29019
rect 8953 28917 8987 28951
rect 11345 28917 11379 28951
rect 12725 28917 12759 28951
rect 14933 28917 14967 28951
rect 37841 28917 37875 28951
rect 42441 28917 42475 28951
rect 8033 28713 8067 28747
rect 9781 28713 9815 28747
rect 14105 28713 14139 28747
rect 15209 28713 15243 28747
rect 18245 28713 18279 28747
rect 19717 28713 19751 28747
rect 29285 28713 29319 28747
rect 33885 28713 33919 28747
rect 37013 28713 37047 28747
rect 38761 28713 38795 28747
rect 5917 28645 5951 28679
rect 28549 28645 28583 28679
rect 44189 28645 44223 28679
rect 3249 28577 3283 28611
rect 7297 28577 7331 28611
rect 7481 28577 7515 28611
rect 9505 28577 9539 28611
rect 10241 28577 10275 28611
rect 10425 28577 10459 28611
rect 11161 28577 11195 28611
rect 11713 28577 11747 28611
rect 12633 28577 12667 28611
rect 28181 28577 28215 28611
rect 29561 28577 29595 28611
rect 32505 28577 32539 28611
rect 32597 28577 32631 28611
rect 33517 28577 33551 28611
rect 33609 28577 33643 28611
rect 42073 28577 42107 28611
rect 44465 28577 44499 28611
rect 44557 28577 44591 28611
rect 4445 28509 4479 28543
rect 4537 28509 4571 28543
rect 7205 28509 7239 28543
rect 8217 28509 8251 28543
rect 10977 28509 11011 28543
rect 11989 28509 12023 28543
rect 12909 28509 12943 28543
rect 14289 28509 14323 28543
rect 14565 28509 14599 28543
rect 18429 28509 18463 28543
rect 19533 28509 19567 28543
rect 21281 28509 21315 28543
rect 21741 28509 21775 28543
rect 26157 28509 26191 28543
rect 27997 28509 28031 28543
rect 28733 28509 28767 28543
rect 34069 28509 34103 28543
rect 37197 28509 37231 28543
rect 41797 28509 41831 28543
rect 41889 28509 41923 28543
rect 43729 28509 43763 28543
rect 44373 28509 44407 28543
rect 44649 28509 44683 28543
rect 45017 28509 45051 28543
rect 45201 28509 45235 28543
rect 4782 28441 4816 28475
rect 9413 28441 9447 28475
rect 10149 28441 10183 28475
rect 15025 28441 15059 28475
rect 15225 28441 15259 28475
rect 20177 28441 20211 28475
rect 20545 28441 20579 28475
rect 26424 28441 26458 28475
rect 29009 28441 29043 28475
rect 29806 28441 29840 28475
rect 33425 28441 33459 28475
rect 37473 28441 37507 28475
rect 38669 28441 38703 28475
rect 43913 28441 43947 28475
rect 2605 28373 2639 28407
rect 2973 28373 3007 28407
rect 3065 28373 3099 28407
rect 4261 28373 4295 28407
rect 6837 28373 6871 28407
rect 8953 28373 8987 28407
rect 9321 28373 9355 28407
rect 10609 28373 10643 28407
rect 11069 28373 11103 28407
rect 14473 28373 14507 28407
rect 15393 28373 15427 28407
rect 21097 28373 21131 28407
rect 21557 28373 21591 28407
rect 27537 28373 27571 28407
rect 27629 28373 27663 28407
rect 28089 28373 28123 28407
rect 30941 28373 30975 28407
rect 32045 28373 32079 28407
rect 32413 28373 32447 28407
rect 33057 28373 33091 28407
rect 37381 28373 37415 28407
rect 42073 28373 42107 28407
rect 44097 28373 44131 28407
rect 45201 28373 45235 28407
rect 11897 28169 11931 28203
rect 12357 28169 12391 28203
rect 18245 28169 18279 28203
rect 21557 28169 21591 28203
rect 21833 28169 21867 28203
rect 26617 28169 26651 28203
rect 27813 28169 27847 28203
rect 28825 28169 28859 28203
rect 29377 28169 29411 28203
rect 29745 28169 29779 28203
rect 29837 28169 29871 28203
rect 31769 28169 31803 28203
rect 33517 28169 33551 28203
rect 39773 28169 39807 28203
rect 41705 28169 41739 28203
rect 42165 28169 42199 28203
rect 42641 28169 42675 28203
rect 44281 28169 44315 28203
rect 44925 28169 44959 28203
rect 46673 28169 46707 28203
rect 12265 28101 12299 28135
rect 13829 28101 13863 28135
rect 14105 28101 14139 28135
rect 14197 28101 14231 28135
rect 15945 28101 15979 28135
rect 17141 28101 17175 28135
rect 21281 28101 21315 28135
rect 22201 28101 22235 28135
rect 32382 28101 32416 28135
rect 39405 28101 39439 28135
rect 42441 28101 42475 28135
rect 43913 28101 43947 28135
rect 44113 28101 44147 28135
rect 44557 28101 44591 28135
rect 2329 28033 2363 28067
rect 2605 28033 2639 28067
rect 2872 28033 2906 28067
rect 4629 28033 4663 28067
rect 4905 28033 4939 28067
rect 7389 28033 7423 28067
rect 7665 28033 7699 28067
rect 12725 28033 12759 28067
rect 14013 28033 14047 28067
rect 14657 28033 14691 28067
rect 14841 28033 14875 28067
rect 14933 28033 14967 28067
rect 15577 28033 15611 28067
rect 16773 28033 16807 28067
rect 18153 28033 18187 28067
rect 18613 28033 18647 28067
rect 19073 28033 19107 28067
rect 19625 28033 19659 28067
rect 20361 28033 20395 28067
rect 22293 28033 22327 28067
rect 26801 28033 26835 28067
rect 27721 28033 27755 28067
rect 29009 28033 29043 28067
rect 30573 28033 30607 28067
rect 31953 28033 31987 28067
rect 38209 28033 38243 28067
rect 39957 28033 39991 28067
rect 40049 28033 40083 28067
rect 40233 28033 40267 28067
rect 40325 28033 40359 28067
rect 41521 28033 41555 28067
rect 41797 28033 41831 28067
rect 43545 28033 43579 28067
rect 44373 28033 44407 28067
rect 44649 28033 44683 28067
rect 44741 28033 44775 28067
rect 45201 28033 45235 28067
rect 45385 28033 45419 28067
rect 45661 28033 45695 28067
rect 46581 28033 46615 28067
rect 12541 27965 12575 27999
rect 14565 27965 14599 27999
rect 15393 27965 15427 27999
rect 15853 27965 15887 27999
rect 16037 27965 16071 27999
rect 20085 27965 20119 27999
rect 22477 27965 22511 27999
rect 23213 27965 23247 27999
rect 23397 27965 23431 27999
rect 24133 27965 24167 27999
rect 24271 27965 24305 27999
rect 24409 27965 24443 27999
rect 25145 27965 25179 27999
rect 27905 27965 27939 27999
rect 30021 27965 30055 27999
rect 30665 27965 30699 27999
rect 30757 27965 30791 27999
rect 32137 27965 32171 27999
rect 33609 27965 33643 27999
rect 38393 27965 38427 27999
rect 41337 27965 41371 27999
rect 41889 27965 41923 27999
rect 45017 27965 45051 27999
rect 13001 27897 13035 27931
rect 13185 27897 13219 27931
rect 23857 27897 23891 27931
rect 25053 27897 25087 27931
rect 25421 27897 25455 27931
rect 39589 27897 39623 27931
rect 43729 27897 43763 27931
rect 2145 27829 2179 27863
rect 3985 27829 4019 27863
rect 7205 27829 7239 27863
rect 7481 27829 7515 27863
rect 16221 27829 16255 27863
rect 18797 27829 18831 27863
rect 19349 27829 19383 27863
rect 19901 27829 19935 27863
rect 25605 27829 25639 27863
rect 27353 27829 27387 27863
rect 30205 27829 30239 27863
rect 33839 27829 33873 27863
rect 38669 27829 38703 27863
rect 41889 27829 41923 27863
rect 42625 27829 42659 27863
rect 42809 27829 42843 27863
rect 44097 27829 44131 27863
rect 45477 27829 45511 27863
rect 3065 27625 3099 27659
rect 3157 27625 3191 27659
rect 5457 27625 5491 27659
rect 6469 27625 6503 27659
rect 14979 27625 15013 27659
rect 17601 27625 17635 27659
rect 22661 27625 22695 27659
rect 28457 27625 28491 27659
rect 29285 27625 29319 27659
rect 31401 27625 31435 27659
rect 37657 27625 37691 27659
rect 45845 27625 45879 27659
rect 8401 27557 8435 27591
rect 12357 27557 12391 27591
rect 18613 27557 18647 27591
rect 18981 27557 19015 27591
rect 19625 27557 19659 27591
rect 22845 27557 22879 27591
rect 26249 27557 26283 27591
rect 34529 27557 34563 27591
rect 40141 27557 40175 27591
rect 40325 27557 40359 27591
rect 41705 27557 41739 27591
rect 46213 27557 46247 27591
rect 1685 27489 1719 27523
rect 4445 27489 4479 27523
rect 6009 27489 6043 27523
rect 7941 27489 7975 27523
rect 10149 27489 10183 27523
rect 10333 27489 10367 27523
rect 10977 27489 11011 27523
rect 11069 27489 11103 27523
rect 12449 27489 12483 27523
rect 14565 27489 14599 27523
rect 14749 27489 14783 27523
rect 16589 27489 16623 27523
rect 24133 27489 24167 27523
rect 26801 27489 26835 27523
rect 29745 27489 29779 27523
rect 30205 27489 30239 27523
rect 30598 27489 30632 27523
rect 30757 27489 30791 27523
rect 32413 27489 32447 27523
rect 32689 27489 32723 27523
rect 33333 27489 33367 27523
rect 33726 27489 33760 27523
rect 35265 27489 35299 27523
rect 38577 27489 38611 27523
rect 41889 27489 41923 27523
rect 45477 27489 45511 27523
rect 1952 27421 1986 27455
rect 3341 27421 3375 27455
rect 4169 27421 4203 27455
rect 5825 27421 5859 27455
rect 6285 27421 6319 27455
rect 8217 27421 8251 27455
rect 16957 27421 16991 27455
rect 17049 27421 17083 27455
rect 18337 27421 18371 27455
rect 18797 27421 18831 27455
rect 19349 27421 19383 27455
rect 19809 27421 19843 27455
rect 21281 27421 21315 27455
rect 21548 27421 21582 27455
rect 23029 27421 23063 27455
rect 23949 27421 23983 27455
rect 24409 27421 24443 27455
rect 24665 27421 24699 27455
rect 26157 27421 26191 27455
rect 27077 27421 27111 27455
rect 28733 27421 28767 27455
rect 29561 27421 29595 27455
rect 30481 27421 30515 27455
rect 32229 27421 32263 27455
rect 32873 27421 32907 27455
rect 33609 27421 33643 27455
rect 33885 27421 33919 27455
rect 35173 27421 35207 27455
rect 37289 27421 37323 27455
rect 37381 27421 37415 27455
rect 38117 27421 38151 27455
rect 38209 27421 38243 27455
rect 38393 27421 38427 27455
rect 38495 27421 38529 27455
rect 38853 27421 38887 27455
rect 40417 27421 40451 27455
rect 40969 27421 41003 27455
rect 41429 27421 41463 27455
rect 45661 27421 45695 27455
rect 46397 27421 46431 27455
rect 7757 27353 7791 27387
rect 11989 27353 12023 27387
rect 14289 27353 14323 27387
rect 16497 27353 16531 27387
rect 17141 27353 17175 27387
rect 17509 27353 17543 27387
rect 20076 27353 20110 27387
rect 23213 27353 23247 27387
rect 23857 27353 23891 27387
rect 27344 27353 27378 27387
rect 29009 27353 29043 27387
rect 32321 27353 32355 27387
rect 35510 27353 35544 27387
rect 36737 27353 36771 27387
rect 36921 27353 36955 27387
rect 37933 27353 37967 27387
rect 39865 27353 39899 27387
rect 41153 27353 41187 27387
rect 3801 27285 3835 27319
rect 4261 27285 4295 27319
rect 5917 27285 5951 27319
rect 7389 27285 7423 27319
rect 7849 27285 7883 27319
rect 9689 27285 9723 27319
rect 10057 27285 10091 27319
rect 10517 27285 10551 27319
rect 10885 27285 10919 27319
rect 21189 27285 21223 27319
rect 23305 27285 23339 27319
rect 23489 27285 23523 27319
rect 25789 27285 25823 27319
rect 25973 27285 26007 27319
rect 26617 27285 26651 27319
rect 26709 27285 26743 27319
rect 28549 27285 28583 27319
rect 31861 27285 31895 27319
rect 34989 27285 35023 27319
rect 36645 27285 36679 27319
rect 37013 27285 37047 27319
rect 37105 27285 37139 27319
rect 37841 27285 37875 27319
rect 40601 27285 40635 27319
rect 41337 27285 41371 27319
rect 4813 27081 4847 27115
rect 11805 27081 11839 27115
rect 11989 27081 12023 27115
rect 12909 27081 12943 27115
rect 19073 27081 19107 27115
rect 21833 27081 21867 27115
rect 28365 27081 28399 27115
rect 35265 27081 35299 27115
rect 35633 27081 35667 27115
rect 38117 27081 38151 27115
rect 38761 27081 38795 27115
rect 40141 27081 40175 27115
rect 41337 27081 41371 27115
rect 46397 27081 46431 27115
rect 8392 27013 8426 27047
rect 11621 27013 11655 27047
rect 11897 27013 11931 27047
rect 12541 27013 12575 27047
rect 12725 27013 12759 27047
rect 15209 27013 15243 27047
rect 15669 27013 15703 27047
rect 16865 27013 16899 27047
rect 17325 27013 17359 27047
rect 18245 27013 18279 27047
rect 18797 27013 18831 27047
rect 21097 27013 21131 27047
rect 22293 27013 22327 27047
rect 27230 27013 27264 27047
rect 1409 26945 1443 26979
rect 4721 26945 4755 26979
rect 6561 26945 6595 26979
rect 6828 26945 6862 26979
rect 8125 26945 8159 26979
rect 9689 26945 9723 26979
rect 10241 26945 10275 26979
rect 10793 26945 10827 26979
rect 12633 26945 12667 26979
rect 13461 26945 13495 26979
rect 13645 26945 13679 26979
rect 14013 26945 14047 26979
rect 15301 26945 15335 26979
rect 17233 26945 17267 26979
rect 17417 26945 17451 26979
rect 17877 26945 17911 26979
rect 18429 26945 18463 26979
rect 18981 26945 19015 26979
rect 19533 26945 19567 26979
rect 20269 26945 20303 26979
rect 21281 26945 21315 26979
rect 21465 26945 21499 26979
rect 21557 26945 21591 26979
rect 22201 26945 22235 26979
rect 23121 26945 23155 26979
rect 23995 26945 24029 26979
rect 25421 26945 25455 26979
rect 25513 26945 25547 26979
rect 25789 26945 25823 26979
rect 25973 26945 26007 26979
rect 26341 26945 26375 26979
rect 26985 26945 27019 26979
rect 29101 26945 29135 26979
rect 29837 26945 29871 26979
rect 32321 26945 32355 26979
rect 33057 26945 33091 26979
rect 33241 26945 33275 26979
rect 34094 26945 34128 26979
rect 35725 26945 35759 26979
rect 36093 26945 36127 26979
rect 36369 26945 36403 26979
rect 38301 26945 38335 26979
rect 38945 26945 38979 26979
rect 39405 26945 39439 26979
rect 39589 26945 39623 26979
rect 39773 26945 39807 26979
rect 40233 26945 40267 26979
rect 41521 26945 41555 26979
rect 41705 26945 41739 26979
rect 41889 26945 41923 26979
rect 42625 26945 42659 26979
rect 42901 26945 42935 26979
rect 43085 26945 43119 26979
rect 43269 26945 43303 26979
rect 45569 26945 45603 26979
rect 45661 26945 45695 26979
rect 46581 26945 46615 26979
rect 4997 26877 5031 26911
rect 12357 26877 12391 26911
rect 13737 26877 13771 26911
rect 15761 26877 15795 26911
rect 16773 26877 16807 26911
rect 19993 26877 20027 26911
rect 22385 26877 22419 26911
rect 22937 26877 22971 26911
rect 23857 26877 23891 26911
rect 24133 26877 24167 26911
rect 25697 26877 25731 26911
rect 28917 26877 28951 26911
rect 29954 26877 29988 26911
rect 30123 26877 30157 26911
rect 33977 26877 34011 26911
rect 34253 26877 34287 26911
rect 35817 26877 35851 26911
rect 39865 26877 39899 26911
rect 41797 26877 41831 26911
rect 42165 26877 42199 26911
rect 42993 26877 43027 26911
rect 45845 26877 45879 26911
rect 7941 26809 7975 26843
rect 9505 26809 9539 26843
rect 23581 26809 23615 26843
rect 29561 26809 29595 26843
rect 33701 26809 33735 26843
rect 39589 26809 39623 26843
rect 41889 26809 41923 26843
rect 41981 26809 42015 26843
rect 43361 26809 43395 26843
rect 45385 26809 45419 26843
rect 46029 26809 46063 26843
rect 1593 26741 1627 26775
rect 4353 26741 4387 26775
rect 9873 26741 9907 26775
rect 10057 26741 10091 26775
rect 10609 26741 10643 26775
rect 12173 26741 12207 26775
rect 13461 26741 13495 26775
rect 19625 26741 19659 26775
rect 24777 26741 24811 26775
rect 25237 26741 25271 26775
rect 30757 26741 30791 26775
rect 32137 26741 32171 26775
rect 34897 26741 34931 26775
rect 37105 26741 37139 26775
rect 39957 26741 39991 26775
rect 40417 26741 40451 26775
rect 2973 26537 3007 26571
rect 6377 26537 6411 26571
rect 7021 26537 7055 26571
rect 12081 26537 12115 26571
rect 12357 26537 12391 26571
rect 13001 26537 13035 26571
rect 14289 26537 14323 26571
rect 18705 26537 18739 26571
rect 33149 26537 33183 26571
rect 35633 26537 35667 26571
rect 38301 26537 38335 26571
rect 38853 26537 38887 26571
rect 46029 26537 46063 26571
rect 46213 26537 46247 26571
rect 46397 26537 46431 26571
rect 46765 26537 46799 26571
rect 7757 26469 7791 26503
rect 12541 26469 12575 26503
rect 13185 26469 13219 26503
rect 13829 26469 13863 26503
rect 15301 26469 15335 26503
rect 20361 26469 20395 26503
rect 20821 26469 20855 26503
rect 21189 26469 21223 26503
rect 23765 26469 23799 26503
rect 26433 26469 26467 26503
rect 30205 26469 30239 26503
rect 42165 26469 42199 26503
rect 4077 26401 4111 26435
rect 4721 26401 4755 26435
rect 4997 26401 5031 26435
rect 5114 26401 5148 26435
rect 5273 26401 5307 26435
rect 8217 26401 8251 26435
rect 8309 26401 8343 26435
rect 9229 26401 9263 26435
rect 10701 26401 10735 26435
rect 15393 26401 15427 26435
rect 15761 26401 15795 26435
rect 16589 26401 16623 26435
rect 30849 26401 30883 26435
rect 42717 26401 42751 26435
rect 43545 26401 43579 26435
rect 1593 26333 1627 26367
rect 3985 26333 4019 26367
rect 4261 26333 4295 26367
rect 6193 26333 6227 26367
rect 7205 26333 7239 26367
rect 9496 26333 9530 26367
rect 10957 26333 10991 26367
rect 12633 26333 12667 26367
rect 13277 26333 13311 26367
rect 14565 26333 14599 26367
rect 14841 26333 14875 26367
rect 14933 26333 14967 26367
rect 17049 26333 17083 26367
rect 17233 26333 17267 26367
rect 17785 26333 17819 26367
rect 18613 26333 18647 26367
rect 19533 26333 19567 26367
rect 20177 26333 20211 26367
rect 20637 26333 20671 26367
rect 21005 26333 21039 26367
rect 30573 26333 30607 26367
rect 31769 26333 31803 26367
rect 32036 26333 32070 26367
rect 35541 26333 35575 26367
rect 38209 26333 38243 26367
rect 38761 26333 38795 26367
rect 41613 26333 41647 26367
rect 41889 26333 41923 26367
rect 41981 26333 42015 26367
rect 42257 26333 42291 26367
rect 42533 26333 42567 26367
rect 42809 26333 42843 26367
rect 42993 26333 43027 26367
rect 43177 26333 43211 26367
rect 43361 26333 43395 26367
rect 45753 26333 45787 26367
rect 46305 26333 46339 26367
rect 1860 26265 1894 26299
rect 5917 26265 5951 26299
rect 8125 26265 8159 26299
rect 12173 26265 12207 26299
rect 13001 26265 13035 26299
rect 13645 26265 13679 26299
rect 14105 26265 14139 26299
rect 14289 26265 14323 26299
rect 16681 26265 16715 26299
rect 17141 26265 17175 26299
rect 17601 26265 17635 26299
rect 19901 26265 19935 26299
rect 23397 26265 23431 26299
rect 26249 26265 26283 26299
rect 30665 26265 30699 26299
rect 41797 26265 41831 26299
rect 3801 26197 3835 26231
rect 10609 26197 10643 26231
rect 12383 26197 12417 26231
rect 13461 26197 13495 26231
rect 13553 26197 13587 26231
rect 23857 26197 23891 26231
rect 38669 26197 38703 26231
rect 39221 26197 39255 26231
rect 2053 25993 2087 26027
rect 2421 25993 2455 26027
rect 2789 25993 2823 26027
rect 2881 25993 2915 26027
rect 13553 25993 13587 26027
rect 17417 25993 17451 26027
rect 23949 25993 23983 26027
rect 46213 25993 46247 26027
rect 5825 25925 5859 25959
rect 13369 25925 13403 25959
rect 36737 25925 36771 25959
rect 2237 25857 2271 25891
rect 3985 25857 4019 25891
rect 4905 25857 4939 25891
rect 5043 25857 5077 25891
rect 7389 25857 7423 25891
rect 8585 25857 8619 25891
rect 9045 25857 9079 25891
rect 9965 25857 9999 25891
rect 11529 25857 11563 25891
rect 13829 25857 13863 25891
rect 14197 25857 14231 25891
rect 14289 25857 14323 25891
rect 14381 25857 14415 25891
rect 15485 25857 15519 25891
rect 17233 25857 17267 25891
rect 17877 25857 17911 25891
rect 18153 25857 18187 25891
rect 19073 25857 19107 25891
rect 23305 25857 23339 25891
rect 23397 25857 23431 25891
rect 23673 25857 23707 25891
rect 23857 25857 23891 25891
rect 25973 25857 26007 25891
rect 33793 25857 33827 25891
rect 36553 25857 36587 25891
rect 36829 25857 36863 25891
rect 39681 25857 39715 25891
rect 42441 25857 42475 25891
rect 42901 25857 42935 25891
rect 43269 25857 43303 25891
rect 43545 25857 43579 25891
rect 44097 25857 44131 25891
rect 44281 25857 44315 25891
rect 44373 25857 44407 25891
rect 45753 25857 45787 25891
rect 3065 25789 3099 25823
rect 4169 25789 4203 25823
rect 5181 25789 5215 25823
rect 7481 25789 7515 25823
rect 7573 25789 7607 25823
rect 9321 25789 9355 25823
rect 10241 25789 10275 25823
rect 11805 25789 11839 25823
rect 12449 25789 12483 25823
rect 12725 25789 12759 25823
rect 15209 25789 15243 25823
rect 23581 25789 23615 25823
rect 33517 25789 33551 25823
rect 42809 25789 42843 25823
rect 43177 25789 43211 25823
rect 4629 25721 4663 25755
rect 7021 25653 7055 25687
rect 8401 25653 8435 25687
rect 13553 25653 13587 25687
rect 14565 25653 14599 25687
rect 18383 25653 18417 25687
rect 19257 25653 19291 25687
rect 23121 25653 23155 25687
rect 26249 25653 26283 25687
rect 36369 25653 36403 25687
rect 39497 25653 39531 25687
rect 42533 25653 42567 25687
rect 43637 25653 43671 25687
rect 44005 25653 44039 25687
rect 44373 25653 44407 25687
rect 46029 25653 46063 25687
rect 5181 25449 5215 25483
rect 14105 25449 14139 25483
rect 21741 25449 21775 25483
rect 37381 25449 37415 25483
rect 12725 25381 12759 25415
rect 21557 25381 21591 25415
rect 24133 25381 24167 25415
rect 26341 25381 26375 25415
rect 37565 25381 37599 25415
rect 39037 25381 39071 25415
rect 45293 25381 45327 25415
rect 7757 25313 7791 25347
rect 7941 25313 7975 25347
rect 9137 25313 9171 25347
rect 12449 25313 12483 25347
rect 14749 25313 14783 25347
rect 15025 25313 15059 25347
rect 15761 25313 15795 25347
rect 15853 25313 15887 25347
rect 16773 25313 16807 25347
rect 16865 25313 16899 25347
rect 21281 25313 21315 25347
rect 36277 25313 36311 25347
rect 37289 25313 37323 25347
rect 40141 25313 40175 25347
rect 43913 25313 43947 25347
rect 46213 25313 46247 25347
rect 1869 25245 1903 25279
rect 3801 25245 3835 25279
rect 4057 25245 4091 25279
rect 6837 25245 6871 25279
rect 7665 25245 7699 25279
rect 9413 25245 9447 25279
rect 12541 25245 12575 25279
rect 14105 25245 14139 25279
rect 14289 25245 14323 25279
rect 16221 25245 16255 25279
rect 16313 25245 16347 25279
rect 16405 25245 16439 25279
rect 17233 25245 17267 25279
rect 17325 25245 17359 25279
rect 17417 25245 17451 25279
rect 17969 25245 18003 25279
rect 18061 25245 18095 25279
rect 18337 25245 18371 25279
rect 23121 25245 23155 25279
rect 23397 25245 23431 25279
rect 27169 25245 27203 25279
rect 31033 25245 31067 25279
rect 33149 25245 33183 25279
rect 34989 25245 35023 25279
rect 36553 25245 36587 25279
rect 37197 25245 37231 25279
rect 37933 25245 37967 25279
rect 38393 25245 38427 25279
rect 38485 25245 38519 25279
rect 38853 25245 38887 25279
rect 40049 25245 40083 25279
rect 40325 25245 40359 25279
rect 44005 25245 44039 25279
rect 44465 25245 44499 25279
rect 44741 25245 44775 25279
rect 45937 25245 45971 25279
rect 2136 25177 2170 25211
rect 26065 25177 26099 25211
rect 33394 25177 33428 25211
rect 39313 25177 39347 25211
rect 44281 25177 44315 25211
rect 45017 25177 45051 25211
rect 3249 25109 3283 25143
rect 6653 25109 6687 25143
rect 7297 25109 7331 25143
rect 12081 25109 12115 25143
rect 17785 25109 17819 25143
rect 26985 25109 27019 25143
rect 30849 25109 30883 25143
rect 34529 25109 34563 25143
rect 34805 25109 34839 25143
rect 39405 25109 39439 25143
rect 39865 25109 39899 25143
rect 40785 25109 40819 25143
rect 45477 25109 45511 25143
rect 2789 24905 2823 24939
rect 19257 24905 19291 24939
rect 33149 24905 33183 24939
rect 37013 24905 37047 24939
rect 41153 24905 41187 24939
rect 44005 24905 44039 24939
rect 2329 24837 2363 24871
rect 9290 24837 9324 24871
rect 23213 24837 23247 24871
rect 30389 24837 30423 24871
rect 30840 24837 30874 24871
rect 38393 24837 38427 24871
rect 1409 24769 1443 24803
rect 2973 24769 3007 24803
rect 7829 24769 7863 24803
rect 12173 24769 12207 24803
rect 12265 24769 12299 24803
rect 16681 24769 16715 24803
rect 18052 24769 18086 24803
rect 19441 24769 19475 24803
rect 22385 24769 22419 24803
rect 24961 24769 24995 24803
rect 25421 24769 25455 24803
rect 25688 24769 25722 24803
rect 27252 24769 27286 24803
rect 30205 24769 30239 24803
rect 30481 24769 30515 24803
rect 32413 24769 32447 24803
rect 33333 24769 33367 24803
rect 34345 24769 34379 24803
rect 34621 24769 34655 24803
rect 36461 24769 36495 24803
rect 36921 24769 36955 24803
rect 38577 24769 38611 24803
rect 38945 24769 38979 24803
rect 39313 24769 39347 24803
rect 39589 24769 39623 24803
rect 40509 24769 40543 24803
rect 40693 24769 40727 24803
rect 40785 24769 40819 24803
rect 40877 24769 40911 24803
rect 41337 24769 41371 24803
rect 41429 24769 41463 24803
rect 43913 24769 43947 24803
rect 44097 24769 44131 24803
rect 44741 24769 44775 24803
rect 46489 24769 46523 24803
rect 2421 24701 2455 24735
rect 2513 24701 2547 24735
rect 7573 24701 7607 24735
rect 9045 24701 9079 24735
rect 11805 24701 11839 24735
rect 16957 24701 16991 24735
rect 17785 24701 17819 24735
rect 19533 24701 19567 24735
rect 19717 24701 19751 24735
rect 20453 24701 20487 24735
rect 20570 24701 20604 24735
rect 20729 24701 20763 24735
rect 22109 24701 22143 24735
rect 26985 24701 27019 24735
rect 29101 24701 29135 24735
rect 30573 24701 30607 24735
rect 33425 24701 33459 24735
rect 33609 24701 33643 24735
rect 34069 24701 34103 24735
rect 34462 24701 34496 24735
rect 39865 24701 39899 24735
rect 41521 24701 41555 24735
rect 41613 24701 41647 24735
rect 1961 24633 1995 24667
rect 20177 24633 20211 24667
rect 23581 24633 23615 24667
rect 29469 24633 29503 24667
rect 41061 24633 41095 24667
rect 44557 24633 44591 24667
rect 1593 24565 1627 24599
rect 8953 24565 8987 24599
rect 10425 24565 10459 24599
rect 12449 24565 12483 24599
rect 19165 24565 19199 24599
rect 21373 24565 21407 24599
rect 23121 24565 23155 24599
rect 23673 24565 23707 24599
rect 24777 24565 24811 24599
rect 26801 24565 26835 24599
rect 28365 24565 28399 24599
rect 29561 24565 29595 24599
rect 30021 24565 30055 24599
rect 31953 24565 31987 24599
rect 32229 24565 32263 24599
rect 35265 24565 35299 24599
rect 39037 24565 39071 24599
rect 39405 24565 39439 24599
rect 46581 24565 46615 24599
rect 7665 24361 7699 24395
rect 12725 24361 12759 24395
rect 14657 24361 14691 24395
rect 18153 24361 18187 24395
rect 21373 24361 21407 24395
rect 22201 24361 22235 24395
rect 26065 24361 26099 24395
rect 27169 24361 27203 24395
rect 30021 24361 30055 24395
rect 30849 24361 30883 24395
rect 33609 24361 33643 24395
rect 39497 24361 39531 24395
rect 40233 24361 40267 24395
rect 42441 24361 42475 24395
rect 46397 24361 46431 24395
rect 12633 24293 12667 24327
rect 21925 24293 21959 24327
rect 41889 24293 41923 24327
rect 42257 24293 42291 24327
rect 45661 24293 45695 24327
rect 5181 24225 5215 24259
rect 6285 24225 6319 24259
rect 13277 24225 13311 24259
rect 16037 24225 16071 24259
rect 18797 24225 18831 24259
rect 19717 24225 19751 24259
rect 20177 24225 20211 24259
rect 20570 24225 20604 24259
rect 20729 24225 20763 24259
rect 22109 24225 22143 24259
rect 22661 24225 22695 24259
rect 26985 24225 27019 24259
rect 27445 24225 27479 24259
rect 28089 24225 28123 24259
rect 28482 24225 28516 24259
rect 31401 24225 31435 24259
rect 34253 24225 34287 24259
rect 35357 24225 35391 24259
rect 39865 24225 39899 24259
rect 42441 24225 42475 24259
rect 42533 24225 42567 24259
rect 43361 24225 43395 24259
rect 6552 24157 6586 24191
rect 7941 24157 7975 24191
rect 11161 24157 11195 24191
rect 11253 24157 11287 24191
rect 13093 24157 13127 24191
rect 14105 24157 14139 24191
rect 14473 24157 14507 24191
rect 14933 24157 14967 24191
rect 15945 24157 15979 24191
rect 18521 24157 18555 24191
rect 19533 24157 19567 24191
rect 20453 24157 20487 24191
rect 22385 24157 22419 24191
rect 22477 24157 22511 24191
rect 22753 24157 22787 24191
rect 23029 24157 23063 24191
rect 23305 24157 23339 24191
rect 24409 24157 24443 24191
rect 24676 24157 24710 24191
rect 26249 24157 26283 24191
rect 26709 24157 26743 24191
rect 26801 24157 26835 24191
rect 27353 24157 27387 24191
rect 27629 24157 27663 24191
rect 28365 24157 28399 24191
rect 28641 24157 28675 24191
rect 29745 24157 29779 24191
rect 29837 24157 29871 24191
rect 30113 24157 30147 24191
rect 31953 24157 31987 24191
rect 32220 24157 32254 24191
rect 33977 24157 34011 24191
rect 35613 24157 35647 24191
rect 36829 24157 36863 24191
rect 38301 24157 38335 24191
rect 38449 24157 38483 24191
rect 38669 24157 38703 24191
rect 38766 24157 38800 24191
rect 39221 24157 39255 24191
rect 40049 24157 40083 24191
rect 41705 24157 41739 24191
rect 41797 24157 41831 24191
rect 41981 24157 42015 24191
rect 42165 24157 42199 24191
rect 42625 24157 42659 24191
rect 43085 24157 43119 24191
rect 43177 24157 43211 24191
rect 43269 24157 43303 24191
rect 45017 24157 45051 24191
rect 45201 24157 45235 24191
rect 45385 24157 45419 24191
rect 45753 24157 45787 24191
rect 45845 24157 45879 24191
rect 46029 24157 46063 24191
rect 46121 24157 46155 24191
rect 46397 24157 46431 24191
rect 46581 24157 46615 24191
rect 4997 24089 5031 24123
rect 11498 24089 11532 24123
rect 16282 24089 16316 24123
rect 21649 24089 21683 24123
rect 22845 24089 22879 24123
rect 24041 24089 24075 24123
rect 29561 24089 29595 24123
rect 31309 24089 31343 24123
rect 37074 24089 37108 24123
rect 38577 24089 38611 24123
rect 42901 24089 42935 24123
rect 45477 24089 45511 24123
rect 46305 24089 46339 24123
rect 4537 24021 4571 24055
rect 4905 24021 4939 24055
rect 7757 24021 7791 24055
rect 10977 24021 11011 24055
rect 13185 24021 13219 24055
rect 14289 24021 14323 24055
rect 15117 24021 15151 24055
rect 15761 24021 15795 24055
rect 17417 24021 17451 24055
rect 18613 24021 18647 24055
rect 23213 24021 23247 24055
rect 24133 24021 24167 24055
rect 25789 24021 25823 24055
rect 26341 24021 26375 24055
rect 29285 24021 29319 24055
rect 31217 24021 31251 24055
rect 33333 24021 33367 24055
rect 34069 24021 34103 24055
rect 36737 24021 36771 24055
rect 38209 24021 38243 24055
rect 38945 24021 38979 24055
rect 39681 24021 39715 24055
rect 41521 24021 41555 24055
rect 45569 24021 45603 24055
rect 12357 23817 12391 23851
rect 12541 23817 12575 23851
rect 13553 23817 13587 23851
rect 16681 23817 16715 23851
rect 17049 23817 17083 23851
rect 25237 23817 25271 23851
rect 27077 23817 27111 23851
rect 29745 23817 29779 23851
rect 32413 23817 32447 23851
rect 32781 23817 32815 23851
rect 35265 23817 35299 23851
rect 35357 23817 35391 23851
rect 35817 23817 35851 23851
rect 40233 23817 40267 23851
rect 41429 23817 41463 23851
rect 41797 23817 41831 23851
rect 42625 23817 42659 23851
rect 44005 23817 44039 23851
rect 44557 23817 44591 23851
rect 14004 23749 14038 23783
rect 17601 23749 17635 23783
rect 24777 23749 24811 23783
rect 27537 23749 27571 23783
rect 32873 23749 32907 23783
rect 39313 23749 39347 23783
rect 41245 23749 41279 23783
rect 42441 23749 42475 23783
rect 2421 23681 2455 23715
rect 5549 23681 5583 23715
rect 9137 23681 9171 23715
rect 12265 23681 12299 23715
rect 13001 23681 13035 23715
rect 13369 23681 13403 23715
rect 13737 23681 13771 23715
rect 15393 23681 15427 23715
rect 18521 23681 18555 23715
rect 19993 23681 20027 23715
rect 21097 23681 21131 23715
rect 21281 23681 21315 23715
rect 21373 23681 21407 23715
rect 25605 23681 25639 23715
rect 27445 23681 27479 23715
rect 28942 23681 28976 23715
rect 30481 23681 30515 23715
rect 34345 23681 34379 23715
rect 35725 23681 35759 23715
rect 36185 23681 36219 23715
rect 38117 23681 38151 23715
rect 38393 23681 38427 23715
rect 39497 23681 39531 23715
rect 39773 23681 39807 23715
rect 39957 23681 39991 23715
rect 40417 23681 40451 23715
rect 40601 23681 40635 23715
rect 40693 23681 40727 23715
rect 41521 23681 41555 23715
rect 41613 23681 41647 23715
rect 41797 23681 41831 23715
rect 42717 23681 42751 23715
rect 43729 23681 43763 23715
rect 43913 23681 43947 23715
rect 44373 23681 44407 23715
rect 44649 23681 44683 23715
rect 45845 23681 45879 23715
rect 46305 23681 46339 23715
rect 4353 23613 4387 23647
rect 4537 23613 4571 23647
rect 5273 23613 5307 23647
rect 5411 23613 5445 23647
rect 6193 23613 6227 23647
rect 9229 23613 9263 23647
rect 9321 23613 9355 23647
rect 12909 23613 12943 23647
rect 17141 23613 17175 23647
rect 17233 23613 17267 23647
rect 25697 23613 25731 23647
rect 25881 23613 25915 23647
rect 27629 23613 27663 23647
rect 27905 23613 27939 23647
rect 28089 23613 28123 23647
rect 28825 23613 28859 23647
rect 29101 23613 29135 23647
rect 33057 23613 33091 23647
rect 33425 23613 33459 23647
rect 33609 23613 33643 23647
rect 34462 23613 34496 23647
rect 34621 23613 34655 23647
rect 35909 23613 35943 23647
rect 36461 23613 36495 23647
rect 44189 23613 44223 23647
rect 45753 23613 45787 23647
rect 46213 23613 46247 23647
rect 4997 23545 5031 23579
rect 15209 23545 15243 23579
rect 17785 23545 17819 23579
rect 18705 23545 18739 23579
rect 20269 23545 20303 23579
rect 20913 23545 20947 23579
rect 25053 23545 25087 23579
rect 28549 23545 28583 23579
rect 34069 23545 34103 23579
rect 39129 23545 39163 23579
rect 39589 23545 39623 23579
rect 39681 23545 39715 23579
rect 40509 23545 40543 23579
rect 42441 23545 42475 23579
rect 44925 23545 44959 23579
rect 45109 23545 45143 23579
rect 46397 23545 46431 23579
rect 2237 23477 2271 23511
rect 8769 23477 8803 23511
rect 13185 23477 13219 23511
rect 15117 23477 15151 23511
rect 30297 23477 30331 23511
rect 41245 23477 41279 23511
rect 13645 23273 13679 23307
rect 14105 23273 14139 23307
rect 31309 23273 31343 23307
rect 35909 23273 35943 23307
rect 39037 23273 39071 23307
rect 46213 23273 46247 23307
rect 3157 23205 3191 23239
rect 17417 23205 17451 23239
rect 22109 23205 22143 23239
rect 22293 23205 22327 23239
rect 36369 23205 36403 23239
rect 41981 23205 42015 23239
rect 44465 23205 44499 23239
rect 45845 23205 45879 23239
rect 46765 23205 46799 23239
rect 4721 23137 4755 23171
rect 5181 23137 5215 23171
rect 5595 23137 5629 23171
rect 6377 23137 6411 23171
rect 14749 23137 14783 23171
rect 21833 23137 21867 23171
rect 23029 23137 23063 23171
rect 33333 23137 33367 23171
rect 36921 23137 36955 23171
rect 42533 23137 42567 23171
rect 42993 23137 43027 23171
rect 43729 23137 43763 23171
rect 1777 23069 1811 23103
rect 2044 23069 2078 23103
rect 4445 23069 4479 23103
rect 4537 23069 4571 23103
rect 5457 23069 5491 23103
rect 5733 23069 5767 23103
rect 8769 23069 8803 23103
rect 8953 23069 8987 23103
rect 15577 23069 15611 23103
rect 15669 23069 15703 23103
rect 15936 23069 15970 23103
rect 17601 23069 17635 23103
rect 17693 23069 17727 23103
rect 22753 23069 22787 23103
rect 22845 23069 22879 23103
rect 23121 23069 23155 23103
rect 23397 23069 23431 23103
rect 23673 23069 23707 23103
rect 29929 23069 29963 23103
rect 30196 23069 30230 23103
rect 33057 23069 33091 23103
rect 36093 23069 36127 23103
rect 36737 23069 36771 23103
rect 38853 23069 38887 23103
rect 42349 23069 42383 23103
rect 42625 23069 42659 23103
rect 42717 23069 42751 23103
rect 43453 23069 43487 23103
rect 43545 23069 43579 23103
rect 43821 23069 43855 23103
rect 43913 23069 43947 23103
rect 44189 23069 44223 23103
rect 44281 23069 44315 23103
rect 44649 23069 44683 23103
rect 44741 23069 44775 23103
rect 45017 23069 45051 23103
rect 45385 23069 45419 23103
rect 45845 23069 45879 23103
rect 46213 23069 46247 23103
rect 46397 23069 46431 23103
rect 46581 23069 46615 23103
rect 9198 23001 9232 23035
rect 11161 23001 11195 23035
rect 13553 23001 13587 23035
rect 14473 23001 14507 23035
rect 17938 23001 17972 23035
rect 23213 23001 23247 23035
rect 42257 23001 42291 23035
rect 44097 23001 44131 23035
rect 4261 22933 4295 22967
rect 8585 22933 8619 22967
rect 10333 22933 10367 22967
rect 11253 22933 11287 22967
rect 14565 22933 14599 22967
rect 15393 22933 15427 22967
rect 17049 22933 17083 22967
rect 19073 22933 19107 22967
rect 22569 22933 22603 22967
rect 23581 22933 23615 22967
rect 36829 22933 36863 22967
rect 42165 22933 42199 22967
rect 42809 22933 42843 22967
rect 42901 22933 42935 22967
rect 43269 22933 43303 22967
rect 3249 22729 3283 22763
rect 3617 22729 3651 22763
rect 4537 22729 4571 22763
rect 6193 22729 6227 22763
rect 8125 22729 8159 22763
rect 8493 22729 8527 22763
rect 8953 22729 8987 22763
rect 11345 22729 11379 22763
rect 16681 22729 16715 22763
rect 18337 22729 18371 22763
rect 21557 22729 21591 22763
rect 22293 22729 22327 22763
rect 23397 22729 23431 22763
rect 27721 22729 27755 22763
rect 29377 22729 29411 22763
rect 30481 22729 30515 22763
rect 30941 22729 30975 22763
rect 38761 22729 38795 22763
rect 3709 22661 3743 22695
rect 5058 22661 5092 22695
rect 11805 22661 11839 22695
rect 17141 22661 17175 22695
rect 38669 22661 38703 22695
rect 2044 22593 2078 22627
rect 4721 22593 4755 22627
rect 8033 22593 8067 22627
rect 8861 22593 8895 22627
rect 9505 22593 9539 22627
rect 11529 22593 11563 22627
rect 12081 22593 12115 22627
rect 12909 22593 12943 22627
rect 13176 22593 13210 22627
rect 14749 22593 14783 22627
rect 16037 22593 16071 22627
rect 17049 22593 17083 22627
rect 18705 22593 18739 22627
rect 22661 22593 22695 22627
rect 24584 22593 24618 22627
rect 27629 22593 27663 22627
rect 28089 22593 28123 22627
rect 30297 22593 30331 22627
rect 30849 22593 30883 22627
rect 37289 22593 37323 22627
rect 38485 22593 38519 22627
rect 38761 22593 38795 22627
rect 39129 22593 39163 22627
rect 42717 22593 42751 22627
rect 42901 22593 42935 22627
rect 1777 22525 1811 22559
rect 3801 22525 3835 22559
rect 4813 22525 4847 22559
rect 8217 22525 8251 22559
rect 9045 22525 9079 22559
rect 9689 22525 9723 22559
rect 10149 22525 10183 22559
rect 10425 22525 10459 22559
rect 10542 22525 10576 22559
rect 10701 22525 10735 22559
rect 14841 22525 14875 22559
rect 14933 22525 14967 22559
rect 17233 22525 17267 22559
rect 18797 22525 18831 22559
rect 18889 22525 18923 22559
rect 19717 22525 19751 22559
rect 19901 22525 19935 22559
rect 20361 22525 20395 22559
rect 20637 22525 20671 22559
rect 20754 22525 20788 22559
rect 20913 22525 20947 22559
rect 21833 22525 21867 22559
rect 22937 22525 22971 22559
rect 24317 22525 24351 22559
rect 27905 22525 27939 22559
rect 28365 22525 28399 22559
rect 29469 22525 29503 22559
rect 29653 22525 29687 22559
rect 31125 22525 31159 22559
rect 37565 22525 37599 22559
rect 42441 22525 42475 22559
rect 12265 22457 12299 22491
rect 14381 22457 14415 22491
rect 22109 22457 22143 22491
rect 23305 22457 23339 22491
rect 3157 22389 3191 22423
rect 7665 22389 7699 22423
rect 14289 22389 14323 22423
rect 16221 22389 16255 22423
rect 22477 22389 22511 22423
rect 25697 22389 25731 22423
rect 27261 22389 27295 22423
rect 29009 22389 29043 22423
rect 30113 22389 30147 22423
rect 39221 22389 39255 22423
rect 42717 22389 42751 22423
rect 2145 22185 2179 22219
rect 5273 22185 5307 22219
rect 5365 22185 5399 22219
rect 8585 22185 8619 22219
rect 13277 22185 13311 22219
rect 17509 22185 17543 22219
rect 23489 22185 23523 22219
rect 31217 22185 31251 22219
rect 34713 22185 34747 22219
rect 38669 22185 38703 22219
rect 38945 22185 38979 22219
rect 20361 22117 20395 22151
rect 42809 22117 42843 22151
rect 3249 22049 3283 22083
rect 3893 22049 3927 22083
rect 6009 22049 6043 22083
rect 7205 22049 7239 22083
rect 9505 22049 9539 22083
rect 10149 22049 10183 22083
rect 10425 22049 10459 22083
rect 10542 22049 10576 22083
rect 19901 22049 19935 22083
rect 20637 22049 20671 22083
rect 20754 22049 20788 22083
rect 20913 22049 20947 22083
rect 21557 22049 21591 22083
rect 23949 22049 23983 22083
rect 24133 22049 24167 22083
rect 24961 22049 24995 22083
rect 25145 22049 25179 22083
rect 25973 22049 26007 22083
rect 26249 22049 26283 22083
rect 31677 22049 31711 22083
rect 31769 22049 31803 22083
rect 35265 22049 35299 22083
rect 37013 22049 37047 22083
rect 38853 22049 38887 22083
rect 1593 21981 1627 22015
rect 2329 21981 2363 22015
rect 2973 21981 3007 22015
rect 4160 21981 4194 22015
rect 5733 21981 5767 22015
rect 7113 21981 7147 22015
rect 9689 21981 9723 22015
rect 10701 21981 10735 22015
rect 11529 21981 11563 22015
rect 13461 21981 13495 22015
rect 14105 21981 14139 22015
rect 16405 21981 16439 22015
rect 17417 21981 17451 22015
rect 19717 21981 19751 22015
rect 22017 21981 22051 22015
rect 24869 21981 24903 22015
rect 25329 21981 25363 22015
rect 25513 21981 25547 22015
rect 26366 21981 26400 22015
rect 26525 21981 26559 22015
rect 27261 21981 27295 22015
rect 28917 21981 28951 22015
rect 29745 21981 29779 22015
rect 30012 21981 30046 22015
rect 35081 21981 35115 22015
rect 35725 21981 35759 22015
rect 36737 21981 36771 22015
rect 37197 21981 37231 22015
rect 37473 21981 37507 22015
rect 39681 21981 39715 22015
rect 39865 21981 39899 22015
rect 40141 21981 40175 22015
rect 42349 21981 42383 22015
rect 42441 21981 42475 22015
rect 42625 21981 42659 22015
rect 42717 21981 42751 22015
rect 42813 21981 42847 22015
rect 43085 21981 43119 22015
rect 7450 21913 7484 21947
rect 17785 21913 17819 21947
rect 22284 21913 22318 21947
rect 27528 21913 27562 21947
rect 38669 21913 38703 21947
rect 39037 21913 39071 21947
rect 42993 21913 43027 21947
rect 1409 21845 1443 21879
rect 2605 21845 2639 21879
rect 3065 21845 3099 21879
rect 5825 21845 5859 21879
rect 6929 21845 6963 21879
rect 11345 21845 11379 21879
rect 11805 21845 11839 21879
rect 14289 21845 14323 21879
rect 16589 21845 16623 21879
rect 18061 21845 18095 21879
rect 23397 21845 23431 21879
rect 23857 21845 23891 21879
rect 24501 21845 24535 21879
rect 27169 21845 27203 21879
rect 28641 21845 28675 21879
rect 28733 21845 28767 21879
rect 31125 21845 31159 21879
rect 31585 21845 31619 21879
rect 35173 21845 35207 21879
rect 35541 21845 35575 21879
rect 36369 21845 36403 21879
rect 36829 21845 36863 21879
rect 38209 21845 38243 21879
rect 39497 21845 39531 21879
rect 40877 21845 40911 21879
rect 42165 21845 42199 21879
rect 8585 21641 8619 21675
rect 10333 21641 10367 21675
rect 10793 21641 10827 21675
rect 21557 21641 21591 21675
rect 24501 21641 24535 21675
rect 26617 21641 26651 21675
rect 27353 21641 27387 21675
rect 27813 21641 27847 21675
rect 32505 21641 32539 21675
rect 32965 21641 32999 21675
rect 36737 21641 36771 21675
rect 36829 21641 36863 21675
rect 38669 21641 38703 21675
rect 19257 21573 19291 21607
rect 24225 21573 24259 21607
rect 27445 21573 27479 21607
rect 28356 21573 28390 21607
rect 35624 21573 35658 21607
rect 37534 21573 37568 21607
rect 7205 21505 7239 21539
rect 7472 21505 7506 21539
rect 10241 21505 10275 21539
rect 10701 21505 10735 21539
rect 15853 21505 15887 21539
rect 18061 21505 18095 21539
rect 18178 21505 18212 21539
rect 18337 21505 18371 21539
rect 21373 21505 21407 21539
rect 21649 21505 21683 21539
rect 22385 21505 22419 21539
rect 22537 21505 22571 21539
rect 22753 21505 22787 21539
rect 23857 21505 23891 21539
rect 24685 21505 24719 21539
rect 24777 21505 24811 21539
rect 25697 21505 25731 21539
rect 25814 21505 25848 21539
rect 25973 21505 26007 21539
rect 27997 21505 28031 21539
rect 28089 21505 28123 21539
rect 32413 21505 32447 21539
rect 32873 21505 32907 21539
rect 33425 21505 33459 21539
rect 35357 21505 35391 21539
rect 37013 21505 37047 21539
rect 39865 21505 39899 21539
rect 41061 21505 41095 21539
rect 42625 21505 42659 21539
rect 43177 21505 43211 21539
rect 43269 21505 43303 21539
rect 46121 21505 46155 21539
rect 10885 21437 10919 21471
rect 16037 21437 16071 21471
rect 17141 21437 17175 21471
rect 17325 21437 17359 21471
rect 22201 21437 22235 21471
rect 24961 21437 24995 21471
rect 27537 21437 27571 21471
rect 33057 21437 33091 21471
rect 33609 21437 33643 21471
rect 34069 21437 34103 21471
rect 34345 21437 34379 21471
rect 34483 21437 34517 21471
rect 34621 21437 34655 21471
rect 37289 21437 37323 21471
rect 40325 21437 40359 21471
rect 42717 21437 42751 21471
rect 42809 21437 42843 21471
rect 42901 21437 42935 21471
rect 17785 21369 17819 21403
rect 18981 21369 19015 21403
rect 19533 21369 19567 21403
rect 21189 21369 21223 21403
rect 22661 21369 22695 21403
rect 25421 21369 25455 21403
rect 26985 21369 27019 21403
rect 29469 21369 29503 21403
rect 43177 21369 43211 21403
rect 10057 21301 10091 21335
rect 19717 21301 19751 21335
rect 32229 21301 32263 21335
rect 35265 21301 35299 21335
rect 39957 21301 39991 21335
rect 41245 21301 41279 21335
rect 42441 21301 42475 21335
rect 45937 21301 45971 21335
rect 7481 21097 7515 21131
rect 11437 21097 11471 21131
rect 13921 21097 13955 21131
rect 20821 21097 20855 21131
rect 21189 21097 21223 21131
rect 34897 21097 34931 21131
rect 38117 21097 38151 21131
rect 43913 21097 43947 21131
rect 46397 21097 46431 21131
rect 46765 21097 46799 21131
rect 11897 21029 11931 21063
rect 33333 21029 33367 21063
rect 45937 21029 45971 21063
rect 3249 20961 3283 20995
rect 10057 20961 10091 20995
rect 12173 20961 12207 20995
rect 17233 20961 17267 20995
rect 17693 20961 17727 20995
rect 18245 20961 18279 20995
rect 20361 20961 20395 20995
rect 34161 20961 34195 20995
rect 34253 20961 34287 20995
rect 44557 20961 44591 20995
rect 44833 20961 44867 20995
rect 45569 20961 45603 20995
rect 45753 20961 45787 20995
rect 2329 20893 2363 20927
rect 4997 20893 5031 20927
rect 7665 20893 7699 20927
rect 10313 20893 10347 20927
rect 11713 20893 11747 20927
rect 11989 20893 12023 20927
rect 12541 20893 12575 20927
rect 14473 20893 14507 20927
rect 15945 20893 15979 20927
rect 17049 20893 17083 20927
rect 17969 20893 18003 20927
rect 18107 20893 18141 20927
rect 20545 20893 20579 20927
rect 20637 20893 20671 20927
rect 20913 20893 20947 20927
rect 21005 20893 21039 20927
rect 31953 20893 31987 20927
rect 32220 20893 32254 20927
rect 33609 20893 33643 20927
rect 37105 20893 37139 20927
rect 37381 20893 37415 20927
rect 39865 20893 39899 20927
rect 40141 20893 40175 20927
rect 43361 20893 43395 20927
rect 43729 20893 43763 20927
rect 44465 20893 44499 20927
rect 46305 20893 46339 20927
rect 5264 20825 5298 20859
rect 12808 20825 12842 20859
rect 14740 20825 14774 20859
rect 34069 20825 34103 20859
rect 34805 20825 34839 20859
rect 43545 20825 43579 20859
rect 43637 20825 43671 20859
rect 2145 20757 2179 20791
rect 2605 20757 2639 20791
rect 2973 20757 3007 20791
rect 3065 20757 3099 20791
rect 6377 20757 6411 20791
rect 15853 20757 15887 20791
rect 16129 20757 16163 20791
rect 18889 20757 18923 20791
rect 33425 20757 33459 20791
rect 33701 20757 33735 20791
rect 40877 20757 40911 20791
rect 3065 20553 3099 20587
rect 12173 20553 12207 20587
rect 13001 20553 13035 20587
rect 13277 20553 13311 20587
rect 13645 20553 13679 20587
rect 14749 20553 14783 20587
rect 15025 20553 15059 20587
rect 15393 20553 15427 20587
rect 16865 20553 16899 20587
rect 18521 20553 18555 20587
rect 19441 20553 19475 20587
rect 32137 20553 32171 20587
rect 35357 20553 35391 20587
rect 43545 20553 43579 20587
rect 46673 20553 46707 20587
rect 1952 20485 1986 20519
rect 3985 20485 4019 20519
rect 8300 20485 8334 20519
rect 17386 20485 17420 20519
rect 21005 20485 21039 20519
rect 29561 20485 29595 20519
rect 30840 20485 30874 20519
rect 38669 20485 38703 20519
rect 45937 20485 45971 20519
rect 1593 20417 1627 20451
rect 3893 20417 3927 20451
rect 5549 20417 5583 20451
rect 7665 20417 7699 20451
rect 9781 20417 9815 20451
rect 10333 20417 10367 20451
rect 11621 20417 11655 20451
rect 13185 20417 13219 20451
rect 14933 20417 14967 20451
rect 15945 20417 15979 20451
rect 17049 20417 17083 20451
rect 17141 20417 17175 20451
rect 18981 20417 19015 20451
rect 20177 20417 20211 20451
rect 20361 20417 20395 20451
rect 20453 20417 20487 20451
rect 20821 20417 20855 20451
rect 23581 20417 23615 20451
rect 29745 20417 29779 20451
rect 29837 20417 29871 20451
rect 30113 20417 30147 20451
rect 30573 20417 30607 20451
rect 32321 20417 32355 20451
rect 33517 20417 33551 20451
rect 33701 20417 33735 20451
rect 34554 20417 34588 20451
rect 34713 20417 34747 20451
rect 38393 20417 38427 20451
rect 38577 20417 38611 20451
rect 38766 20417 38800 20451
rect 41061 20417 41095 20451
rect 41153 20417 41187 20451
rect 41337 20417 41371 20451
rect 41429 20417 41463 20451
rect 42165 20417 42199 20451
rect 42441 20417 42475 20451
rect 42625 20417 42659 20451
rect 42717 20417 42751 20451
rect 42993 20417 43027 20451
rect 43361 20417 43395 20451
rect 43545 20417 43579 20451
rect 46213 20417 46247 20451
rect 46489 20417 46523 20451
rect 1685 20349 1719 20383
rect 4077 20349 4111 20383
rect 4353 20349 4387 20383
rect 4537 20349 4571 20383
rect 5273 20349 5307 20383
rect 5411 20349 5445 20383
rect 6377 20349 6411 20383
rect 6653 20349 6687 20383
rect 8033 20349 8067 20383
rect 12541 20349 12575 20383
rect 12633 20349 12667 20383
rect 13737 20349 13771 20383
rect 13829 20349 13863 20383
rect 15485 20349 15519 20383
rect 15669 20349 15703 20383
rect 30021 20349 30055 20383
rect 34161 20349 34195 20383
rect 34437 20349 34471 20383
rect 41889 20349 41923 20383
rect 41981 20349 42015 20383
rect 42073 20349 42107 20383
rect 42809 20349 42843 20383
rect 45293 20349 45327 20383
rect 45477 20349 45511 20383
rect 4997 20281 5031 20315
rect 10609 20281 10643 20315
rect 16129 20281 16163 20315
rect 19257 20281 19291 20315
rect 19993 20281 20027 20315
rect 38945 20281 38979 20315
rect 46029 20281 46063 20315
rect 1409 20213 1443 20247
rect 3525 20213 3559 20247
rect 6193 20213 6227 20247
rect 7849 20213 7883 20247
rect 9413 20213 9447 20247
rect 9965 20213 9999 20247
rect 11713 20213 11747 20247
rect 12817 20213 12851 20247
rect 23397 20213 23431 20247
rect 31953 20213 31987 20247
rect 40877 20213 40911 20247
rect 41705 20213 41739 20247
rect 42441 20213 42475 20247
rect 43177 20213 43211 20247
rect 3065 20009 3099 20043
rect 17601 20009 17635 20043
rect 24409 20009 24443 20043
rect 30941 20009 30975 20043
rect 31401 20009 31435 20043
rect 34529 20009 34563 20043
rect 38761 20009 38795 20043
rect 41521 20009 41555 20043
rect 43177 20009 43211 20043
rect 43361 20009 43395 20043
rect 45937 20009 45971 20043
rect 46213 20009 46247 20043
rect 5181 19941 5215 19975
rect 8677 19941 8711 19975
rect 26249 19941 26283 19975
rect 27537 19941 27571 19975
rect 30849 19941 30883 19975
rect 38117 19941 38151 19975
rect 5457 19873 5491 19907
rect 5574 19873 5608 19907
rect 5733 19873 5767 19907
rect 6929 19873 6963 19907
rect 7113 19873 7147 19907
rect 18061 19873 18095 19907
rect 18245 19873 18279 19907
rect 20177 19873 20211 19907
rect 22845 19873 22879 19907
rect 24869 19873 24903 19907
rect 24961 19873 24995 19907
rect 26642 19873 26676 19907
rect 28181 19873 28215 19907
rect 29561 19873 29595 19907
rect 30481 19873 30515 19907
rect 32045 19873 32079 19907
rect 1685 19805 1719 19839
rect 1952 19805 1986 19839
rect 4169 19805 4203 19839
rect 4537 19805 4571 19839
rect 4721 19805 4755 19839
rect 6837 19805 6871 19839
rect 8493 19805 8527 19839
rect 15301 19805 15335 19839
rect 17233 19805 17267 19839
rect 17969 19805 18003 19839
rect 20085 19805 20119 19839
rect 20453 19805 20487 19839
rect 23112 19805 23146 19839
rect 25605 19805 25639 19839
rect 25789 19805 25823 19839
rect 26525 19805 26559 19839
rect 26801 19805 26835 19839
rect 29193 19805 29227 19839
rect 29837 19805 29871 19839
rect 31769 19805 31803 19839
rect 33149 19805 33183 19839
rect 33416 19805 33450 19839
rect 37565 19805 37599 19839
rect 37749 19805 37783 19839
rect 37841 19805 37875 19839
rect 37938 19805 37972 19839
rect 38669 19805 38703 19839
rect 41521 19805 41555 19839
rect 41705 19805 41739 19839
rect 43269 19805 43303 19839
rect 43453 19805 43487 19839
rect 44557 19805 44591 19839
rect 44649 19805 44683 19839
rect 45753 19805 45787 19839
rect 12541 19737 12575 19771
rect 12909 19737 12943 19771
rect 27997 19737 28031 19771
rect 42809 19737 42843 19771
rect 42993 19737 43027 19771
rect 3985 19669 4019 19703
rect 6377 19669 6411 19703
rect 6469 19669 6503 19703
rect 15485 19669 15519 19703
rect 17417 19669 17451 19703
rect 19901 19669 19935 19703
rect 21189 19669 21223 19703
rect 24225 19669 24259 19703
rect 24777 19669 24811 19703
rect 27445 19669 27479 19703
rect 27905 19669 27939 19703
rect 29285 19669 29319 19703
rect 31861 19669 31895 19703
rect 44189 19669 44223 19703
rect 44833 19669 44867 19703
rect 1593 19465 1627 19499
rect 2605 19465 2639 19499
rect 2973 19465 3007 19499
rect 3065 19465 3099 19499
rect 4905 19465 4939 19499
rect 5365 19465 5399 19499
rect 10517 19465 10551 19499
rect 11713 19465 11747 19499
rect 15393 19465 15427 19499
rect 18153 19465 18187 19499
rect 20177 19465 20211 19499
rect 22661 19465 22695 19499
rect 26985 19465 27019 19499
rect 30849 19465 30883 19499
rect 37933 19465 37967 19499
rect 39589 19465 39623 19499
rect 43545 19465 43579 19499
rect 3792 19397 3826 19431
rect 20637 19397 20671 19431
rect 22753 19397 22787 19431
rect 25688 19397 25722 19431
rect 27528 19397 27562 19431
rect 31493 19397 31527 19431
rect 1409 19329 1443 19363
rect 3525 19329 3559 19363
rect 5549 19329 5583 19363
rect 10425 19329 10459 19363
rect 11529 19329 11563 19363
rect 13093 19329 13127 19363
rect 15761 19329 15795 19363
rect 15853 19329 15887 19363
rect 18337 19329 18371 19363
rect 20545 19329 20579 19363
rect 25421 19329 25455 19363
rect 27169 19329 27203 19363
rect 27261 19329 27295 19363
rect 28917 19329 28951 19363
rect 29009 19329 29043 19363
rect 29276 19329 29310 19363
rect 30665 19329 30699 19363
rect 30941 19329 30975 19363
rect 31401 19329 31435 19363
rect 35909 19329 35943 19363
rect 37841 19329 37875 19363
rect 38117 19329 38151 19363
rect 38393 19329 38427 19363
rect 38853 19329 38887 19363
rect 40233 19329 40267 19363
rect 40509 19329 40543 19363
rect 40693 19329 40727 19363
rect 40877 19329 40911 19363
rect 41429 19329 41463 19363
rect 43085 19329 43119 19363
rect 44281 19329 44315 19363
rect 3249 19261 3283 19295
rect 15945 19261 15979 19295
rect 20821 19261 20855 19295
rect 22937 19261 22971 19295
rect 23121 19261 23155 19295
rect 23305 19261 23339 19295
rect 24041 19261 24075 19295
rect 24158 19261 24192 19295
rect 24317 19261 24351 19295
rect 30481 19261 30515 19295
rect 31585 19261 31619 19295
rect 33517 19261 33551 19295
rect 33701 19261 33735 19295
rect 34161 19261 34195 19295
rect 34437 19261 34471 19295
rect 34554 19261 34588 19295
rect 34713 19261 34747 19295
rect 38577 19261 38611 19295
rect 41521 19261 41555 19295
rect 42257 19261 42291 19295
rect 44373 19261 44407 19295
rect 44649 19261 44683 19295
rect 23765 19193 23799 19227
rect 28641 19193 28675 19227
rect 28733 19193 28767 19227
rect 31033 19193 31067 19227
rect 37657 19193 37691 19227
rect 38209 19193 38243 19227
rect 38301 19193 38335 19227
rect 40601 19193 40635 19227
rect 12909 19125 12943 19159
rect 22293 19125 22327 19159
rect 24961 19125 24995 19159
rect 26801 19125 26835 19159
rect 30389 19125 30423 19159
rect 35357 19125 35391 19159
rect 35725 19125 35759 19159
rect 43177 19125 43211 19159
rect 16681 18921 16715 18955
rect 24041 18921 24075 18955
rect 27445 18921 27479 18955
rect 29193 18921 29227 18955
rect 38301 18921 38335 18955
rect 40417 18921 40451 18955
rect 41337 18921 41371 18955
rect 10333 18853 10367 18887
rect 11161 18853 11195 18887
rect 15485 18853 15519 18887
rect 19073 18853 19107 18887
rect 20085 18853 20119 18887
rect 21373 18853 21407 18887
rect 38945 18853 38979 18887
rect 40325 18853 40359 18887
rect 41521 18853 41555 18887
rect 11437 18785 11471 18819
rect 11713 18785 11747 18819
rect 14841 18785 14875 18819
rect 17693 18785 17727 18819
rect 19809 18785 19843 18819
rect 20729 18785 20763 18819
rect 21766 18785 21800 18819
rect 21925 18785 21959 18819
rect 24869 18785 24903 18819
rect 24961 18785 24995 18819
rect 25513 18785 25547 18819
rect 25697 18785 25731 18819
rect 26157 18785 26191 18819
rect 26433 18785 26467 18819
rect 27353 18785 27387 18819
rect 27905 18785 27939 18819
rect 28089 18785 28123 18819
rect 30113 18785 30147 18819
rect 31861 18785 31895 18819
rect 41429 18785 41463 18819
rect 44097 18785 44131 18819
rect 6929 18717 6963 18751
rect 8953 18717 8987 18751
rect 10517 18717 10551 18751
rect 10701 18717 10735 18751
rect 11554 18717 11588 18751
rect 12541 18717 12575 18751
rect 12808 18717 12842 18751
rect 14289 18717 14323 18751
rect 15025 18717 15059 18751
rect 15761 18717 15795 18751
rect 15899 18717 15933 18751
rect 16037 18717 16071 18751
rect 17509 18717 17543 18751
rect 19625 18717 19659 18751
rect 20269 18717 20303 18751
rect 20545 18717 20579 18751
rect 20913 18717 20947 18751
rect 21649 18717 21683 18751
rect 22661 18717 22695 18751
rect 26571 18717 26605 18751
rect 26709 18717 26743 18751
rect 27813 18717 27847 18751
rect 29377 18717 29411 18751
rect 30021 18717 30055 18751
rect 31769 18717 31803 18751
rect 33701 18717 33735 18751
rect 33977 18717 34011 18751
rect 35449 18717 35483 18751
rect 35716 18717 35750 18751
rect 36921 18717 36955 18751
rect 38393 18717 38427 18751
rect 38761 18717 38795 18751
rect 40049 18717 40083 18751
rect 40187 18717 40221 18751
rect 40509 18717 40543 18751
rect 40910 18717 40944 18751
rect 41521 18717 41555 18751
rect 41705 18717 41739 18751
rect 44189 18717 44223 18751
rect 44557 18717 44591 18751
rect 44741 18717 44775 18751
rect 46121 18717 46155 18751
rect 7174 18649 7208 18683
rect 9198 18649 9232 18683
rect 12357 18649 12391 18683
rect 17325 18649 17359 18683
rect 17960 18649 17994 18683
rect 22906 18649 22940 18683
rect 29929 18649 29963 18683
rect 32106 18649 32140 18683
rect 37166 18649 37200 18683
rect 8309 18581 8343 18615
rect 13921 18581 13955 18615
rect 14105 18581 14139 18615
rect 19257 18581 19291 18615
rect 19717 18581 19751 18615
rect 20453 18581 20487 18615
rect 22569 18581 22603 18615
rect 24409 18581 24443 18615
rect 24777 18581 24811 18615
rect 29561 18581 29595 18615
rect 31585 18581 31619 18615
rect 33241 18581 33275 18615
rect 36829 18581 36863 18615
rect 38577 18581 38611 18615
rect 40785 18581 40819 18615
rect 40969 18581 41003 18615
rect 44833 18581 44867 18615
rect 45937 18581 45971 18615
rect 6377 18377 6411 18411
rect 6653 18377 6687 18411
rect 8309 18377 8343 18411
rect 14473 18377 14507 18411
rect 16405 18377 16439 18411
rect 18337 18377 18371 18411
rect 18705 18377 18739 18411
rect 20223 18377 20257 18411
rect 21925 18377 21959 18411
rect 24869 18377 24903 18411
rect 31125 18377 31159 18411
rect 32137 18377 32171 18411
rect 32505 18377 32539 18411
rect 32597 18377 32631 18411
rect 35725 18377 35759 18411
rect 36185 18377 36219 18411
rect 36645 18377 36679 18411
rect 37289 18377 37323 18411
rect 37657 18377 37691 18411
rect 41337 18377 41371 18411
rect 44097 18377 44131 18411
rect 2697 18309 2731 18343
rect 7174 18309 7208 18343
rect 10210 18309 10244 18343
rect 13360 18309 13394 18343
rect 36093 18309 36127 18343
rect 40601 18309 40635 18343
rect 40877 18309 40911 18343
rect 46305 18309 46339 18343
rect 2145 18241 2179 18275
rect 3065 18241 3099 18275
rect 4701 18241 4735 18275
rect 6561 18241 6595 18275
rect 6837 18241 6871 18275
rect 8861 18241 8895 18275
rect 9873 18241 9907 18275
rect 11897 18241 11931 18275
rect 13093 18241 13127 18275
rect 15761 18241 15795 18275
rect 16937 18241 16971 18275
rect 18153 18241 18187 18275
rect 18889 18241 18923 18275
rect 22109 18241 22143 18275
rect 23029 18241 23063 18275
rect 23949 18241 23983 18275
rect 24087 18241 24121 18275
rect 29469 18241 29503 18275
rect 30481 18241 30515 18275
rect 33701 18241 33735 18275
rect 34554 18241 34588 18275
rect 36829 18241 36863 18275
rect 40785 18241 40819 18275
rect 41005 18241 41039 18275
rect 41337 18241 41371 18275
rect 41797 18241 41831 18275
rect 42441 18241 42475 18275
rect 43821 18241 43855 18275
rect 45017 18241 45051 18275
rect 45845 18241 45879 18275
rect 2237 18173 2271 18207
rect 2421 18173 2455 18207
rect 4445 18173 4479 18207
rect 6929 18173 6963 18207
rect 8585 18173 8619 18207
rect 9965 18173 9999 18207
rect 11989 18173 12023 18207
rect 12081 18173 12115 18207
rect 14565 18173 14599 18207
rect 14749 18173 14783 18207
rect 15485 18173 15519 18207
rect 15623 18173 15657 18207
rect 16681 18173 16715 18207
rect 19993 18173 20027 18207
rect 23213 18173 23247 18207
rect 24225 18173 24259 18207
rect 29285 18173 29319 18207
rect 30205 18173 30239 18207
rect 30322 18173 30356 18207
rect 32689 18173 32723 18207
rect 33517 18173 33551 18207
rect 34437 18173 34471 18207
rect 34713 18173 34747 18207
rect 36277 18173 36311 18207
rect 37749 18173 37783 18207
rect 37841 18173 37875 18207
rect 40693 18173 40727 18207
rect 41153 18173 41187 18207
rect 41705 18173 41739 18207
rect 42073 18173 42107 18207
rect 42901 18173 42935 18207
rect 44097 18173 44131 18207
rect 44925 18173 44959 18207
rect 45385 18173 45419 18207
rect 45661 18173 45695 18207
rect 1777 18105 1811 18139
rect 9689 18105 9723 18139
rect 11529 18105 11563 18139
rect 15209 18105 15243 18139
rect 23673 18105 23707 18139
rect 29929 18105 29963 18139
rect 34161 18105 34195 18139
rect 41889 18105 41923 18139
rect 5825 18037 5859 18071
rect 11345 18037 11379 18071
rect 18061 18037 18095 18071
rect 35357 18037 35391 18071
rect 41981 18037 42015 18071
rect 42533 18037 42567 18071
rect 43913 18037 43947 18071
rect 2973 17833 3007 17867
rect 3893 17833 3927 17867
rect 6285 17833 6319 17867
rect 7573 17833 7607 17867
rect 8585 17833 8619 17867
rect 8953 17833 8987 17867
rect 13093 17833 13127 17867
rect 16313 17833 16347 17867
rect 16589 17833 16623 17867
rect 20545 17833 20579 17867
rect 45845 17833 45879 17867
rect 46213 17833 46247 17867
rect 6009 17765 6043 17799
rect 28641 17765 28675 17799
rect 30481 17765 30515 17799
rect 31677 17765 31711 17799
rect 38393 17765 38427 17799
rect 4353 17697 4387 17731
rect 4813 17697 4847 17731
rect 8125 17697 8159 17731
rect 9505 17697 9539 17731
rect 10517 17697 10551 17731
rect 10977 17697 11011 17731
rect 13645 17697 13679 17731
rect 14381 17697 14415 17731
rect 17233 17697 17267 17731
rect 29101 17697 29135 17731
rect 29193 17697 29227 17731
rect 29837 17697 29871 17731
rect 30021 17697 30055 17731
rect 30757 17697 30791 17731
rect 35265 17697 35299 17731
rect 1593 17629 1627 17663
rect 3341 17629 3375 17663
rect 4077 17629 4111 17663
rect 4169 17629 4203 17663
rect 5089 17629 5123 17663
rect 5227 17629 5261 17663
rect 5365 17629 5399 17663
rect 6193 17629 6227 17663
rect 7021 17629 7055 17663
rect 7941 17629 7975 17663
rect 8769 17629 8803 17663
rect 9321 17629 9355 17663
rect 10333 17629 10367 17663
rect 11253 17629 11287 17663
rect 11370 17629 11404 17663
rect 11529 17629 11563 17663
rect 12173 17629 12207 17663
rect 13461 17629 13495 17663
rect 14105 17629 14139 17663
rect 15393 17629 15427 17663
rect 15669 17629 15703 17663
rect 16497 17629 16531 17663
rect 16957 17629 16991 17663
rect 23213 17629 23247 17663
rect 26617 17629 26651 17663
rect 29745 17629 29779 17663
rect 30874 17629 30908 17663
rect 31033 17629 31067 17663
rect 37841 17629 37875 17663
rect 38214 17629 38248 17663
rect 38669 17629 38703 17663
rect 44189 17629 44223 17663
rect 44281 17629 44315 17663
rect 44373 17629 44407 17663
rect 44557 17629 44591 17663
rect 45753 17629 45787 17663
rect 46397 17629 46431 17663
rect 46765 17629 46799 17663
rect 1860 17561 1894 17595
rect 17049 17561 17083 17595
rect 20453 17561 20487 17595
rect 35081 17561 35115 17595
rect 38025 17561 38059 17595
rect 38117 17561 38151 17595
rect 39681 17561 39715 17595
rect 3157 17493 3191 17527
rect 7205 17493 7239 17527
rect 8033 17493 8067 17527
rect 9413 17493 9447 17527
rect 13553 17493 13587 17527
rect 23029 17493 23063 17527
rect 26433 17493 26467 17527
rect 29009 17493 29043 17527
rect 29561 17493 29595 17527
rect 34713 17493 34747 17527
rect 35173 17493 35207 17527
rect 43913 17493 43947 17527
rect 1409 17289 1443 17323
rect 6745 17289 6779 17323
rect 7481 17289 7515 17323
rect 7849 17289 7883 17323
rect 14197 17289 14231 17323
rect 14565 17289 14599 17323
rect 14657 17289 14691 17323
rect 21281 17289 21315 17323
rect 24041 17289 24075 17323
rect 25881 17289 25915 17323
rect 26341 17289 26375 17323
rect 28365 17289 28399 17323
rect 29929 17289 29963 17323
rect 33425 17289 33459 17323
rect 38301 17289 38335 17323
rect 40141 17289 40175 17323
rect 42533 17289 42567 17323
rect 42625 17289 42659 17323
rect 44557 17289 44591 17323
rect 22928 17221 22962 17255
rect 24768 17221 24802 17255
rect 27230 17221 27264 17255
rect 28816 17221 28850 17255
rect 31585 17221 31619 17255
rect 40601 17221 40635 17255
rect 1593 17153 1627 17187
rect 2320 17153 2354 17187
rect 4353 17153 4387 17187
rect 6561 17153 6595 17187
rect 7941 17153 7975 17187
rect 19257 17153 19291 17187
rect 20545 17153 20579 17187
rect 21557 17153 21591 17187
rect 22661 17153 22695 17187
rect 24501 17153 24535 17187
rect 31677 17153 31711 17187
rect 34345 17153 34379 17187
rect 35449 17153 35483 17187
rect 37565 17153 37599 17187
rect 38577 17153 38611 17187
rect 38669 17153 38703 17187
rect 38853 17153 38887 17187
rect 38945 17153 38979 17187
rect 39957 17153 39991 17187
rect 40233 17153 40267 17187
rect 40785 17153 40819 17187
rect 40969 17153 41003 17187
rect 42441 17153 42475 17187
rect 44097 17153 44131 17187
rect 44741 17153 44775 17187
rect 45293 17153 45327 17187
rect 45385 17153 45419 17187
rect 2053 17085 2087 17119
rect 4169 17085 4203 17119
rect 5089 17085 5123 17119
rect 5227 17085 5261 17119
rect 5365 17085 5399 17119
rect 8033 17085 8067 17119
rect 14749 17085 14783 17119
rect 18061 17085 18095 17119
rect 18245 17085 18279 17119
rect 18981 17085 19015 17119
rect 19119 17085 19153 17119
rect 20269 17085 20303 17119
rect 26433 17085 26467 17119
rect 26617 17085 26651 17119
rect 26985 17085 27019 17119
rect 28549 17085 28583 17119
rect 31861 17085 31895 17119
rect 33517 17085 33551 17119
rect 33609 17085 33643 17119
rect 37289 17085 37323 17119
rect 41061 17085 41095 17119
rect 42809 17085 42843 17119
rect 45017 17085 45051 17119
rect 45569 17085 45603 17119
rect 4813 17017 4847 17051
rect 6009 17017 6043 17051
rect 18705 17017 18739 17051
rect 34575 17017 34609 17051
rect 39957 17017 39991 17051
rect 44925 17017 44959 17051
rect 3433 16949 3467 16983
rect 19901 16949 19935 16983
rect 21557 16949 21591 16983
rect 25973 16949 26007 16983
rect 31217 16949 31251 16983
rect 33057 16949 33091 16983
rect 35265 16949 35299 16983
rect 38393 16949 38427 16983
rect 42533 16949 42567 16983
rect 44189 16949 44223 16983
rect 45477 16949 45511 16983
rect 2513 16745 2547 16779
rect 5089 16745 5123 16779
rect 12633 16745 12667 16779
rect 18337 16745 18371 16779
rect 20361 16745 20395 16779
rect 20821 16745 20855 16779
rect 23213 16745 23247 16779
rect 24869 16745 24903 16779
rect 26433 16745 26467 16779
rect 32137 16745 32171 16779
rect 34345 16745 34379 16779
rect 43453 16745 43487 16779
rect 44741 16745 44775 16779
rect 45017 16745 45051 16779
rect 13369 16677 13403 16711
rect 20085 16677 20119 16711
rect 20269 16677 20303 16711
rect 40785 16677 40819 16711
rect 41981 16677 42015 16711
rect 44557 16677 44591 16711
rect 4353 16609 4387 16643
rect 5733 16609 5767 16643
rect 9413 16609 9447 16643
rect 12357 16609 12391 16643
rect 12449 16609 12483 16643
rect 13093 16609 13127 16643
rect 13185 16609 13219 16643
rect 15577 16609 15611 16643
rect 23673 16609 23707 16643
rect 23857 16609 23891 16643
rect 26893 16609 26927 16643
rect 27077 16609 27111 16643
rect 32965 16609 32999 16643
rect 34713 16609 34747 16643
rect 38025 16609 38059 16643
rect 42625 16609 42659 16643
rect 43361 16609 43395 16643
rect 45109 16609 45143 16643
rect 45661 16609 45695 16643
rect 45937 16609 45971 16643
rect 2697 16541 2731 16575
rect 4169 16541 4203 16575
rect 5457 16541 5491 16575
rect 14841 16541 14875 16575
rect 16957 16541 16991 16575
rect 19809 16541 19843 16575
rect 20545 16541 20579 16575
rect 20637 16541 20671 16575
rect 20913 16541 20947 16575
rect 23581 16541 23615 16575
rect 25053 16541 25087 16575
rect 26801 16541 26835 16575
rect 30757 16541 30791 16575
rect 32873 16541 32907 16575
rect 37105 16541 37139 16575
rect 37289 16541 37323 16575
rect 38301 16541 38335 16575
rect 38485 16541 38519 16575
rect 38853 16541 38887 16575
rect 40049 16541 40083 16575
rect 40233 16541 40267 16575
rect 40417 16541 40451 16575
rect 40693 16541 40727 16575
rect 40877 16541 40911 16575
rect 40969 16541 41003 16575
rect 41245 16541 41279 16575
rect 41337 16541 41371 16575
rect 41981 16541 42015 16575
rect 42165 16541 42199 16575
rect 42349 16541 42383 16575
rect 42533 16541 42567 16575
rect 42809 16541 42843 16575
rect 42993 16541 43027 16575
rect 43177 16541 43211 16575
rect 43637 16541 43671 16575
rect 43821 16541 43855 16575
rect 45017 16541 45051 16575
rect 9680 16473 9714 16507
rect 17224 16473 17258 16507
rect 31024 16473 31058 16507
rect 33210 16473 33244 16507
rect 34958 16473 34992 16507
rect 40325 16473 40359 16507
rect 41521 16473 41555 16507
rect 43545 16473 43579 16507
rect 44281 16473 44315 16507
rect 45753 16473 45787 16507
rect 3801 16405 3835 16439
rect 4261 16405 4295 16439
rect 5549 16405 5583 16439
rect 10793 16405 10827 16439
rect 11989 16405 12023 16439
rect 12725 16405 12759 16439
rect 14657 16405 14691 16439
rect 14933 16405 14967 16439
rect 15301 16405 15335 16439
rect 15393 16405 15427 16439
rect 32689 16405 32723 16439
rect 36093 16405 36127 16439
rect 38945 16405 38979 16439
rect 40509 16405 40543 16439
rect 43269 16405 43303 16439
rect 43729 16405 43763 16439
rect 45385 16405 45419 16439
rect 3709 16201 3743 16235
rect 4169 16201 4203 16235
rect 10701 16201 10735 16235
rect 11805 16201 11839 16235
rect 13553 16201 13587 16235
rect 13921 16201 13955 16235
rect 17233 16201 17267 16235
rect 17509 16201 17543 16235
rect 17969 16201 18003 16235
rect 21189 16201 21223 16235
rect 28089 16201 28123 16235
rect 31125 16201 31159 16235
rect 33517 16201 33551 16235
rect 34069 16201 34103 16235
rect 35725 16201 35759 16235
rect 40049 16201 40083 16235
rect 42901 16201 42935 16235
rect 45385 16201 45419 16235
rect 7021 16133 7055 16167
rect 10609 16133 10643 16167
rect 12326 16133 12360 16167
rect 14013 16133 14047 16167
rect 23489 16133 23523 16167
rect 23857 16133 23891 16167
rect 34612 16133 34646 16167
rect 2329 16065 2363 16099
rect 2596 16065 2630 16099
rect 4261 16065 4295 16099
rect 6561 16065 6595 16099
rect 9965 16065 9999 16099
rect 10885 16065 10919 16099
rect 11989 16065 12023 16099
rect 14473 16065 14507 16099
rect 14740 16065 14774 16099
rect 16221 16065 16255 16099
rect 17417 16065 17451 16099
rect 17877 16065 17911 16099
rect 18521 16065 18555 16099
rect 19374 16065 19408 16099
rect 21373 16065 21407 16099
rect 21557 16065 21591 16099
rect 21649 16065 21683 16099
rect 22385 16065 22419 16099
rect 22477 16065 22511 16099
rect 22753 16065 22787 16099
rect 23029 16065 23063 16099
rect 23121 16065 23155 16099
rect 23397 16065 23431 16099
rect 23673 16065 23707 16099
rect 23949 16065 23983 16099
rect 24869 16065 24903 16099
rect 24961 16065 24995 16099
rect 25237 16065 25271 16099
rect 26525 16065 26559 16099
rect 27077 16065 27111 16099
rect 27905 16065 27939 16099
rect 28273 16065 28307 16099
rect 29009 16065 29043 16099
rect 31309 16065 31343 16099
rect 32137 16065 32171 16099
rect 32404 16065 32438 16099
rect 34253 16065 34287 16099
rect 34345 16065 34379 16099
rect 37565 16065 37599 16099
rect 39589 16065 39623 16099
rect 40141 16065 40175 16099
rect 40785 16065 40819 16099
rect 41245 16065 41279 16099
rect 42533 16065 42567 16099
rect 42717 16065 42751 16099
rect 42993 16065 43027 16099
rect 45017 16065 45051 16099
rect 45753 16065 45787 16099
rect 46489 16065 46523 16099
rect 4445 15997 4479 16031
rect 7113 15997 7147 16031
rect 7205 15997 7239 16031
rect 8769 15997 8803 16031
rect 8953 15997 8987 16031
rect 9689 15997 9723 16031
rect 9806 15997 9840 16031
rect 12081 15997 12115 16031
rect 14105 15997 14139 16031
rect 18061 15997 18095 16031
rect 18337 15997 18371 16031
rect 19257 15997 19291 16031
rect 19533 15997 19567 16031
rect 24133 15997 24167 16031
rect 24685 15997 24719 16031
rect 37289 15997 37323 16031
rect 40693 15997 40727 16031
rect 41337 15997 41371 16031
rect 43085 15997 43119 16031
rect 43269 15997 43303 16031
rect 45109 15997 45143 16031
rect 45477 15997 45511 16031
rect 6653 15929 6687 15963
rect 9413 15929 9447 15963
rect 13461 15929 13495 15963
rect 15853 15929 15887 15963
rect 18981 15929 19015 15963
rect 20177 15929 20211 15963
rect 24409 15929 24443 15963
rect 24593 15929 24627 15963
rect 25145 15929 25179 15963
rect 27353 15929 27387 15963
rect 38301 15929 38335 15963
rect 39773 15929 39807 15963
rect 3801 15861 3835 15895
rect 6377 15861 6411 15895
rect 16313 15861 16347 15895
rect 22201 15861 22235 15895
rect 22661 15861 22695 15895
rect 22845 15861 22879 15895
rect 23305 15861 23339 15895
rect 26709 15861 26743 15895
rect 28457 15861 28491 15895
rect 29193 15861 29227 15895
rect 43177 15861 43211 15895
rect 46673 15861 46707 15895
rect 2789 15657 2823 15691
rect 10793 15657 10827 15691
rect 22109 15657 22143 15691
rect 32413 15657 32447 15691
rect 34713 15657 34747 15691
rect 36369 15657 36403 15691
rect 37933 15657 37967 15691
rect 46213 15657 46247 15691
rect 7205 15589 7239 15623
rect 8033 15589 8067 15623
rect 14565 15589 14599 15623
rect 17141 15589 17175 15623
rect 17509 15589 17543 15623
rect 20361 15589 20395 15623
rect 21557 15589 21591 15623
rect 21925 15589 21959 15623
rect 31585 15589 31619 15623
rect 4813 15521 4847 15555
rect 8585 15521 8619 15555
rect 9137 15521 9171 15555
rect 9597 15521 9631 15555
rect 9873 15521 9907 15555
rect 10149 15521 10183 15555
rect 12173 15521 12207 15555
rect 14841 15521 14875 15555
rect 18061 15521 18095 15555
rect 19901 15521 19935 15555
rect 20637 15521 20671 15555
rect 20913 15521 20947 15555
rect 29561 15521 29595 15555
rect 32137 15521 32171 15555
rect 35265 15521 35299 15555
rect 39589 15521 39623 15555
rect 40049 15521 40083 15555
rect 45569 15521 45603 15555
rect 2973 15453 3007 15487
rect 4537 15453 4571 15487
rect 5733 15453 5767 15487
rect 5825 15453 5859 15487
rect 7941 15453 7975 15487
rect 8401 15453 8435 15487
rect 8953 15453 8987 15487
rect 9990 15453 10024 15487
rect 14749 15453 14783 15487
rect 17417 15453 17451 15487
rect 17969 15453 18003 15487
rect 19717 15453 19751 15487
rect 20754 15453 20788 15487
rect 21649 15453 21683 15487
rect 26065 15453 26099 15487
rect 29377 15453 29411 15487
rect 32597 15453 32631 15487
rect 35081 15453 35115 15487
rect 35173 15453 35207 15487
rect 36185 15453 36219 15487
rect 36921 15453 36955 15487
rect 37197 15453 37231 15487
rect 40325 15453 40359 15487
rect 45293 15453 45327 15487
rect 46397 15453 46431 15487
rect 6070 15385 6104 15419
rect 8493 15385 8527 15419
rect 12440 15385 12474 15419
rect 15086 15385 15120 15419
rect 16957 15385 16991 15419
rect 17877 15385 17911 15419
rect 26332 15385 26366 15419
rect 29806 15385 29840 15419
rect 39405 15385 39439 15419
rect 4169 15317 4203 15351
rect 4629 15317 4663 15351
rect 5549 15317 5583 15351
rect 7757 15317 7791 15351
rect 13553 15317 13587 15351
rect 16221 15317 16255 15351
rect 17233 15317 17267 15351
rect 27445 15317 27479 15351
rect 29193 15317 29227 15351
rect 30941 15317 30975 15351
rect 31953 15317 31987 15351
rect 32045 15317 32079 15351
rect 4813 15113 4847 15147
rect 9321 15113 9355 15147
rect 9781 15113 9815 15147
rect 12541 15113 12575 15147
rect 12817 15113 12851 15147
rect 13185 15113 13219 15147
rect 15301 15113 15335 15147
rect 15669 15113 15703 15147
rect 18337 15113 18371 15147
rect 21557 15113 21591 15147
rect 23121 15113 23155 15147
rect 26341 15113 26375 15147
rect 26985 15113 27019 15147
rect 29285 15113 29319 15147
rect 29653 15113 29687 15147
rect 42533 15113 42567 15147
rect 45661 15113 45695 15147
rect 6622 15045 6656 15079
rect 8186 15045 8220 15079
rect 10149 15045 10183 15079
rect 10241 15045 10275 15079
rect 13277 15045 13311 15079
rect 15761 15045 15795 15079
rect 17224 15045 17258 15079
rect 21097 15045 21131 15079
rect 3433 14977 3467 15011
rect 3700 14977 3734 15011
rect 7941 14977 7975 15011
rect 12725 14977 12759 15011
rect 16957 14977 16991 15011
rect 19349 14977 19383 15011
rect 20085 14977 20119 15011
rect 20361 14977 20395 15011
rect 26525 14977 26559 15011
rect 27353 14977 27387 15011
rect 29193 14977 29227 15011
rect 33793 14977 33827 15011
rect 35541 14977 35575 15011
rect 38853 14977 38887 15011
rect 38945 14977 38979 15011
rect 39129 14977 39163 15011
rect 39313 14977 39347 15011
rect 39405 14977 39439 15011
rect 41337 14977 41371 15011
rect 42717 14977 42751 15011
rect 43177 14977 43211 15011
rect 43361 14977 43395 15011
rect 43729 14977 43763 15011
rect 43821 14977 43855 15011
rect 44005 14977 44039 15011
rect 45201 14977 45235 15011
rect 6377 14909 6411 14943
rect 10425 14909 10459 14943
rect 13461 14909 13495 14943
rect 15945 14909 15979 14943
rect 19165 14909 19199 14943
rect 20223 14909 20257 14943
rect 22661 14909 22695 14943
rect 27445 14909 27479 14943
rect 27537 14909 27571 14943
rect 29745 14909 29779 14943
rect 29837 14909 29871 14943
rect 35817 14909 35851 14943
rect 39865 14909 39899 14943
rect 19809 14841 19843 14875
rect 21005 14841 21039 14875
rect 21373 14841 21407 14875
rect 23029 14841 23063 14875
rect 39037 14841 39071 14875
rect 43637 14841 43671 14875
rect 7757 14773 7791 14807
rect 29009 14773 29043 14807
rect 33977 14773 34011 14807
rect 38669 14773 38703 14807
rect 39681 14773 39715 14807
rect 41153 14773 41187 14807
rect 43913 14773 43947 14807
rect 45477 14773 45511 14807
rect 3893 14569 3927 14603
rect 6561 14569 6595 14603
rect 24409 14569 24443 14603
rect 27813 14569 27847 14603
rect 28641 14569 28675 14603
rect 30665 14569 30699 14603
rect 31493 14569 31527 14603
rect 37197 14569 37231 14603
rect 38025 14569 38059 14603
rect 40233 14569 40267 14603
rect 41245 14569 41279 14603
rect 41981 14569 42015 14603
rect 42165 14569 42199 14603
rect 43821 14569 43855 14603
rect 7113 14433 7147 14467
rect 18521 14433 18555 14467
rect 19901 14433 19935 14467
rect 22293 14433 22327 14467
rect 25053 14433 25087 14467
rect 26617 14433 26651 14467
rect 27010 14433 27044 14467
rect 28549 14433 28583 14467
rect 29101 14433 29135 14467
rect 29193 14433 29227 14467
rect 31217 14433 31251 14467
rect 32045 14433 32079 14467
rect 33885 14433 33919 14467
rect 38209 14433 38243 14467
rect 40601 14433 40635 14467
rect 1409 14365 1443 14399
rect 4077 14365 4111 14399
rect 7021 14365 7055 14399
rect 12265 14365 12299 14399
rect 15853 14365 15887 14399
rect 18245 14365 18279 14399
rect 20177 14365 20211 14399
rect 20913 14365 20947 14399
rect 25605 14365 25639 14399
rect 25973 14365 26007 14399
rect 26157 14365 26191 14399
rect 26893 14365 26927 14399
rect 27169 14365 27203 14399
rect 28365 14365 28399 14399
rect 29561 14365 29595 14399
rect 33609 14365 33643 14399
rect 35817 14365 35851 14399
rect 38301 14365 38335 14399
rect 39865 14365 39899 14399
rect 40049 14365 40083 14399
rect 40877 14365 40911 14399
rect 40974 14365 41008 14399
rect 41153 14365 41187 14399
rect 41705 14365 41739 14399
rect 43177 14365 43211 14399
rect 43545 14365 43579 14399
rect 6929 14297 6963 14331
rect 12449 14297 12483 14331
rect 16129 14297 16163 14331
rect 23305 14297 23339 14331
rect 23673 14297 23707 14331
rect 29009 14297 29043 14331
rect 31125 14297 31159 14331
rect 36084 14297 36118 14331
rect 38025 14297 38059 14331
rect 38393 14297 38427 14331
rect 40601 14297 40635 14331
rect 40785 14297 40819 14331
rect 1593 14229 1627 14263
rect 21005 14229 21039 14263
rect 21741 14229 21775 14263
rect 22109 14229 22143 14263
rect 22201 14229 22235 14263
rect 24777 14229 24811 14263
rect 24869 14229 24903 14263
rect 25421 14229 25455 14263
rect 29791 14229 29825 14263
rect 31033 14229 31067 14263
rect 31861 14229 31895 14263
rect 31953 14229 31987 14263
rect 41613 14229 41647 14263
rect 43269 14229 43303 14263
rect 44005 14229 44039 14263
rect 21097 14025 21131 14059
rect 28825 14025 28859 14059
rect 31585 14025 31619 14059
rect 32137 14025 32171 14059
rect 32505 14025 32539 14059
rect 35265 14025 35299 14059
rect 35449 14025 35483 14059
rect 37657 14025 37691 14059
rect 37749 14025 37783 14059
rect 40141 14025 40175 14059
rect 41613 14025 41647 14059
rect 42993 14025 43027 14059
rect 44005 14025 44039 14059
rect 10241 13957 10275 13991
rect 13277 13957 13311 13991
rect 22569 13957 22603 13991
rect 25412 13957 25446 13991
rect 35970 13957 36004 13991
rect 7113 13889 7147 13923
rect 9505 13889 9539 13923
rect 12541 13889 12575 13923
rect 12633 13889 12667 13923
rect 13461 13889 13495 13923
rect 15301 13889 15335 13923
rect 19717 13889 19751 13923
rect 19984 13889 20018 13923
rect 23397 13889 23431 13923
rect 25145 13889 25179 13923
rect 28181 13889 28215 13923
rect 29285 13889 29319 13923
rect 30665 13889 30699 13923
rect 30782 13889 30816 13923
rect 30941 13889 30975 13923
rect 31953 13889 31987 13923
rect 32597 13889 32631 13923
rect 34621 13889 34655 13923
rect 35633 13889 35667 13923
rect 40325 13889 40359 13923
rect 41153 13889 41187 13923
rect 42809 13889 42843 13923
rect 43085 13889 43119 13923
rect 43453 13889 43487 13923
rect 44189 13889 44223 13923
rect 45017 13889 45051 13923
rect 12173 13821 12207 13855
rect 12817 13821 12851 13855
rect 26985 13821 27019 13855
rect 27169 13821 27203 13855
rect 27905 13821 27939 13855
rect 28022 13821 28056 13855
rect 29377 13821 29411 13855
rect 29561 13821 29595 13855
rect 29745 13821 29779 13855
rect 29929 13821 29963 13855
rect 32689 13821 32723 13855
rect 33425 13821 33459 13855
rect 33609 13821 33643 13855
rect 34069 13821 34103 13855
rect 34345 13821 34379 13855
rect 34462 13821 34496 13855
rect 35725 13821 35759 13855
rect 37841 13821 37875 13855
rect 40969 13821 41003 13855
rect 43269 13821 43303 13855
rect 22753 13753 22787 13787
rect 27629 13753 27663 13787
rect 30389 13753 30423 13787
rect 6929 13685 6963 13719
rect 9321 13685 9355 13719
rect 10333 13685 10367 13719
rect 15117 13685 15151 13719
rect 23581 13685 23615 13719
rect 26525 13685 26559 13719
rect 28917 13685 28951 13719
rect 31769 13685 31803 13719
rect 37105 13685 37139 13719
rect 37289 13685 37323 13719
rect 42809 13685 42843 13719
rect 43637 13685 43671 13719
rect 45293 13685 45327 13719
rect 45477 13685 45511 13719
rect 9045 13481 9079 13515
rect 20269 13481 20303 13515
rect 21465 13481 21499 13515
rect 24225 13481 24259 13515
rect 25513 13481 25547 13515
rect 28825 13481 28859 13515
rect 31769 13481 31803 13515
rect 33241 13481 33275 13515
rect 36185 13481 36219 13515
rect 20729 13413 20763 13447
rect 29101 13413 29135 13447
rect 30573 13413 30607 13447
rect 33517 13413 33551 13447
rect 42993 13413 43027 13447
rect 6469 13345 6503 13379
rect 9321 13345 9355 13379
rect 14749 13345 14783 13379
rect 23029 13345 23063 13379
rect 23581 13345 23615 13379
rect 25053 13345 25087 13379
rect 26157 13345 26191 13379
rect 30113 13345 30147 13379
rect 30849 13345 30883 13379
rect 30966 13345 31000 13379
rect 31125 13345 31159 13379
rect 31861 13345 31895 13379
rect 34253 13345 34287 13379
rect 34345 13345 34379 13379
rect 36829 13345 36863 13379
rect 4445 13277 4479 13311
rect 9229 13277 9263 13311
rect 10977 13277 11011 13311
rect 11713 13277 11747 13311
rect 11805 13277 11839 13311
rect 14657 13277 14691 13311
rect 15016 13277 15050 13311
rect 16865 13277 16899 13311
rect 20453 13277 20487 13311
rect 20913 13277 20947 13311
rect 21189 13277 21223 13311
rect 22385 13277 22419 13311
rect 22569 13277 22603 13311
rect 23305 13277 23339 13311
rect 23422 13277 23456 13311
rect 24869 13277 24903 13311
rect 25881 13277 25915 13311
rect 27445 13277 27479 13311
rect 29285 13277 29319 13311
rect 29929 13277 29963 13311
rect 32117 13277 32151 13311
rect 33701 13277 33735 13311
rect 34713 13277 34747 13311
rect 34969 13277 35003 13311
rect 36553 13277 36587 13311
rect 37381 13277 37415 13311
rect 43177 13277 43211 13311
rect 43269 13277 43303 13311
rect 45477 13277 45511 13311
rect 46489 13277 46523 13311
rect 6736 13209 6770 13243
rect 9588 13209 9622 13243
rect 12050 13209 12084 13243
rect 17110 13209 17144 13243
rect 21373 13209 21407 13243
rect 25973 13209 26007 13243
rect 27712 13209 27746 13243
rect 34161 13209 34195 13243
rect 42993 13209 43027 13243
rect 4261 13141 4295 13175
rect 7849 13141 7883 13175
rect 10701 13141 10735 13175
rect 10793 13141 10827 13175
rect 11529 13141 11563 13175
rect 13185 13141 13219 13175
rect 14473 13141 14507 13175
rect 16129 13141 16163 13175
rect 18245 13141 18279 13175
rect 21097 13141 21131 13175
rect 24409 13141 24443 13175
rect 24777 13141 24811 13175
rect 33793 13141 33827 13175
rect 36093 13141 36127 13175
rect 36645 13141 36679 13175
rect 37473 13141 37507 13175
rect 45293 13141 45327 13175
rect 46673 13141 46707 13175
rect 5181 12937 5215 12971
rect 10425 12937 10459 12971
rect 10793 12937 10827 12971
rect 13461 12937 13495 12971
rect 13829 12937 13863 12971
rect 15761 12937 15795 12971
rect 16129 12937 16163 12971
rect 16865 12937 16899 12971
rect 19073 12937 19107 12971
rect 19441 12937 19475 12971
rect 24869 12937 24903 12971
rect 30205 12937 30239 12971
rect 35081 12937 35115 12971
rect 36093 12937 36127 12971
rect 39681 12937 39715 12971
rect 42809 12937 42843 12971
rect 3976 12869 4010 12903
rect 9220 12869 9254 12903
rect 10885 12869 10919 12903
rect 19901 12869 19935 12903
rect 1501 12801 1535 12835
rect 5549 12801 5583 12835
rect 6377 12801 6411 12835
rect 8953 12801 8987 12835
rect 11529 12801 11563 12835
rect 11713 12801 11747 12835
rect 12725 12801 12759 12835
rect 14289 12801 14323 12835
rect 14556 12801 14590 12835
rect 17049 12801 17083 12835
rect 17325 12801 17359 12835
rect 18178 12801 18212 12835
rect 18337 12801 18371 12835
rect 19533 12801 19567 12835
rect 20913 12801 20947 12835
rect 21097 12801 21131 12835
rect 21189 12801 21223 12835
rect 25145 12801 25179 12835
rect 27905 12801 27939 12835
rect 29092 12801 29126 12835
rect 33241 12801 33275 12835
rect 34161 12801 34195 12835
rect 34299 12801 34333 12835
rect 36277 12801 36311 12835
rect 39221 12801 39255 12835
rect 39405 12801 39439 12835
rect 39497 12801 39531 12835
rect 39589 12801 39623 12835
rect 39773 12801 39807 12835
rect 40417 12801 40451 12835
rect 45109 12801 45143 12835
rect 1685 12733 1719 12767
rect 3709 12733 3743 12767
rect 5641 12733 5675 12767
rect 5825 12733 5859 12767
rect 6561 12733 6595 12767
rect 7297 12733 7331 12767
rect 7414 12733 7448 12767
rect 7573 12733 7607 12767
rect 10977 12733 11011 12767
rect 12449 12733 12483 12767
rect 12587 12733 12621 12767
rect 13921 12733 13955 12767
rect 14013 12733 14047 12767
rect 16221 12733 16255 12767
rect 16405 12733 16439 12767
rect 17141 12733 17175 12767
rect 17785 12733 17819 12767
rect 18061 12733 18095 12767
rect 19625 12733 19659 12767
rect 23029 12733 23063 12767
rect 23213 12733 23247 12767
rect 23949 12733 23983 12767
rect 24066 12733 24100 12767
rect 24225 12733 24259 12767
rect 28825 12733 28859 12767
rect 33425 12733 33459 12767
rect 34437 12733 34471 12767
rect 40509 12733 40543 12767
rect 40785 12733 40819 12767
rect 42993 12733 43027 12767
rect 43085 12733 43119 12767
rect 43177 12733 43211 12767
rect 44925 12733 44959 12767
rect 5089 12665 5123 12699
rect 7021 12665 7055 12699
rect 12173 12665 12207 12699
rect 18981 12665 19015 12699
rect 20177 12665 20211 12699
rect 23673 12665 23707 12699
rect 27721 12665 27755 12699
rect 33885 12665 33919 12699
rect 39221 12665 39255 12699
rect 8217 12597 8251 12631
rect 10333 12597 10367 12631
rect 13369 12597 13403 12631
rect 15669 12597 15703 12631
rect 20361 12597 20395 12631
rect 20729 12597 20763 12631
rect 24961 12597 24995 12631
rect 45293 12597 45327 12631
rect 5181 12393 5215 12427
rect 7757 12393 7791 12427
rect 9689 12393 9723 12427
rect 14565 12393 14599 12427
rect 19717 12393 19751 12427
rect 25789 12393 25823 12427
rect 39129 12393 39163 12427
rect 39589 12393 39623 12427
rect 40049 12393 40083 12427
rect 41613 12393 41647 12427
rect 43453 12393 43487 12427
rect 7665 12325 7699 12359
rect 12265 12325 12299 12359
rect 23029 12325 23063 12359
rect 26157 12325 26191 12359
rect 30021 12325 30055 12359
rect 36461 12325 36495 12359
rect 38669 12325 38703 12359
rect 41245 12325 41279 12359
rect 3801 12257 3835 12291
rect 6009 12257 6043 12291
rect 6469 12257 6503 12291
rect 6745 12257 6779 12291
rect 6883 12257 6917 12291
rect 8401 12257 8435 12291
rect 10241 12257 10275 12291
rect 11621 12257 11655 12291
rect 11805 12257 11839 12291
rect 12541 12257 12575 12291
rect 12658 12257 12692 12291
rect 15117 12257 15151 12291
rect 16957 12257 16991 12291
rect 17141 12257 17175 12291
rect 17601 12257 17635 12291
rect 17877 12257 17911 12291
rect 18015 12257 18049 12291
rect 18153 12257 18187 12291
rect 23765 12257 23799 12291
rect 27721 12257 27755 12291
rect 38945 12257 38979 12291
rect 41429 12257 41463 12291
rect 43085 12257 43119 12291
rect 5825 12189 5859 12223
rect 7021 12189 7055 12223
rect 8125 12189 8159 12223
rect 10057 12189 10091 12223
rect 12817 12189 12851 12223
rect 14933 12189 14967 12223
rect 19441 12189 19475 12223
rect 19533 12189 19567 12223
rect 19809 12189 19843 12223
rect 19901 12189 19935 12223
rect 20177 12189 20211 12223
rect 21649 12189 21683 12223
rect 24409 12189 24443 12223
rect 24676 12189 24710 12223
rect 29837 12189 29871 12223
rect 32505 12189 32539 12223
rect 35909 12189 35943 12223
rect 36185 12189 36219 12223
rect 36329 12189 36363 12223
rect 38393 12189 38427 12223
rect 38577 12189 38611 12223
rect 39037 12189 39071 12223
rect 39313 12189 39347 12223
rect 39865 12189 39899 12223
rect 40049 12189 40083 12223
rect 41153 12189 41187 12223
rect 41797 12189 41831 12223
rect 42257 12189 42291 12223
rect 42441 12189 42475 12223
rect 42809 12189 42843 12223
rect 43729 12189 43763 12223
rect 43821 12189 43855 12223
rect 43913 12189 43947 12223
rect 44097 12189 44131 12223
rect 44189 12189 44223 12223
rect 44465 12189 44499 12223
rect 44557 12189 44591 12223
rect 4068 12121 4102 12155
rect 15025 12121 15059 12155
rect 16681 12121 16715 12155
rect 19257 12121 19291 12155
rect 21916 12121 21950 12155
rect 23581 12121 23615 12155
rect 25881 12121 25915 12155
rect 27445 12121 27479 12155
rect 36093 12121 36127 12155
rect 44373 12121 44407 12155
rect 8217 12053 8251 12087
rect 10149 12053 10183 12087
rect 13461 12053 13495 12087
rect 16773 12053 16807 12087
rect 18797 12053 18831 12087
rect 20913 12053 20947 12087
rect 23121 12053 23155 12087
rect 23489 12053 23523 12087
rect 26341 12053 26375 12087
rect 27077 12053 27111 12087
rect 27537 12053 27571 12087
rect 32689 12053 32723 12087
rect 38853 12053 38887 12087
rect 40233 12053 40267 12087
rect 41429 12053 41463 12087
rect 44741 12053 44775 12087
rect 4169 11849 4203 11883
rect 4813 11849 4847 11883
rect 5181 11849 5215 11883
rect 10425 11849 10459 11883
rect 10885 11849 10919 11883
rect 22017 11849 22051 11883
rect 23397 11849 23431 11883
rect 26617 11849 26651 11883
rect 30389 11849 30423 11883
rect 33425 11849 33459 11883
rect 34253 11849 34287 11883
rect 38025 11849 38059 11883
rect 41613 11849 41647 11883
rect 42257 11849 42291 11883
rect 42625 11849 42659 11883
rect 6837 11781 6871 11815
rect 23489 11781 23523 11815
rect 27230 11781 27264 11815
rect 31585 11781 31619 11815
rect 31677 11781 31711 11815
rect 33333 11781 33367 11815
rect 38739 11781 38773 11815
rect 39129 11781 39163 11815
rect 4353 11713 4387 11747
rect 5273 11713 5307 11747
rect 6009 11713 6043 11747
rect 6745 11713 6779 11747
rect 9045 11713 9079 11747
rect 9312 11713 9346 11747
rect 10977 11713 11011 11747
rect 22201 11713 22235 11747
rect 26801 11713 26835 11747
rect 26985 11713 27019 11747
rect 29377 11713 29411 11747
rect 29469 11713 29503 11747
rect 29745 11713 29779 11747
rect 30205 11713 30239 11747
rect 30481 11713 30515 11747
rect 32229 11713 32263 11747
rect 32597 11713 32631 11747
rect 34161 11713 34195 11747
rect 37565 11713 37599 11747
rect 38117 11713 38151 11747
rect 38301 11713 38335 11747
rect 39037 11713 39071 11747
rect 39313 11713 39347 11747
rect 41521 11713 41555 11747
rect 41797 11713 41831 11747
rect 43361 11713 43395 11747
rect 43545 11713 43579 11747
rect 44097 11713 44131 11747
rect 5457 11645 5491 11679
rect 7021 11645 7055 11679
rect 11069 11645 11103 11679
rect 23673 11645 23707 11679
rect 30021 11645 30055 11679
rect 31769 11645 31803 11679
rect 33609 11645 33643 11679
rect 34345 11645 34379 11679
rect 38209 11645 38243 11679
rect 38669 11645 38703 11679
rect 38853 11645 38887 11679
rect 42441 11645 42475 11679
rect 42809 11645 42843 11679
rect 43269 11645 43303 11679
rect 43453 11645 43487 11679
rect 44005 11645 44039 11679
rect 44465 11645 44499 11679
rect 6377 11577 6411 11611
rect 29193 11577 29227 11611
rect 38945 11577 38979 11611
rect 5825 11509 5859 11543
rect 10517 11509 10551 11543
rect 23029 11509 23063 11543
rect 28365 11509 28399 11543
rect 29653 11509 29687 11543
rect 31217 11509 31251 11543
rect 32965 11509 32999 11543
rect 33793 11509 33827 11543
rect 37841 11509 37875 11543
rect 39497 11509 39531 11543
rect 41889 11509 41923 11543
rect 42993 11509 43027 11543
rect 43085 11509 43119 11543
rect 6745 11305 6779 11339
rect 9413 11305 9447 11339
rect 13553 11305 13587 11339
rect 23857 11305 23891 11339
rect 26525 11305 26559 11339
rect 30021 11305 30055 11339
rect 32229 11305 32263 11339
rect 34161 11305 34195 11339
rect 38209 11305 38243 11339
rect 39037 11305 39071 11339
rect 42809 11305 42843 11339
rect 43361 11305 43395 11339
rect 15485 11237 15519 11271
rect 20085 11237 20119 11271
rect 25145 11237 25179 11271
rect 25881 11237 25915 11271
rect 26341 11237 26375 11271
rect 29929 11237 29963 11271
rect 32505 11237 32539 11271
rect 36645 11237 36679 11271
rect 39497 11237 39531 11271
rect 44281 11237 44315 11271
rect 5365 11169 5399 11203
rect 10977 11169 11011 11203
rect 12909 11169 12943 11203
rect 14473 11169 14507 11203
rect 14565 11169 14599 11203
rect 16129 11169 16163 11203
rect 18153 11169 18187 11203
rect 19809 11169 19843 11203
rect 24869 11169 24903 11203
rect 26065 11169 26099 11203
rect 29561 11169 29595 11203
rect 35633 11169 35667 11203
rect 43913 11169 43947 11203
rect 5632 11101 5666 11135
rect 9597 11101 9631 11135
rect 13277 11101 13311 11135
rect 13369 11101 13403 11135
rect 15393 11101 15427 11135
rect 15945 11101 15979 11135
rect 17969 11101 18003 11135
rect 22477 11101 22511 11135
rect 25605 11101 25639 11135
rect 25697 11101 25731 11135
rect 25973 11101 26007 11135
rect 26801 11101 26835 11135
rect 27077 11101 27111 11135
rect 30849 11101 30883 11135
rect 32689 11101 32723 11135
rect 32781 11101 32815 11135
rect 33037 11101 33071 11135
rect 34437 11101 34471 11135
rect 35909 11101 35943 11135
rect 37749 11101 37783 11135
rect 37933 11101 37967 11135
rect 38209 11101 38243 11135
rect 38393 11101 38427 11135
rect 38761 11101 38795 11135
rect 38853 11101 38887 11135
rect 39129 11101 39163 11135
rect 39221 11101 39255 11135
rect 39359 11101 39393 11135
rect 39681 11101 39715 11135
rect 42533 11101 42567 11135
rect 42717 11101 42751 11135
rect 42993 11101 43027 11135
rect 43269 11101 43303 11135
rect 43545 11101 43579 11135
rect 43821 11101 43855 11135
rect 44097 11101 44131 11135
rect 10885 11033 10919 11067
rect 14105 11033 14139 11067
rect 14749 11033 14783 11067
rect 17877 11033 17911 11067
rect 22744 11033 22778 11067
rect 25421 11033 25455 11067
rect 26617 11033 26651 11067
rect 26985 11033 27019 11067
rect 31116 11033 31150 11067
rect 38117 11033 38151 11067
rect 10425 10965 10459 10999
rect 10793 10965 10827 10999
rect 15209 10965 15243 10999
rect 15853 10965 15887 10999
rect 17509 10965 17543 10999
rect 20269 10965 20303 10999
rect 25329 10965 25363 10999
rect 34253 10965 34287 10999
rect 38577 10965 38611 10999
rect 39589 10965 39623 10999
rect 42717 10965 42751 10999
rect 43177 10965 43211 10999
rect 43729 10965 43763 10999
rect 6745 10761 6779 10795
rect 7113 10761 7147 10795
rect 10977 10761 11011 10795
rect 14105 10761 14139 10795
rect 14565 10761 14599 10795
rect 16313 10761 16347 10795
rect 21189 10761 21223 10795
rect 22845 10761 22879 10795
rect 30481 10761 30515 10795
rect 31217 10761 31251 10795
rect 34621 10761 34655 10795
rect 36737 10761 36771 10795
rect 38301 10761 38335 10795
rect 39129 10761 39163 10795
rect 40601 10761 40635 10795
rect 41245 10761 41279 10795
rect 43361 10761 43395 10795
rect 43653 10761 43687 10795
rect 15200 10693 15234 10727
rect 19717 10693 19751 10727
rect 33508 10693 33542 10727
rect 40233 10693 40267 10727
rect 42809 10693 42843 10727
rect 42993 10693 43027 10727
rect 43453 10693 43487 10727
rect 6561 10625 6595 10659
rect 8702 10625 8736 10659
rect 8861 10625 8895 10659
rect 9853 10625 9887 10659
rect 12725 10625 12759 10659
rect 14013 10625 14047 10659
rect 14473 10625 14507 10659
rect 14933 10625 14967 10659
rect 17325 10625 17359 10659
rect 17785 10625 17819 10659
rect 18061 10625 18095 10659
rect 18914 10625 18948 10659
rect 19073 10625 19107 10659
rect 20453 10625 20487 10659
rect 23029 10625 23063 10659
rect 28641 10625 28675 10659
rect 29678 10625 29712 10659
rect 29837 10625 29871 10659
rect 31401 10625 31435 10659
rect 33241 10625 33275 10659
rect 35725 10625 35759 10659
rect 36001 10625 36035 10659
rect 37933 10625 37967 10659
rect 38117 10625 38151 10659
rect 38393 10625 38427 10659
rect 38485 10625 38519 10659
rect 38761 10625 38795 10659
rect 38945 10625 38979 10659
rect 40049 10625 40083 10659
rect 40325 10625 40359 10659
rect 40417 10625 40451 10659
rect 40693 10625 40727 10659
rect 41061 10625 41095 10659
rect 42717 10625 42751 10659
rect 42901 10625 42935 10659
rect 43177 10625 43211 10659
rect 46489 10625 46523 10659
rect 7205 10557 7239 10591
rect 7389 10557 7423 10591
rect 7665 10557 7699 10591
rect 7849 10557 7883 10591
rect 8309 10557 8343 10591
rect 8585 10557 8619 10591
rect 9597 10557 9631 10591
rect 11529 10557 11563 10591
rect 11713 10557 11747 10591
rect 12173 10557 12207 10591
rect 12449 10557 12483 10591
rect 12587 10557 12621 10591
rect 14749 10557 14783 10591
rect 17509 10557 17543 10591
rect 17877 10557 17911 10591
rect 18797 10557 18831 10591
rect 20177 10557 20211 10591
rect 28825 10557 28859 10591
rect 29285 10557 29319 10591
rect 29561 10557 29595 10591
rect 38669 10557 38703 10591
rect 17601 10489 17635 10523
rect 18521 10489 18555 10523
rect 38577 10489 38611 10523
rect 40049 10489 40083 10523
rect 40417 10489 40451 10523
rect 43821 10489 43855 10523
rect 6377 10421 6411 10455
rect 9505 10421 9539 10455
rect 13369 10421 13403 10455
rect 13829 10421 13863 10455
rect 43637 10421 43671 10455
rect 46673 10421 46707 10455
rect 7665 10217 7699 10251
rect 9229 10217 9263 10251
rect 13921 10217 13955 10251
rect 18337 10217 18371 10251
rect 20085 10217 20119 10251
rect 20545 10217 20579 10251
rect 20729 10217 20763 10251
rect 40785 10217 40819 10251
rect 11897 10149 11931 10183
rect 15485 10149 15519 10183
rect 22661 10149 22695 10183
rect 27537 10149 27571 10183
rect 30205 10149 30239 10183
rect 31493 10149 31527 10183
rect 37289 10149 37323 10183
rect 42717 10149 42751 10183
rect 6193 10081 6227 10115
rect 8125 10081 8159 10115
rect 8217 10081 8251 10115
rect 11253 10081 11287 10115
rect 11437 10081 11471 10115
rect 12311 10081 12345 10115
rect 13277 10081 13311 10115
rect 13645 10081 13679 10115
rect 14105 10081 14139 10115
rect 21189 10081 21223 10115
rect 22017 10081 22051 10115
rect 23121 10081 23155 10115
rect 27813 10081 27847 10115
rect 29561 10081 29595 10115
rect 30481 10081 30515 10115
rect 30757 10081 30791 10115
rect 32045 10081 32079 10115
rect 35173 10081 35207 10115
rect 36277 10081 36311 10115
rect 39681 10081 39715 10115
rect 42901 10081 42935 10115
rect 6101 10013 6135 10047
rect 9413 10013 9447 10047
rect 9689 10013 9723 10047
rect 9781 10013 9815 10047
rect 12173 10013 12207 10047
rect 12449 10013 12483 10047
rect 13737 10013 13771 10047
rect 14361 10013 14395 10047
rect 16957 10013 16991 10047
rect 17224 10013 17258 10047
rect 20269 10013 20303 10047
rect 20361 10013 20395 10047
rect 20637 10013 20671 10047
rect 20913 10013 20947 10047
rect 21005 10013 21039 10047
rect 21281 10013 21315 10047
rect 21649 10013 21683 10047
rect 21909 10007 21943 10041
rect 22201 10013 22235 10047
rect 22477 10013 22511 10047
rect 22845 10013 22879 10047
rect 22937 10013 22971 10047
rect 23213 10013 23247 10047
rect 27721 10013 27755 10047
rect 29745 10013 29779 10047
rect 30598 10013 30632 10047
rect 35449 10013 35483 10047
rect 36553 10013 36587 10047
rect 39405 10013 39439 10047
rect 39497 10013 39531 10047
rect 39865 10013 39899 10047
rect 40141 10013 40175 10047
rect 41061 10013 41095 10047
rect 41153 10013 41187 10047
rect 41245 10013 41279 10047
rect 41429 10013 41463 10047
rect 42625 10013 42659 10047
rect 42993 10013 43027 10047
rect 43177 10013 43211 10047
rect 1501 9945 1535 9979
rect 2237 9945 2271 9979
rect 6438 9945 6472 9979
rect 8033 9945 8067 9979
rect 10026 9945 10060 9979
rect 13093 9945 13127 9979
rect 28058 9945 28092 9979
rect 31401 9945 31435 9979
rect 31861 9945 31895 9979
rect 1593 9877 1627 9911
rect 5917 9877 5951 9911
rect 7573 9877 7607 9911
rect 9505 9877 9539 9911
rect 11161 9877 11195 9911
rect 21465 9877 21499 9911
rect 21833 9877 21867 9911
rect 22385 9877 22419 9911
rect 29193 9877 29227 9911
rect 31953 9877 31987 9911
rect 36185 9877 36219 9911
rect 39681 9877 39715 9911
rect 42901 9877 42935 9911
rect 43177 9877 43211 9911
rect 7757 9673 7791 9707
rect 28457 9673 28491 9707
rect 28917 9673 28951 9707
rect 30757 9673 30791 9707
rect 6622 9605 6656 9639
rect 10057 9605 10091 9639
rect 19717 9605 19751 9639
rect 19809 9605 19843 9639
rect 20821 9605 20855 9639
rect 25881 9605 25915 9639
rect 28825 9605 28859 9639
rect 42257 9605 42291 9639
rect 8125 9537 8159 9571
rect 8861 9537 8895 9571
rect 17877 9537 17911 9571
rect 18061 9537 18095 9571
rect 18797 9537 18831 9571
rect 18914 9537 18948 9571
rect 19073 9537 19107 9571
rect 24041 9537 24075 9571
rect 25237 9537 25271 9571
rect 26801 9537 26835 9571
rect 27241 9537 27275 9571
rect 31125 9537 31159 9571
rect 36185 9537 36219 9571
rect 38393 9537 38427 9571
rect 38577 9537 38611 9571
rect 40325 9537 40359 9571
rect 40417 9537 40451 9571
rect 40601 9537 40635 9571
rect 41245 9537 41279 9571
rect 42625 9537 42659 9571
rect 43453 9537 43487 9571
rect 6377 9469 6411 9503
rect 7941 9469 7975 9503
rect 8978 9469 9012 9503
rect 9137 9469 9171 9503
rect 20269 9469 20303 9503
rect 21281 9469 21315 9503
rect 24225 9469 24259 9503
rect 24961 9469 24995 9503
rect 25099 9469 25133 9503
rect 26985 9469 27019 9503
rect 29009 9469 29043 9503
rect 31217 9469 31251 9503
rect 31401 9469 31435 9503
rect 32229 9469 32263 9503
rect 32505 9469 32539 9503
rect 35909 9469 35943 9503
rect 40141 9469 40175 9503
rect 40509 9469 40543 9503
rect 42533 9469 42567 9503
rect 43085 9469 43119 9503
rect 43269 9469 43303 9503
rect 43361 9469 43395 9503
rect 43545 9469 43579 9503
rect 8585 9401 8619 9435
rect 18521 9401 18555 9435
rect 20085 9401 20119 9435
rect 21097 9401 21131 9435
rect 24685 9401 24719 9435
rect 26617 9401 26651 9435
rect 42993 9401 43027 9435
rect 9781 9333 9815 9367
rect 10149 9333 10183 9367
rect 28365 9333 28399 9367
rect 36921 9333 36955 9367
rect 38393 9333 38427 9367
rect 26341 9129 26375 9163
rect 27261 9129 27295 9163
rect 36737 9129 36771 9163
rect 38485 9129 38519 9163
rect 42717 9129 42751 9163
rect 10609 9061 10643 9095
rect 13185 9061 13219 9095
rect 21465 9061 21499 9095
rect 21649 9061 21683 9095
rect 22845 9061 22879 9095
rect 30389 9061 30423 9095
rect 11161 8993 11195 9027
rect 13737 8993 13771 9027
rect 15853 8993 15887 9027
rect 16589 8993 16623 9027
rect 21189 8993 21223 9027
rect 22201 8993 22235 9027
rect 24409 8993 24443 9027
rect 24593 8993 24627 9027
rect 25053 8993 25087 9027
rect 25329 8993 25363 9027
rect 26985 8993 27019 9027
rect 27721 8993 27755 9027
rect 27813 8993 27847 9027
rect 30941 8993 30975 9027
rect 10977 8925 11011 8959
rect 21925 8925 21959 8959
rect 22017 8925 22051 8959
rect 22293 8925 22327 8959
rect 22569 8925 22603 8959
rect 22661 8925 22695 8959
rect 22937 8925 22971 8959
rect 24225 8925 24259 8959
rect 25446 8925 25480 8959
rect 25605 8925 25639 8959
rect 26709 8925 26743 8959
rect 27629 8925 27663 8959
rect 32137 8925 32171 8959
rect 36185 8925 36219 8959
rect 36369 8925 36403 8959
rect 36461 8925 36495 8959
rect 36558 8925 36592 8959
rect 37473 8925 37507 8959
rect 37749 8925 37783 8959
rect 39681 8925 39715 8959
rect 42717 8925 42751 8959
rect 42901 8925 42935 8959
rect 42993 8925 43027 8959
rect 13645 8857 13679 8891
rect 16405 8857 16439 8891
rect 32404 8857 32438 8891
rect 38669 8857 38703 8891
rect 11069 8789 11103 8823
rect 13553 8789 13587 8823
rect 15209 8789 15243 8823
rect 15577 8789 15611 8823
rect 15669 8789 15703 8823
rect 16037 8789 16071 8823
rect 16497 8789 16531 8823
rect 21741 8789 21775 8823
rect 22385 8789 22419 8823
rect 24041 8789 24075 8823
rect 26249 8789 26283 8823
rect 26801 8789 26835 8823
rect 30757 8789 30791 8823
rect 30849 8789 30883 8823
rect 33517 8789 33551 8823
rect 38761 8789 38795 8823
rect 8401 8585 8435 8619
rect 14013 8585 14047 8619
rect 14657 8585 14691 8619
rect 16313 8585 16347 8619
rect 18981 8585 19015 8619
rect 20913 8585 20947 8619
rect 22293 8585 22327 8619
rect 26065 8585 26099 8619
rect 31309 8585 31343 8619
rect 32321 8585 32355 8619
rect 34805 8585 34839 8619
rect 38025 8585 38059 8619
rect 39865 8585 39899 8619
rect 15178 8517 15212 8551
rect 24930 8517 24964 8551
rect 36001 8517 36035 8551
rect 38752 8517 38786 8551
rect 7941 8449 7975 8483
rect 8493 8449 8527 8483
rect 10701 8449 10735 8483
rect 12909 8449 12943 8483
rect 13921 8449 13955 8483
rect 14841 8449 14875 8483
rect 18178 8449 18212 8483
rect 21833 8449 21867 8483
rect 23121 8449 23155 8483
rect 30665 8449 30699 8483
rect 32505 8449 32539 8483
rect 34161 8449 34195 8483
rect 37657 8449 37691 8483
rect 37913 8449 37947 8483
rect 38209 8449 38243 8483
rect 46213 8449 46247 8483
rect 8585 8381 8619 8415
rect 12633 8381 12667 8415
rect 14197 8381 14231 8415
rect 14933 8381 14967 8415
rect 17141 8381 17175 8415
rect 17325 8381 17359 8415
rect 18061 8381 18095 8415
rect 18337 8381 18371 8415
rect 19073 8381 19107 8415
rect 19257 8381 19291 8415
rect 19993 8381 20027 8415
rect 20110 8381 20144 8415
rect 20269 8381 20303 8415
rect 24685 8381 24719 8415
rect 29469 8381 29503 8415
rect 29653 8381 29687 8415
rect 30113 8381 30147 8415
rect 30389 8381 30423 8415
rect 30527 8381 30561 8415
rect 32965 8381 32999 8415
rect 33149 8381 33183 8415
rect 33885 8381 33919 8415
rect 34002 8381 34036 8415
rect 38117 8381 38151 8415
rect 38485 8381 38519 8415
rect 45937 8381 45971 8415
rect 8033 8313 8067 8347
rect 13553 8313 13587 8347
rect 17785 8313 17819 8347
rect 19717 8313 19751 8347
rect 22109 8313 22143 8347
rect 33609 8313 33643 8347
rect 36185 8313 36219 8347
rect 7757 8245 7791 8279
rect 10517 8245 10551 8279
rect 22937 8245 22971 8279
rect 37473 8245 37507 8279
rect 8953 8041 8987 8075
rect 11621 8041 11655 8075
rect 11713 8041 11747 8075
rect 13921 8041 13955 8075
rect 17141 8041 17175 8075
rect 19073 8041 19107 8075
rect 21097 8041 21131 8075
rect 31401 8041 31435 8075
rect 31861 8041 31895 8075
rect 34529 8041 34563 8075
rect 36645 8041 36679 8075
rect 38669 8041 38703 8075
rect 8769 7973 8803 8007
rect 17877 7973 17911 8007
rect 24961 7973 24995 8007
rect 9413 7905 9447 7939
rect 9597 7905 9631 7939
rect 10241 7905 10275 7939
rect 12265 7905 12299 7939
rect 15025 7905 15059 7939
rect 17233 7905 17267 7939
rect 18153 7905 18187 7939
rect 18270 7905 18304 7939
rect 18429 7905 18463 7939
rect 19257 7905 19291 7939
rect 19441 7905 19475 7939
rect 19901 7905 19935 7939
rect 20294 7905 20328 7939
rect 20453 7905 20487 7939
rect 25513 7905 25547 7939
rect 28089 7905 28123 7939
rect 29561 7905 29595 7939
rect 30205 7905 30239 7939
rect 30598 7905 30632 7939
rect 32505 7905 32539 7939
rect 32873 7905 32907 7939
rect 33333 7905 33367 7939
rect 33609 7905 33643 7939
rect 35265 7905 35299 7939
rect 7297 7837 7331 7871
rect 7389 7837 7423 7871
rect 10508 7837 10542 7871
rect 12081 7837 12115 7871
rect 12541 7837 12575 7871
rect 14289 7837 14323 7871
rect 14565 7837 14599 7871
rect 15761 7837 15795 7871
rect 17417 7837 17451 7871
rect 20177 7837 20211 7871
rect 22569 7837 22603 7871
rect 22836 7837 22870 7871
rect 25329 7837 25363 7871
rect 27905 7837 27939 7871
rect 29745 7837 29779 7871
rect 30481 7837 30515 7871
rect 30757 7837 30791 7871
rect 32229 7837 32263 7871
rect 32689 7837 32723 7871
rect 33726 7837 33760 7871
rect 33885 7837 33919 7871
rect 35173 7837 35207 7871
rect 38577 7837 38611 7871
rect 38761 7837 38795 7871
rect 7634 7769 7668 7803
rect 12173 7769 12207 7803
rect 12808 7769 12842 7803
rect 14841 7769 14875 7803
rect 16028 7769 16062 7803
rect 27997 7769 28031 7803
rect 35510 7769 35544 7803
rect 7113 7701 7147 7735
rect 9321 7701 9355 7735
rect 14105 7701 14139 7735
rect 14381 7701 14415 7735
rect 23949 7701 23983 7735
rect 25421 7701 25455 7735
rect 27537 7701 27571 7735
rect 32321 7701 32355 7735
rect 34989 7701 35023 7735
rect 8861 7497 8895 7531
rect 11345 7497 11379 7531
rect 11897 7497 11931 7531
rect 11989 7497 12023 7531
rect 13829 7497 13863 7531
rect 15945 7497 15979 7531
rect 18061 7497 18095 7531
rect 20913 7497 20947 7531
rect 22017 7497 22051 7531
rect 23121 7497 23155 7531
rect 23489 7497 23523 7531
rect 28733 7497 28767 7531
rect 29193 7497 29227 7531
rect 31769 7497 31803 7531
rect 35909 7497 35943 7531
rect 36369 7497 36403 7531
rect 7748 7429 7782 7463
rect 12716 7429 12750 7463
rect 17969 7429 18003 7463
rect 19625 7429 19659 7463
rect 22385 7429 22419 7463
rect 22477 7429 22511 7463
rect 27506 7429 27540 7463
rect 30113 7429 30147 7463
rect 32382 7429 32416 7463
rect 36277 7429 36311 7463
rect 1501 7361 1535 7395
rect 10232 7361 10266 7395
rect 16129 7361 16163 7395
rect 19073 7361 19107 7395
rect 19533 7361 19567 7395
rect 21281 7361 21315 7395
rect 21373 7361 21407 7395
rect 24317 7361 24351 7395
rect 26801 7361 26835 7395
rect 27169 7361 27203 7395
rect 29101 7361 29135 7395
rect 31953 7361 31987 7395
rect 32137 7361 32171 7395
rect 33977 7361 34011 7395
rect 34437 7361 34471 7395
rect 34693 7361 34727 7395
rect 7481 7293 7515 7327
rect 9965 7293 9999 7327
rect 12081 7293 12115 7327
rect 12449 7293 12483 7327
rect 19809 7293 19843 7327
rect 19993 7293 20027 7327
rect 20269 7293 20303 7327
rect 21465 7293 21499 7327
rect 22661 7293 22695 7327
rect 23581 7293 23615 7327
rect 23765 7293 23799 7327
rect 24593 7293 24627 7327
rect 27261 7293 27295 7327
rect 29285 7293 29319 7327
rect 30205 7293 30239 7327
rect 30297 7293 30331 7327
rect 34069 7293 34103 7327
rect 34253 7293 34287 7327
rect 36553 7293 36587 7327
rect 18889 7225 18923 7259
rect 26617 7225 26651 7259
rect 28641 7225 28675 7259
rect 1593 7157 1627 7191
rect 11529 7157 11563 7191
rect 19165 7157 19199 7191
rect 26985 7157 27019 7191
rect 29745 7157 29779 7191
rect 33517 7157 33551 7191
rect 33609 7157 33643 7191
rect 35817 7157 35851 7191
rect 10425 6953 10459 6987
rect 20637 6953 20671 6987
rect 28549 6953 28583 6987
rect 32045 6953 32079 6987
rect 33977 6885 34011 6919
rect 15209 6817 15243 6851
rect 15602 6817 15636 6851
rect 15761 6817 15795 6851
rect 17877 6817 17911 6851
rect 24685 6817 24719 6851
rect 29745 6817 29779 6851
rect 32505 6817 32539 6851
rect 32597 6817 32631 6851
rect 10609 6749 10643 6783
rect 14565 6749 14599 6783
rect 14749 6749 14783 6783
rect 15485 6749 15519 6783
rect 19073 6749 19107 6783
rect 19257 6749 19291 6783
rect 27169 6749 27203 6783
rect 27425 6749 27459 6783
rect 30021 6749 30055 6783
rect 30849 6749 30883 6783
rect 32413 6749 32447 6783
rect 33793 6749 33827 6783
rect 34345 6749 34379 6783
rect 16405 6681 16439 6715
rect 19502 6681 19536 6715
rect 24952 6681 24986 6715
rect 17325 6613 17359 6647
rect 17693 6613 17727 6647
rect 17785 6613 17819 6647
rect 18889 6613 18923 6647
rect 26065 6613 26099 6647
rect 30665 6613 30699 6647
rect 34161 6613 34195 6647
rect 18153 6409 18187 6443
rect 23673 6409 23707 6443
rect 25605 6409 25639 6443
rect 26525 6409 26559 6443
rect 31217 6409 31251 6443
rect 19226 6341 19260 6375
rect 30104 6341 30138 6375
rect 13185 6273 13219 6307
rect 14013 6273 14047 6307
rect 15531 6273 15565 6307
rect 15669 6273 15703 6307
rect 16773 6273 16807 6307
rect 17040 6273 17074 6307
rect 18889 6273 18923 6307
rect 20821 6273 20855 6307
rect 21833 6273 21867 6307
rect 24225 6273 24259 6307
rect 24492 6273 24526 6307
rect 26065 6273 26099 6307
rect 26157 6273 26191 6307
rect 26709 6273 26743 6307
rect 28917 6273 28951 6307
rect 29837 6273 29871 6307
rect 31493 6273 31527 6307
rect 14105 6205 14139 6239
rect 14289 6205 14323 6239
rect 14473 6205 14507 6239
rect 14657 6205 14691 6239
rect 15393 6205 15427 6239
rect 18981 6205 19015 6239
rect 20913 6205 20947 6239
rect 21005 6205 21039 6239
rect 22017 6205 22051 6239
rect 22477 6205 22511 6239
rect 22753 6205 22787 6239
rect 22870 6205 22904 6239
rect 23029 6205 23063 6239
rect 26341 6205 26375 6239
rect 29193 6205 29227 6239
rect 15117 6137 15151 6171
rect 18705 6137 18739 6171
rect 20453 6137 20487 6171
rect 25697 6137 25731 6171
rect 13001 6069 13035 6103
rect 13645 6069 13679 6103
rect 16313 6069 16347 6103
rect 20361 6069 20395 6103
rect 31309 6069 31343 6103
rect 14105 5865 14139 5899
rect 17141 5865 17175 5899
rect 23489 5865 23523 5899
rect 24501 5865 24535 5899
rect 31033 5865 31067 5899
rect 13921 5797 13955 5831
rect 25697 5797 25731 5831
rect 14565 5729 14599 5763
rect 14749 5729 14783 5763
rect 19257 5729 19291 5763
rect 19533 5729 19567 5763
rect 21833 5729 21867 5763
rect 22293 5729 22327 5763
rect 22686 5729 22720 5763
rect 22845 5729 22879 5763
rect 26249 5729 26283 5763
rect 29653 5729 29687 5763
rect 12541 5661 12575 5695
rect 17325 5661 17359 5695
rect 21649 5661 21683 5695
rect 22569 5661 22603 5695
rect 24685 5661 24719 5695
rect 29920 5661 29954 5695
rect 35265 5661 35299 5695
rect 46397 5661 46431 5695
rect 12808 5593 12842 5627
rect 24869 5593 24903 5627
rect 25053 5593 25087 5627
rect 26065 5593 26099 5627
rect 14473 5525 14507 5559
rect 26157 5525 26191 5559
rect 35081 5525 35115 5559
rect 46673 5525 46707 5559
rect 18061 5321 18095 5355
rect 21465 5321 21499 5355
rect 23397 5321 23431 5355
rect 26801 5321 26835 5355
rect 27813 5321 27847 5355
rect 29653 5321 29687 5355
rect 33977 5321 34011 5355
rect 11897 5253 11931 5287
rect 12716 5253 12750 5287
rect 22262 5253 22296 5287
rect 30021 5253 30055 5287
rect 35072 5253 35106 5287
rect 1409 5185 1443 5219
rect 9965 5185 9999 5219
rect 10232 5185 10266 5219
rect 14105 5185 14139 5219
rect 16681 5185 16715 5219
rect 16948 5185 16982 5219
rect 19165 5185 19199 5219
rect 21649 5185 21683 5219
rect 26157 5185 26191 5219
rect 27721 5185 27755 5219
rect 11989 5117 12023 5151
rect 12173 5117 12207 5151
rect 12449 5117 12483 5151
rect 22017 5117 22051 5151
rect 24961 5117 24995 5151
rect 25145 5117 25179 5151
rect 25881 5117 25915 5151
rect 26019 5117 26053 5151
rect 27997 5117 28031 5151
rect 30113 5117 30147 5151
rect 30205 5117 30239 5151
rect 32137 5117 32171 5151
rect 32321 5117 32355 5151
rect 33057 5117 33091 5151
rect 33174 5117 33208 5151
rect 33333 5117 33367 5151
rect 34805 5117 34839 5151
rect 13829 5049 13863 5083
rect 25605 5049 25639 5083
rect 32781 5049 32815 5083
rect 1593 4981 1627 5015
rect 11345 4981 11379 5015
rect 11529 4981 11563 5015
rect 13921 4981 13955 5015
rect 19257 4981 19291 5015
rect 27353 4981 27387 5015
rect 36185 4981 36219 5015
rect 10701 4777 10735 4811
rect 17233 4777 17267 4811
rect 22477 4777 22511 4811
rect 33977 4777 34011 4811
rect 35081 4777 35115 4811
rect 26249 4709 26283 4743
rect 27445 4709 27479 4743
rect 28917 4709 28951 4743
rect 29009 4709 29043 4743
rect 29561 4709 29595 4743
rect 32781 4709 32815 4743
rect 15393 4641 15427 4675
rect 18337 4641 18371 4675
rect 19901 4641 19935 4675
rect 23121 4641 23155 4675
rect 25605 4641 25639 4675
rect 25789 4641 25823 4675
rect 26525 4641 26559 4675
rect 26801 4641 26835 4675
rect 30113 4641 30147 4675
rect 32137 4641 32171 4675
rect 33057 4641 33091 4675
rect 35725 4641 35759 4675
rect 10885 4573 10919 4607
rect 15577 4573 15611 4607
rect 15853 4573 15887 4607
rect 17417 4573 17451 4607
rect 18061 4573 18095 4607
rect 18153 4573 18187 4607
rect 22845 4573 22879 4607
rect 26642 4573 26676 4607
rect 27537 4573 27571 4607
rect 29193 4573 29227 4607
rect 29929 4573 29963 4607
rect 32045 4573 32079 4607
rect 32321 4573 32355 4607
rect 33174 4573 33208 4607
rect 33333 4573 33367 4607
rect 35449 4573 35483 4607
rect 35541 4573 35575 4607
rect 38301 4573 38335 4607
rect 15209 4505 15243 4539
rect 19625 4505 19659 4539
rect 22937 4505 22971 4539
rect 27782 4505 27816 4539
rect 14749 4437 14783 4471
rect 15117 4437 15151 4471
rect 17693 4437 17727 4471
rect 19257 4437 19291 4471
rect 19717 4437 19751 4471
rect 30021 4437 30055 4471
rect 31861 4437 31895 4471
rect 18429 4233 18463 4267
rect 20085 4233 20119 4267
rect 22201 4233 22235 4267
rect 24961 4233 24995 4267
rect 17509 4165 17543 4199
rect 33026 4165 33060 4199
rect 38108 4165 38142 4199
rect 14372 4097 14406 4131
rect 17049 4097 17083 4131
rect 18613 4097 18647 4131
rect 18961 4097 18995 4131
rect 21281 4097 21315 4131
rect 23949 4097 23983 4131
rect 26157 4097 26191 4131
rect 27537 4097 27571 4131
rect 28641 4097 28675 4131
rect 28908 4097 28942 4131
rect 31033 4097 31067 4131
rect 32781 4097 32815 4131
rect 37841 4097 37875 4131
rect 14105 4029 14139 4063
rect 17601 4029 17635 4063
rect 17785 4029 17819 4063
rect 18705 4029 18739 4063
rect 22293 4029 22327 4063
rect 22477 4029 22511 4063
rect 25053 4029 25087 4063
rect 25145 4029 25179 4063
rect 15485 3961 15519 3995
rect 17141 3961 17175 3995
rect 21833 3961 21867 3995
rect 27353 3961 27387 3995
rect 30021 3961 30055 3995
rect 39221 3961 39255 3995
rect 16865 3893 16899 3927
rect 21097 3893 21131 3927
rect 23765 3893 23799 3927
rect 24593 3893 24627 3927
rect 25973 3893 26007 3927
rect 30849 3893 30883 3927
rect 34161 3893 34195 3927
rect 14565 3689 14599 3723
rect 18245 3689 18279 3723
rect 22201 3689 22235 3723
rect 23489 3689 23523 3723
rect 25789 3689 25823 3723
rect 32597 3689 32631 3723
rect 18153 3621 18187 3655
rect 22293 3621 22327 3655
rect 31861 3621 31895 3655
rect 15669 3553 15703 3587
rect 18797 3553 18831 3587
rect 20453 3553 20487 3587
rect 20637 3553 20671 3587
rect 22753 3553 22787 3587
rect 22845 3553 22879 3587
rect 24133 3553 24167 3587
rect 25973 3553 26007 3587
rect 30021 3553 30055 3587
rect 30205 3553 30239 3587
rect 30481 3553 30515 3587
rect 33241 3553 33275 3587
rect 33885 3553 33919 3587
rect 34069 3553 34103 3587
rect 35265 3553 35299 3587
rect 14473 3485 14507 3519
rect 14749 3485 14783 3519
rect 15393 3485 15427 3519
rect 16681 3485 16715 3519
rect 16773 3485 16807 3519
rect 18613 3485 18647 3519
rect 19901 3485 19935 3519
rect 20821 3485 20855 3519
rect 21088 3485 21122 3519
rect 23305 3485 23339 3519
rect 23949 3485 23983 3519
rect 24409 3485 24443 3519
rect 26229 3485 26263 3519
rect 27629 3485 27663 3519
rect 29929 3485 29963 3519
rect 30748 3485 30782 3519
rect 32137 3485 32171 3519
rect 33793 3485 33827 3519
rect 35081 3485 35115 3519
rect 17018 3417 17052 3451
rect 20361 3417 20395 3451
rect 23857 3417 23891 3451
rect 24676 3417 24710 3451
rect 33057 3417 33091 3451
rect 14289 3349 14323 3383
rect 15025 3349 15059 3383
rect 15485 3349 15519 3383
rect 16497 3349 16531 3383
rect 18705 3349 18739 3383
rect 19717 3349 19751 3383
rect 19993 3349 20027 3383
rect 22661 3349 22695 3383
rect 23121 3349 23155 3383
rect 27353 3349 27387 3383
rect 29561 3349 29595 3383
rect 31953 3349 31987 3383
rect 32965 3349 32999 3383
rect 33425 3349 33459 3383
rect 34713 3349 34747 3383
rect 35173 3349 35207 3383
rect 15669 3145 15703 3179
rect 18061 3145 18095 3179
rect 20913 3145 20947 3179
rect 23213 3145 23247 3179
rect 24869 3145 24903 3179
rect 24961 3145 24995 3179
rect 25789 3145 25823 3179
rect 30297 3145 30331 3179
rect 31033 3145 31067 3179
rect 31401 3145 31435 3179
rect 33517 3145 33551 3179
rect 34989 3145 35023 3179
rect 46673 3145 46707 3179
rect 14534 3077 14568 3111
rect 22100 3077 22134 3111
rect 23756 3077 23790 3111
rect 26157 3077 26191 3111
rect 27344 3077 27378 3111
rect 31493 3077 31527 3111
rect 32382 3077 32416 3111
rect 1501 3009 1535 3043
rect 16681 3009 16715 3043
rect 16948 3009 16982 3043
rect 19533 3009 19567 3043
rect 19800 3009 19834 3043
rect 21833 3009 21867 3043
rect 25145 3009 25179 3043
rect 27077 3009 27111 3043
rect 28917 3009 28951 3043
rect 29184 3009 29218 3043
rect 32137 3009 32171 3043
rect 33865 3009 33899 3043
rect 46581 3009 46615 3043
rect 14289 2941 14323 2975
rect 23489 2941 23523 2975
rect 26249 2941 26283 2975
rect 26341 2941 26375 2975
rect 31677 2941 31711 2975
rect 33609 2941 33643 2975
rect 2237 2873 2271 2907
rect 1593 2805 1627 2839
rect 28457 2805 28491 2839
rect 6561 2601 6595 2635
rect 14335 2601 14369 2635
rect 23305 2601 23339 2635
rect 39405 2601 39439 2635
rect 2421 2533 2455 2567
rect 9413 2465 9447 2499
rect 25513 2465 25547 2499
rect 42717 2465 42751 2499
rect 45937 2465 45971 2499
rect 46213 2465 46247 2499
rect 1409 2397 1443 2431
rect 2237 2397 2271 2431
rect 4629 2397 4663 2431
rect 6745 2397 6779 2431
rect 9137 2397 9171 2431
rect 11713 2397 11747 2431
rect 14105 2397 14139 2431
rect 16681 2397 16715 2431
rect 16957 2397 16991 2431
rect 18797 2397 18831 2431
rect 21005 2397 21039 2431
rect 23489 2397 23523 2431
rect 25237 2397 25271 2431
rect 27813 2397 27847 2431
rect 29377 2397 29411 2431
rect 32321 2397 32355 2431
rect 33609 2397 33643 2431
rect 34897 2397 34931 2431
rect 37473 2397 37507 2431
rect 39589 2397 39623 2431
rect 42441 2397 42475 2431
rect 44557 2397 44591 2431
rect 45845 2397 45879 2431
rect 2053 2329 2087 2363
rect 20821 2329 20855 2363
rect 30297 2329 30331 2363
rect 1593 2261 1627 2295
rect 4813 2261 4847 2295
rect 11897 2261 11931 2295
rect 18981 2261 19015 2295
rect 27997 2261 28031 2295
rect 29193 2261 29227 2295
rect 30389 2261 30423 2295
rect 32505 2261 32539 2295
rect 33425 2261 33459 2295
rect 35081 2261 35115 2295
rect 37657 2261 37691 2295
rect 44741 2261 44775 2295
rect 45661 2261 45695 2295
<< metal1 >>
rect 6086 48016 6092 48068
rect 6144 48056 6150 48068
rect 32122 48056 32128 48068
rect 6144 48028 32128 48056
rect 6144 48016 6150 48028
rect 32122 48016 32128 48028
rect 32180 48016 32186 48068
rect 1104 47898 47104 47920
rect 1104 47846 4874 47898
rect 4926 47846 4938 47898
rect 4990 47846 5002 47898
rect 5054 47846 5066 47898
rect 5118 47846 5130 47898
rect 5182 47846 35594 47898
rect 35646 47846 35658 47898
rect 35710 47846 35722 47898
rect 35774 47846 35786 47898
rect 35838 47846 35850 47898
rect 35902 47846 47104 47898
rect 1104 47824 47104 47846
rect 1762 47744 1768 47796
rect 1820 47744 1826 47796
rect 3234 47744 3240 47796
rect 3292 47784 3298 47796
rect 3513 47787 3571 47793
rect 3513 47784 3525 47787
rect 3292 47756 3525 47784
rect 3292 47744 3298 47756
rect 3513 47753 3525 47756
rect 3559 47753 3571 47787
rect 3513 47747 3571 47753
rect 6086 47744 6092 47796
rect 6144 47744 6150 47796
rect 10594 47744 10600 47796
rect 10652 47744 10658 47796
rect 13170 47744 13176 47796
rect 13228 47744 13234 47796
rect 15746 47744 15752 47796
rect 15804 47744 15810 47796
rect 17402 47744 17408 47796
rect 17460 47784 17466 47796
rect 17497 47787 17555 47793
rect 17497 47784 17509 47787
rect 17460 47756 17509 47784
rect 17460 47744 17466 47756
rect 17497 47753 17509 47756
rect 17543 47753 17555 47787
rect 17497 47747 17555 47753
rect 17957 47787 18015 47793
rect 17957 47753 17969 47787
rect 18003 47784 18015 47787
rect 18003 47756 18828 47784
rect 18003 47753 18015 47756
rect 17957 47747 18015 47753
rect 5994 47676 6000 47728
rect 6052 47676 6058 47728
rect 1673 47651 1731 47657
rect 1673 47617 1685 47651
rect 1719 47648 1731 47651
rect 2314 47648 2320 47660
rect 1719 47620 2320 47648
rect 1719 47617 1731 47620
rect 1673 47611 1731 47617
rect 2314 47608 2320 47620
rect 2372 47608 2378 47660
rect 3050 47608 3056 47660
rect 3108 47648 3114 47660
rect 3329 47651 3387 47657
rect 3329 47648 3341 47651
rect 3108 47620 3341 47648
rect 3108 47608 3114 47620
rect 3329 47617 3341 47620
rect 3375 47617 3387 47651
rect 3329 47611 3387 47617
rect 8662 47608 8668 47660
rect 8720 47608 8726 47660
rect 10226 47608 10232 47660
rect 10284 47648 10290 47660
rect 10413 47651 10471 47657
rect 10413 47648 10425 47651
rect 10284 47620 10425 47648
rect 10284 47608 10290 47620
rect 10413 47617 10425 47620
rect 10459 47617 10471 47651
rect 10413 47611 10471 47617
rect 12989 47651 13047 47657
rect 12989 47617 13001 47651
rect 13035 47617 13047 47651
rect 12989 47611 13047 47617
rect 13004 47580 13032 47611
rect 15194 47608 15200 47660
rect 15252 47648 15258 47660
rect 15565 47651 15623 47657
rect 15565 47648 15577 47651
rect 15252 47620 15577 47648
rect 15252 47608 15258 47620
rect 15565 47617 15577 47620
rect 15611 47617 15623 47651
rect 15565 47611 15623 47617
rect 17310 47608 17316 47660
rect 17368 47608 17374 47660
rect 18248 47657 18276 47756
rect 18800 47716 18828 47756
rect 19978 47744 19984 47796
rect 20036 47784 20042 47796
rect 20349 47787 20407 47793
rect 20349 47784 20361 47787
rect 20036 47756 20361 47784
rect 20036 47744 20042 47756
rect 20349 47753 20361 47756
rect 20395 47753 20407 47787
rect 20349 47747 20407 47753
rect 22554 47744 22560 47796
rect 22612 47784 22618 47796
rect 22833 47787 22891 47793
rect 22833 47784 22845 47787
rect 22612 47756 22845 47784
rect 22612 47744 22618 47756
rect 22833 47753 22845 47756
rect 22879 47753 22891 47787
rect 22833 47747 22891 47753
rect 28994 47744 29000 47796
rect 29052 47784 29058 47796
rect 29273 47787 29331 47793
rect 29273 47784 29285 47787
rect 29052 47756 29285 47784
rect 29052 47744 29058 47756
rect 29273 47753 29285 47756
rect 29319 47753 29331 47787
rect 29273 47747 29331 47753
rect 31754 47744 31760 47796
rect 31812 47784 31818 47796
rect 32309 47787 32367 47793
rect 32309 47784 32321 47787
rect 31812 47756 32321 47784
rect 31812 47744 31818 47756
rect 32309 47753 32321 47756
rect 32355 47753 32367 47787
rect 32309 47747 32367 47753
rect 34422 47744 34428 47796
rect 34480 47744 34486 47796
rect 36078 47744 36084 47796
rect 36136 47784 36142 47796
rect 36357 47787 36415 47793
rect 36357 47784 36369 47787
rect 36136 47756 36369 47784
rect 36136 47744 36142 47756
rect 36357 47753 36369 47756
rect 36403 47753 36415 47787
rect 36357 47747 36415 47753
rect 41414 47744 41420 47796
rect 41472 47784 41478 47796
rect 41509 47787 41567 47793
rect 41509 47784 41521 47787
rect 41472 47756 41521 47784
rect 41472 47744 41478 47756
rect 41509 47753 41521 47756
rect 41555 47753 41567 47787
rect 41509 47747 41567 47753
rect 18800 47688 26924 47716
rect 18233 47651 18291 47657
rect 18233 47617 18245 47651
rect 18279 47617 18291 47651
rect 18233 47611 18291 47617
rect 18340 47620 18644 47648
rect 18340 47580 18368 47620
rect 13004 47552 18368 47580
rect 18616 47580 18644 47620
rect 19242 47608 19248 47660
rect 19300 47648 19306 47660
rect 19337 47651 19395 47657
rect 19337 47648 19349 47651
rect 19300 47620 19349 47648
rect 19300 47608 19306 47620
rect 19337 47617 19349 47620
rect 19383 47617 19395 47651
rect 19337 47611 19395 47617
rect 20165 47651 20223 47657
rect 20165 47617 20177 47651
rect 20211 47648 20223 47651
rect 20346 47648 20352 47660
rect 20211 47620 20352 47648
rect 20211 47617 20223 47620
rect 20165 47611 20223 47617
rect 20346 47608 20352 47620
rect 20404 47608 20410 47660
rect 22649 47651 22707 47657
rect 22649 47617 22661 47651
rect 22695 47648 22707 47651
rect 23198 47648 23204 47660
rect 22695 47620 23204 47648
rect 22695 47617 22707 47620
rect 22649 47611 22707 47617
rect 23198 47608 23204 47620
rect 23256 47608 23262 47660
rect 24578 47608 24584 47660
rect 24636 47608 24642 47660
rect 18616 47552 24808 47580
rect 8481 47515 8539 47521
rect 8481 47481 8493 47515
rect 8527 47512 8539 47515
rect 24780 47512 24808 47552
rect 24854 47540 24860 47592
rect 24912 47540 24918 47592
rect 26896 47580 26924 47688
rect 27246 47676 27252 47728
rect 27304 47676 27310 47728
rect 28258 47676 28264 47728
rect 28316 47716 28322 47728
rect 38378 47716 38384 47728
rect 28316 47688 38384 47716
rect 28316 47676 28322 47688
rect 38378 47676 38384 47688
rect 38436 47676 38442 47728
rect 27338 47608 27344 47660
rect 27396 47648 27402 47660
rect 29089 47651 29147 47657
rect 29089 47648 29101 47651
rect 27396 47620 29101 47648
rect 27396 47608 27402 47620
rect 29089 47617 29101 47620
rect 29135 47617 29147 47651
rect 29089 47611 29147 47617
rect 32214 47608 32220 47660
rect 32272 47608 32278 47660
rect 34241 47651 34299 47657
rect 34241 47617 34253 47651
rect 34287 47648 34299 47651
rect 34330 47648 34336 47660
rect 34287 47620 34336 47648
rect 34287 47617 34299 47620
rect 34241 47611 34299 47617
rect 34330 47608 34336 47620
rect 34388 47608 34394 47660
rect 36173 47651 36231 47657
rect 36173 47617 36185 47651
rect 36219 47648 36231 47651
rect 36906 47648 36912 47660
rect 36219 47620 36912 47648
rect 36219 47617 36231 47620
rect 36173 47611 36231 47617
rect 36906 47608 36912 47620
rect 36964 47608 36970 47660
rect 38654 47608 38660 47660
rect 38712 47648 38718 47660
rect 38933 47651 38991 47657
rect 38933 47648 38945 47651
rect 38712 47620 38945 47648
rect 38712 47608 38718 47620
rect 38933 47617 38945 47620
rect 38979 47617 38991 47651
rect 38933 47611 38991 47617
rect 41417 47651 41475 47657
rect 41417 47617 41429 47651
rect 41463 47617 41475 47651
rect 41417 47611 41475 47617
rect 32398 47580 32404 47592
rect 26896 47552 32404 47580
rect 32398 47540 32404 47552
rect 32456 47540 32462 47592
rect 36446 47540 36452 47592
rect 36504 47580 36510 47592
rect 41432 47580 41460 47611
rect 43254 47608 43260 47660
rect 43312 47608 43318 47660
rect 45830 47608 45836 47660
rect 45888 47608 45894 47660
rect 45922 47608 45928 47660
rect 45980 47608 45986 47660
rect 36504 47552 41460 47580
rect 36504 47540 36510 47552
rect 42886 47540 42892 47592
rect 42944 47580 42950 47592
rect 43533 47583 43591 47589
rect 43533 47580 43545 47583
rect 42944 47552 43545 47580
rect 42944 47540 42950 47552
rect 43533 47549 43545 47552
rect 43579 47549 43591 47583
rect 43533 47543 43591 47549
rect 46198 47540 46204 47592
rect 46256 47540 46262 47592
rect 27154 47512 27160 47524
rect 8527 47484 22094 47512
rect 24780 47484 27160 47512
rect 8527 47481 8539 47484
rect 8481 47475 8539 47481
rect 18230 47404 18236 47456
rect 18288 47444 18294 47456
rect 18463 47447 18521 47453
rect 18463 47444 18475 47447
rect 18288 47416 18475 47444
rect 18288 47404 18294 47416
rect 18463 47413 18475 47416
rect 18509 47413 18521 47447
rect 18463 47407 18521 47413
rect 19426 47404 19432 47456
rect 19484 47404 19490 47456
rect 22066 47444 22094 47484
rect 27154 47472 27160 47484
rect 27212 47472 27218 47524
rect 27430 47472 27436 47524
rect 27488 47472 27494 47524
rect 31386 47444 31392 47456
rect 22066 47416 31392 47444
rect 31386 47404 31392 47416
rect 31444 47404 31450 47456
rect 31478 47404 31484 47456
rect 31536 47444 31542 47456
rect 33502 47444 33508 47456
rect 31536 47416 33508 47444
rect 31536 47404 31542 47416
rect 33502 47404 33508 47416
rect 33560 47404 33566 47456
rect 38749 47447 38807 47453
rect 38749 47413 38761 47447
rect 38795 47444 38807 47447
rect 38838 47444 38844 47456
rect 38795 47416 38844 47444
rect 38795 47413 38807 47416
rect 38749 47407 38807 47413
rect 38838 47404 38844 47416
rect 38896 47404 38902 47456
rect 45646 47404 45652 47456
rect 45704 47404 45710 47456
rect 1104 47354 47104 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 47104 47354
rect 1104 47280 47104 47302
rect 3050 47200 3056 47252
rect 3108 47200 3114 47252
rect 17310 47200 17316 47252
rect 17368 47240 17374 47252
rect 20625 47243 20683 47249
rect 20625 47240 20637 47243
rect 17368 47212 20637 47240
rect 17368 47200 17374 47212
rect 20625 47209 20637 47212
rect 20671 47240 20683 47243
rect 20671 47212 25452 47240
rect 20671 47209 20683 47212
rect 20625 47203 20683 47209
rect 1118 47132 1124 47184
rect 1176 47172 1182 47184
rect 2133 47175 2191 47181
rect 2133 47172 2145 47175
rect 1176 47144 2145 47172
rect 1176 47132 1182 47144
rect 2133 47141 2145 47144
rect 2179 47141 2191 47175
rect 2133 47135 2191 47141
rect 17773 47107 17831 47113
rect 17773 47073 17785 47107
rect 17819 47104 17831 47107
rect 17862 47104 17868 47116
rect 17819 47076 17868 47104
rect 17819 47073 17831 47076
rect 17773 47067 17831 47073
rect 17862 47064 17868 47076
rect 17920 47064 17926 47116
rect 20254 47064 20260 47116
rect 20312 47104 20318 47116
rect 21729 47107 21787 47113
rect 21729 47104 21741 47107
rect 20312 47076 21741 47104
rect 20312 47064 20318 47076
rect 21729 47073 21741 47076
rect 21775 47073 21787 47107
rect 25424 47104 25452 47212
rect 25682 47200 25688 47252
rect 25740 47240 25746 47252
rect 25777 47243 25835 47249
rect 25777 47240 25789 47243
rect 25740 47212 25789 47240
rect 25740 47200 25746 47212
rect 25777 47209 25789 47212
rect 25823 47240 25835 47243
rect 27249 47243 27307 47249
rect 25823 47212 27200 47240
rect 25823 47209 25835 47212
rect 25777 47203 25835 47209
rect 27172 47172 27200 47212
rect 27249 47209 27261 47243
rect 27295 47240 27307 47243
rect 27338 47240 27344 47252
rect 27295 47212 27344 47240
rect 27295 47209 27307 47212
rect 27249 47203 27307 47209
rect 27338 47200 27344 47212
rect 27396 47200 27402 47252
rect 29178 47200 29184 47252
rect 29236 47240 29242 47252
rect 29917 47243 29975 47249
rect 29917 47240 29929 47243
rect 29236 47212 29929 47240
rect 29236 47200 29242 47212
rect 29917 47209 29929 47212
rect 29963 47240 29975 47243
rect 30098 47240 30104 47252
rect 29963 47212 30104 47240
rect 29963 47209 29975 47212
rect 29917 47203 29975 47209
rect 30098 47200 30104 47212
rect 30156 47200 30162 47252
rect 32214 47240 32220 47252
rect 30208 47212 32220 47240
rect 27172 47144 29684 47172
rect 27341 47107 27399 47113
rect 25424 47076 26004 47104
rect 21729 47067 21787 47073
rect 1673 47039 1731 47045
rect 1673 47005 1685 47039
rect 1719 47036 1731 47039
rect 1946 47036 1952 47048
rect 1719 47008 1952 47036
rect 1719 47005 1731 47008
rect 1673 46999 1731 47005
rect 1946 46996 1952 47008
rect 2004 46996 2010 47048
rect 3237 47039 3295 47045
rect 3237 47005 3249 47039
rect 3283 47036 3295 47039
rect 4617 47039 4675 47045
rect 4617 47036 4629 47039
rect 3283 47008 4629 47036
rect 3283 47005 3295 47008
rect 3237 46999 3295 47005
rect 4617 47005 4629 47008
rect 4663 47036 4675 47039
rect 11330 47036 11336 47048
rect 4663 47008 11336 47036
rect 4663 47005 4675 47008
rect 4617 46999 4675 47005
rect 11330 46996 11336 47008
rect 11388 46996 11394 47048
rect 18141 47039 18199 47045
rect 18141 47005 18153 47039
rect 18187 47005 18199 47039
rect 18141 46999 18199 47005
rect 4884 46971 4942 46977
rect 4884 46937 4896 46971
rect 4930 46937 4942 46971
rect 18156 46968 18184 46999
rect 18230 46996 18236 47048
rect 18288 46996 18294 47048
rect 18414 46996 18420 47048
rect 18472 47036 18478 47048
rect 18509 47039 18567 47045
rect 18509 47036 18521 47039
rect 18472 47008 18521 47036
rect 18472 46996 18478 47008
rect 18509 47005 18521 47008
rect 18555 47036 18567 47039
rect 19242 47036 19248 47048
rect 18555 47008 19248 47036
rect 18555 47005 18567 47008
rect 18509 46999 18567 47005
rect 19242 46996 19248 47008
rect 19300 46996 19306 47048
rect 21085 47039 21143 47045
rect 21085 47005 21097 47039
rect 21131 47036 21143 47039
rect 21358 47036 21364 47048
rect 21131 47008 21364 47036
rect 21131 47005 21143 47008
rect 21085 46999 21143 47005
rect 21358 46996 21364 47008
rect 21416 46996 21422 47048
rect 21744 47036 21772 47067
rect 23474 47036 23480 47048
rect 21744 47008 23480 47036
rect 23474 46996 23480 47008
rect 23532 46996 23538 47048
rect 24213 47039 24271 47045
rect 24213 47005 24225 47039
rect 24259 47005 24271 47039
rect 24213 46999 24271 47005
rect 19490 46971 19548 46977
rect 19490 46968 19502 46971
rect 18156 46940 19502 46968
rect 4884 46931 4942 46937
rect 19490 46937 19502 46940
rect 19536 46937 19548 46971
rect 19490 46931 19548 46937
rect 4798 46860 4804 46912
rect 4856 46900 4862 46912
rect 4908 46900 4936 46931
rect 20346 46928 20352 46980
rect 20404 46968 20410 46980
rect 21996 46971 22054 46977
rect 20404 46940 21036 46968
rect 20404 46928 20410 46940
rect 4856 46872 4936 46900
rect 4856 46860 4862 46872
rect 5994 46860 6000 46912
rect 6052 46860 6058 46912
rect 17126 46860 17132 46912
rect 17184 46860 17190 46912
rect 17494 46860 17500 46912
rect 17552 46860 17558 46912
rect 17586 46860 17592 46912
rect 17644 46860 17650 46912
rect 20898 46860 20904 46912
rect 20956 46860 20962 46912
rect 21008 46900 21036 46940
rect 21996 46937 22008 46971
rect 22042 46968 22054 46971
rect 22370 46968 22376 46980
rect 22042 46940 22376 46968
rect 22042 46937 22054 46940
rect 21996 46931 22054 46937
rect 22370 46928 22376 46940
rect 22428 46928 22434 46980
rect 24228 46968 24256 46999
rect 24394 46996 24400 47048
rect 24452 47036 24458 47048
rect 25869 47039 25927 47045
rect 25869 47036 25881 47039
rect 24452 47008 25881 47036
rect 24452 46996 24458 47008
rect 25869 47005 25881 47008
rect 25915 47005 25927 47039
rect 25976 47036 26004 47076
rect 27341 47073 27353 47107
rect 27387 47104 27399 47107
rect 27387 47076 27936 47104
rect 27387 47073 27399 47076
rect 27341 47067 27399 47073
rect 27908 47048 27936 47076
rect 28258 47064 28264 47116
rect 28316 47064 28322 47116
rect 29656 47104 29684 47144
rect 29822 47132 29828 47184
rect 29880 47172 29886 47184
rect 30009 47175 30067 47181
rect 30009 47172 30021 47175
rect 29880 47144 30021 47172
rect 29880 47132 29886 47144
rect 30009 47141 30021 47144
rect 30055 47141 30067 47175
rect 30009 47135 30067 47141
rect 30208 47104 30236 47212
rect 32214 47200 32220 47212
rect 32272 47200 32278 47252
rect 31113 47175 31171 47181
rect 31113 47141 31125 47175
rect 31159 47172 31171 47175
rect 31938 47172 31944 47184
rect 31159 47144 31944 47172
rect 31159 47141 31171 47144
rect 31113 47135 31171 47141
rect 31938 47132 31944 47144
rect 31996 47132 32002 47184
rect 29196 47076 29592 47104
rect 29656 47076 30236 47104
rect 26694 47036 26700 47048
rect 25976 47008 26700 47036
rect 25869 46999 25927 47005
rect 24642 46971 24700 46977
rect 24642 46968 24654 46971
rect 24228 46940 24654 46968
rect 24642 46937 24654 46940
rect 24688 46937 24700 46971
rect 25884 46968 25912 46999
rect 26694 46996 26700 47008
rect 26752 46996 26758 47048
rect 27062 46996 27068 47048
rect 27120 47036 27126 47048
rect 27617 47039 27675 47045
rect 27617 47036 27629 47039
rect 27120 47008 27629 47036
rect 27120 46996 27126 47008
rect 27617 47005 27629 47008
rect 27663 47005 27675 47039
rect 27617 46999 27675 47005
rect 27890 46996 27896 47048
rect 27948 47036 27954 47048
rect 29196 47045 29224 47076
rect 29564 47045 29592 47076
rect 31386 47064 31392 47116
rect 31444 47104 31450 47116
rect 31573 47107 31631 47113
rect 31573 47104 31585 47107
rect 31444 47076 31585 47104
rect 31444 47064 31450 47076
rect 31573 47073 31585 47076
rect 31619 47073 31631 47107
rect 31573 47067 31631 47073
rect 31757 47107 31815 47113
rect 31757 47073 31769 47107
rect 31803 47073 31815 47107
rect 33318 47104 33324 47116
rect 31757 47067 31815 47073
rect 31956 47076 33324 47104
rect 28537 47039 28595 47045
rect 28537 47036 28549 47039
rect 27948 47008 28549 47036
rect 27948 46996 27954 47008
rect 28537 47005 28549 47008
rect 28583 47005 28595 47039
rect 28537 46999 28595 47005
rect 29181 47039 29239 47045
rect 29181 47005 29193 47039
rect 29227 47005 29239 47039
rect 29181 46999 29239 47005
rect 29365 47039 29423 47045
rect 29365 47005 29377 47039
rect 29411 47005 29423 47039
rect 29365 46999 29423 47005
rect 29549 47039 29607 47045
rect 29549 47005 29561 47039
rect 29595 47036 29607 47039
rect 29595 47008 29960 47036
rect 29595 47005 29607 47008
rect 29549 46999 29607 47005
rect 26142 46977 26148 46980
rect 25884 46940 26096 46968
rect 24642 46931 24700 46937
rect 22922 46900 22928 46912
rect 21008 46872 22928 46900
rect 22922 46860 22928 46872
rect 22980 46860 22986 46912
rect 23109 46903 23167 46909
rect 23109 46869 23121 46903
rect 23155 46900 23167 46903
rect 23198 46900 23204 46912
rect 23155 46872 23204 46900
rect 23155 46869 23167 46872
rect 23109 46863 23167 46869
rect 23198 46860 23204 46872
rect 23256 46860 23262 46912
rect 26068 46900 26096 46940
rect 26136 46931 26148 46977
rect 26142 46928 26148 46931
rect 26200 46928 26206 46980
rect 28350 46928 28356 46980
rect 28408 46968 28414 46980
rect 29380 46968 29408 46999
rect 29733 46971 29791 46977
rect 29733 46968 29745 46971
rect 28408 46940 29745 46968
rect 28408 46928 28414 46940
rect 29733 46937 29745 46940
rect 29779 46937 29791 46971
rect 29733 46931 29791 46937
rect 27062 46900 27068 46912
rect 26068 46872 27068 46900
rect 27062 46860 27068 46872
rect 27120 46860 27126 46912
rect 29270 46860 29276 46912
rect 29328 46860 29334 46912
rect 29932 46900 29960 47008
rect 30098 46996 30104 47048
rect 30156 47036 30162 47048
rect 30193 47039 30251 47045
rect 30193 47036 30205 47039
rect 30156 47008 30205 47036
rect 30156 46996 30162 47008
rect 30193 47005 30205 47008
rect 30239 47005 30251 47039
rect 30193 46999 30251 47005
rect 30282 46996 30288 47048
rect 30340 46996 30346 47048
rect 31478 46996 31484 47048
rect 31536 46996 31542 47048
rect 30006 46928 30012 46980
rect 30064 46928 30070 46980
rect 31496 46968 31524 46996
rect 30116 46940 31524 46968
rect 31772 46968 31800 47067
rect 31956 47045 31984 47076
rect 33318 47064 33324 47076
rect 33376 47064 33382 47116
rect 31941 47039 31999 47045
rect 31941 47005 31953 47039
rect 31987 47005 31999 47039
rect 31941 46999 31999 47005
rect 32214 46996 32220 47048
rect 32272 46996 32278 47048
rect 32876 47008 34928 47036
rect 31772 46940 31984 46968
rect 30116 46900 30144 46940
rect 29932 46872 30144 46900
rect 31956 46900 31984 46940
rect 32876 46900 32904 47008
rect 33502 46928 33508 46980
rect 33560 46968 33566 46980
rect 33597 46971 33655 46977
rect 33597 46968 33609 46971
rect 33560 46940 33609 46968
rect 33560 46928 33566 46940
rect 33597 46937 33609 46940
rect 33643 46937 33655 46971
rect 34900 46968 34928 47008
rect 34974 46996 34980 47048
rect 35032 46996 35038 47048
rect 46753 47039 46811 47045
rect 46753 47005 46765 47039
rect 46799 47036 46811 47039
rect 47670 47036 47676 47048
rect 46799 47008 47676 47036
rect 46799 47005 46811 47008
rect 46753 46999 46811 47005
rect 47670 46996 47676 47008
rect 47728 46996 47734 47048
rect 35434 46968 35440 46980
rect 34900 46940 35440 46968
rect 33597 46931 33655 46937
rect 35434 46928 35440 46940
rect 35492 46928 35498 46980
rect 31956 46872 32904 46900
rect 34790 46860 34796 46912
rect 34848 46860 34854 46912
rect 46566 46860 46572 46912
rect 46624 46860 46630 46912
rect 1104 46810 47104 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 35594 46810
rect 35646 46758 35658 46810
rect 35710 46758 35722 46810
rect 35774 46758 35786 46810
rect 35838 46758 35850 46810
rect 35902 46758 47104 46810
rect 1104 46736 47104 46758
rect 1302 46656 1308 46708
rect 1360 46696 1366 46708
rect 1581 46699 1639 46705
rect 1581 46696 1593 46699
rect 1360 46668 1593 46696
rect 1360 46656 1366 46668
rect 1581 46665 1593 46668
rect 1627 46665 1639 46699
rect 1581 46659 1639 46665
rect 17494 46656 17500 46708
rect 17552 46696 17558 46708
rect 18049 46699 18107 46705
rect 18049 46696 18061 46699
rect 17552 46668 18061 46696
rect 17552 46656 17558 46668
rect 18049 46665 18061 46668
rect 18095 46665 18107 46699
rect 18049 46659 18107 46665
rect 19613 46699 19671 46705
rect 19613 46665 19625 46699
rect 19659 46696 19671 46699
rect 20254 46696 20260 46708
rect 19659 46668 20260 46696
rect 19659 46665 19671 46668
rect 19613 46659 19671 46665
rect 20254 46656 20260 46668
rect 20312 46656 20318 46708
rect 20530 46656 20536 46708
rect 20588 46696 20594 46708
rect 21545 46699 21603 46705
rect 21545 46696 21557 46699
rect 20588 46668 21557 46696
rect 20588 46656 20594 46668
rect 21545 46665 21557 46668
rect 21591 46665 21603 46699
rect 21545 46659 21603 46665
rect 22370 46656 22376 46708
rect 22428 46656 22434 46708
rect 25133 46699 25191 46705
rect 25133 46696 25145 46699
rect 22756 46668 25145 46696
rect 1489 46631 1547 46637
rect 1489 46597 1501 46631
rect 1535 46628 1547 46631
rect 5994 46628 6000 46640
rect 1535 46600 6000 46628
rect 1535 46597 1547 46600
rect 1489 46591 1547 46597
rect 5994 46588 6000 46600
rect 6052 46628 6058 46640
rect 20432 46631 20490 46637
rect 6052 46600 18644 46628
rect 6052 46588 6058 46600
rect 4798 46520 4804 46572
rect 4856 46560 4862 46572
rect 16942 46569 16948 46572
rect 5077 46563 5135 46569
rect 5077 46560 5089 46563
rect 4856 46532 5089 46560
rect 4856 46520 4862 46532
rect 5077 46529 5089 46532
rect 5123 46529 5135 46563
rect 5077 46523 5135 46529
rect 16936 46523 16948 46569
rect 16942 46520 16948 46523
rect 17000 46520 17006 46572
rect 17954 46520 17960 46572
rect 18012 46560 18018 46572
rect 18489 46563 18547 46569
rect 18489 46560 18501 46563
rect 18012 46532 18501 46560
rect 18012 46520 18018 46532
rect 18489 46529 18501 46532
rect 18535 46529 18547 46563
rect 18616 46560 18644 46600
rect 20432 46597 20444 46631
rect 20478 46628 20490 46631
rect 20898 46628 20904 46640
rect 20478 46600 20904 46628
rect 20478 46597 20490 46600
rect 20432 46591 20490 46597
rect 20898 46588 20904 46600
rect 20956 46588 20962 46640
rect 22756 46628 22784 46668
rect 25133 46665 25145 46668
rect 25179 46665 25191 46699
rect 25133 46659 25191 46665
rect 26513 46699 26571 46705
rect 26513 46665 26525 46699
rect 26559 46696 26571 46699
rect 27338 46696 27344 46708
rect 26559 46668 27344 46696
rect 26559 46665 26571 46668
rect 26513 46659 26571 46665
rect 23385 46631 23443 46637
rect 23385 46628 23397 46631
rect 22066 46600 22784 46628
rect 22848 46600 23397 46628
rect 22066 46560 22094 46600
rect 18616 46532 22094 46560
rect 22557 46563 22615 46569
rect 18489 46523 18547 46529
rect 22557 46529 22569 46563
rect 22603 46560 22615 46563
rect 22738 46560 22744 46572
rect 22603 46532 22744 46560
rect 22603 46529 22615 46532
rect 22557 46523 22615 46529
rect 22738 46520 22744 46532
rect 22796 46520 22802 46572
rect 22848 46569 22876 46600
rect 23385 46597 23397 46600
rect 23431 46597 23443 46631
rect 25148 46628 25176 46659
rect 27338 46656 27344 46668
rect 27396 46656 27402 46708
rect 29270 46656 29276 46708
rect 29328 46696 29334 46708
rect 30282 46696 30288 46708
rect 29328 46668 30288 46696
rect 29328 46656 29334 46668
rect 30282 46656 30288 46668
rect 30340 46656 30346 46708
rect 32125 46699 32183 46705
rect 32125 46665 32137 46699
rect 32171 46696 32183 46699
rect 32214 46696 32220 46708
rect 32171 46668 32220 46696
rect 32171 46665 32183 46668
rect 32125 46659 32183 46665
rect 32214 46656 32220 46668
rect 32272 46656 32278 46708
rect 34974 46656 34980 46708
rect 35032 46696 35038 46708
rect 35437 46699 35495 46705
rect 35437 46696 35449 46699
rect 35032 46668 35449 46696
rect 35032 46656 35038 46668
rect 35437 46665 35449 46668
rect 35483 46665 35495 46699
rect 35437 46659 35495 46665
rect 26421 46631 26479 46637
rect 25148 46600 25820 46628
rect 23385 46591 23443 46597
rect 22833 46563 22891 46569
rect 22833 46529 22845 46563
rect 22879 46529 22891 46563
rect 22833 46523 22891 46529
rect 23014 46520 23020 46572
rect 23072 46520 23078 46572
rect 23106 46520 23112 46572
rect 23164 46520 23170 46572
rect 23474 46520 23480 46572
rect 23532 46520 23538 46572
rect 23744 46563 23802 46569
rect 23744 46529 23756 46563
rect 23790 46560 23802 46563
rect 25314 46560 25320 46572
rect 23790 46532 25320 46560
rect 23790 46529 23802 46532
rect 23744 46523 23802 46529
rect 25314 46520 25320 46532
rect 25372 46520 25378 46572
rect 25501 46563 25559 46569
rect 25501 46529 25513 46563
rect 25547 46529 25559 46563
rect 25501 46523 25559 46529
rect 16669 46495 16727 46501
rect 16669 46461 16681 46495
rect 16715 46461 16727 46495
rect 16669 46455 16727 46461
rect 15654 46316 15660 46368
rect 15712 46356 15718 46368
rect 16684 46356 16712 46455
rect 17678 46452 17684 46504
rect 17736 46492 17742 46504
rect 18233 46495 18291 46501
rect 18233 46492 18245 46495
rect 17736 46464 18245 46492
rect 17736 46452 17742 46464
rect 18233 46461 18245 46464
rect 18279 46461 18291 46495
rect 18233 46455 18291 46461
rect 20162 46452 20168 46504
rect 20220 46452 20226 46504
rect 22646 46452 22652 46504
rect 22704 46492 22710 46504
rect 23201 46495 23259 46501
rect 23201 46492 23213 46495
rect 22704 46464 23213 46492
rect 22704 46452 22710 46464
rect 23201 46461 23213 46464
rect 23247 46461 23259 46495
rect 23201 46455 23259 46461
rect 23290 46452 23296 46504
rect 23348 46492 23354 46504
rect 23385 46495 23443 46501
rect 23385 46492 23397 46495
rect 23348 46464 23397 46492
rect 23348 46452 23354 46464
rect 23385 46461 23397 46464
rect 23431 46461 23443 46495
rect 25516 46492 25544 46523
rect 25682 46520 25688 46572
rect 25740 46520 25746 46572
rect 25792 46569 25820 46600
rect 26421 46597 26433 46631
rect 26467 46628 26479 46631
rect 28534 46628 28540 46640
rect 26467 46600 28540 46628
rect 26467 46597 26479 46600
rect 26421 46591 26479 46597
rect 28534 46588 28540 46600
rect 28592 46588 28598 46640
rect 34232 46631 34290 46637
rect 30208 46600 31754 46628
rect 25777 46563 25835 46569
rect 25777 46529 25789 46563
rect 25823 46529 25835 46563
rect 25777 46523 25835 46529
rect 26973 46563 27031 46569
rect 26973 46529 26985 46563
rect 27019 46560 27031 46563
rect 27062 46560 27068 46572
rect 27019 46532 27068 46560
rect 27019 46529 27031 46532
rect 26973 46523 27031 46529
rect 27062 46520 27068 46532
rect 27120 46520 27126 46572
rect 27246 46569 27252 46572
rect 27240 46523 27252 46569
rect 27246 46520 27252 46523
rect 27304 46520 27310 46572
rect 29641 46563 29699 46569
rect 29641 46560 29653 46563
rect 29012 46532 29653 46560
rect 29012 46501 29040 46532
rect 29641 46529 29653 46532
rect 29687 46529 29699 46563
rect 29641 46523 29699 46529
rect 29822 46520 29828 46572
rect 29880 46520 29886 46572
rect 30208 46569 30236 46600
rect 30193 46563 30251 46569
rect 30193 46529 30205 46563
rect 30239 46529 30251 46563
rect 30193 46523 30251 46529
rect 30282 46520 30288 46572
rect 30340 46560 30346 46572
rect 30449 46563 30507 46569
rect 30449 46560 30461 46563
rect 30340 46532 30461 46560
rect 30340 46520 30346 46532
rect 30449 46529 30461 46532
rect 30495 46529 30507 46563
rect 30449 46523 30507 46529
rect 23385 46455 23443 46461
rect 24872 46464 25544 46492
rect 26697 46495 26755 46501
rect 22741 46427 22799 46433
rect 22741 46393 22753 46427
rect 22787 46424 22799 46427
rect 23308 46424 23336 46452
rect 22787 46396 23336 46424
rect 22787 46393 22799 46396
rect 22741 46387 22799 46393
rect 19426 46356 19432 46368
rect 15712 46328 19432 46356
rect 15712 46316 15718 46328
rect 19426 46316 19432 46328
rect 19484 46316 19490 46368
rect 22922 46316 22928 46368
rect 22980 46356 22986 46368
rect 24872 46365 24900 46464
rect 26697 46461 26709 46495
rect 26743 46492 26755 46495
rect 28997 46495 29055 46501
rect 26743 46464 27016 46492
rect 26743 46461 26755 46464
rect 26697 46455 26755 46461
rect 25961 46427 26019 46433
rect 25961 46393 25973 46427
rect 26007 46424 26019 46427
rect 26878 46424 26884 46436
rect 26007 46396 26884 46424
rect 26007 46393 26019 46396
rect 25961 46387 26019 46393
rect 26878 46384 26884 46396
rect 26936 46384 26942 46436
rect 24857 46359 24915 46365
rect 24857 46356 24869 46359
rect 22980 46328 24869 46356
rect 22980 46316 22986 46328
rect 24857 46325 24869 46328
rect 24903 46325 24915 46359
rect 24857 46319 24915 46325
rect 25777 46359 25835 46365
rect 25777 46325 25789 46359
rect 25823 46356 25835 46359
rect 25866 46356 25872 46368
rect 25823 46328 25872 46356
rect 25823 46325 25835 46328
rect 25777 46319 25835 46325
rect 25866 46316 25872 46328
rect 25924 46316 25930 46368
rect 26053 46359 26111 46365
rect 26053 46325 26065 46359
rect 26099 46356 26111 46359
rect 26326 46356 26332 46368
rect 26099 46328 26332 46356
rect 26099 46325 26111 46328
rect 26053 46319 26111 46325
rect 26326 46316 26332 46328
rect 26384 46316 26390 46368
rect 26988 46356 27016 46464
rect 28997 46461 29009 46495
rect 29043 46461 29055 46495
rect 28997 46455 29055 46461
rect 29178 46452 29184 46504
rect 29236 46452 29242 46504
rect 29270 46452 29276 46504
rect 29328 46452 29334 46504
rect 29365 46495 29423 46501
rect 29365 46461 29377 46495
rect 29411 46461 29423 46495
rect 29365 46455 29423 46461
rect 29380 46424 29408 46455
rect 29454 46452 29460 46504
rect 29512 46452 29518 46504
rect 31726 46492 31754 46600
rect 34232 46597 34244 46631
rect 34278 46628 34290 46631
rect 34790 46628 34796 46640
rect 34278 46600 34796 46628
rect 34278 46597 34290 46600
rect 34232 46591 34290 46597
rect 34790 46588 34796 46600
rect 34848 46588 34854 46640
rect 31938 46520 31944 46572
rect 31996 46560 32002 46572
rect 32309 46563 32367 46569
rect 32309 46560 32321 46563
rect 31996 46532 32321 46560
rect 31996 46520 32002 46532
rect 32309 46529 32321 46532
rect 32355 46529 32367 46563
rect 35710 46560 35716 46572
rect 32309 46523 32367 46529
rect 33060 46532 35716 46560
rect 33060 46501 33088 46532
rect 35710 46520 35716 46532
rect 35768 46520 35774 46572
rect 35802 46520 35808 46572
rect 35860 46520 35866 46572
rect 35897 46563 35955 46569
rect 35897 46529 35909 46563
rect 35943 46560 35955 46563
rect 36725 46563 36783 46569
rect 35943 46532 36676 46560
rect 35943 46529 35955 46532
rect 35897 46523 35955 46529
rect 33045 46495 33103 46501
rect 33045 46492 33057 46495
rect 31726 46464 33057 46492
rect 33045 46461 33057 46464
rect 33091 46461 33103 46495
rect 33045 46455 33103 46461
rect 33318 46452 33324 46504
rect 33376 46492 33382 46504
rect 33965 46495 34023 46501
rect 33965 46492 33977 46495
rect 33376 46464 33977 46492
rect 33376 46452 33382 46464
rect 33965 46461 33977 46464
rect 34011 46461 34023 46495
rect 33965 46455 34023 46461
rect 35434 46452 35440 46504
rect 35492 46492 35498 46504
rect 35989 46495 36047 46501
rect 35989 46492 36001 46495
rect 35492 46464 36001 46492
rect 35492 46452 35498 46464
rect 35989 46461 36001 46464
rect 36035 46461 36047 46495
rect 36648 46492 36676 46532
rect 36725 46529 36737 46563
rect 36771 46560 36783 46563
rect 37274 46560 37280 46572
rect 36771 46532 37280 46560
rect 36771 46529 36783 46532
rect 36725 46523 36783 46529
rect 37274 46520 37280 46532
rect 37332 46520 37338 46572
rect 45646 46492 45652 46504
rect 36648 46464 45652 46492
rect 35989 46455 36047 46461
rect 29546 46424 29552 46436
rect 29380 46396 29552 46424
rect 29546 46384 29552 46396
rect 29604 46424 29610 46436
rect 30006 46424 30012 46436
rect 29604 46396 30012 46424
rect 29604 46384 29610 46396
rect 30006 46384 30012 46396
rect 30064 46384 30070 46436
rect 36004 46424 36032 46455
rect 45646 46452 45652 46464
rect 45704 46452 45710 46504
rect 37366 46424 37372 46436
rect 36004 46396 37372 46424
rect 37366 46384 37372 46396
rect 37424 46384 37430 46436
rect 27338 46356 27344 46368
rect 26988 46328 27344 46356
rect 27338 46316 27344 46328
rect 27396 46316 27402 46368
rect 27614 46316 27620 46368
rect 27672 46356 27678 46368
rect 28350 46356 28356 46368
rect 27672 46328 28356 46356
rect 27672 46316 27678 46328
rect 28350 46316 28356 46328
rect 28408 46356 28414 46368
rect 28626 46356 28632 46368
rect 28408 46328 28632 46356
rect 28408 46316 28414 46328
rect 28626 46316 28632 46328
rect 28684 46316 28690 46368
rect 29638 46316 29644 46368
rect 29696 46316 29702 46368
rect 30834 46316 30840 46368
rect 30892 46356 30898 46368
rect 31573 46359 31631 46365
rect 31573 46356 31585 46359
rect 30892 46328 31585 46356
rect 30892 46316 30898 46328
rect 31573 46325 31585 46328
rect 31619 46325 31631 46359
rect 31573 46319 31631 46325
rect 35342 46316 35348 46368
rect 35400 46316 35406 46368
rect 36354 46316 36360 46368
rect 36412 46356 36418 46368
rect 36541 46359 36599 46365
rect 36541 46356 36553 46359
rect 36412 46328 36553 46356
rect 36412 46316 36418 46328
rect 36541 46325 36553 46328
rect 36587 46325 36599 46359
rect 36541 46319 36599 46325
rect 1104 46266 47104 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 47104 46266
rect 1104 46192 47104 46214
rect 16942 46112 16948 46164
rect 17000 46112 17006 46164
rect 21174 46112 21180 46164
rect 21232 46112 21238 46164
rect 21358 46112 21364 46164
rect 21416 46112 21422 46164
rect 22646 46112 22652 46164
rect 22704 46152 22710 46164
rect 23017 46155 23075 46161
rect 23017 46152 23029 46155
rect 22704 46124 23029 46152
rect 22704 46112 22710 46124
rect 23017 46121 23029 46124
rect 23063 46121 23075 46155
rect 23017 46115 23075 46121
rect 25314 46112 25320 46164
rect 25372 46112 25378 46164
rect 26142 46112 26148 46164
rect 26200 46112 26206 46164
rect 27246 46112 27252 46164
rect 27304 46152 27310 46164
rect 27341 46155 27399 46161
rect 27341 46152 27353 46155
rect 27304 46124 27353 46152
rect 27304 46112 27310 46124
rect 27341 46121 27353 46124
rect 27387 46121 27399 46155
rect 27341 46115 27399 46121
rect 27706 46112 27712 46164
rect 27764 46152 27770 46164
rect 28166 46152 28172 46164
rect 27764 46124 28172 46152
rect 27764 46112 27770 46124
rect 28166 46112 28172 46124
rect 28224 46152 28230 46164
rect 30101 46155 30159 46161
rect 28224 46124 29408 46152
rect 28224 46112 28230 46124
rect 17405 46087 17463 46093
rect 17405 46053 17417 46087
rect 17451 46084 17463 46087
rect 18046 46084 18052 46096
rect 17451 46056 18052 46084
rect 17451 46053 17463 46056
rect 17405 46047 17463 46053
rect 18046 46044 18052 46056
rect 18104 46044 18110 46096
rect 17862 45976 17868 46028
rect 17920 46016 17926 46028
rect 17957 46019 18015 46025
rect 17957 46016 17969 46019
rect 17920 45988 17969 46016
rect 17920 45976 17926 45988
rect 17957 45985 17969 45988
rect 18003 45985 18015 46019
rect 17957 45979 18015 45985
rect 18233 46019 18291 46025
rect 18233 45985 18245 46019
rect 18279 46016 18291 46019
rect 19426 46016 19432 46028
rect 18279 45988 19432 46016
rect 18279 45985 18291 45988
rect 18233 45979 18291 45985
rect 19426 45976 19432 45988
rect 19484 45976 19490 46028
rect 20165 46019 20223 46025
rect 20165 45985 20177 46019
rect 20211 46016 20223 46019
rect 20211 45988 22508 46016
rect 20211 45985 20223 45988
rect 20165 45979 20223 45985
rect 17126 45908 17132 45960
rect 17184 45908 17190 45960
rect 17494 45908 17500 45960
rect 17552 45948 17558 45960
rect 17773 45951 17831 45957
rect 17773 45948 17785 45951
rect 17552 45920 17785 45948
rect 17552 45908 17558 45920
rect 17773 45917 17785 45920
rect 17819 45917 17831 45951
rect 17773 45911 17831 45917
rect 18509 45951 18567 45957
rect 18509 45917 18521 45951
rect 18555 45917 18567 45951
rect 18509 45911 18567 45917
rect 17678 45840 17684 45892
rect 17736 45880 17742 45892
rect 18524 45880 18552 45911
rect 20346 45908 20352 45960
rect 20404 45908 20410 45960
rect 20625 45951 20683 45957
rect 20625 45917 20637 45951
rect 20671 45917 20683 45951
rect 20625 45911 20683 45917
rect 20809 45951 20867 45957
rect 20809 45917 20821 45951
rect 20855 45948 20867 45951
rect 20898 45948 20904 45960
rect 20855 45920 20904 45948
rect 20855 45917 20867 45920
rect 20809 45911 20867 45917
rect 20640 45880 20668 45911
rect 20898 45908 20904 45920
rect 20956 45908 20962 45960
rect 17736 45852 18552 45880
rect 19996 45852 20668 45880
rect 21177 45883 21235 45889
rect 17736 45840 17742 45852
rect 19996 45824 20024 45852
rect 21177 45849 21189 45883
rect 21223 45880 21235 45883
rect 21223 45852 21680 45880
rect 21223 45849 21235 45852
rect 21177 45843 21235 45849
rect 15930 45772 15936 45824
rect 15988 45812 15994 45824
rect 17586 45812 17592 45824
rect 15988 45784 17592 45812
rect 15988 45772 15994 45784
rect 17586 45772 17592 45784
rect 17644 45812 17650 45824
rect 17865 45815 17923 45821
rect 17865 45812 17877 45815
rect 17644 45784 17877 45812
rect 17644 45772 17650 45784
rect 17865 45781 17877 45784
rect 17911 45812 17923 45815
rect 19978 45812 19984 45824
rect 17911 45784 19984 45812
rect 17911 45781 17923 45784
rect 17865 45775 17923 45781
rect 19978 45772 19984 45784
rect 20036 45772 20042 45824
rect 20162 45772 20168 45824
rect 20220 45812 20226 45824
rect 20530 45812 20536 45824
rect 20220 45784 20536 45812
rect 20220 45772 20226 45784
rect 20530 45772 20536 45784
rect 20588 45772 20594 45824
rect 21652 45812 21680 45852
rect 22370 45812 22376 45824
rect 21652 45784 22376 45812
rect 22370 45772 22376 45784
rect 22428 45772 22434 45824
rect 22480 45812 22508 45988
rect 22557 45951 22615 45957
rect 22557 45917 22569 45951
rect 22603 45948 22615 45951
rect 22664 45948 22692 46112
rect 22738 46044 22744 46096
rect 22796 46084 22802 46096
rect 23106 46084 23112 46096
rect 22796 46056 23112 46084
rect 22796 46044 22802 46056
rect 23106 46044 23112 46056
rect 23164 46044 23170 46096
rect 23290 46044 23296 46096
rect 23348 46084 23354 46096
rect 28629 46087 28687 46093
rect 28629 46084 28641 46087
rect 23348 46056 28641 46084
rect 23348 46044 23354 46056
rect 28629 46053 28641 46056
rect 28675 46053 28687 46087
rect 28629 46047 28687 46053
rect 22925 46019 22983 46025
rect 22925 45985 22937 46019
rect 22971 46016 22983 46019
rect 22971 45988 23520 46016
rect 22971 45985 22983 45988
rect 22925 45979 22983 45985
rect 22603 45920 22692 45948
rect 22603 45917 22615 45920
rect 22557 45911 22615 45917
rect 22738 45908 22744 45960
rect 22796 45908 22802 45960
rect 23017 45951 23075 45957
rect 23017 45917 23029 45951
rect 23063 45948 23075 45951
rect 23106 45948 23112 45960
rect 23063 45920 23112 45948
rect 23063 45917 23075 45920
rect 23017 45911 23075 45917
rect 23106 45908 23112 45920
rect 23164 45908 23170 45960
rect 23198 45908 23204 45960
rect 23256 45908 23262 45960
rect 23290 45908 23296 45960
rect 23348 45908 23354 45960
rect 23492 45957 23520 45988
rect 23566 45976 23572 46028
rect 23624 46016 23630 46028
rect 24673 46019 24731 46025
rect 24673 46016 24685 46019
rect 23624 45988 24685 46016
rect 23624 45976 23630 45988
rect 24673 45985 24685 45988
rect 24719 45985 24731 46019
rect 27709 46019 27767 46025
rect 24673 45979 24731 45985
rect 25608 45988 26280 46016
rect 25608 45960 25636 45988
rect 23477 45951 23535 45957
rect 23477 45917 23489 45951
rect 23523 45917 23535 45951
rect 23477 45911 23535 45917
rect 24394 45908 24400 45960
rect 24452 45908 24458 45960
rect 25590 45908 25596 45960
rect 25648 45908 25654 45960
rect 25774 45908 25780 45960
rect 25832 45908 25838 45960
rect 25958 45908 25964 45960
rect 26016 45908 26022 45960
rect 26053 45951 26111 45957
rect 26053 45917 26065 45951
rect 26099 45917 26111 45951
rect 26053 45911 26111 45917
rect 26068 45880 26096 45911
rect 22848 45852 26096 45880
rect 26252 45880 26280 45988
rect 27709 45985 27721 46019
rect 27755 46016 27767 46019
rect 28258 46016 28264 46028
rect 27755 45988 28264 46016
rect 27755 45985 27767 45988
rect 27709 45979 27767 45985
rect 28258 45976 28264 45988
rect 28316 45976 28322 46028
rect 28445 46019 28503 46025
rect 28445 45985 28457 46019
rect 28491 46016 28503 46019
rect 29270 46016 29276 46028
rect 28491 45988 29276 46016
rect 28491 45985 28503 45988
rect 28445 45979 28503 45985
rect 29270 45976 29276 45988
rect 29328 45976 29334 46028
rect 29380 46016 29408 46124
rect 30101 46121 30113 46155
rect 30147 46152 30159 46155
rect 30282 46152 30288 46164
rect 30147 46124 30288 46152
rect 30147 46121 30159 46124
rect 30101 46115 30159 46121
rect 30282 46112 30288 46124
rect 30340 46112 30346 46164
rect 29454 46044 29460 46096
rect 29512 46084 29518 46096
rect 30469 46087 30527 46093
rect 30469 46084 30481 46087
rect 29512 46056 30481 46084
rect 29512 46044 29518 46056
rect 30469 46053 30481 46056
rect 30515 46053 30527 46087
rect 30469 46047 30527 46053
rect 30377 46019 30435 46025
rect 30377 46016 30389 46019
rect 29380 45988 30389 46016
rect 30377 45985 30389 45988
rect 30423 46016 30435 46019
rect 33226 46016 33232 46028
rect 30423 45988 33232 46016
rect 30423 45985 30435 45988
rect 30377 45979 30435 45985
rect 33226 45976 33232 45988
rect 33284 45976 33290 46028
rect 35434 45976 35440 46028
rect 35492 46016 35498 46028
rect 35710 46016 35716 46028
rect 35492 45988 35716 46016
rect 35492 45976 35498 45988
rect 35710 45976 35716 45988
rect 35768 46016 35774 46028
rect 36081 46019 36139 46025
rect 36081 46016 36093 46019
rect 35768 45988 36093 46016
rect 35768 45976 35774 45988
rect 36081 45985 36093 45988
rect 36127 45985 36139 46019
rect 36081 45979 36139 45985
rect 26326 45908 26332 45960
rect 26384 45908 26390 45960
rect 27154 45908 27160 45960
rect 27212 45948 27218 45960
rect 27522 45948 27528 45960
rect 27212 45920 27528 45948
rect 27212 45908 27218 45920
rect 27522 45908 27528 45920
rect 27580 45908 27586 45960
rect 27614 45908 27620 45960
rect 27672 45908 27678 45960
rect 27801 45951 27859 45957
rect 27801 45917 27813 45951
rect 27847 45917 27859 45951
rect 27801 45911 27859 45917
rect 27816 45880 27844 45911
rect 27982 45908 27988 45960
rect 28040 45908 28046 45960
rect 28905 45951 28963 45957
rect 28905 45917 28917 45951
rect 28951 45948 28963 45951
rect 29178 45948 29184 45960
rect 28951 45920 29184 45948
rect 28951 45917 28963 45920
rect 28905 45911 28963 45917
rect 29178 45908 29184 45920
rect 29236 45908 29242 45960
rect 30285 45951 30343 45957
rect 30285 45917 30297 45951
rect 30331 45948 30343 45951
rect 30466 45948 30472 45960
rect 30331 45920 30472 45948
rect 30331 45917 30343 45920
rect 30285 45911 30343 45917
rect 30466 45908 30472 45920
rect 30524 45908 30530 45960
rect 30558 45908 30564 45960
rect 30616 45908 30622 45960
rect 30745 45951 30803 45957
rect 30745 45917 30757 45951
rect 30791 45917 30803 45951
rect 30745 45911 30803 45917
rect 28350 45880 28356 45892
rect 26252 45852 28356 45880
rect 22848 45812 22876 45852
rect 28350 45840 28356 45852
rect 28408 45880 28414 45892
rect 30760 45880 30788 45911
rect 30834 45908 30840 45960
rect 30892 45908 30898 45960
rect 33045 45951 33103 45957
rect 33045 45917 33057 45951
rect 33091 45948 33103 45951
rect 33505 45951 33563 45957
rect 33505 45948 33517 45951
rect 33091 45920 33517 45948
rect 33091 45917 33103 45920
rect 33045 45911 33103 45917
rect 33505 45917 33517 45920
rect 33551 45917 33563 45951
rect 33505 45911 33563 45917
rect 33134 45880 33140 45892
rect 28408 45852 30788 45880
rect 31036 45852 33140 45880
rect 28408 45840 28414 45852
rect 22480 45784 22876 45812
rect 22922 45772 22928 45824
rect 22980 45812 22986 45824
rect 23385 45815 23443 45821
rect 23385 45812 23397 45815
rect 22980 45784 23397 45812
rect 22980 45772 22986 45784
rect 23385 45781 23397 45784
rect 23431 45781 23443 45815
rect 23385 45775 23443 45781
rect 25685 45815 25743 45821
rect 25685 45781 25697 45815
rect 25731 45812 25743 45815
rect 27614 45812 27620 45824
rect 25731 45784 27620 45812
rect 25731 45781 25743 45784
rect 25685 45775 25743 45781
rect 27614 45772 27620 45784
rect 27672 45772 27678 45824
rect 28813 45815 28871 45821
rect 28813 45781 28825 45815
rect 28859 45812 28871 45815
rect 29546 45812 29552 45824
rect 28859 45784 29552 45812
rect 28859 45781 28871 45784
rect 28813 45775 28871 45781
rect 29546 45772 29552 45784
rect 29604 45772 29610 45824
rect 30374 45772 30380 45824
rect 30432 45812 30438 45824
rect 30650 45812 30656 45824
rect 30432 45784 30656 45812
rect 30432 45772 30438 45784
rect 30650 45772 30656 45784
rect 30708 45812 30714 45824
rect 31036 45821 31064 45852
rect 33134 45840 33140 45852
rect 33192 45880 33198 45892
rect 33229 45883 33287 45889
rect 33229 45880 33241 45883
rect 33192 45852 33241 45880
rect 33192 45840 33198 45852
rect 33229 45849 33241 45852
rect 33275 45849 33287 45883
rect 33520 45880 33548 45911
rect 33686 45908 33692 45960
rect 33744 45908 33750 45960
rect 34790 45908 34796 45960
rect 34848 45948 34854 45960
rect 35342 45948 35348 45960
rect 34848 45920 35348 45948
rect 34848 45908 34854 45920
rect 35342 45908 35348 45920
rect 35400 45908 35406 45960
rect 36354 45957 36360 45960
rect 36348 45948 36360 45957
rect 36315 45920 36360 45948
rect 36348 45911 36360 45920
rect 36354 45908 36360 45911
rect 36412 45908 36418 45960
rect 33520 45852 36768 45880
rect 33229 45843 33287 45849
rect 36740 45824 36768 45852
rect 31021 45815 31079 45821
rect 31021 45812 31033 45815
rect 30708 45784 31033 45812
rect 30708 45772 30714 45784
rect 31021 45781 31033 45784
rect 31067 45781 31079 45815
rect 31021 45775 31079 45781
rect 33410 45772 33416 45824
rect 33468 45772 33474 45824
rect 33686 45772 33692 45824
rect 33744 45772 33750 45824
rect 34422 45772 34428 45824
rect 34480 45812 34486 45824
rect 34885 45815 34943 45821
rect 34885 45812 34897 45815
rect 34480 45784 34897 45812
rect 34480 45772 34486 45784
rect 34885 45781 34897 45784
rect 34931 45812 34943 45815
rect 35802 45812 35808 45824
rect 34931 45784 35808 45812
rect 34931 45781 34943 45784
rect 34885 45775 34943 45781
rect 35802 45772 35808 45784
rect 35860 45772 35866 45824
rect 36722 45772 36728 45824
rect 36780 45812 36786 45824
rect 37461 45815 37519 45821
rect 37461 45812 37473 45815
rect 36780 45784 37473 45812
rect 36780 45772 36786 45784
rect 37461 45781 37473 45784
rect 37507 45781 37519 45815
rect 37461 45775 37519 45781
rect 1104 45722 47104 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 35594 45722
rect 35646 45670 35658 45722
rect 35710 45670 35722 45722
rect 35774 45670 35786 45722
rect 35838 45670 35850 45722
rect 35902 45670 47104 45722
rect 1104 45648 47104 45670
rect 20898 45568 20904 45620
rect 20956 45608 20962 45620
rect 25958 45608 25964 45620
rect 20956 45580 25964 45608
rect 20956 45568 20962 45580
rect 25958 45568 25964 45580
rect 26016 45568 26022 45620
rect 27982 45568 27988 45620
rect 28040 45608 28046 45620
rect 28445 45611 28503 45617
rect 28445 45608 28457 45611
rect 28040 45580 28457 45608
rect 28040 45568 28046 45580
rect 28445 45577 28457 45580
rect 28491 45577 28503 45611
rect 28445 45571 28503 45577
rect 28626 45568 28632 45620
rect 28684 45608 28690 45620
rect 28810 45608 28816 45620
rect 28684 45580 28816 45608
rect 28684 45568 28690 45580
rect 28810 45568 28816 45580
rect 28868 45608 28874 45620
rect 28868 45580 29859 45608
rect 28868 45568 28874 45580
rect 22370 45500 22376 45552
rect 22428 45540 22434 45552
rect 22830 45540 22836 45552
rect 22428 45512 22836 45540
rect 22428 45500 22434 45512
rect 22830 45500 22836 45512
rect 22888 45540 22894 45552
rect 23290 45540 23296 45552
rect 22888 45512 23296 45540
rect 22888 45500 22894 45512
rect 23290 45500 23296 45512
rect 23348 45500 23354 45552
rect 29638 45540 29644 45552
rect 29012 45512 29644 45540
rect 16850 45432 16856 45484
rect 16908 45472 16914 45484
rect 17037 45475 17095 45481
rect 17037 45472 17049 45475
rect 16908 45444 17049 45472
rect 16908 45432 16914 45444
rect 17037 45441 17049 45444
rect 17083 45441 17095 45475
rect 17862 45472 17868 45484
rect 17037 45435 17095 45441
rect 17328 45444 17868 45472
rect 17328 45416 17356 45444
rect 17862 45432 17868 45444
rect 17920 45432 17926 45484
rect 18046 45432 18052 45484
rect 18104 45432 18110 45484
rect 19978 45432 19984 45484
rect 20036 45432 20042 45484
rect 20162 45432 20168 45484
rect 20220 45432 20226 45484
rect 28629 45475 28687 45481
rect 28629 45441 28641 45475
rect 28675 45441 28687 45475
rect 28629 45435 28687 45441
rect 17126 45364 17132 45416
rect 17184 45364 17190 45416
rect 17310 45364 17316 45416
rect 17368 45364 17374 45416
rect 28644 45404 28672 45435
rect 28718 45432 28724 45484
rect 28776 45432 28782 45484
rect 28813 45475 28871 45481
rect 28813 45441 28825 45475
rect 28859 45472 28871 45475
rect 28902 45472 28908 45484
rect 28859 45444 28908 45472
rect 28859 45441 28871 45444
rect 28813 45435 28871 45441
rect 28902 45432 28908 45444
rect 28960 45432 28966 45484
rect 29012 45481 29040 45512
rect 29638 45500 29644 45512
rect 29696 45500 29702 45552
rect 28997 45475 29055 45481
rect 28997 45441 29009 45475
rect 29043 45441 29055 45475
rect 28997 45435 29055 45441
rect 29089 45475 29147 45481
rect 29089 45441 29101 45475
rect 29135 45472 29147 45475
rect 29270 45472 29276 45484
rect 29135 45444 29276 45472
rect 29135 45441 29147 45444
rect 29089 45435 29147 45441
rect 29270 45432 29276 45444
rect 29328 45432 29334 45484
rect 29181 45407 29239 45413
rect 29181 45404 29193 45407
rect 28644 45376 29193 45404
rect 29181 45373 29193 45376
rect 29227 45373 29239 45407
rect 29181 45367 29239 45373
rect 29362 45364 29368 45416
rect 29420 45364 29426 45416
rect 29454 45364 29460 45416
rect 29512 45364 29518 45416
rect 29549 45407 29607 45413
rect 29549 45373 29561 45407
rect 29595 45373 29607 45407
rect 29549 45367 29607 45373
rect 29641 45407 29699 45413
rect 29641 45373 29653 45407
rect 29687 45404 29699 45407
rect 29831 45404 29859 45580
rect 30558 45568 30564 45620
rect 30616 45608 30622 45620
rect 31665 45611 31723 45617
rect 31665 45608 31677 45611
rect 30616 45580 31677 45608
rect 30616 45568 30622 45580
rect 31665 45577 31677 45580
rect 31711 45577 31723 45611
rect 31665 45571 31723 45577
rect 33134 45568 33140 45620
rect 33192 45608 33198 45620
rect 33686 45608 33692 45620
rect 33192 45580 33692 45608
rect 33192 45568 33198 45580
rect 33686 45568 33692 45580
rect 33744 45608 33750 45620
rect 33781 45611 33839 45617
rect 33781 45608 33793 45611
rect 33744 45580 33793 45608
rect 33744 45568 33750 45580
rect 33781 45577 33793 45580
rect 33827 45577 33839 45611
rect 33781 45571 33839 45577
rect 37645 45611 37703 45617
rect 37645 45577 37657 45611
rect 37691 45608 37703 45611
rect 38102 45608 38108 45620
rect 37691 45580 38108 45608
rect 37691 45577 37703 45580
rect 37645 45571 37703 45577
rect 38102 45568 38108 45580
rect 38160 45568 38166 45620
rect 33410 45540 33416 45552
rect 30760 45512 32720 45540
rect 29687 45376 29859 45404
rect 29687 45373 29699 45376
rect 29641 45367 29699 45373
rect 17865 45339 17923 45345
rect 17865 45305 17877 45339
rect 17911 45336 17923 45339
rect 17954 45336 17960 45348
rect 17911 45308 17960 45336
rect 17911 45305 17923 45308
rect 17865 45299 17923 45305
rect 17954 45296 17960 45308
rect 18012 45296 18018 45348
rect 29086 45296 29092 45348
rect 29144 45336 29150 45348
rect 29564 45336 29592 45367
rect 30374 45364 30380 45416
rect 30432 45364 30438 45416
rect 30558 45364 30564 45416
rect 30616 45404 30622 45416
rect 30653 45407 30711 45413
rect 30653 45404 30665 45407
rect 30616 45376 30665 45404
rect 30616 45364 30622 45376
rect 30653 45373 30665 45376
rect 30699 45373 30711 45407
rect 30653 45367 30711 45373
rect 29144 45308 29592 45336
rect 29144 45296 29150 45308
rect 29730 45296 29736 45348
rect 29788 45336 29794 45348
rect 30760 45336 30788 45512
rect 31110 45432 31116 45484
rect 31168 45472 31174 45484
rect 31297 45475 31355 45481
rect 31297 45472 31309 45475
rect 31168 45444 31309 45472
rect 31168 45432 31174 45444
rect 31297 45441 31309 45444
rect 31343 45441 31355 45475
rect 31297 45435 31355 45441
rect 31757 45475 31815 45481
rect 31757 45441 31769 45475
rect 31803 45472 31815 45475
rect 32582 45472 32588 45484
rect 31803 45444 32588 45472
rect 31803 45441 31815 45444
rect 31757 45435 31815 45441
rect 32582 45432 32588 45444
rect 32640 45432 32646 45484
rect 32692 45404 32720 45512
rect 32784 45512 33416 45540
rect 32784 45481 32812 45512
rect 33410 45500 33416 45512
rect 33468 45500 33474 45552
rect 33597 45543 33655 45549
rect 33597 45509 33609 45543
rect 33643 45540 33655 45543
rect 34790 45540 34796 45552
rect 33643 45512 34796 45540
rect 33643 45509 33655 45512
rect 33597 45503 33655 45509
rect 32769 45475 32827 45481
rect 32769 45441 32781 45475
rect 32815 45441 32827 45475
rect 32769 45435 32827 45441
rect 32950 45432 32956 45484
rect 33008 45432 33014 45484
rect 33045 45475 33103 45481
rect 33045 45441 33057 45475
rect 33091 45441 33103 45475
rect 33045 45435 33103 45441
rect 33137 45475 33195 45481
rect 33137 45441 33149 45475
rect 33183 45472 33195 45475
rect 33612 45472 33640 45503
rect 34790 45500 34796 45512
rect 34848 45500 34854 45552
rect 36722 45500 36728 45552
rect 36780 45500 36786 45552
rect 37366 45500 37372 45552
rect 37424 45540 37430 45552
rect 37424 45512 37872 45540
rect 37424 45500 37430 45512
rect 33183 45444 33640 45472
rect 33689 45475 33747 45481
rect 33183 45441 33195 45444
rect 33137 45435 33195 45441
rect 33689 45441 33701 45475
rect 33735 45441 33747 45475
rect 33689 45435 33747 45441
rect 33060 45404 33088 45435
rect 33704 45404 33732 45435
rect 37844 45413 37872 45512
rect 46750 45432 46756 45484
rect 46808 45432 46814 45484
rect 32692 45376 33732 45404
rect 37737 45407 37795 45413
rect 37737 45373 37749 45407
rect 37783 45373 37795 45407
rect 37737 45367 37795 45373
rect 37829 45407 37887 45413
rect 37829 45373 37841 45407
rect 37875 45373 37887 45407
rect 37829 45367 37887 45373
rect 29788 45308 30788 45336
rect 29788 45296 29794 45308
rect 37274 45296 37280 45348
rect 37332 45296 37338 45348
rect 37752 45336 37780 45367
rect 46569 45339 46627 45345
rect 46569 45336 46581 45339
rect 37752 45308 46581 45336
rect 46569 45305 46581 45308
rect 46615 45305 46627 45339
rect 46569 45299 46627 45305
rect 15562 45228 15568 45280
rect 15620 45268 15626 45280
rect 16669 45271 16727 45277
rect 16669 45268 16681 45271
rect 15620 45240 16681 45268
rect 15620 45228 15626 45240
rect 16669 45237 16681 45240
rect 16715 45237 16727 45271
rect 16669 45231 16727 45237
rect 20073 45271 20131 45277
rect 20073 45237 20085 45271
rect 20119 45268 20131 45271
rect 21358 45268 21364 45280
rect 20119 45240 21364 45268
rect 20119 45237 20131 45240
rect 20073 45231 20131 45237
rect 21358 45228 21364 45240
rect 21416 45228 21422 45280
rect 28258 45228 28264 45280
rect 28316 45268 28322 45280
rect 29178 45268 29184 45280
rect 28316 45240 29184 45268
rect 28316 45228 28322 45240
rect 29178 45228 29184 45240
rect 29236 45228 29242 45280
rect 29454 45228 29460 45280
rect 29512 45268 29518 45280
rect 30558 45268 30564 45280
rect 29512 45240 30564 45268
rect 29512 45228 29518 45240
rect 30558 45228 30564 45240
rect 30616 45228 30622 45280
rect 31018 45228 31024 45280
rect 31076 45268 31082 45280
rect 31435 45271 31493 45277
rect 31435 45268 31447 45271
rect 31076 45240 31447 45268
rect 31076 45228 31082 45240
rect 31435 45237 31447 45240
rect 31481 45237 31493 45271
rect 31435 45231 31493 45237
rect 31570 45228 31576 45280
rect 31628 45228 31634 45280
rect 32306 45228 32312 45280
rect 32364 45268 32370 45280
rect 33321 45271 33379 45277
rect 33321 45268 33333 45271
rect 32364 45240 33333 45268
rect 32364 45228 32370 45240
rect 33321 45237 33333 45240
rect 33367 45237 33379 45271
rect 33321 45231 33379 45237
rect 33962 45228 33968 45280
rect 34020 45228 34026 45280
rect 37001 45271 37059 45277
rect 37001 45237 37013 45271
rect 37047 45268 37059 45271
rect 38102 45268 38108 45280
rect 37047 45240 38108 45268
rect 37047 45237 37059 45240
rect 37001 45231 37059 45237
rect 38102 45228 38108 45240
rect 38160 45228 38166 45280
rect 1104 45178 47104 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 47104 45178
rect 1104 45104 47104 45126
rect 17126 45024 17132 45076
rect 17184 45064 17190 45076
rect 20622 45064 20628 45076
rect 17184 45036 20628 45064
rect 17184 45024 17190 45036
rect 16393 44999 16451 45005
rect 16393 44965 16405 44999
rect 16439 44996 16451 44999
rect 16850 44996 16856 45008
rect 16439 44968 16856 44996
rect 16439 44965 16451 44968
rect 16393 44959 16451 44965
rect 16850 44956 16856 44968
rect 16908 44956 16914 45008
rect 17236 44996 17264 45036
rect 20622 45024 20628 45036
rect 20680 45024 20686 45076
rect 20809 45067 20867 45073
rect 20809 45033 20821 45067
rect 20855 45064 20867 45067
rect 21174 45064 21180 45076
rect 20855 45036 21180 45064
rect 20855 45033 20867 45036
rect 20809 45027 20867 45033
rect 21174 45024 21180 45036
rect 21232 45024 21238 45076
rect 22738 45024 22744 45076
rect 22796 45064 22802 45076
rect 23293 45067 23351 45073
rect 23293 45064 23305 45067
rect 22796 45036 23305 45064
rect 22796 45024 22802 45036
rect 23293 45033 23305 45036
rect 23339 45033 23351 45067
rect 23293 45027 23351 45033
rect 25501 45067 25559 45073
rect 25501 45033 25513 45067
rect 25547 45064 25559 45067
rect 25774 45064 25780 45076
rect 25547 45036 25780 45064
rect 25547 45033 25559 45036
rect 25501 45027 25559 45033
rect 25774 45024 25780 45036
rect 25832 45064 25838 45076
rect 27706 45064 27712 45076
rect 25832 45036 27712 45064
rect 25832 45024 25838 45036
rect 27706 45024 27712 45036
rect 27764 45024 27770 45076
rect 27982 45024 27988 45076
rect 28040 45064 28046 45076
rect 28040 45036 28856 45064
rect 28040 45024 28046 45036
rect 20714 44996 20720 45008
rect 16960 44968 17264 44996
rect 20272 44968 20720 44996
rect 16574 44888 16580 44940
rect 16632 44928 16638 44940
rect 16960 44937 16988 44968
rect 16945 44931 17003 44937
rect 16945 44928 16957 44931
rect 16632 44900 16957 44928
rect 16632 44888 16638 44900
rect 16945 44897 16957 44900
rect 16991 44897 17003 44931
rect 16945 44891 17003 44897
rect 17129 44931 17187 44937
rect 17129 44897 17141 44931
rect 17175 44928 17187 44931
rect 17310 44928 17316 44940
rect 17175 44900 17316 44928
rect 17175 44897 17187 44900
rect 17129 44891 17187 44897
rect 17310 44888 17316 44900
rect 17368 44888 17374 44940
rect 20272 44928 20300 44968
rect 20714 44956 20720 44968
rect 20772 44956 20778 45008
rect 20898 44956 20904 45008
rect 20956 44956 20962 45008
rect 21266 44956 21272 45008
rect 21324 44996 21330 45008
rect 25685 44999 25743 45005
rect 21324 44968 22048 44996
rect 21324 44956 21330 44968
rect 22020 44937 22048 44968
rect 25685 44965 25697 44999
rect 25731 44965 25743 44999
rect 25685 44959 25743 44965
rect 22005 44931 22063 44937
rect 20180 44900 20300 44928
rect 20548 44900 21404 44928
rect 13722 44820 13728 44872
rect 13780 44860 13786 44872
rect 15013 44863 15071 44869
rect 15013 44860 15025 44863
rect 13780 44832 15025 44860
rect 13780 44820 13786 44832
rect 15013 44829 15025 44832
rect 15059 44860 15071 44863
rect 15654 44860 15660 44872
rect 15059 44832 15660 44860
rect 15059 44829 15071 44832
rect 15013 44823 15071 44829
rect 15654 44820 15660 44832
rect 15712 44820 15718 44872
rect 16850 44820 16856 44872
rect 16908 44820 16914 44872
rect 20180 44869 20208 44900
rect 20165 44863 20223 44869
rect 20165 44829 20177 44863
rect 20211 44829 20223 44863
rect 20165 44823 20223 44829
rect 20258 44863 20316 44869
rect 20258 44829 20270 44863
rect 20304 44829 20316 44863
rect 20258 44823 20316 44829
rect 20395 44863 20453 44869
rect 20395 44829 20407 44863
rect 20441 44860 20453 44863
rect 20548 44860 20576 44900
rect 21376 44872 21404 44900
rect 22005 44897 22017 44931
rect 22051 44897 22063 44931
rect 22005 44891 22063 44897
rect 22097 44931 22155 44937
rect 22097 44897 22109 44931
rect 22143 44928 22155 44931
rect 22646 44928 22652 44940
rect 22143 44900 22652 44928
rect 22143 44897 22155 44900
rect 22097 44891 22155 44897
rect 22646 44888 22652 44900
rect 22704 44888 22710 44940
rect 23198 44928 23204 44940
rect 22940 44900 23204 44928
rect 20441 44832 20576 44860
rect 20441 44829 20453 44832
rect 20395 44823 20453 44829
rect 15280 44795 15338 44801
rect 15280 44761 15292 44795
rect 15326 44792 15338 44795
rect 15378 44792 15384 44804
rect 15326 44764 15384 44792
rect 15326 44761 15338 44764
rect 15280 44755 15338 44761
rect 15378 44752 15384 44764
rect 15436 44752 15442 44804
rect 16482 44684 16488 44736
rect 16540 44684 16546 44736
rect 20272 44724 20300 44823
rect 20622 44820 20628 44872
rect 20680 44869 20686 44872
rect 20680 44823 20688 44869
rect 20680 44820 20686 44823
rect 21174 44820 21180 44872
rect 21232 44820 21238 44872
rect 21269 44863 21327 44869
rect 21269 44829 21281 44863
rect 21315 44829 21327 44863
rect 21269 44823 21327 44829
rect 20530 44752 20536 44804
rect 20588 44752 20594 44804
rect 21082 44752 21088 44804
rect 21140 44792 21146 44804
rect 21284 44792 21312 44823
rect 21358 44820 21364 44872
rect 21416 44820 21422 44872
rect 21542 44820 21548 44872
rect 21600 44820 21606 44872
rect 22186 44820 22192 44872
rect 22244 44820 22250 44872
rect 22278 44820 22284 44872
rect 22336 44820 22342 44872
rect 22554 44820 22560 44872
rect 22612 44860 22618 44872
rect 22940 44869 22968 44900
rect 23198 44888 23204 44900
rect 23256 44888 23262 44940
rect 23290 44888 23296 44940
rect 23348 44928 23354 44940
rect 25700 44928 25728 44959
rect 28626 44956 28632 45008
rect 28684 44956 28690 45008
rect 23348 44900 25728 44928
rect 23348 44888 23354 44900
rect 26694 44888 26700 44940
rect 26752 44888 26758 44940
rect 26881 44931 26939 44937
rect 26881 44897 26893 44931
rect 26927 44928 26939 44931
rect 28442 44928 28448 44940
rect 26927 44900 28448 44928
rect 26927 44897 26939 44900
rect 26881 44891 26939 44897
rect 28442 44888 28448 44900
rect 28500 44888 28506 44940
rect 28828 44928 28856 45036
rect 28902 45024 28908 45076
rect 28960 45064 28966 45076
rect 29362 45064 29368 45076
rect 28960 45036 29368 45064
rect 28960 45024 28966 45036
rect 29362 45024 29368 45036
rect 29420 45064 29426 45076
rect 30466 45064 30472 45076
rect 29420 45036 30472 45064
rect 29420 45024 29426 45036
rect 30466 45024 30472 45036
rect 30524 45064 30530 45076
rect 30837 45067 30895 45073
rect 30837 45064 30849 45067
rect 30524 45036 30849 45064
rect 30524 45024 30530 45036
rect 30837 45033 30849 45036
rect 30883 45033 30895 45067
rect 30837 45027 30895 45033
rect 31018 45024 31024 45076
rect 31076 45024 31082 45076
rect 31110 45024 31116 45076
rect 31168 45024 31174 45076
rect 32493 45067 32551 45073
rect 32493 45033 32505 45067
rect 32539 45033 32551 45067
rect 32493 45027 32551 45033
rect 28994 44956 29000 45008
rect 29052 44996 29058 45008
rect 29822 44996 29828 45008
rect 29052 44968 29828 44996
rect 29052 44956 29058 44968
rect 29822 44956 29828 44968
rect 29880 44956 29886 45008
rect 30377 44999 30435 45005
rect 30377 44965 30389 44999
rect 30423 44996 30435 44999
rect 31570 44996 31576 45008
rect 30423 44968 31576 44996
rect 30423 44965 30435 44968
rect 30377 44959 30435 44965
rect 31570 44956 31576 44968
rect 31628 44956 31634 45008
rect 32508 44996 32536 45027
rect 32582 45024 32588 45076
rect 32640 45064 32646 45076
rect 32953 45067 33011 45073
rect 32953 45064 32965 45067
rect 32640 45036 32965 45064
rect 32640 45024 32646 45036
rect 32953 45033 32965 45036
rect 32999 45033 33011 45067
rect 32953 45027 33011 45033
rect 34790 44996 34796 45008
rect 31726 44968 34796 44996
rect 31726 44928 31754 44968
rect 34790 44956 34796 44968
rect 34848 44956 34854 45008
rect 28828 44900 31754 44928
rect 32674 44888 32680 44940
rect 32732 44928 32738 44940
rect 33962 44928 33968 44940
rect 32732 44900 33968 44928
rect 32732 44888 32738 44900
rect 33962 44888 33968 44900
rect 34020 44888 34026 44940
rect 22925 44863 22983 44869
rect 22925 44860 22937 44863
rect 22612 44832 22937 44860
rect 22612 44820 22618 44832
rect 22925 44829 22937 44832
rect 22971 44829 22983 44863
rect 22925 44823 22983 44829
rect 23106 44820 23112 44872
rect 23164 44820 23170 44872
rect 25590 44860 25596 44872
rect 25548 44835 25596 44860
rect 25547 44829 25596 44835
rect 21140 44764 21312 44792
rect 21140 44752 21146 44764
rect 25314 44752 25320 44804
rect 25372 44752 25378 44804
rect 25547 44795 25559 44829
rect 25593 44820 25596 44829
rect 25648 44820 25654 44872
rect 25774 44820 25780 44872
rect 25832 44820 25838 44872
rect 26602 44820 26608 44872
rect 26660 44820 26666 44872
rect 26786 44820 26792 44872
rect 26844 44820 26850 44872
rect 27617 44863 27675 44869
rect 27617 44829 27629 44863
rect 27663 44829 27675 44863
rect 27617 44823 27675 44829
rect 25593 44795 25605 44820
rect 25547 44789 25605 44795
rect 26418 44752 26424 44804
rect 26476 44752 26482 44804
rect 27632 44792 27660 44823
rect 27798 44820 27804 44872
rect 27856 44860 27862 44872
rect 28169 44863 28227 44869
rect 28169 44860 28181 44863
rect 27856 44832 28181 44860
rect 27856 44820 27862 44832
rect 28169 44829 28181 44832
rect 28215 44860 28227 44863
rect 28537 44863 28595 44869
rect 28215 44832 28488 44860
rect 28215 44829 28227 44832
rect 28169 44823 28227 44829
rect 27982 44792 27988 44804
rect 27632 44764 27988 44792
rect 27982 44752 27988 44764
rect 28040 44752 28046 44804
rect 28258 44752 28264 44804
rect 28316 44792 28322 44804
rect 28353 44795 28411 44801
rect 28353 44792 28365 44795
rect 28316 44764 28365 44792
rect 28316 44752 28322 44764
rect 28353 44761 28365 44764
rect 28399 44761 28411 44795
rect 28460 44792 28488 44832
rect 28537 44829 28549 44863
rect 28583 44857 28595 44863
rect 28626 44857 28632 44872
rect 28583 44829 28632 44857
rect 28537 44823 28595 44829
rect 28626 44820 28632 44829
rect 28684 44820 28690 44872
rect 28810 44820 28816 44872
rect 28868 44860 28874 44872
rect 28905 44863 28963 44869
rect 28905 44860 28917 44863
rect 28868 44832 28917 44860
rect 28868 44820 28874 44832
rect 28905 44829 28917 44832
rect 28951 44829 28963 44863
rect 28905 44823 28963 44829
rect 29178 44820 29184 44872
rect 29236 44820 29242 44872
rect 29362 44820 29368 44872
rect 29420 44860 29426 44872
rect 30377 44863 30435 44869
rect 29420 44832 30052 44860
rect 29420 44820 29426 44832
rect 29454 44792 29460 44804
rect 28460 44764 29460 44792
rect 28353 44755 28411 44761
rect 29454 44752 29460 44764
rect 29512 44752 29518 44804
rect 20346 44724 20352 44736
rect 20272 44696 20352 44724
rect 20346 44684 20352 44696
rect 20404 44684 20410 44736
rect 21818 44684 21824 44736
rect 21876 44684 21882 44736
rect 25682 44684 25688 44736
rect 25740 44724 25746 44736
rect 25961 44727 26019 44733
rect 25961 44724 25973 44727
rect 25740 44696 25973 44724
rect 25740 44684 25746 44696
rect 25961 44693 25973 44696
rect 26007 44693 26019 44727
rect 25961 44687 26019 44693
rect 27706 44684 27712 44736
rect 27764 44684 27770 44736
rect 28626 44684 28632 44736
rect 28684 44684 28690 44736
rect 28721 44727 28779 44733
rect 28721 44693 28733 44727
rect 28767 44724 28779 44727
rect 29086 44724 29092 44736
rect 28767 44696 29092 44724
rect 28767 44693 28779 44696
rect 28721 44687 28779 44693
rect 29086 44684 29092 44696
rect 29144 44684 29150 44736
rect 29270 44684 29276 44736
rect 29328 44724 29334 44736
rect 29914 44724 29920 44736
rect 29328 44696 29920 44724
rect 29328 44684 29334 44696
rect 29914 44684 29920 44696
rect 29972 44684 29978 44736
rect 30024 44724 30052 44832
rect 30377 44829 30389 44863
rect 30423 44860 30435 44863
rect 30466 44860 30472 44872
rect 30423 44832 30472 44860
rect 30423 44829 30435 44832
rect 30377 44823 30435 44829
rect 30466 44820 30472 44832
rect 30524 44820 30530 44872
rect 30558 44820 30564 44872
rect 30616 44820 30622 44872
rect 31294 44820 31300 44872
rect 31352 44820 31358 44872
rect 31573 44863 31631 44869
rect 31573 44829 31585 44863
rect 31619 44860 31631 44863
rect 31662 44860 31668 44872
rect 31619 44832 31668 44860
rect 31619 44829 31631 44832
rect 31573 44823 31631 44829
rect 31662 44820 31668 44832
rect 31720 44820 31726 44872
rect 31757 44863 31815 44869
rect 31757 44829 31769 44863
rect 31803 44860 31815 44863
rect 31803 44832 31837 44860
rect 31803 44829 31815 44832
rect 31757 44823 31815 44829
rect 30098 44752 30104 44804
rect 30156 44792 30162 44804
rect 30576 44792 30604 44820
rect 30653 44795 30711 44801
rect 30653 44792 30665 44795
rect 30156 44764 30665 44792
rect 30156 44752 30162 44764
rect 30653 44761 30665 44764
rect 30699 44761 30711 44795
rect 31772 44792 31800 44823
rect 32306 44820 32312 44872
rect 32364 44820 32370 44872
rect 32769 44863 32827 44869
rect 32769 44829 32781 44863
rect 32815 44860 32827 44863
rect 32950 44860 32956 44872
rect 32815 44832 32956 44860
rect 32815 44829 32827 44832
rect 32769 44823 32827 44829
rect 32950 44820 32956 44832
rect 33008 44820 33014 44872
rect 38838 44820 38844 44872
rect 38896 44820 38902 44872
rect 33318 44792 33324 44804
rect 30653 44755 30711 44761
rect 30760 44764 33324 44792
rect 30760 44724 30788 44764
rect 33318 44752 33324 44764
rect 33376 44752 33382 44804
rect 30024 44696 30788 44724
rect 30863 44727 30921 44733
rect 30863 44693 30875 44727
rect 30909 44724 30921 44727
rect 31294 44724 31300 44736
rect 30909 44696 31300 44724
rect 30909 44693 30921 44696
rect 30863 44687 30921 44693
rect 31294 44684 31300 44696
rect 31352 44684 31358 44736
rect 38286 44684 38292 44736
rect 38344 44724 38350 44736
rect 39025 44727 39083 44733
rect 39025 44724 39037 44727
rect 38344 44696 39037 44724
rect 38344 44684 38350 44696
rect 39025 44693 39037 44696
rect 39071 44693 39083 44727
rect 39025 44687 39083 44693
rect 1104 44634 47104 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 35594 44634
rect 35646 44582 35658 44634
rect 35710 44582 35722 44634
rect 35774 44582 35786 44634
rect 35838 44582 35850 44634
rect 35902 44582 47104 44634
rect 1104 44560 47104 44582
rect 15378 44480 15384 44532
rect 15436 44480 15442 44532
rect 16853 44523 16911 44529
rect 16853 44489 16865 44523
rect 16899 44489 16911 44523
rect 16853 44483 16911 44489
rect 20073 44523 20131 44529
rect 20073 44489 20085 44523
rect 20119 44520 20131 44523
rect 20346 44520 20352 44532
rect 20119 44492 20352 44520
rect 20119 44489 20131 44492
rect 20073 44483 20131 44489
rect 2682 44412 2688 44464
rect 2740 44452 2746 44464
rect 16868 44452 16896 44483
rect 20346 44480 20352 44492
rect 20404 44520 20410 44532
rect 21542 44520 21548 44532
rect 20404 44492 21548 44520
rect 20404 44480 20410 44492
rect 21542 44480 21548 44492
rect 21600 44480 21606 44532
rect 22278 44480 22284 44532
rect 22336 44520 22342 44532
rect 27709 44523 27767 44529
rect 27709 44520 27721 44523
rect 22336 44492 27721 44520
rect 22336 44480 22342 44492
rect 27709 44489 27721 44492
rect 27755 44489 27767 44523
rect 27709 44483 27767 44489
rect 28629 44523 28687 44529
rect 28629 44489 28641 44523
rect 28675 44520 28687 44523
rect 29270 44520 29276 44532
rect 28675 44492 29276 44520
rect 28675 44489 28687 44492
rect 28629 44483 28687 44489
rect 29270 44480 29276 44492
rect 29328 44480 29334 44532
rect 29454 44480 29460 44532
rect 29512 44520 29518 44532
rect 31754 44520 31760 44532
rect 29512 44492 31760 44520
rect 29512 44480 29518 44492
rect 31754 44480 31760 44492
rect 31812 44520 31818 44532
rect 32950 44520 32956 44532
rect 31812 44492 32956 44520
rect 31812 44480 31818 44492
rect 32950 44480 32956 44492
rect 33008 44480 33014 44532
rect 33226 44480 33232 44532
rect 33284 44520 33290 44532
rect 33321 44523 33379 44529
rect 33321 44520 33333 44523
rect 33284 44492 33333 44520
rect 33284 44480 33290 44492
rect 33321 44489 33333 44492
rect 33367 44520 33379 44523
rect 34238 44520 34244 44532
rect 33367 44492 34244 44520
rect 33367 44489 33379 44492
rect 33321 44483 33379 44489
rect 34238 44480 34244 44492
rect 34296 44480 34302 44532
rect 36357 44523 36415 44529
rect 36357 44489 36369 44523
rect 36403 44520 36415 44523
rect 36446 44520 36452 44532
rect 36403 44492 36452 44520
rect 36403 44489 36415 44492
rect 36357 44483 36415 44489
rect 36446 44480 36452 44492
rect 36504 44480 36510 44532
rect 37366 44480 37372 44532
rect 37424 44520 37430 44532
rect 37461 44523 37519 44529
rect 37461 44520 37473 44523
rect 37424 44492 37473 44520
rect 37424 44480 37430 44492
rect 37461 44489 37473 44492
rect 37507 44489 37519 44523
rect 37461 44483 37519 44489
rect 38378 44480 38384 44532
rect 38436 44480 38442 44532
rect 17650 44455 17708 44461
rect 17650 44452 17662 44455
rect 2740 44424 12434 44452
rect 16868 44424 17662 44452
rect 2740 44412 2746 44424
rect 1394 44344 1400 44396
rect 1452 44344 1458 44396
rect 12406 44316 12434 44424
rect 17650 44421 17662 44424
rect 17696 44421 17708 44455
rect 21818 44452 21824 44464
rect 17650 44415 17708 44421
rect 20640 44424 21824 44452
rect 15562 44344 15568 44396
rect 15620 44344 15626 44396
rect 16482 44344 16488 44396
rect 16540 44384 16546 44396
rect 17037 44387 17095 44393
rect 17037 44384 17049 44387
rect 16540 44356 17049 44384
rect 16540 44344 16546 44356
rect 17037 44353 17049 44356
rect 17083 44353 17095 44387
rect 17037 44347 17095 44353
rect 17328 44356 19656 44384
rect 17328 44316 17356 44356
rect 12406 44288 17356 44316
rect 17405 44319 17463 44325
rect 17405 44285 17417 44319
rect 17451 44285 17463 44319
rect 19628 44316 19656 44356
rect 19702 44344 19708 44396
rect 19760 44344 19766 44396
rect 19889 44387 19947 44393
rect 19889 44353 19901 44387
rect 19935 44384 19947 44387
rect 20162 44384 20168 44396
rect 19935 44356 20168 44384
rect 19935 44353 19947 44356
rect 19889 44347 19947 44353
rect 19904 44316 19932 44347
rect 20162 44344 20168 44356
rect 20220 44344 20226 44396
rect 20640 44393 20668 44424
rect 21818 44412 21824 44424
rect 21876 44412 21882 44464
rect 22738 44412 22744 44464
rect 22796 44452 22802 44464
rect 22925 44455 22983 44461
rect 22925 44452 22937 44455
rect 22796 44424 22937 44452
rect 22796 44412 22802 44424
rect 22925 44421 22937 44424
rect 22971 44421 22983 44455
rect 22925 44415 22983 44421
rect 23014 44412 23020 44464
rect 23072 44412 23078 44464
rect 23217 44455 23275 44461
rect 23217 44452 23229 44455
rect 23124 44424 23229 44452
rect 20625 44387 20683 44393
rect 20625 44353 20637 44387
rect 20671 44353 20683 44387
rect 20625 44347 20683 44353
rect 20714 44344 20720 44396
rect 20772 44384 20778 44396
rect 20809 44387 20867 44393
rect 20809 44384 20821 44387
rect 20772 44356 20821 44384
rect 20772 44344 20778 44356
rect 20809 44353 20821 44356
rect 20855 44384 20867 44387
rect 21082 44384 21088 44396
rect 20855 44356 21088 44384
rect 20855 44353 20867 44356
rect 20809 44347 20867 44353
rect 21082 44344 21088 44356
rect 21140 44344 21146 44396
rect 22186 44344 22192 44396
rect 22244 44384 22250 44396
rect 22281 44387 22339 44393
rect 22281 44384 22293 44387
rect 22244 44356 22293 44384
rect 22244 44344 22250 44356
rect 22281 44353 22293 44356
rect 22327 44353 22339 44387
rect 22281 44347 22339 44353
rect 22649 44387 22707 44393
rect 22649 44353 22661 44387
rect 22695 44384 22707 44387
rect 22830 44384 22836 44396
rect 22695 44356 22836 44384
rect 22695 44353 22707 44356
rect 22649 44347 22707 44353
rect 22830 44344 22836 44356
rect 22888 44344 22894 44396
rect 19628 44288 19932 44316
rect 20180 44316 20208 44344
rect 20180 44288 22324 44316
rect 17405 44279 17463 44285
rect 934 44208 940 44260
rect 992 44248 998 44260
rect 1581 44251 1639 44257
rect 1581 44248 1593 44251
rect 992 44220 1593 44248
rect 992 44208 998 44220
rect 1581 44217 1593 44220
rect 1627 44217 1639 44251
rect 1581 44211 1639 44217
rect 17034 44140 17040 44192
rect 17092 44180 17098 44192
rect 17420 44180 17448 44279
rect 22296 44260 22324 44288
rect 22094 44208 22100 44260
rect 22152 44208 22158 44260
rect 22278 44208 22284 44260
rect 22336 44208 22342 44260
rect 22646 44208 22652 44260
rect 22704 44248 22710 44260
rect 23124 44248 23152 44424
rect 23217 44421 23229 44424
rect 23263 44421 23275 44455
rect 23217 44415 23275 44421
rect 25314 44412 25320 44464
rect 25372 44452 25378 44464
rect 29362 44452 29368 44464
rect 25372 44424 29368 44452
rect 25372 44412 25378 44424
rect 25406 44344 25412 44396
rect 25464 44344 25470 44396
rect 25593 44387 25651 44393
rect 25593 44353 25605 44387
rect 25639 44353 25651 44387
rect 25593 44347 25651 44353
rect 25608 44316 25636 44347
rect 25682 44344 25688 44396
rect 25740 44384 25746 44396
rect 25777 44387 25835 44393
rect 25777 44384 25789 44387
rect 25740 44356 25789 44384
rect 25740 44344 25746 44356
rect 25777 44353 25789 44356
rect 25823 44353 25835 44387
rect 25777 44347 25835 44353
rect 26418 44344 26424 44396
rect 26476 44384 26482 44396
rect 26970 44384 26976 44396
rect 26476 44356 26976 44384
rect 26476 44344 26482 44356
rect 26970 44344 26976 44356
rect 27028 44384 27034 44396
rect 27172 44393 27200 44424
rect 29362 44412 29368 44424
rect 29420 44412 29426 44464
rect 29733 44455 29791 44461
rect 29472 44424 29684 44452
rect 27065 44387 27123 44393
rect 27065 44384 27077 44387
rect 27028 44356 27077 44384
rect 27028 44344 27034 44356
rect 27065 44353 27077 44356
rect 27111 44353 27123 44387
rect 27065 44347 27123 44353
rect 27157 44387 27215 44393
rect 27157 44353 27169 44387
rect 27203 44353 27215 44387
rect 27157 44347 27215 44353
rect 27525 44387 27583 44393
rect 27525 44353 27537 44387
rect 27571 44384 27583 44387
rect 27798 44384 27804 44396
rect 27571 44356 27804 44384
rect 27571 44353 27583 44356
rect 27525 44347 27583 44353
rect 27798 44344 27804 44356
rect 27856 44344 27862 44396
rect 28537 44387 28595 44393
rect 28537 44353 28549 44387
rect 28583 44384 28595 44387
rect 28994 44384 29000 44396
rect 28583 44356 29000 44384
rect 28583 44353 28595 44356
rect 28537 44347 28595 44353
rect 28994 44344 29000 44356
rect 29052 44344 29058 44396
rect 29086 44344 29092 44396
rect 29144 44384 29150 44396
rect 29472 44384 29500 44424
rect 29144 44356 29500 44384
rect 29549 44387 29607 44393
rect 29144 44344 29150 44356
rect 29549 44353 29561 44387
rect 29595 44353 29607 44387
rect 29656 44384 29684 44424
rect 29733 44421 29745 44455
rect 29779 44452 29791 44455
rect 30098 44452 30104 44464
rect 29779 44424 30104 44452
rect 29779 44421 29791 44424
rect 29733 44415 29791 44421
rect 30098 44412 30104 44424
rect 30156 44412 30162 44464
rect 35244 44455 35302 44461
rect 35244 44421 35256 44455
rect 35290 44452 35302 44455
rect 35342 44452 35348 44464
rect 35290 44424 35348 44452
rect 35290 44421 35302 44424
rect 35244 44415 35302 44421
rect 35342 44412 35348 44424
rect 35400 44412 35406 44464
rect 35434 44412 35440 44464
rect 35492 44452 35498 44464
rect 38838 44452 38844 44464
rect 35492 44424 38844 44452
rect 35492 44412 35498 44424
rect 38838 44412 38844 44424
rect 38896 44412 38902 44464
rect 29825 44387 29883 44393
rect 29825 44384 29837 44387
rect 29656 44356 29837 44384
rect 29549 44347 29607 44353
rect 29825 44353 29837 44356
rect 29871 44384 29883 44387
rect 30282 44384 30288 44396
rect 29871 44356 30288 44384
rect 29871 44353 29883 44356
rect 29825 44347 29883 44353
rect 25961 44319 26019 44325
rect 25961 44316 25973 44319
rect 25608 44288 25973 44316
rect 25961 44285 25973 44288
rect 26007 44316 26019 44319
rect 26510 44316 26516 44328
rect 26007 44288 26516 44316
rect 26007 44285 26019 44288
rect 25961 44279 26019 44285
rect 26510 44276 26516 44288
rect 26568 44316 26574 44328
rect 28813 44319 28871 44325
rect 28813 44316 28825 44319
rect 26568 44288 28825 44316
rect 26568 44276 26574 44288
rect 28813 44285 28825 44288
rect 28859 44316 28871 44319
rect 28902 44316 28908 44328
rect 28859 44288 28908 44316
rect 28859 44285 28871 44288
rect 28813 44279 28871 44285
rect 28902 44276 28908 44288
rect 28960 44276 28966 44328
rect 29564 44316 29592 44347
rect 30282 44344 30288 44356
rect 30340 44344 30346 44396
rect 33229 44387 33287 44393
rect 33229 44353 33241 44387
rect 33275 44384 33287 44387
rect 33318 44384 33324 44396
rect 33275 44356 33324 44384
rect 33275 44353 33287 44356
rect 33229 44347 33287 44353
rect 33318 44344 33324 44356
rect 33376 44344 33382 44396
rect 33505 44387 33563 44393
rect 33505 44353 33517 44387
rect 33551 44384 33563 44387
rect 34790 44384 34796 44396
rect 33551 44356 34796 44384
rect 33551 44353 33563 44356
rect 33505 44347 33563 44353
rect 34790 44344 34796 44356
rect 34848 44344 34854 44396
rect 34977 44387 35035 44393
rect 34977 44353 34989 44387
rect 35023 44384 35035 44387
rect 35452 44384 35480 44412
rect 35023 44356 35480 44384
rect 35023 44353 35035 44356
rect 34977 44347 35035 44353
rect 37274 44344 37280 44396
rect 37332 44344 37338 44396
rect 38286 44344 38292 44396
rect 38344 44344 38350 44396
rect 38470 44344 38476 44396
rect 38528 44384 38534 44396
rect 38657 44387 38715 44393
rect 38657 44384 38669 44387
rect 38528 44356 38669 44384
rect 38528 44344 38534 44356
rect 38657 44353 38669 44356
rect 38703 44384 38715 44387
rect 39761 44387 39819 44393
rect 39761 44384 39773 44387
rect 38703 44356 39773 44384
rect 38703 44353 38715 44356
rect 38657 44347 38715 44353
rect 39761 44353 39773 44356
rect 39807 44353 39819 44387
rect 39761 44347 39819 44353
rect 29730 44316 29736 44328
rect 29564 44288 29736 44316
rect 22704 44220 23152 44248
rect 25501 44251 25559 44257
rect 22704 44208 22710 44220
rect 25501 44217 25513 44251
rect 25547 44248 25559 44251
rect 26418 44248 26424 44260
rect 25547 44220 26424 44248
rect 25547 44217 25559 44220
rect 25501 44211 25559 44217
rect 26418 44208 26424 44220
rect 26476 44208 26482 44260
rect 28169 44251 28227 44257
rect 28169 44248 28181 44251
rect 26528 44220 28181 44248
rect 17770 44180 17776 44192
rect 17092 44152 17776 44180
rect 17092 44140 17098 44152
rect 17770 44140 17776 44152
rect 17828 44140 17834 44192
rect 18785 44183 18843 44189
rect 18785 44149 18797 44183
rect 18831 44180 18843 44183
rect 19978 44180 19984 44192
rect 18831 44152 19984 44180
rect 18831 44149 18843 44152
rect 18785 44143 18843 44149
rect 19978 44140 19984 44152
rect 20036 44140 20042 44192
rect 20530 44140 20536 44192
rect 20588 44180 20594 44192
rect 20625 44183 20683 44189
rect 20625 44180 20637 44183
rect 20588 44152 20637 44180
rect 20588 44140 20594 44152
rect 20625 44149 20637 44152
rect 20671 44149 20683 44183
rect 20625 44143 20683 44149
rect 23201 44183 23259 44189
rect 23201 44149 23213 44183
rect 23247 44180 23259 44183
rect 23290 44180 23296 44192
rect 23247 44152 23296 44180
rect 23247 44149 23259 44152
rect 23201 44143 23259 44149
rect 23290 44140 23296 44152
rect 23348 44140 23354 44192
rect 23382 44140 23388 44192
rect 23440 44140 23446 44192
rect 25958 44140 25964 44192
rect 26016 44180 26022 44192
rect 26528 44180 26556 44220
rect 28169 44217 28181 44220
rect 28215 44217 28227 44251
rect 28169 44211 28227 44217
rect 28718 44208 28724 44260
rect 28776 44248 28782 44260
rect 29656 44248 29684 44288
rect 29730 44276 29736 44288
rect 29788 44276 29794 44328
rect 29914 44276 29920 44328
rect 29972 44316 29978 44328
rect 31294 44316 31300 44328
rect 29972 44288 31300 44316
rect 29972 44276 29978 44288
rect 31294 44276 31300 44288
rect 31352 44316 31358 44328
rect 33781 44319 33839 44325
rect 31352 44288 31754 44316
rect 31352 44276 31358 44288
rect 28776 44220 29684 44248
rect 31726 44248 31754 44288
rect 33781 44285 33793 44319
rect 33827 44316 33839 44319
rect 34514 44316 34520 44328
rect 33827 44288 34520 44316
rect 33827 44285 33839 44288
rect 33781 44279 33839 44285
rect 33796 44248 33824 44279
rect 34514 44276 34520 44288
rect 34572 44276 34578 44328
rect 31726 44220 33824 44248
rect 28776 44208 28782 44220
rect 26016 44152 26556 44180
rect 27525 44183 27583 44189
rect 26016 44140 26022 44152
rect 27525 44149 27537 44183
rect 27571 44180 27583 44183
rect 27982 44180 27988 44192
rect 27571 44152 27988 44180
rect 27571 44149 27583 44152
rect 27525 44143 27583 44149
rect 27982 44140 27988 44152
rect 28040 44140 28046 44192
rect 28074 44140 28080 44192
rect 28132 44180 28138 44192
rect 29086 44180 29092 44192
rect 28132 44152 29092 44180
rect 28132 44140 28138 44152
rect 29086 44140 29092 44152
rect 29144 44140 29150 44192
rect 29822 44140 29828 44192
rect 29880 44140 29886 44192
rect 32398 44140 32404 44192
rect 32456 44180 32462 44192
rect 38304 44180 38332 44344
rect 38378 44276 38384 44328
rect 38436 44316 38442 44328
rect 39022 44316 39028 44328
rect 38436 44288 39028 44316
rect 38436 44276 38442 44288
rect 39022 44276 39028 44288
rect 39080 44316 39086 44328
rect 39485 44319 39543 44325
rect 39485 44316 39497 44319
rect 39080 44288 39497 44316
rect 39080 44276 39086 44288
rect 39485 44285 39497 44288
rect 39531 44285 39543 44319
rect 39485 44279 39543 44285
rect 32456 44152 38332 44180
rect 32456 44140 32462 44152
rect 1104 44090 47104 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 47104 44090
rect 1104 44016 47104 44038
rect 4614 43936 4620 43988
rect 4672 43976 4678 43988
rect 19702 43976 19708 43988
rect 4672 43948 6914 43976
rect 4672 43936 4678 43948
rect 6886 43908 6914 43948
rect 16224 43948 19708 43976
rect 15930 43908 15936 43920
rect 6886 43880 15936 43908
rect 15930 43868 15936 43880
rect 15988 43868 15994 43920
rect 16224 43840 16252 43948
rect 19702 43936 19708 43948
rect 19760 43936 19766 43988
rect 20165 43979 20223 43985
rect 20165 43945 20177 43979
rect 20211 43976 20223 43979
rect 21266 43976 21272 43988
rect 20211 43948 21272 43976
rect 20211 43945 20223 43948
rect 20165 43939 20223 43945
rect 21266 43936 21272 43948
rect 21324 43936 21330 43988
rect 22557 43979 22615 43985
rect 22557 43945 22569 43979
rect 22603 43976 22615 43979
rect 23014 43976 23020 43988
rect 22603 43948 23020 43976
rect 22603 43945 22615 43948
rect 22557 43939 22615 43945
rect 23014 43936 23020 43948
rect 23072 43936 23078 43988
rect 23106 43936 23112 43988
rect 23164 43976 23170 43988
rect 24213 43979 24271 43985
rect 24213 43976 24225 43979
rect 23164 43948 24225 43976
rect 23164 43936 23170 43948
rect 24213 43945 24225 43948
rect 24259 43945 24271 43979
rect 24213 43939 24271 43945
rect 17954 43868 17960 43920
rect 18012 43908 18018 43920
rect 19150 43908 19156 43920
rect 18012 43880 19156 43908
rect 18012 43868 18018 43880
rect 19150 43868 19156 43880
rect 19208 43908 19214 43920
rect 19208 43880 20300 43908
rect 19208 43868 19214 43880
rect 20272 43849 20300 43880
rect 21358 43868 21364 43920
rect 21416 43908 21422 43920
rect 22646 43908 22652 43920
rect 21416 43880 22652 43908
rect 21416 43868 21422 43880
rect 22646 43868 22652 43880
rect 22704 43868 22710 43920
rect 22830 43868 22836 43920
rect 22888 43868 22894 43920
rect 20257 43843 20315 43849
rect 6886 43812 16252 43840
rect 16684 43812 17080 43840
rect 6886 43772 6914 43812
rect 3896 43744 6914 43772
rect 15105 43775 15163 43781
rect 3234 43664 3240 43716
rect 3292 43704 3298 43716
rect 3896 43713 3924 43744
rect 15105 43741 15117 43775
rect 15151 43772 15163 43775
rect 15470 43772 15476 43784
rect 15151 43744 15476 43772
rect 15151 43741 15163 43744
rect 15105 43735 15163 43741
rect 15470 43732 15476 43744
rect 15528 43772 15534 43784
rect 16684 43772 16712 43812
rect 15528 43744 16712 43772
rect 15528 43732 15534 43744
rect 16758 43732 16764 43784
rect 16816 43772 16822 43784
rect 16853 43775 16911 43781
rect 16853 43772 16865 43775
rect 16816 43744 16865 43772
rect 16816 43732 16822 43744
rect 16853 43741 16865 43744
rect 16899 43741 16911 43775
rect 16853 43735 16911 43741
rect 16942 43732 16948 43784
rect 17000 43732 17006 43784
rect 17052 43772 17080 43812
rect 18892 43812 19564 43840
rect 18892 43781 18920 43812
rect 18877 43775 18935 43781
rect 18877 43772 18889 43775
rect 17052 43744 18889 43772
rect 18877 43741 18889 43744
rect 18923 43741 18935 43775
rect 18877 43735 18935 43741
rect 19058 43732 19064 43784
rect 19116 43772 19122 43784
rect 19536 43781 19564 43812
rect 20257 43809 20269 43843
rect 20303 43809 20315 43843
rect 22848 43840 22876 43868
rect 20257 43803 20315 43809
rect 21928 43812 22876 43840
rect 24228 43840 24256 43939
rect 25774 43936 25780 43988
rect 25832 43976 25838 43988
rect 26145 43979 26203 43985
rect 26145 43976 26157 43979
rect 25832 43948 26157 43976
rect 25832 43936 25838 43948
rect 26145 43945 26157 43948
rect 26191 43976 26203 43979
rect 26191 43948 30696 43976
rect 26191 43945 26203 43948
rect 26145 43939 26203 43945
rect 24302 43868 24308 43920
rect 24360 43908 24366 43920
rect 30190 43908 30196 43920
rect 24360 43880 24808 43908
rect 24360 43868 24366 43880
rect 24780 43849 24808 43880
rect 26344 43880 30196 43908
rect 24765 43843 24823 43849
rect 24228 43812 24348 43840
rect 20530 43781 20536 43784
rect 19337 43775 19395 43781
rect 19337 43772 19349 43775
rect 19116 43744 19349 43772
rect 19116 43732 19122 43744
rect 19337 43741 19349 43744
rect 19383 43741 19395 43775
rect 19337 43735 19395 43741
rect 19521 43775 19579 43781
rect 19521 43741 19533 43775
rect 19567 43741 19579 43775
rect 19521 43735 19579 43741
rect 19705 43775 19763 43781
rect 19705 43741 19717 43775
rect 19751 43772 19763 43775
rect 20524 43772 20536 43781
rect 19751 43744 20024 43772
rect 20491 43744 20536 43772
rect 19751 43741 19763 43744
rect 19705 43735 19763 43741
rect 3881 43707 3939 43713
rect 3881 43704 3893 43707
rect 3292 43676 3893 43704
rect 3292 43664 3298 43676
rect 3881 43673 3893 43676
rect 3927 43673 3939 43707
rect 3881 43667 3939 43673
rect 4249 43707 4307 43713
rect 4249 43673 4261 43707
rect 4295 43704 4307 43707
rect 4614 43704 4620 43716
rect 4295 43676 4620 43704
rect 4295 43673 4307 43676
rect 4249 43667 4307 43673
rect 4614 43664 4620 43676
rect 4672 43664 4678 43716
rect 19996 43713 20024 43744
rect 20524 43735 20536 43744
rect 20530 43732 20536 43735
rect 20588 43732 20594 43784
rect 21928 43781 21956 43812
rect 21913 43775 21971 43781
rect 21913 43741 21925 43775
rect 21959 43741 21971 43775
rect 21913 43735 21971 43741
rect 22006 43775 22064 43781
rect 22006 43741 22018 43775
rect 22052 43772 22064 43775
rect 22094 43772 22100 43784
rect 22052 43744 22100 43772
rect 22052 43741 22064 43744
rect 22006 43735 22064 43741
rect 22094 43732 22100 43744
rect 22152 43732 22158 43784
rect 22186 43732 22192 43784
rect 22244 43732 22250 43784
rect 22419 43775 22477 43781
rect 22419 43741 22431 43775
rect 22465 43772 22477 43775
rect 22465 43744 22692 43772
rect 22465 43741 22477 43744
rect 22419 43735 22477 43741
rect 17190 43707 17248 43713
rect 17190 43704 17202 43707
rect 16684 43676 17202 43704
rect 15289 43639 15347 43645
rect 15289 43605 15301 43639
rect 15335 43636 15347 43639
rect 16022 43636 16028 43648
rect 15335 43608 16028 43636
rect 15335 43605 15347 43608
rect 15289 43599 15347 43605
rect 16022 43596 16028 43608
rect 16080 43636 16086 43648
rect 16574 43636 16580 43648
rect 16080 43608 16580 43636
rect 16080 43596 16086 43608
rect 16574 43596 16580 43608
rect 16632 43596 16638 43648
rect 16684 43645 16712 43676
rect 17190 43673 17202 43676
rect 17236 43673 17248 43707
rect 17190 43667 17248 43673
rect 18969 43707 19027 43713
rect 18969 43673 18981 43707
rect 19015 43704 19027 43707
rect 19797 43707 19855 43713
rect 19797 43704 19809 43707
rect 19015 43676 19809 43704
rect 19015 43673 19027 43676
rect 18969 43667 19027 43673
rect 19797 43673 19809 43676
rect 19843 43673 19855 43707
rect 19797 43667 19855 43673
rect 19981 43707 20039 43713
rect 19981 43673 19993 43707
rect 20027 43704 20039 43707
rect 21174 43704 21180 43716
rect 20027 43676 21180 43704
rect 20027 43673 20039 43676
rect 19981 43667 20039 43673
rect 21174 43664 21180 43676
rect 21232 43664 21238 43716
rect 21726 43664 21732 43716
rect 21784 43704 21790 43716
rect 22204 43704 22232 43732
rect 21784 43676 22232 43704
rect 22281 43707 22339 43713
rect 21784 43664 21790 43676
rect 22281 43673 22293 43707
rect 22327 43704 22339 43707
rect 22554 43704 22560 43716
rect 22327 43676 22560 43704
rect 22327 43673 22339 43676
rect 22281 43667 22339 43673
rect 16669 43639 16727 43645
rect 16669 43605 16681 43639
rect 16715 43605 16727 43639
rect 16669 43599 16727 43605
rect 18322 43596 18328 43648
rect 18380 43596 18386 43648
rect 19058 43596 19064 43648
rect 19116 43636 19122 43648
rect 20622 43636 20628 43648
rect 19116 43608 20628 43636
rect 19116 43596 19122 43608
rect 20622 43596 20628 43608
rect 20680 43636 20686 43648
rect 21637 43639 21695 43645
rect 21637 43636 21649 43639
rect 20680 43608 21649 43636
rect 20680 43596 20686 43608
rect 21637 43605 21649 43608
rect 21683 43636 21695 43639
rect 21818 43636 21824 43648
rect 21683 43608 21824 43636
rect 21683 43605 21695 43608
rect 21637 43599 21695 43605
rect 21818 43596 21824 43608
rect 21876 43596 21882 43648
rect 22186 43596 22192 43648
rect 22244 43636 22250 43648
rect 22296 43636 22324 43667
rect 22554 43664 22560 43676
rect 22612 43664 22618 43716
rect 22664 43648 22692 43744
rect 22738 43732 22744 43784
rect 22796 43772 22802 43784
rect 22833 43775 22891 43781
rect 22833 43772 22845 43775
rect 22796 43744 22845 43772
rect 22796 43732 22802 43744
rect 22833 43741 22845 43744
rect 22879 43772 22891 43775
rect 23474 43772 23480 43784
rect 22879 43744 23480 43772
rect 22879 43741 22891 43744
rect 22833 43735 22891 43741
rect 23474 43732 23480 43744
rect 23532 43772 23538 43784
rect 24210 43772 24216 43784
rect 23532 43744 24216 43772
rect 23532 43732 23538 43744
rect 24210 43732 24216 43744
rect 24268 43732 24274 43784
rect 24320 43774 24348 43812
rect 24765 43809 24777 43843
rect 24811 43809 24823 43843
rect 24765 43803 24823 43809
rect 24403 43775 24461 43781
rect 24403 43774 24415 43775
rect 24320 43746 24415 43774
rect 24403 43741 24415 43746
rect 24449 43741 24461 43775
rect 26344 43772 26372 43880
rect 30190 43868 30196 43880
rect 30248 43868 30254 43920
rect 27982 43840 27988 43852
rect 26528 43812 27988 43840
rect 24403 43735 24461 43741
rect 24964 43744 26372 43772
rect 23100 43707 23158 43713
rect 23100 43673 23112 43707
rect 23146 43704 23158 43707
rect 24964 43704 24992 43744
rect 26418 43732 26424 43784
rect 26476 43732 26482 43784
rect 23146 43676 24992 43704
rect 25032 43707 25090 43713
rect 23146 43673 23158 43676
rect 23100 43667 23158 43673
rect 25032 43673 25044 43707
rect 25078 43704 25090 43707
rect 25498 43704 25504 43716
rect 25078 43676 25504 43704
rect 25078 43673 25090 43676
rect 25032 43667 25090 43673
rect 25498 43664 25504 43676
rect 25556 43664 25562 43716
rect 26234 43664 26240 43716
rect 26292 43664 26298 43716
rect 26528 43704 26556 43812
rect 27982 43800 27988 43812
rect 28040 43800 28046 43852
rect 28166 43800 28172 43852
rect 28224 43800 28230 43852
rect 28258 43800 28264 43852
rect 28316 43800 28322 43852
rect 28813 43843 28871 43849
rect 28813 43840 28825 43843
rect 28552 43812 28825 43840
rect 26970 43732 26976 43784
rect 27028 43732 27034 43784
rect 27154 43732 27160 43784
rect 27212 43732 27218 43784
rect 28074 43732 28080 43784
rect 28132 43732 28138 43784
rect 28350 43732 28356 43784
rect 28408 43732 28414 43784
rect 28552 43781 28580 43812
rect 28813 43809 28825 43812
rect 28859 43809 28871 43843
rect 28813 43803 28871 43809
rect 29273 43843 29331 43849
rect 29273 43809 29285 43843
rect 29319 43840 29331 43843
rect 29549 43843 29607 43849
rect 29549 43840 29561 43843
rect 29319 43812 29561 43840
rect 29319 43809 29331 43812
rect 29273 43803 29331 43809
rect 29549 43809 29561 43812
rect 29595 43809 29607 43843
rect 29549 43803 29607 43809
rect 29822 43800 29828 43852
rect 29880 43800 29886 43852
rect 29914 43800 29920 43852
rect 29972 43800 29978 43852
rect 30006 43800 30012 43852
rect 30064 43800 30070 43852
rect 28537 43775 28595 43781
rect 28537 43741 28549 43775
rect 28583 43741 28595 43775
rect 28537 43735 28595 43741
rect 28626 43732 28632 43784
rect 28684 43772 28690 43784
rect 28997 43775 29055 43781
rect 28997 43772 29009 43775
rect 28684 43744 29009 43772
rect 28684 43732 28690 43744
rect 28997 43741 29009 43744
rect 29043 43741 29055 43775
rect 28997 43735 29055 43741
rect 29086 43732 29092 43784
rect 29144 43732 29150 43784
rect 29178 43732 29184 43784
rect 29236 43732 29242 43784
rect 29733 43775 29791 43781
rect 29733 43741 29745 43775
rect 29779 43772 29791 43775
rect 30193 43775 30251 43781
rect 30193 43772 30205 43775
rect 29779 43744 30205 43772
rect 29779 43741 29791 43744
rect 29733 43735 29791 43741
rect 30193 43741 30205 43744
rect 30239 43741 30251 43775
rect 30193 43735 30251 43741
rect 30377 43775 30435 43781
rect 30377 43741 30389 43775
rect 30423 43772 30435 43775
rect 30466 43772 30472 43784
rect 30423 43744 30472 43772
rect 30423 43741 30435 43744
rect 30377 43735 30435 43741
rect 30466 43732 30472 43744
rect 30524 43732 30530 43784
rect 30668 43781 30696 43948
rect 33318 43936 33324 43988
rect 33376 43976 33382 43988
rect 33781 43979 33839 43985
rect 33781 43976 33793 43979
rect 33376 43948 33793 43976
rect 33376 43936 33382 43948
rect 33781 43945 33793 43948
rect 33827 43945 33839 43979
rect 33781 43939 33839 43945
rect 35069 43979 35127 43985
rect 35069 43945 35081 43979
rect 35115 43976 35127 43979
rect 35342 43976 35348 43988
rect 35115 43948 35348 43976
rect 35115 43945 35127 43948
rect 35069 43939 35127 43945
rect 35342 43936 35348 43948
rect 35400 43936 35406 43988
rect 36446 43976 36452 43988
rect 35544 43948 36452 43976
rect 34882 43868 34888 43920
rect 34940 43908 34946 43920
rect 35437 43911 35495 43917
rect 35437 43908 35449 43911
rect 34940 43880 35449 43908
rect 34940 43868 34946 43880
rect 35437 43877 35449 43880
rect 35483 43877 35495 43911
rect 35437 43871 35495 43877
rect 35544 43840 35572 43948
rect 36446 43936 36452 43948
rect 36504 43936 36510 43988
rect 37274 43936 37280 43988
rect 37332 43976 37338 43988
rect 37461 43979 37519 43985
rect 37461 43976 37473 43979
rect 37332 43948 37473 43976
rect 37332 43936 37338 43948
rect 37461 43945 37473 43948
rect 37507 43945 37519 43979
rect 38838 43976 38844 43988
rect 37461 43939 37519 43945
rect 38212 43948 38844 43976
rect 35268 43812 35572 43840
rect 30653 43775 30711 43781
rect 30653 43741 30665 43775
rect 30699 43741 30711 43775
rect 30653 43735 30711 43741
rect 32030 43732 32036 43784
rect 32088 43772 32094 43784
rect 35268 43781 35296 43812
rect 35986 43800 35992 43852
rect 36044 43800 36050 43852
rect 32401 43775 32459 43781
rect 32401 43772 32413 43775
rect 32088 43744 32413 43772
rect 32088 43732 32094 43744
rect 32401 43741 32413 43744
rect 32447 43741 32459 43775
rect 32401 43735 32459 43741
rect 35253 43775 35311 43781
rect 35253 43741 35265 43775
rect 35299 43741 35311 43775
rect 35253 43735 35311 43741
rect 35342 43732 35348 43784
rect 35400 43732 35406 43784
rect 35529 43775 35587 43781
rect 35529 43741 35541 43775
rect 35575 43741 35587 43775
rect 35529 43735 35587 43741
rect 35713 43775 35771 43781
rect 35713 43741 35725 43775
rect 35759 43772 35771 43775
rect 36004 43772 36032 43800
rect 35759 43744 36032 43772
rect 36081 43775 36139 43781
rect 35759 43741 35771 43744
rect 35713 43735 35771 43741
rect 36081 43741 36093 43775
rect 36127 43772 36139 43775
rect 37274 43772 37280 43784
rect 36127 43744 37280 43772
rect 36127 43741 36139 43744
rect 36081 43735 36139 43741
rect 28077 43729 28135 43732
rect 26344 43676 26556 43704
rect 26605 43707 26663 43713
rect 22244 43608 22324 43636
rect 22244 43596 22250 43608
rect 22646 43596 22652 43648
rect 22704 43636 22710 43648
rect 24581 43639 24639 43645
rect 24581 43636 24593 43639
rect 22704 43608 24593 43636
rect 22704 43596 22710 43608
rect 24581 43605 24593 43608
rect 24627 43636 24639 43639
rect 26344 43636 26372 43676
rect 26605 43673 26617 43707
rect 26651 43704 26663 43707
rect 27706 43704 27712 43716
rect 26651 43676 27712 43704
rect 26651 43673 26663 43676
rect 26605 43667 26663 43673
rect 27706 43664 27712 43676
rect 27764 43664 27770 43716
rect 30561 43707 30619 43713
rect 28736 43676 28994 43704
rect 24627 43608 26372 43636
rect 26513 43639 26571 43645
rect 24627 43605 24639 43608
rect 24581 43599 24639 43605
rect 26513 43605 26525 43639
rect 26559 43636 26571 43639
rect 26694 43636 26700 43648
rect 26559 43608 26700 43636
rect 26559 43605 26571 43608
rect 26513 43599 26571 43605
rect 26694 43596 26700 43608
rect 26752 43596 26758 43648
rect 26786 43596 26792 43648
rect 26844 43596 26850 43648
rect 27614 43596 27620 43648
rect 27672 43636 27678 43648
rect 27893 43639 27951 43645
rect 27893 43636 27905 43639
rect 27672 43608 27905 43636
rect 27672 43596 27678 43608
rect 27893 43605 27905 43608
rect 27939 43605 27951 43639
rect 27893 43599 27951 43605
rect 27982 43596 27988 43648
rect 28040 43636 28046 43648
rect 28736 43636 28764 43676
rect 28040 43608 28764 43636
rect 28966 43648 28994 43676
rect 30561 43673 30573 43707
rect 30607 43704 30619 43707
rect 30834 43704 30840 43716
rect 30607 43676 30840 43704
rect 30607 43673 30619 43676
rect 30561 43667 30619 43673
rect 30834 43664 30840 43676
rect 30892 43664 30898 43716
rect 32668 43707 32726 43713
rect 32668 43673 32680 43707
rect 32714 43704 32726 43707
rect 33594 43704 33600 43716
rect 32714 43676 33600 43704
rect 32714 43673 32726 43676
rect 32668 43667 32726 43673
rect 33594 43664 33600 43676
rect 33652 43664 33658 43716
rect 34698 43664 34704 43716
rect 34756 43704 34762 43716
rect 35434 43704 35440 43716
rect 34756 43676 35440 43704
rect 34756 43664 34762 43676
rect 35434 43664 35440 43676
rect 35492 43704 35498 43716
rect 35544 43704 35572 43735
rect 37274 43732 37280 43744
rect 37332 43732 37338 43784
rect 37476 43772 37504 43939
rect 38212 43849 38240 43948
rect 38838 43936 38844 43948
rect 38896 43936 38902 43988
rect 38197 43843 38255 43849
rect 38197 43809 38209 43843
rect 38243 43809 38255 43843
rect 40405 43843 40463 43849
rect 40405 43840 40417 43843
rect 38197 43803 38255 43809
rect 39224 43812 40417 43840
rect 37553 43775 37611 43781
rect 37553 43772 37565 43775
rect 37476 43744 37565 43772
rect 37553 43741 37565 43744
rect 37599 43741 37611 43775
rect 39224 43772 39252 43812
rect 40405 43809 40417 43812
rect 40451 43809 40463 43843
rect 40405 43803 40463 43809
rect 37553 43735 37611 43741
rect 38396 43744 39252 43772
rect 40313 43775 40371 43781
rect 35492 43676 35572 43704
rect 35492 43664 35498 43676
rect 35986 43664 35992 43716
rect 36044 43704 36050 43716
rect 36326 43707 36384 43713
rect 36326 43704 36338 43707
rect 36044 43676 36338 43704
rect 36044 43664 36050 43676
rect 36326 43673 36338 43676
rect 36372 43673 36384 43707
rect 36326 43667 36384 43673
rect 37826 43664 37832 43716
rect 37884 43704 37890 43716
rect 38396 43704 38424 43744
rect 40313 43741 40325 43775
rect 40359 43772 40371 43775
rect 46566 43772 46572 43784
rect 40359 43744 46572 43772
rect 40359 43741 40371 43744
rect 40313 43735 40371 43741
rect 46566 43732 46572 43744
rect 46624 43732 46630 43784
rect 37884 43676 38424 43704
rect 38464 43707 38522 43713
rect 37884 43664 37890 43676
rect 38464 43673 38476 43707
rect 38510 43704 38522 43707
rect 38746 43704 38752 43716
rect 38510 43676 38752 43704
rect 38510 43673 38522 43676
rect 38464 43667 38522 43673
rect 38746 43664 38752 43676
rect 38804 43664 38810 43716
rect 40221 43707 40279 43713
rect 40221 43704 40233 43707
rect 39592 43676 40233 43704
rect 28966 43608 29000 43648
rect 28040 43596 28046 43608
rect 28994 43596 29000 43608
rect 29052 43596 29058 43648
rect 29086 43596 29092 43648
rect 29144 43636 29150 43648
rect 30374 43636 30380 43648
rect 29144 43608 30380 43636
rect 29144 43596 29150 43608
rect 30374 43596 30380 43608
rect 30432 43596 30438 43648
rect 30742 43596 30748 43648
rect 30800 43636 30806 43648
rect 38102 43636 38108 43648
rect 30800 43608 38108 43636
rect 30800 43596 30806 43608
rect 38102 43596 38108 43608
rect 38160 43596 38166 43648
rect 39206 43596 39212 43648
rect 39264 43636 39270 43648
rect 39592 43645 39620 43676
rect 40221 43673 40233 43676
rect 40267 43673 40279 43707
rect 40221 43667 40279 43673
rect 39577 43639 39635 43645
rect 39577 43636 39589 43639
rect 39264 43608 39589 43636
rect 39264 43596 39270 43608
rect 39577 43605 39589 43608
rect 39623 43605 39635 43639
rect 39577 43599 39635 43605
rect 39850 43596 39856 43648
rect 39908 43596 39914 43648
rect 1104 43546 47104 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 35594 43546
rect 35646 43494 35658 43546
rect 35710 43494 35722 43546
rect 35774 43494 35786 43546
rect 35838 43494 35850 43546
rect 35902 43494 47104 43546
rect 1104 43472 47104 43494
rect 13449 43435 13507 43441
rect 13449 43401 13461 43435
rect 13495 43401 13507 43435
rect 13449 43395 13507 43401
rect 15105 43435 15163 43441
rect 15105 43401 15117 43435
rect 15151 43432 15163 43435
rect 15194 43432 15200 43444
rect 15151 43404 15200 43432
rect 15151 43401 15163 43404
rect 15105 43395 15163 43401
rect 13464 43364 13492 43395
rect 15194 43392 15200 43404
rect 15252 43392 15258 43444
rect 16301 43435 16359 43441
rect 16301 43401 16313 43435
rect 16347 43401 16359 43435
rect 16301 43395 16359 43401
rect 13970 43367 14028 43373
rect 13970 43364 13982 43367
rect 13464 43336 13982 43364
rect 13970 43333 13982 43336
rect 14016 43333 14028 43367
rect 16316 43364 16344 43395
rect 16758 43392 16764 43444
rect 16816 43432 16822 43444
rect 18141 43435 18199 43441
rect 18141 43432 18153 43435
rect 16816 43404 18153 43432
rect 16816 43392 16822 43404
rect 18141 43401 18153 43404
rect 18187 43401 18199 43435
rect 18141 43395 18199 43401
rect 21269 43435 21327 43441
rect 21269 43401 21281 43435
rect 21315 43432 21327 43435
rect 21637 43435 21695 43441
rect 21637 43432 21649 43435
rect 21315 43404 21649 43432
rect 21315 43401 21327 43404
rect 21269 43395 21327 43401
rect 21637 43401 21649 43404
rect 21683 43432 21695 43435
rect 21726 43432 21732 43444
rect 21683 43404 21732 43432
rect 21683 43401 21695 43404
rect 21637 43395 21695 43401
rect 21726 43392 21732 43404
rect 21784 43392 21790 43444
rect 22094 43432 22100 43444
rect 21836 43404 22100 43432
rect 16914 43367 16972 43373
rect 16914 43364 16926 43367
rect 16316 43336 16926 43364
rect 13970 43327 14028 43333
rect 16914 43333 16926 43336
rect 16960 43333 16972 43367
rect 16914 43327 16972 43333
rect 17034 43324 17040 43376
rect 17092 43324 17098 43376
rect 18601 43367 18659 43373
rect 18601 43333 18613 43367
rect 18647 43364 18659 43367
rect 19702 43364 19708 43376
rect 18647 43336 19708 43364
rect 18647 43333 18659 43336
rect 18601 43327 18659 43333
rect 19702 43324 19708 43336
rect 19760 43324 19766 43376
rect 20162 43324 20168 43376
rect 20220 43364 20226 43376
rect 20533 43367 20591 43373
rect 20533 43364 20545 43367
rect 20220 43336 20545 43364
rect 20220 43324 20226 43336
rect 20533 43333 20545 43336
rect 20579 43333 20591 43367
rect 20533 43327 20591 43333
rect 20717 43367 20775 43373
rect 20717 43333 20729 43367
rect 20763 43364 20775 43367
rect 21836 43364 21864 43404
rect 22094 43392 22100 43404
rect 22152 43392 22158 43444
rect 24121 43435 24179 43441
rect 24121 43401 24133 43435
rect 24167 43401 24179 43435
rect 24121 43395 24179 43401
rect 20763 43336 21864 43364
rect 20763 43333 20775 43336
rect 20717 43327 20775 43333
rect 13633 43299 13691 43305
rect 13633 43265 13645 43299
rect 13679 43296 13691 43299
rect 15102 43296 15108 43308
rect 13679 43268 15108 43296
rect 13679 43265 13691 43268
rect 13633 43259 13691 43265
rect 15102 43256 15108 43268
rect 15160 43256 15166 43308
rect 16485 43299 16543 43305
rect 16485 43265 16497 43299
rect 16531 43296 16543 43299
rect 16574 43296 16580 43308
rect 16531 43268 16580 43296
rect 16531 43265 16543 43268
rect 16485 43259 16543 43265
rect 16574 43256 16580 43268
rect 16632 43256 16638 43308
rect 16669 43299 16727 43305
rect 16669 43265 16681 43299
rect 16715 43296 16727 43299
rect 17052 43296 17080 43324
rect 16715 43268 17080 43296
rect 16715 43265 16727 43268
rect 16669 43259 16727 43265
rect 17310 43256 17316 43308
rect 17368 43296 17374 43308
rect 17368 43268 17724 43296
rect 17368 43256 17374 43268
rect 13722 43188 13728 43240
rect 13780 43188 13786 43240
rect 17696 43228 17724 43268
rect 18322 43256 18328 43308
rect 18380 43296 18386 43308
rect 18509 43299 18567 43305
rect 18509 43296 18521 43299
rect 18380 43268 18521 43296
rect 18380 43256 18386 43268
rect 18509 43265 18521 43268
rect 18555 43296 18567 43299
rect 19610 43296 19616 43308
rect 18555 43268 19616 43296
rect 18555 43265 18567 43268
rect 18509 43259 18567 43265
rect 19610 43256 19616 43268
rect 19668 43256 19674 43308
rect 20346 43256 20352 43308
rect 20404 43256 20410 43308
rect 18693 43231 18751 43237
rect 18693 43228 18705 43231
rect 17696 43200 18705 43228
rect 18693 43197 18705 43200
rect 18739 43197 18751 43231
rect 20548 43228 20576 43327
rect 21910 43324 21916 43376
rect 21968 43364 21974 43376
rect 24136 43364 24164 43395
rect 25498 43392 25504 43444
rect 25556 43392 25562 43444
rect 26234 43392 26240 43444
rect 26292 43432 26298 43444
rect 26421 43435 26479 43441
rect 26421 43432 26433 43435
rect 26292 43404 26433 43432
rect 26292 43392 26298 43404
rect 26421 43401 26433 43404
rect 26467 43401 26479 43435
rect 26421 43395 26479 43401
rect 26602 43392 26608 43444
rect 26660 43432 26666 43444
rect 27433 43435 27491 43441
rect 27433 43432 27445 43435
rect 26660 43404 27445 43432
rect 26660 43392 26666 43404
rect 27433 43401 27445 43404
rect 27479 43401 27491 43435
rect 30282 43432 30288 43444
rect 27433 43395 27491 43401
rect 29472 43404 30288 43432
rect 26786 43364 26792 43376
rect 21968 43336 24164 43364
rect 25884 43336 26792 43364
rect 21968 43324 21974 43336
rect 21085 43299 21143 43305
rect 21085 43265 21097 43299
rect 21131 43296 21143 43299
rect 21266 43296 21272 43308
rect 21131 43268 21272 43296
rect 21131 43265 21143 43268
rect 21085 43259 21143 43265
rect 21266 43256 21272 43268
rect 21324 43256 21330 43308
rect 21358 43256 21364 43308
rect 21416 43256 21422 43308
rect 21450 43256 21456 43308
rect 21508 43256 21514 43308
rect 21637 43299 21695 43305
rect 21637 43265 21649 43299
rect 21683 43265 21695 43299
rect 21637 43259 21695 43265
rect 21821 43299 21879 43305
rect 21821 43265 21833 43299
rect 21867 43296 21879 43299
rect 22097 43299 22155 43305
rect 21867 43268 22048 43296
rect 21867 43265 21879 43268
rect 21821 43259 21879 43265
rect 21652 43228 21680 43259
rect 21910 43228 21916 43240
rect 20548 43200 21916 43228
rect 18693 43191 18751 43197
rect 21910 43188 21916 43200
rect 21968 43188 21974 43240
rect 22020 43228 22048 43268
rect 22097 43265 22109 43299
rect 22143 43296 22155 43299
rect 22278 43296 22284 43308
rect 22143 43268 22284 43296
rect 22143 43265 22155 43268
rect 22097 43259 22155 43265
rect 22278 43256 22284 43268
rect 22336 43256 22342 43308
rect 22554 43256 22560 43308
rect 22612 43296 22618 43308
rect 22997 43299 23055 43305
rect 22997 43296 23009 43299
rect 22612 43268 23009 43296
rect 22612 43256 22618 43268
rect 22997 43265 23009 43268
rect 23043 43265 23055 43299
rect 22997 43259 23055 43265
rect 25590 43256 25596 43308
rect 25648 43296 25654 43308
rect 25884 43305 25912 43336
rect 26786 43324 26792 43336
rect 26844 43324 26850 43376
rect 26878 43324 26884 43376
rect 26936 43364 26942 43376
rect 26973 43367 27031 43373
rect 26973 43364 26985 43367
rect 26936 43336 26985 43364
rect 26936 43324 26942 43336
rect 26973 43333 26985 43336
rect 27019 43333 27031 43367
rect 28166 43364 28172 43376
rect 26973 43327 27031 43333
rect 27080 43336 28172 43364
rect 25685 43299 25743 43305
rect 25685 43296 25697 43299
rect 25648 43268 25697 43296
rect 25648 43256 25654 43268
rect 25685 43265 25697 43268
rect 25731 43265 25743 43299
rect 25685 43259 25743 43265
rect 25869 43299 25927 43305
rect 25869 43265 25881 43299
rect 25915 43265 25927 43299
rect 25869 43259 25927 43265
rect 25958 43256 25964 43308
rect 26016 43256 26022 43308
rect 26050 43256 26056 43308
rect 26108 43256 26114 43308
rect 26237 43299 26295 43305
rect 26237 43265 26249 43299
rect 26283 43296 26295 43299
rect 26510 43296 26516 43308
rect 26283 43268 26516 43296
rect 26283 43265 26295 43268
rect 26237 43259 26295 43265
rect 26510 43256 26516 43268
rect 26568 43256 26574 43308
rect 26694 43256 26700 43308
rect 26752 43296 26758 43308
rect 27080 43296 27108 43336
rect 28166 43324 28172 43336
rect 28224 43324 28230 43376
rect 26752 43268 27108 43296
rect 26752 43256 26758 43268
rect 27246 43256 27252 43308
rect 27304 43256 27310 43308
rect 29365 43299 29423 43305
rect 29365 43265 29377 43299
rect 29411 43296 29423 43299
rect 29472 43296 29500 43404
rect 30282 43392 30288 43404
rect 30340 43392 30346 43444
rect 30374 43392 30380 43444
rect 30432 43392 30438 43444
rect 30650 43392 30656 43444
rect 30708 43392 30714 43444
rect 34790 43392 34796 43444
rect 34848 43392 34854 43444
rect 34882 43392 34888 43444
rect 34940 43432 34946 43444
rect 35713 43435 35771 43441
rect 34940 43404 35664 43432
rect 34940 43392 34946 43404
rect 29546 43324 29552 43376
rect 29604 43364 29610 43376
rect 29641 43367 29699 43373
rect 29641 43364 29653 43367
rect 29604 43336 29653 43364
rect 29604 43324 29610 43336
rect 29641 43333 29653 43336
rect 29687 43333 29699 43367
rect 29641 43327 29699 43333
rect 30469 43367 30527 43373
rect 30469 43333 30481 43367
rect 30515 43364 30527 43367
rect 30834 43364 30840 43376
rect 30515 43336 30840 43364
rect 30515 43333 30527 43336
rect 30469 43327 30527 43333
rect 30834 43324 30840 43336
rect 30892 43324 30898 43376
rect 33680 43367 33738 43373
rect 33680 43333 33692 43367
rect 33726 43364 33738 43367
rect 35636 43364 35664 43404
rect 35713 43401 35725 43435
rect 35759 43432 35771 43435
rect 35986 43432 35992 43444
rect 35759 43404 35992 43432
rect 35759 43401 35771 43404
rect 35713 43395 35771 43401
rect 35986 43392 35992 43404
rect 36044 43392 36050 43444
rect 36078 43392 36084 43444
rect 36136 43432 36142 43444
rect 37366 43432 37372 43444
rect 36136 43404 37372 43432
rect 36136 43392 36142 43404
rect 37366 43392 37372 43404
rect 37424 43392 37430 43444
rect 37642 43392 37648 43444
rect 37700 43432 37706 43444
rect 38562 43432 38568 43444
rect 37700 43404 38568 43432
rect 37700 43392 37706 43404
rect 38562 43392 38568 43404
rect 38620 43392 38626 43444
rect 38746 43392 38752 43444
rect 38804 43392 38810 43444
rect 40402 43392 40408 43444
rect 40460 43392 40466 43444
rect 39850 43364 39856 43376
rect 33726 43336 35204 43364
rect 35636 43336 36124 43364
rect 33726 43333 33738 43336
rect 33680 43327 33738 43333
rect 29411 43268 29500 43296
rect 29411 43265 29423 43268
rect 29365 43259 29423 43265
rect 29730 43256 29736 43308
rect 29788 43256 29794 43308
rect 29826 43299 29884 43305
rect 29826 43265 29838 43299
rect 29872 43265 29884 43299
rect 29826 43259 29884 43265
rect 22186 43228 22192 43240
rect 22020 43200 22192 43228
rect 22186 43188 22192 43200
rect 22244 43188 22250 43240
rect 22296 43228 22324 43256
rect 22649 43231 22707 43237
rect 22649 43228 22661 43231
rect 22296 43200 22661 43228
rect 22649 43197 22661 43200
rect 22695 43197 22707 43231
rect 22649 43191 22707 43197
rect 22738 43188 22744 43240
rect 22796 43188 22802 43240
rect 27065 43231 27123 43237
rect 27065 43228 27077 43231
rect 24688 43200 27077 43228
rect 21082 43120 21088 43172
rect 21140 43120 21146 43172
rect 22281 43163 22339 43169
rect 22281 43129 22293 43163
rect 22327 43129 22339 43163
rect 22281 43123 22339 43129
rect 18046 43052 18052 43104
rect 18104 43052 18110 43104
rect 21818 43052 21824 43104
rect 21876 43052 21882 43104
rect 22296 43092 22324 43123
rect 24688 43092 24716 43200
rect 27065 43197 27077 43200
rect 27111 43197 27123 43231
rect 27065 43191 27123 43197
rect 29546 43188 29552 43240
rect 29604 43228 29610 43240
rect 29641 43231 29699 43237
rect 29641 43228 29653 43231
rect 29604 43200 29653 43228
rect 29604 43188 29610 43200
rect 29641 43197 29653 43200
rect 29687 43228 29699 43231
rect 29840 43228 29868 43259
rect 29914 43256 29920 43308
rect 29972 43296 29978 43308
rect 30009 43299 30067 43305
rect 30009 43296 30021 43299
rect 29972 43268 30021 43296
rect 29972 43256 29978 43268
rect 30009 43265 30021 43268
rect 30055 43265 30067 43299
rect 30009 43259 30067 43265
rect 30098 43256 30104 43308
rect 30156 43256 30162 43308
rect 30239 43299 30297 43305
rect 30239 43265 30251 43299
rect 30285 43296 30297 43299
rect 30285 43268 30420 43296
rect 30285 43265 30297 43268
rect 30239 43259 30297 43265
rect 30392 43228 30420 43268
rect 30742 43256 30748 43308
rect 30800 43256 30806 43308
rect 32030 43256 32036 43308
rect 32088 43296 32094 43308
rect 33410 43296 33416 43308
rect 32088 43268 33416 43296
rect 32088 43256 32094 43268
rect 33410 43256 33416 43268
rect 33468 43256 33474 43308
rect 34698 43256 34704 43308
rect 34756 43296 34762 43308
rect 34885 43299 34943 43305
rect 34885 43296 34897 43299
rect 34756 43268 34897 43296
rect 34756 43256 34762 43268
rect 34885 43265 34897 43268
rect 34931 43265 34943 43299
rect 34885 43259 34943 43265
rect 35066 43256 35072 43308
rect 35124 43256 35130 43308
rect 35176 43296 35204 43336
rect 35176 43268 35388 43296
rect 30760 43228 30788 43256
rect 29687 43200 29868 43228
rect 30116 43200 30788 43228
rect 29687 43197 29699 43200
rect 29641 43191 29699 43197
rect 29457 43163 29515 43169
rect 29457 43129 29469 43163
rect 29503 43160 29515 43163
rect 30006 43160 30012 43172
rect 29503 43132 30012 43160
rect 29503 43129 29515 43132
rect 29457 43123 29515 43129
rect 30006 43120 30012 43132
rect 30064 43120 30070 43172
rect 22296 43064 24716 43092
rect 27062 43052 27068 43104
rect 27120 43052 27126 43104
rect 28534 43052 28540 43104
rect 28592 43092 28598 43104
rect 30116 43092 30144 43200
rect 34514 43188 34520 43240
rect 34572 43228 34578 43240
rect 35161 43231 35219 43237
rect 35161 43228 35173 43231
rect 34572 43200 35173 43228
rect 34572 43188 34578 43200
rect 35161 43197 35173 43200
rect 35207 43197 35219 43231
rect 35161 43191 35219 43197
rect 35253 43231 35311 43237
rect 35253 43197 35265 43231
rect 35299 43197 35311 43231
rect 35253 43191 35311 43197
rect 34606 43120 34612 43172
rect 34664 43160 34670 43172
rect 35268 43160 35296 43191
rect 34664 43132 35296 43160
rect 35360 43160 35388 43268
rect 35434 43256 35440 43308
rect 35492 43256 35498 43308
rect 35986 43256 35992 43308
rect 36044 43256 36050 43308
rect 36096 43305 36124 43336
rect 38948 43336 39856 43364
rect 36081 43299 36139 43305
rect 36081 43265 36093 43299
rect 36127 43265 36139 43299
rect 36081 43259 36139 43265
rect 36173 43299 36231 43305
rect 36173 43265 36185 43299
rect 36219 43265 36231 43299
rect 36173 43259 36231 43265
rect 35526 43188 35532 43240
rect 35584 43228 35590 43240
rect 36188 43228 36216 43259
rect 36262 43256 36268 43308
rect 36320 43296 36326 43308
rect 36357 43299 36415 43305
rect 36357 43296 36369 43299
rect 36320 43268 36369 43296
rect 36320 43256 36326 43268
rect 36357 43265 36369 43268
rect 36403 43265 36415 43299
rect 36357 43259 36415 43265
rect 36725 43299 36783 43305
rect 36725 43265 36737 43299
rect 36771 43296 36783 43299
rect 36771 43268 37320 43296
rect 36771 43265 36783 43268
rect 36725 43259 36783 43265
rect 35584 43200 36216 43228
rect 35584 43188 35590 43200
rect 37292 43169 37320 43268
rect 37366 43256 37372 43308
rect 37424 43296 37430 43308
rect 38948 43305 38976 43336
rect 39850 43324 39856 43336
rect 39908 43324 39914 43376
rect 38933 43299 38991 43305
rect 37424 43268 37872 43296
rect 37424 43256 37430 43268
rect 37734 43188 37740 43240
rect 37792 43188 37798 43240
rect 37844 43237 37872 43268
rect 38933 43265 38945 43299
rect 38979 43265 38991 43299
rect 38933 43259 38991 43265
rect 39292 43299 39350 43305
rect 39292 43265 39304 43299
rect 39338 43296 39350 43299
rect 39574 43296 39580 43308
rect 39338 43268 39580 43296
rect 39338 43265 39350 43268
rect 39292 43259 39350 43265
rect 39574 43256 39580 43268
rect 39632 43256 39638 43308
rect 45830 43256 45836 43308
rect 45888 43296 45894 43308
rect 46477 43299 46535 43305
rect 46477 43296 46489 43299
rect 45888 43268 46489 43296
rect 45888 43256 45894 43268
rect 46477 43265 46489 43268
rect 46523 43265 46535 43299
rect 46477 43259 46535 43265
rect 37829 43231 37887 43237
rect 37829 43197 37841 43231
rect 37875 43197 37887 43231
rect 37829 43191 37887 43197
rect 38838 43188 38844 43240
rect 38896 43228 38902 43240
rect 39025 43231 39083 43237
rect 39025 43228 39037 43231
rect 38896 43200 39037 43228
rect 38896 43188 38902 43200
rect 39025 43197 39037 43200
rect 39071 43197 39083 43231
rect 39025 43191 39083 43197
rect 35621 43163 35679 43169
rect 35621 43160 35633 43163
rect 35360 43132 35633 43160
rect 34664 43120 34670 43132
rect 35621 43129 35633 43132
rect 35667 43129 35679 43163
rect 35621 43123 35679 43129
rect 37277 43163 37335 43169
rect 37277 43129 37289 43163
rect 37323 43129 37335 43163
rect 37277 43123 37335 43129
rect 28592 43064 30144 43092
rect 28592 43052 28598 43064
rect 30374 43052 30380 43104
rect 30432 43092 30438 43104
rect 30469 43095 30527 43101
rect 30469 43092 30481 43095
rect 30432 43064 30481 43092
rect 30432 43052 30438 43064
rect 30469 43061 30481 43064
rect 30515 43061 30527 43095
rect 30469 43055 30527 43061
rect 34514 43052 34520 43104
rect 34572 43092 34578 43104
rect 35986 43092 35992 43104
rect 34572 43064 35992 43092
rect 34572 43052 34578 43064
rect 35986 43052 35992 43064
rect 36044 43052 36050 43104
rect 36538 43052 36544 43104
rect 36596 43052 36602 43104
rect 40402 43052 40408 43104
rect 40460 43092 40466 43104
rect 46474 43092 46480 43104
rect 40460 43064 46480 43092
rect 40460 43052 40466 43064
rect 46474 43052 46480 43064
rect 46532 43052 46538 43104
rect 46658 43052 46664 43104
rect 46716 43052 46722 43104
rect 1104 43002 47104 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 47104 43002
rect 1104 42928 47104 42950
rect 15470 42848 15476 42900
rect 15528 42848 15534 42900
rect 16574 42848 16580 42900
rect 16632 42848 16638 42900
rect 17310 42848 17316 42900
rect 17368 42888 17374 42900
rect 17589 42891 17647 42897
rect 17589 42888 17601 42891
rect 17368 42860 17601 42888
rect 17368 42848 17374 42860
rect 17589 42857 17601 42860
rect 17635 42857 17647 42891
rect 17589 42851 17647 42857
rect 22554 42848 22560 42900
rect 22612 42848 22618 42900
rect 29917 42891 29975 42897
rect 29917 42857 29929 42891
rect 29963 42888 29975 42891
rect 30006 42888 30012 42900
rect 29963 42860 30012 42888
rect 29963 42857 29975 42860
rect 29917 42851 29975 42857
rect 30006 42848 30012 42860
rect 30064 42848 30070 42900
rect 35253 42891 35311 42897
rect 35253 42857 35265 42891
rect 35299 42888 35311 42891
rect 35434 42888 35440 42900
rect 35299 42860 35440 42888
rect 35299 42857 35311 42860
rect 35253 42851 35311 42857
rect 35434 42848 35440 42860
rect 35492 42848 35498 42900
rect 39574 42848 39580 42900
rect 39632 42848 39638 42900
rect 13722 42712 13728 42764
rect 13780 42752 13786 42764
rect 14093 42755 14151 42761
rect 14093 42752 14105 42755
rect 13780 42724 14105 42752
rect 13780 42712 13786 42724
rect 14093 42721 14105 42724
rect 14139 42721 14151 42755
rect 14093 42715 14151 42721
rect 15194 42712 15200 42764
rect 15252 42752 15258 42764
rect 16025 42755 16083 42761
rect 16025 42752 16037 42755
rect 15252 42724 16037 42752
rect 15252 42712 15258 42724
rect 16025 42721 16037 42724
rect 16071 42721 16083 42755
rect 16025 42715 16083 42721
rect 16206 42712 16212 42764
rect 16264 42712 16270 42764
rect 17221 42755 17279 42761
rect 17221 42721 17233 42755
rect 17267 42752 17279 42755
rect 17328 42752 17356 42848
rect 22646 42820 22652 42832
rect 19720 42792 22652 42820
rect 19720 42764 19748 42792
rect 22646 42780 22652 42792
rect 22704 42780 22710 42832
rect 29178 42780 29184 42832
rect 29236 42820 29242 42832
rect 30101 42823 30159 42829
rect 30101 42820 30113 42823
rect 29236 42792 30113 42820
rect 29236 42780 29242 42792
rect 30101 42789 30113 42792
rect 30147 42789 30159 42823
rect 30101 42783 30159 42789
rect 30190 42780 30196 42832
rect 30248 42820 30254 42832
rect 36538 42820 36544 42832
rect 30248 42792 36544 42820
rect 30248 42780 30254 42792
rect 36538 42780 36544 42792
rect 36596 42780 36602 42832
rect 17267 42724 17356 42752
rect 17267 42721 17279 42724
rect 17221 42715 17279 42721
rect 19702 42712 19708 42764
rect 19760 42712 19766 42764
rect 19886 42712 19892 42764
rect 19944 42712 19950 42764
rect 26970 42712 26976 42764
rect 27028 42712 27034 42764
rect 29365 42755 29423 42761
rect 29365 42721 29377 42755
rect 29411 42752 29423 42755
rect 30466 42752 30472 42764
rect 29411 42724 30472 42752
rect 29411 42721 29423 42724
rect 29365 42715 29423 42721
rect 16945 42687 17003 42693
rect 16945 42653 16957 42687
rect 16991 42684 17003 42687
rect 18046 42684 18052 42696
rect 16991 42656 18052 42684
rect 16991 42653 17003 42656
rect 16945 42647 17003 42653
rect 18046 42644 18052 42656
rect 18104 42644 18110 42696
rect 19610 42644 19616 42696
rect 19668 42644 19674 42696
rect 22741 42687 22799 42693
rect 22741 42653 22753 42687
rect 22787 42684 22799 42687
rect 23382 42684 23388 42696
rect 22787 42656 23388 42684
rect 22787 42653 22799 42656
rect 22741 42647 22799 42653
rect 23382 42644 23388 42656
rect 23440 42644 23446 42696
rect 27240 42687 27298 42693
rect 27240 42653 27252 42687
rect 27286 42684 27298 42687
rect 27614 42684 27620 42696
rect 27286 42656 27620 42684
rect 27286 42653 27298 42656
rect 27240 42647 27298 42653
rect 27614 42644 27620 42656
rect 27672 42644 27678 42696
rect 29454 42644 29460 42696
rect 29512 42684 29518 42696
rect 29549 42687 29607 42693
rect 29549 42684 29561 42687
rect 29512 42656 29561 42684
rect 29512 42644 29518 42656
rect 29549 42653 29561 42656
rect 29595 42653 29607 42687
rect 29549 42647 29607 42653
rect 29917 42687 29975 42693
rect 29917 42653 29929 42687
rect 29963 42684 29975 42687
rect 30282 42684 30288 42696
rect 29963 42656 30288 42684
rect 29963 42653 29975 42656
rect 29917 42647 29975 42653
rect 30282 42644 30288 42656
rect 30340 42644 30346 42696
rect 30392 42693 30420 42724
rect 30466 42712 30472 42724
rect 30524 42712 30530 42764
rect 30377 42687 30435 42693
rect 30377 42653 30389 42687
rect 30423 42653 30435 42687
rect 30377 42647 30435 42653
rect 31665 42687 31723 42693
rect 31665 42653 31677 42687
rect 31711 42684 31723 42687
rect 32122 42684 32128 42696
rect 31711 42656 32128 42684
rect 31711 42653 31723 42656
rect 31665 42647 31723 42653
rect 32122 42644 32128 42656
rect 32180 42644 32186 42696
rect 32769 42687 32827 42693
rect 32769 42653 32781 42687
rect 32815 42653 32827 42687
rect 32769 42647 32827 42653
rect 13262 42576 13268 42628
rect 13320 42616 13326 42628
rect 14338 42619 14396 42625
rect 14338 42616 14350 42619
rect 13320 42588 14350 42616
rect 13320 42576 13326 42588
rect 14338 42585 14350 42588
rect 14384 42585 14396 42619
rect 14338 42579 14396 42585
rect 15102 42576 15108 42628
rect 15160 42616 15166 42628
rect 17497 42619 17555 42625
rect 15160 42588 15608 42616
rect 15160 42576 15166 42588
rect 15580 42557 15608 42588
rect 17497 42585 17509 42619
rect 17543 42616 17555 42619
rect 17586 42616 17592 42628
rect 17543 42588 17592 42616
rect 17543 42585 17555 42588
rect 17497 42579 17555 42585
rect 17586 42576 17592 42588
rect 17644 42616 17650 42628
rect 20438 42616 20444 42628
rect 17644 42588 20444 42616
rect 17644 42576 17650 42588
rect 20438 42576 20444 42588
rect 20496 42576 20502 42628
rect 25866 42576 25872 42628
rect 25924 42616 25930 42628
rect 28810 42616 28816 42628
rect 25924 42588 28816 42616
rect 25924 42576 25930 42588
rect 28810 42576 28816 42588
rect 28868 42576 28874 42628
rect 29181 42619 29239 42625
rect 29181 42585 29193 42619
rect 29227 42616 29239 42619
rect 29227 42588 29500 42616
rect 29227 42585 29239 42588
rect 29181 42579 29239 42585
rect 15565 42551 15623 42557
rect 15565 42517 15577 42551
rect 15611 42517 15623 42551
rect 15565 42511 15623 42517
rect 15838 42508 15844 42560
rect 15896 42548 15902 42560
rect 15933 42551 15991 42557
rect 15933 42548 15945 42551
rect 15896 42520 15945 42548
rect 15896 42508 15902 42520
rect 15933 42517 15945 42520
rect 15979 42548 15991 42551
rect 17037 42551 17095 42557
rect 17037 42548 17049 42551
rect 15979 42520 17049 42548
rect 15979 42517 15991 42520
rect 15933 42511 15991 42517
rect 17037 42517 17049 42520
rect 17083 42548 17095 42551
rect 19058 42548 19064 42560
rect 17083 42520 19064 42548
rect 17083 42517 17095 42520
rect 17037 42511 17095 42517
rect 19058 42508 19064 42520
rect 19116 42508 19122 42560
rect 19242 42508 19248 42560
rect 19300 42508 19306 42560
rect 19702 42508 19708 42560
rect 19760 42548 19766 42560
rect 28353 42551 28411 42557
rect 28353 42548 28365 42551
rect 19760 42520 28365 42548
rect 19760 42508 19766 42520
rect 28353 42517 28365 42520
rect 28399 42548 28411 42551
rect 29196 42548 29224 42579
rect 28399 42520 29224 42548
rect 29472 42548 29500 42588
rect 30190 42576 30196 42628
rect 30248 42576 30254 42628
rect 32784 42616 32812 42647
rect 32950 42644 32956 42696
rect 33008 42644 33014 42696
rect 33045 42687 33103 42693
rect 33045 42653 33057 42687
rect 33091 42684 33103 42687
rect 35066 42684 35072 42696
rect 33091 42656 35072 42684
rect 33091 42653 33103 42656
rect 33045 42647 33103 42653
rect 35066 42644 35072 42656
rect 35124 42644 35130 42696
rect 35161 42687 35219 42693
rect 35161 42653 35173 42687
rect 35207 42653 35219 42687
rect 35161 42647 35219 42653
rect 34146 42616 34152 42628
rect 32784 42588 34152 42616
rect 34146 42576 34152 42588
rect 34204 42576 34210 42628
rect 35176 42616 35204 42647
rect 37274 42644 37280 42696
rect 37332 42684 37338 42696
rect 37461 42687 37519 42693
rect 37461 42684 37473 42687
rect 37332 42656 37473 42684
rect 37332 42644 37338 42656
rect 37461 42653 37473 42656
rect 37507 42684 37519 42687
rect 38286 42684 38292 42696
rect 37507 42656 38292 42684
rect 37507 42653 37519 42656
rect 37461 42647 37519 42653
rect 38286 42644 38292 42656
rect 38344 42684 38350 42696
rect 38470 42684 38476 42696
rect 38344 42656 38476 42684
rect 38344 42644 38350 42656
rect 38470 42644 38476 42656
rect 38528 42644 38534 42696
rect 35986 42616 35992 42628
rect 35176 42588 35992 42616
rect 35986 42576 35992 42588
rect 36044 42616 36050 42628
rect 37706 42619 37764 42625
rect 37706 42616 37718 42619
rect 36044 42588 37718 42616
rect 36044 42576 36050 42588
rect 37706 42585 37718 42588
rect 37752 42585 37764 42619
rect 37706 42579 37764 42585
rect 29546 42548 29552 42560
rect 29472 42520 29552 42548
rect 28399 42517 28411 42520
rect 28353 42511 28411 42517
rect 29546 42508 29552 42520
rect 29604 42508 29610 42560
rect 29914 42508 29920 42560
rect 29972 42548 29978 42560
rect 30561 42551 30619 42557
rect 30561 42548 30573 42551
rect 29972 42520 30573 42548
rect 29972 42508 29978 42520
rect 30561 42517 30573 42520
rect 30607 42517 30619 42551
rect 30561 42511 30619 42517
rect 30834 42508 30840 42560
rect 30892 42548 30898 42560
rect 31481 42551 31539 42557
rect 31481 42548 31493 42551
rect 30892 42520 31493 42548
rect 30892 42508 30898 42520
rect 31481 42517 31493 42520
rect 31527 42517 31539 42551
rect 31481 42511 31539 42517
rect 32582 42508 32588 42560
rect 32640 42508 32646 42560
rect 38838 42508 38844 42560
rect 38896 42508 38902 42560
rect 1104 42458 47104 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 35594 42458
rect 35646 42406 35658 42458
rect 35710 42406 35722 42458
rect 35774 42406 35786 42458
rect 35838 42406 35850 42458
rect 35902 42406 47104 42458
rect 1104 42384 47104 42406
rect 13262 42304 13268 42356
rect 13320 42304 13326 42356
rect 15838 42304 15844 42356
rect 15896 42304 15902 42356
rect 18046 42304 18052 42356
rect 18104 42344 18110 42356
rect 18969 42347 19027 42353
rect 18969 42344 18981 42347
rect 18104 42316 18981 42344
rect 18104 42304 18110 42316
rect 18969 42313 18981 42316
rect 19015 42313 19027 42347
rect 18969 42307 19027 42313
rect 19058 42304 19064 42356
rect 19116 42344 19122 42356
rect 21450 42344 21456 42356
rect 19116 42316 21456 42344
rect 19116 42304 19122 42316
rect 21450 42304 21456 42316
rect 21508 42304 21514 42356
rect 22021 42316 31616 42344
rect 1394 42236 1400 42288
rect 1452 42276 1458 42288
rect 22021 42276 22049 42316
rect 1452 42248 22049 42276
rect 1452 42236 1458 42248
rect 29454 42236 29460 42288
rect 29512 42236 29518 42288
rect 30006 42236 30012 42288
rect 30064 42236 30070 42288
rect 31588 42276 31616 42316
rect 31662 42304 31668 42356
rect 31720 42344 31726 42356
rect 31941 42347 31999 42353
rect 31941 42344 31953 42347
rect 31720 42316 31953 42344
rect 31720 42304 31726 42316
rect 31941 42313 31953 42316
rect 31987 42313 31999 42347
rect 31941 42307 31999 42313
rect 32950 42304 32956 42356
rect 33008 42344 33014 42356
rect 33505 42347 33563 42353
rect 33505 42344 33517 42347
rect 33008 42316 33517 42344
rect 33008 42304 33014 42316
rect 33505 42313 33517 42316
rect 33551 42313 33563 42347
rect 33505 42307 33563 42313
rect 33594 42304 33600 42356
rect 33652 42304 33658 42356
rect 32392 42279 32450 42285
rect 30576 42248 31524 42276
rect 31588 42248 32352 42276
rect 12710 42168 12716 42220
rect 12768 42208 12774 42220
rect 13449 42211 13507 42217
rect 13449 42208 13461 42211
rect 12768 42180 13461 42208
rect 12768 42168 12774 42180
rect 13449 42177 13461 42180
rect 13495 42177 13507 42211
rect 13449 42171 13507 42177
rect 13538 42168 13544 42220
rect 13596 42208 13602 42220
rect 13981 42211 14039 42217
rect 13981 42208 13993 42211
rect 13596 42180 13993 42208
rect 13596 42168 13602 42180
rect 13981 42177 13993 42180
rect 14027 42177 14039 42211
rect 13981 42171 14039 42177
rect 15657 42211 15715 42217
rect 15657 42177 15669 42211
rect 15703 42208 15715 42211
rect 15703 42180 17080 42208
rect 15703 42177 15715 42180
rect 15657 42171 15715 42177
rect 13722 42100 13728 42152
rect 13780 42100 13786 42152
rect 15105 42075 15163 42081
rect 15105 42041 15117 42075
rect 15151 42072 15163 42075
rect 15672 42072 15700 42171
rect 15151 42044 15700 42072
rect 17052 42072 17080 42180
rect 19242 42168 19248 42220
rect 19300 42208 19306 42220
rect 19613 42211 19671 42217
rect 19613 42208 19625 42211
rect 19300 42180 19625 42208
rect 19300 42168 19306 42180
rect 19613 42177 19625 42180
rect 19659 42177 19671 42211
rect 19613 42171 19671 42177
rect 29365 42211 29423 42217
rect 29365 42177 29377 42211
rect 29411 42208 29423 42211
rect 29411 42180 29500 42208
rect 29411 42177 29423 42180
rect 29365 42171 29423 42177
rect 19153 42143 19211 42149
rect 19153 42109 19165 42143
rect 19199 42140 19211 42143
rect 19886 42140 19892 42152
rect 19199 42112 19892 42140
rect 19199 42109 19211 42112
rect 19153 42103 19211 42109
rect 19886 42100 19892 42112
rect 19944 42100 19950 42152
rect 20346 42072 20352 42084
rect 17052 42044 20352 42072
rect 15151 42041 15163 42044
rect 15105 42035 15163 42041
rect 20346 42032 20352 42044
rect 20404 42032 20410 42084
rect 20438 42032 20444 42084
rect 20496 42072 20502 42084
rect 26878 42072 26884 42084
rect 20496 42044 26884 42072
rect 20496 42032 20502 42044
rect 26878 42032 26884 42044
rect 26936 42032 26942 42084
rect 29472 42072 29500 42180
rect 29546 42168 29552 42220
rect 29604 42168 29610 42220
rect 29914 42168 29920 42220
rect 29972 42168 29978 42220
rect 30576 42217 30604 42248
rect 30834 42217 30840 42220
rect 30101 42211 30159 42217
rect 30101 42177 30113 42211
rect 30147 42177 30159 42211
rect 30101 42171 30159 42177
rect 30561 42211 30619 42217
rect 30561 42177 30573 42211
rect 30607 42177 30619 42211
rect 30828 42208 30840 42217
rect 30795 42180 30840 42208
rect 30561 42171 30619 42177
rect 30828 42171 30840 42180
rect 29564 42140 29592 42168
rect 30116 42140 30144 42171
rect 30834 42168 30840 42171
rect 30892 42168 30898 42220
rect 31496 42208 31524 42248
rect 32324 42208 32352 42248
rect 32392 42245 32404 42279
rect 32438 42276 32450 42279
rect 32582 42276 32588 42288
rect 32438 42248 32588 42276
rect 32438 42245 32450 42248
rect 32392 42239 32450 42245
rect 32582 42236 32588 42248
rect 32640 42236 32646 42288
rect 34238 42236 34244 42288
rect 34296 42236 34302 42288
rect 33873 42211 33931 42217
rect 31496 42180 31616 42208
rect 32324 42180 33732 42208
rect 29564 42112 30144 42140
rect 31588 42140 31616 42180
rect 32030 42140 32036 42152
rect 31588 42112 32036 42140
rect 32030 42100 32036 42112
rect 32088 42140 32094 42152
rect 32125 42143 32183 42149
rect 32125 42140 32137 42143
rect 32088 42112 32137 42140
rect 32088 42100 32094 42112
rect 32125 42109 32137 42112
rect 32171 42109 32183 42143
rect 32125 42103 32183 42109
rect 30190 42072 30196 42084
rect 29472 42044 30196 42072
rect 30190 42032 30196 42044
rect 30248 42032 30254 42084
rect 18601 42007 18659 42013
rect 18601 41973 18613 42007
rect 18647 42004 18659 42007
rect 19058 42004 19064 42016
rect 18647 41976 19064 42004
rect 18647 41973 18659 41976
rect 18601 41967 18659 41973
rect 19058 41964 19064 41976
rect 19116 41964 19122 42016
rect 19429 42007 19487 42013
rect 19429 41973 19441 42007
rect 19475 42004 19487 42007
rect 19518 42004 19524 42016
rect 19475 41976 19524 42004
rect 19475 41973 19487 41976
rect 19429 41967 19487 41973
rect 19518 41964 19524 41976
rect 19576 41964 19582 42016
rect 21634 41964 21640 42016
rect 21692 42004 21698 42016
rect 31662 42004 31668 42016
rect 21692 41976 31668 42004
rect 21692 41964 21698 41976
rect 31662 41964 31668 41976
rect 31720 41964 31726 42016
rect 33704 42004 33732 42180
rect 33873 42177 33885 42211
rect 33919 42208 33931 42211
rect 34698 42208 34704 42220
rect 33919 42180 34704 42208
rect 33919 42177 33931 42180
rect 33873 42171 33931 42177
rect 34698 42168 34704 42180
rect 34756 42168 34762 42220
rect 35342 42168 35348 42220
rect 35400 42168 35406 42220
rect 33781 42143 33839 42149
rect 33781 42109 33793 42143
rect 33827 42109 33839 42143
rect 33781 42103 33839 42109
rect 34149 42143 34207 42149
rect 34149 42109 34161 42143
rect 34195 42140 34207 42143
rect 34238 42140 34244 42152
rect 34195 42112 34244 42140
rect 34195 42109 34207 42112
rect 34149 42103 34207 42109
rect 33796 42072 33824 42103
rect 34238 42100 34244 42112
rect 34296 42100 34302 42152
rect 35066 42100 35072 42152
rect 35124 42140 35130 42152
rect 35437 42143 35495 42149
rect 35437 42140 35449 42143
rect 35124 42112 35449 42140
rect 35124 42100 35130 42112
rect 35437 42109 35449 42112
rect 35483 42140 35495 42143
rect 35618 42140 35624 42152
rect 35483 42112 35624 42140
rect 35483 42109 35495 42112
rect 35437 42103 35495 42109
rect 35618 42100 35624 42112
rect 35676 42100 35682 42152
rect 35713 42075 35771 42081
rect 35713 42072 35725 42075
rect 33796 42044 35725 42072
rect 35713 42041 35725 42044
rect 35759 42041 35771 42075
rect 35713 42035 35771 42041
rect 35434 42004 35440 42016
rect 33704 41976 35440 42004
rect 35434 41964 35440 41976
rect 35492 41964 35498 42016
rect 35529 42007 35587 42013
rect 35529 41973 35541 42007
rect 35575 42004 35587 42007
rect 37090 42004 37096 42016
rect 35575 41976 37096 42004
rect 35575 41973 35587 41976
rect 35529 41967 35587 41973
rect 37090 41964 37096 41976
rect 37148 41964 37154 42016
rect 1104 41914 47104 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 47104 41914
rect 1104 41840 47104 41862
rect 13449 41803 13507 41809
rect 13449 41769 13461 41803
rect 13495 41800 13507 41803
rect 13538 41800 13544 41812
rect 13495 41772 13544 41800
rect 13495 41769 13507 41772
rect 13449 41763 13507 41769
rect 13538 41760 13544 41772
rect 13596 41760 13602 41812
rect 19886 41760 19892 41812
rect 19944 41800 19950 41812
rect 19944 41772 31754 41800
rect 19944 41760 19950 41772
rect 20625 41735 20683 41741
rect 20625 41701 20637 41735
rect 20671 41732 20683 41735
rect 21266 41732 21272 41744
rect 20671 41704 21272 41732
rect 20671 41701 20683 41704
rect 20625 41695 20683 41701
rect 21266 41692 21272 41704
rect 21324 41692 21330 41744
rect 31726 41732 31754 41772
rect 32122 41760 32128 41812
rect 32180 41760 32186 41812
rect 32508 41772 32812 41800
rect 32508 41732 32536 41772
rect 31726 41704 32536 41732
rect 32784 41732 32812 41772
rect 32858 41760 32864 41812
rect 32916 41800 32922 41812
rect 32916 41772 34836 41800
rect 32916 41760 32922 41772
rect 33134 41732 33140 41744
rect 32784 41704 33140 41732
rect 33134 41692 33140 41704
rect 33192 41692 33198 41744
rect 34514 41732 34520 41744
rect 34256 41704 34520 41732
rect 11330 41624 11336 41676
rect 11388 41624 11394 41676
rect 17034 41624 17040 41676
rect 17092 41664 17098 41676
rect 17405 41667 17463 41673
rect 17405 41664 17417 41667
rect 17092 41636 17417 41664
rect 17092 41624 17098 41636
rect 17405 41633 17417 41636
rect 17451 41633 17463 41667
rect 17405 41627 17463 41633
rect 19150 41624 19156 41676
rect 19208 41664 19214 41676
rect 19245 41667 19303 41673
rect 19245 41664 19257 41667
rect 19208 41636 19257 41664
rect 19208 41624 19214 41636
rect 19245 41633 19257 41636
rect 19291 41633 19303 41667
rect 32674 41664 32680 41676
rect 19245 41627 19303 41633
rect 31956 41636 32680 41664
rect 1394 41556 1400 41608
rect 1452 41596 1458 41608
rect 1949 41599 2007 41605
rect 1949 41596 1961 41599
rect 1452 41568 1961 41596
rect 1452 41556 1458 41568
rect 1949 41565 1961 41568
rect 1995 41565 2007 41599
rect 1949 41559 2007 41565
rect 11057 41599 11115 41605
rect 11057 41565 11069 41599
rect 11103 41565 11115 41599
rect 11057 41559 11115 41565
rect 934 41420 940 41472
rect 992 41460 998 41472
rect 1581 41463 1639 41469
rect 1581 41460 1593 41463
rect 992 41432 1593 41460
rect 992 41420 998 41432
rect 1581 41429 1593 41432
rect 1627 41429 1639 41463
rect 11072 41460 11100 41559
rect 12894 41556 12900 41608
rect 12952 41596 12958 41608
rect 13633 41599 13691 41605
rect 13633 41596 13645 41599
rect 12952 41568 13645 41596
rect 12952 41556 12958 41568
rect 13633 41565 13645 41568
rect 13679 41565 13691 41599
rect 13633 41559 13691 41565
rect 17129 41599 17187 41605
rect 17129 41565 17141 41599
rect 17175 41596 17187 41599
rect 17310 41596 17316 41608
rect 17175 41568 17316 41596
rect 17175 41565 17187 41568
rect 17129 41559 17187 41565
rect 17310 41556 17316 41568
rect 17368 41556 17374 41608
rect 19058 41556 19064 41608
rect 19116 41556 19122 41608
rect 19518 41605 19524 41608
rect 19512 41596 19524 41605
rect 19479 41568 19524 41596
rect 19512 41559 19524 41568
rect 19518 41556 19524 41559
rect 19576 41556 19582 41608
rect 20898 41556 20904 41608
rect 20956 41556 20962 41608
rect 21818 41556 21824 41608
rect 21876 41596 21882 41608
rect 22097 41599 22155 41605
rect 22097 41596 22109 41599
rect 21876 41568 22109 41596
rect 21876 41556 21882 41568
rect 22097 41565 22109 41568
rect 22143 41565 22155 41599
rect 22097 41559 22155 41565
rect 24302 41556 24308 41608
rect 24360 41596 24366 41608
rect 24397 41599 24455 41605
rect 24397 41596 24409 41599
rect 24360 41568 24409 41596
rect 24360 41556 24366 41568
rect 24397 41565 24409 41568
rect 24443 41565 24455 41599
rect 24397 41559 24455 41565
rect 26878 41556 26884 41608
rect 26936 41596 26942 41608
rect 31846 41596 31852 41608
rect 26936 41568 31852 41596
rect 26936 41556 26942 41568
rect 31846 41556 31852 41568
rect 31904 41556 31910 41608
rect 23934 41488 23940 41540
rect 23992 41528 23998 41540
rect 24642 41531 24700 41537
rect 24642 41528 24654 41531
rect 23992 41500 24654 41528
rect 23992 41488 23998 41500
rect 24642 41497 24654 41500
rect 24688 41497 24700 41531
rect 24642 41491 24700 41497
rect 27338 41488 27344 41540
rect 27396 41528 27402 41540
rect 27982 41528 27988 41540
rect 27396 41500 27988 41528
rect 27396 41488 27402 41500
rect 27982 41488 27988 41500
rect 28040 41488 28046 41540
rect 29914 41488 29920 41540
rect 29972 41528 29978 41540
rect 31205 41531 31263 41537
rect 31205 41528 31217 41531
rect 29972 41500 31217 41528
rect 29972 41488 29978 41500
rect 31205 41497 31217 41500
rect 31251 41528 31263 41531
rect 31570 41528 31576 41540
rect 31251 41500 31576 41528
rect 31251 41497 31263 41500
rect 31205 41491 31263 41497
rect 31570 41488 31576 41500
rect 31628 41488 31634 41540
rect 31662 41488 31668 41540
rect 31720 41528 31726 41540
rect 31956 41528 31984 41636
rect 32674 41624 32680 41636
rect 32732 41624 32738 41676
rect 32769 41667 32827 41673
rect 32769 41633 32781 41667
rect 32815 41664 32827 41667
rect 34256 41664 34284 41704
rect 34514 41692 34520 41704
rect 34572 41692 34578 41744
rect 34808 41732 34836 41772
rect 34882 41760 34888 41812
rect 34940 41760 34946 41812
rect 35158 41760 35164 41812
rect 35216 41760 35222 41812
rect 35434 41760 35440 41812
rect 35492 41800 35498 41812
rect 36722 41800 36728 41812
rect 35492 41772 36728 41800
rect 35492 41760 35498 41772
rect 36722 41760 36728 41772
rect 36780 41800 36786 41812
rect 37185 41803 37243 41809
rect 37185 41800 37197 41803
rect 36780 41772 37197 41800
rect 36780 41760 36786 41772
rect 37185 41769 37197 41772
rect 37231 41800 37243 41803
rect 37642 41800 37648 41812
rect 37231 41772 37648 41800
rect 37231 41769 37243 41772
rect 37185 41763 37243 41769
rect 37642 41760 37648 41772
rect 37700 41760 37706 41812
rect 38749 41803 38807 41809
rect 38749 41769 38761 41803
rect 38795 41800 38807 41803
rect 38838 41800 38844 41812
rect 38795 41772 38844 41800
rect 38795 41769 38807 41772
rect 38749 41763 38807 41769
rect 38838 41760 38844 41772
rect 38896 41760 38902 41812
rect 36633 41735 36691 41741
rect 36633 41732 36645 41735
rect 34808 41704 36645 41732
rect 36633 41701 36645 41704
rect 36679 41701 36691 41735
rect 36633 41695 36691 41701
rect 34790 41664 34796 41676
rect 32815 41636 34284 41664
rect 34348 41636 34796 41664
rect 32815 41633 32827 41636
rect 32769 41627 32827 41633
rect 32030 41556 32036 41608
rect 32088 41596 32094 41608
rect 32953 41599 33011 41605
rect 32953 41596 32965 41599
rect 32088 41568 32965 41596
rect 32088 41556 32094 41568
rect 32953 41565 32965 41568
rect 32999 41596 33011 41599
rect 33318 41596 33324 41608
rect 32999 41568 33324 41596
rect 32999 41565 33011 41568
rect 32953 41559 33011 41565
rect 33318 41556 33324 41568
rect 33376 41556 33382 41608
rect 34348 41605 34376 41636
rect 34790 41624 34796 41636
rect 34848 41624 34854 41676
rect 34885 41667 34943 41673
rect 34885 41633 34897 41667
rect 34931 41664 34943 41667
rect 35342 41664 35348 41676
rect 34931 41636 35348 41664
rect 34931 41633 34943 41636
rect 34885 41627 34943 41633
rect 35342 41624 35348 41636
rect 35400 41624 35406 41676
rect 35897 41667 35955 41673
rect 35897 41633 35909 41667
rect 35943 41664 35955 41667
rect 36354 41664 36360 41676
rect 35943 41636 36360 41664
rect 35943 41633 35955 41636
rect 35897 41627 35955 41633
rect 36354 41624 36360 41636
rect 36412 41624 36418 41676
rect 34333 41599 34391 41605
rect 34333 41565 34345 41599
rect 34379 41565 34391 41599
rect 34333 41559 34391 41565
rect 34517 41599 34575 41605
rect 34517 41565 34529 41599
rect 34563 41596 34575 41599
rect 34563 41568 34928 41596
rect 34563 41565 34575 41568
rect 34517 41559 34575 41565
rect 34348 41528 34376 41559
rect 31720 41500 31984 41528
rect 32048 41500 32444 41528
rect 34348 41500 34560 41528
rect 31720 41488 31726 41500
rect 18046 41460 18052 41472
rect 11072 41432 18052 41460
rect 1581 41423 1639 41429
rect 18046 41420 18052 41432
rect 18104 41420 18110 41472
rect 18874 41420 18880 41472
rect 18932 41420 18938 41472
rect 20714 41420 20720 41472
rect 20772 41420 20778 41472
rect 21913 41463 21971 41469
rect 21913 41429 21925 41463
rect 21959 41460 21971 41463
rect 22094 41460 22100 41472
rect 21959 41432 22100 41460
rect 21959 41429 21971 41432
rect 21913 41423 21971 41429
rect 22094 41420 22100 41432
rect 22152 41420 22158 41472
rect 24486 41420 24492 41472
rect 24544 41460 24550 41472
rect 25777 41463 25835 41469
rect 25777 41460 25789 41463
rect 24544 41432 25789 41460
rect 24544 41420 24550 41432
rect 25777 41429 25789 41432
rect 25823 41429 25835 41463
rect 25777 41423 25835 41429
rect 30190 41420 30196 41472
rect 30248 41460 30254 41472
rect 31481 41463 31539 41469
rect 31481 41460 31493 41463
rect 30248 41432 31493 41460
rect 30248 41420 30254 41432
rect 31481 41429 31493 41432
rect 31527 41460 31539 41463
rect 32048 41460 32076 41500
rect 32416 41472 32444 41500
rect 31527 41432 32076 41460
rect 31527 41429 31539 41432
rect 31481 41423 31539 41429
rect 32398 41420 32404 41472
rect 32456 41460 32462 41472
rect 32493 41463 32551 41469
rect 32493 41460 32505 41463
rect 32456 41432 32505 41460
rect 32456 41420 32462 41432
rect 32493 41429 32505 41432
rect 32539 41429 32551 41463
rect 32493 41423 32551 41429
rect 32582 41420 32588 41472
rect 32640 41420 32646 41472
rect 34422 41420 34428 41472
rect 34480 41420 34486 41472
rect 34532 41460 34560 41500
rect 34606 41488 34612 41540
rect 34664 41528 34670 41540
rect 34701 41531 34759 41537
rect 34701 41528 34713 41531
rect 34664 41500 34713 41528
rect 34664 41488 34670 41500
rect 34701 41497 34713 41500
rect 34747 41528 34759 41531
rect 34790 41528 34796 41540
rect 34747 41500 34796 41528
rect 34747 41497 34759 41500
rect 34701 41491 34759 41497
rect 34790 41488 34796 41500
rect 34848 41488 34854 41540
rect 34900 41528 34928 41568
rect 34974 41556 34980 41608
rect 35032 41596 35038 41608
rect 35032 41568 35388 41596
rect 35032 41556 35038 41568
rect 35066 41528 35072 41540
rect 34900 41500 35072 41528
rect 35066 41488 35072 41500
rect 35124 41488 35130 41540
rect 35253 41531 35311 41537
rect 35253 41497 35265 41531
rect 35299 41497 35311 41531
rect 35360 41528 35388 41568
rect 35434 41556 35440 41608
rect 35492 41596 35498 41608
rect 35529 41599 35587 41605
rect 35529 41596 35541 41599
rect 35492 41568 35541 41596
rect 35492 41556 35498 41568
rect 35529 41565 35541 41568
rect 35575 41565 35587 41599
rect 35529 41559 35587 41565
rect 35621 41599 35679 41605
rect 35621 41565 35633 41599
rect 35667 41596 35679 41599
rect 35710 41596 35716 41608
rect 35667 41568 35716 41596
rect 35667 41565 35679 41568
rect 35621 41559 35679 41565
rect 35710 41556 35716 41568
rect 35768 41556 35774 41608
rect 35989 41599 36047 41605
rect 35989 41565 36001 41599
rect 36035 41565 36047 41599
rect 36648 41596 36676 41695
rect 37001 41599 37059 41605
rect 37001 41596 37013 41599
rect 36648 41568 37013 41596
rect 35989 41559 36047 41565
rect 37001 41565 37013 41568
rect 37047 41565 37059 41599
rect 37001 41559 37059 41565
rect 36004 41528 36032 41559
rect 35360 41500 36032 41528
rect 38565 41531 38623 41537
rect 35253 41491 35311 41497
rect 35268 41460 35296 41491
rect 35636 41472 35664 41500
rect 38565 41497 38577 41531
rect 38611 41528 38623 41531
rect 39390 41528 39396 41540
rect 38611 41500 39396 41528
rect 38611 41497 38623 41500
rect 38565 41491 38623 41497
rect 39390 41488 39396 41500
rect 39448 41488 39454 41540
rect 34532 41432 35296 41460
rect 35342 41420 35348 41472
rect 35400 41460 35406 41472
rect 35526 41460 35532 41472
rect 35400 41432 35532 41460
rect 35400 41420 35406 41432
rect 35526 41420 35532 41432
rect 35584 41420 35590 41472
rect 35618 41420 35624 41472
rect 35676 41420 35682 41472
rect 35713 41463 35771 41469
rect 35713 41429 35725 41463
rect 35759 41460 35771 41463
rect 35986 41460 35992 41472
rect 35759 41432 35992 41460
rect 35759 41429 35771 41432
rect 35713 41423 35771 41429
rect 35986 41420 35992 41432
rect 36044 41460 36050 41472
rect 36446 41460 36452 41472
rect 36044 41432 36452 41460
rect 36044 41420 36050 41432
rect 36446 41420 36452 41432
rect 36504 41420 36510 41472
rect 38654 41420 38660 41472
rect 38712 41460 38718 41472
rect 38765 41463 38823 41469
rect 38765 41460 38777 41463
rect 38712 41432 38777 41460
rect 38712 41420 38718 41432
rect 38765 41429 38777 41432
rect 38811 41429 38823 41463
rect 38765 41423 38823 41429
rect 38930 41420 38936 41472
rect 38988 41420 38994 41472
rect 1104 41370 47104 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 35594 41370
rect 35646 41318 35658 41370
rect 35710 41318 35722 41370
rect 35774 41318 35786 41370
rect 35838 41318 35850 41370
rect 35902 41318 47104 41370
rect 1104 41296 47104 41318
rect 10042 41216 10048 41268
rect 10100 41256 10106 41268
rect 10100 41228 23888 41256
rect 10100 41216 10106 41228
rect 11330 41188 11336 41200
rect 11072 41160 11336 41188
rect 11072 41129 11100 41160
rect 11330 41148 11336 41160
rect 11388 41188 11394 41200
rect 11609 41191 11667 41197
rect 11609 41188 11621 41191
rect 11388 41160 11621 41188
rect 11388 41148 11394 41160
rect 11609 41157 11621 41160
rect 11655 41157 11667 41191
rect 11609 41151 11667 41157
rect 17402 41148 17408 41200
rect 17460 41188 17466 41200
rect 18414 41188 18420 41200
rect 17460 41160 18420 41188
rect 17460 41148 17466 41160
rect 18414 41148 18420 41160
rect 18472 41188 18478 41200
rect 18472 41160 18828 41188
rect 18472 41148 18478 41160
rect 11057 41123 11115 41129
rect 11057 41089 11069 41123
rect 11103 41089 11115 41123
rect 11057 41083 11115 41089
rect 12158 41080 12164 41132
rect 12216 41120 12222 41132
rect 12805 41123 12863 41129
rect 12805 41120 12817 41123
rect 12216 41092 12817 41120
rect 12216 41080 12222 41092
rect 12805 41089 12817 41092
rect 12851 41089 12863 41123
rect 12805 41083 12863 41089
rect 12897 41123 12955 41129
rect 12897 41089 12909 41123
rect 12943 41120 12955 41123
rect 13630 41120 13636 41132
rect 12943 41092 13636 41120
rect 12943 41089 12955 41092
rect 12897 41083 12955 41089
rect 13630 41080 13636 41092
rect 13688 41080 13694 41132
rect 14458 41129 14464 41132
rect 14452 41083 14464 41129
rect 14458 41080 14464 41083
rect 14516 41080 14522 41132
rect 16942 41080 16948 41132
rect 17000 41080 17006 41132
rect 17304 41123 17362 41129
rect 17304 41089 17316 41123
rect 17350 41120 17362 41123
rect 18598 41120 18604 41132
rect 17350 41092 18604 41120
rect 17350 41089 17362 41092
rect 17304 41083 17362 41089
rect 18598 41080 18604 41092
rect 18656 41080 18662 41132
rect 18800 41129 18828 41160
rect 18874 41148 18880 41200
rect 18932 41188 18938 41200
rect 19030 41191 19088 41197
rect 19030 41188 19042 41191
rect 18932 41160 19042 41188
rect 18932 41148 18938 41160
rect 19030 41157 19042 41160
rect 19076 41157 19088 41191
rect 19030 41151 19088 41157
rect 20524 41191 20582 41197
rect 20524 41157 20536 41191
rect 20570 41188 20582 41191
rect 20714 41188 20720 41200
rect 20570 41160 20720 41188
rect 20570 41157 20582 41160
rect 20524 41151 20582 41157
rect 20714 41148 20720 41160
rect 20772 41148 20778 41200
rect 22094 41197 22100 41200
rect 22088 41151 22100 41197
rect 22152 41188 22158 41200
rect 23860 41188 23888 41228
rect 23934 41216 23940 41268
rect 23992 41216 23998 41268
rect 26050 41256 26056 41268
rect 24044 41228 26056 41256
rect 24044 41188 24072 41228
rect 26050 41216 26056 41228
rect 26108 41216 26114 41268
rect 34606 41216 34612 41268
rect 34664 41256 34670 41268
rect 34882 41256 34888 41268
rect 34664 41228 34888 41256
rect 34664 41216 34670 41228
rect 34882 41216 34888 41228
rect 34940 41216 34946 41268
rect 34977 41259 35035 41265
rect 34977 41225 34989 41259
rect 35023 41256 35035 41259
rect 35066 41256 35072 41268
rect 35023 41228 35072 41256
rect 35023 41225 35035 41228
rect 34977 41219 35035 41225
rect 35066 41216 35072 41228
rect 35124 41256 35130 41268
rect 35342 41256 35348 41268
rect 35124 41228 35348 41256
rect 35124 41216 35130 41228
rect 35342 41216 35348 41228
rect 35400 41216 35406 41268
rect 37369 41259 37427 41265
rect 37369 41225 37381 41259
rect 37415 41225 37427 41259
rect 37369 41219 37427 41225
rect 37476 41228 39528 41256
rect 22152 41160 22188 41188
rect 23860 41160 24072 41188
rect 22094 41148 22100 41151
rect 22152 41148 22158 41160
rect 24210 41148 24216 41200
rect 24268 41188 24274 41200
rect 24734 41191 24792 41197
rect 24734 41188 24746 41191
rect 24268 41160 24746 41188
rect 24268 41148 24274 41160
rect 24734 41157 24746 41160
rect 24780 41157 24792 41191
rect 24734 41151 24792 41157
rect 34146 41148 34152 41200
rect 34204 41188 34210 41200
rect 36078 41188 36084 41200
rect 34204 41160 35480 41188
rect 34204 41148 34210 41160
rect 18785 41123 18843 41129
rect 18785 41089 18797 41123
rect 18831 41089 18843 41123
rect 18785 41083 18843 41089
rect 20257 41123 20315 41129
rect 20257 41089 20269 41123
rect 20303 41120 20315 41123
rect 20303 41092 23980 41120
rect 20303 41089 20315 41092
rect 20257 41083 20315 41089
rect 13081 41055 13139 41061
rect 13081 41021 13093 41055
rect 13127 41052 13139 41055
rect 13262 41052 13268 41064
rect 13127 41024 13268 41052
rect 13127 41021 13139 41024
rect 13081 41015 13139 41021
rect 13262 41012 13268 41024
rect 13320 41012 13326 41064
rect 13998 41012 14004 41064
rect 14056 41052 14062 41064
rect 14185 41055 14243 41061
rect 14185 41052 14197 41055
rect 14056 41024 14197 41052
rect 14056 41012 14062 41024
rect 14185 41021 14197 41024
rect 14231 41021 14243 41055
rect 14185 41015 14243 41021
rect 17034 41012 17040 41064
rect 17092 41012 17098 41064
rect 21726 41012 21732 41064
rect 21784 41052 21790 41064
rect 21836 41061 21864 41092
rect 21821 41055 21879 41061
rect 21821 41052 21833 41055
rect 21784 41024 21833 41052
rect 21784 41012 21790 41024
rect 21821 41021 21833 41024
rect 21867 41021 21879 41055
rect 23952 41052 23980 41092
rect 24026 41080 24032 41132
rect 24084 41120 24090 41132
rect 24121 41123 24179 41129
rect 24121 41120 24133 41123
rect 24084 41092 24133 41120
rect 24084 41080 24090 41092
rect 24121 41089 24133 41092
rect 24167 41089 24179 41123
rect 24121 41083 24179 41089
rect 24394 41080 24400 41132
rect 24452 41080 24458 41132
rect 33686 41080 33692 41132
rect 33744 41120 33750 41132
rect 33965 41123 34023 41129
rect 33965 41120 33977 41123
rect 33744 41092 33977 41120
rect 33744 41080 33750 41092
rect 33965 41089 33977 41092
rect 34011 41120 34023 41123
rect 34422 41120 34428 41132
rect 34011 41092 34428 41120
rect 34011 41089 34023 41092
rect 33965 41083 34023 41089
rect 34422 41080 34428 41092
rect 34480 41080 34486 41132
rect 34974 41080 34980 41132
rect 35032 41120 35038 41132
rect 35253 41123 35311 41129
rect 35253 41120 35265 41123
rect 35032 41092 35265 41120
rect 35032 41080 35038 41092
rect 35253 41089 35265 41092
rect 35299 41089 35311 41123
rect 35253 41083 35311 41089
rect 24302 41052 24308 41064
rect 23952 41024 24308 41052
rect 21821 41015 21879 41021
rect 24302 41012 24308 41024
rect 24360 41052 24366 41064
rect 24489 41055 24547 41061
rect 24489 41052 24501 41055
rect 24360 41024 24501 41052
rect 24360 41012 24366 41024
rect 24489 41021 24501 41024
rect 24535 41021 24547 41055
rect 24489 41015 24547 41021
rect 27798 41012 27804 41064
rect 27856 41052 27862 41064
rect 27893 41055 27951 41061
rect 27893 41052 27905 41055
rect 27856 41024 27905 41052
rect 27856 41012 27862 41024
rect 27893 41021 27905 41024
rect 27939 41021 27951 41055
rect 27893 41015 27951 41021
rect 28169 41055 28227 41061
rect 28169 41021 28181 41055
rect 28215 41052 28227 41055
rect 28442 41052 28448 41064
rect 28215 41024 28448 41052
rect 28215 41021 28227 41024
rect 28169 41015 28227 41021
rect 28442 41012 28448 41024
rect 28500 41012 28506 41064
rect 34790 41012 34796 41064
rect 34848 41012 34854 41064
rect 35268 41052 35296 41083
rect 35342 41080 35348 41132
rect 35400 41080 35406 41132
rect 35452 41129 35480 41160
rect 35728 41160 36084 41188
rect 35437 41123 35495 41129
rect 35437 41089 35449 41123
rect 35483 41089 35495 41123
rect 35437 41083 35495 41089
rect 35526 41080 35532 41132
rect 35584 41120 35590 41132
rect 35728 41129 35756 41160
rect 36078 41148 36084 41160
rect 36136 41148 36142 41200
rect 36173 41191 36231 41197
rect 36173 41157 36185 41191
rect 36219 41188 36231 41191
rect 36722 41188 36728 41200
rect 36219 41160 36728 41188
rect 36219 41157 36231 41160
rect 36173 41151 36231 41157
rect 36722 41148 36728 41160
rect 36780 41148 36786 41200
rect 36998 41148 37004 41200
rect 37056 41188 37062 41200
rect 37384 41188 37412 41219
rect 37056 41160 37412 41188
rect 37056 41148 37062 41160
rect 35621 41123 35679 41129
rect 35621 41120 35633 41123
rect 35584 41092 35633 41120
rect 35584 41080 35590 41092
rect 35621 41089 35633 41092
rect 35667 41089 35679 41123
rect 35621 41083 35679 41089
rect 35713 41123 35771 41129
rect 35713 41089 35725 41123
rect 35759 41089 35771 41123
rect 35713 41083 35771 41089
rect 35897 41123 35955 41129
rect 35897 41089 35909 41123
rect 35943 41120 35955 41123
rect 36909 41123 36967 41129
rect 36909 41120 36921 41123
rect 35943 41092 36921 41120
rect 35943 41089 35955 41092
rect 35897 41083 35955 41089
rect 36909 41089 36921 41092
rect 36955 41089 36967 41123
rect 36909 41083 36967 41089
rect 37274 41080 37280 41132
rect 37332 41080 37338 41132
rect 35802 41052 35808 41064
rect 35268 41024 35808 41052
rect 35802 41012 35808 41024
rect 35860 41012 35866 41064
rect 36633 41055 36691 41061
rect 36633 41021 36645 41055
rect 36679 41021 36691 41055
rect 36633 41015 36691 41021
rect 36725 41055 36783 41061
rect 36725 41021 36737 41055
rect 36771 41052 36783 41055
rect 36814 41052 36820 41064
rect 36771 41024 36820 41052
rect 36771 41021 36783 41024
rect 36725 41015 36783 41021
rect 10686 40944 10692 40996
rect 10744 40984 10750 40996
rect 12437 40987 12495 40993
rect 12437 40984 12449 40987
rect 10744 40956 12449 40984
rect 10744 40944 10750 40956
rect 12437 40953 12449 40956
rect 12483 40953 12495 40987
rect 12437 40947 12495 40953
rect 21634 40944 21640 40996
rect 21692 40944 21698 40996
rect 24210 40944 24216 40996
rect 24268 40944 24274 40996
rect 34422 40944 34428 40996
rect 34480 40984 34486 40996
rect 34808 40984 34836 41012
rect 34480 40956 34836 40984
rect 34480 40944 34486 40956
rect 35342 40944 35348 40996
rect 35400 40984 35406 40996
rect 36173 40987 36231 40993
rect 35400 40956 35848 40984
rect 35400 40944 35406 40956
rect 10778 40876 10784 40928
rect 10836 40916 10842 40928
rect 10873 40919 10931 40925
rect 10873 40916 10885 40919
rect 10836 40888 10885 40916
rect 10836 40876 10842 40888
rect 10873 40885 10885 40888
rect 10919 40885 10931 40919
rect 10873 40879 10931 40885
rect 11514 40876 11520 40928
rect 11572 40916 11578 40928
rect 11701 40919 11759 40925
rect 11701 40916 11713 40919
rect 11572 40888 11713 40916
rect 11572 40876 11578 40888
rect 11701 40885 11713 40888
rect 11747 40885 11759 40919
rect 11701 40879 11759 40885
rect 15378 40876 15384 40928
rect 15436 40916 15442 40928
rect 15565 40919 15623 40925
rect 15565 40916 15577 40919
rect 15436 40888 15577 40916
rect 15436 40876 15442 40888
rect 15565 40885 15577 40888
rect 15611 40885 15623 40919
rect 15565 40879 15623 40885
rect 16574 40876 16580 40928
rect 16632 40916 16638 40928
rect 16761 40919 16819 40925
rect 16761 40916 16773 40919
rect 16632 40888 16773 40916
rect 16632 40876 16638 40888
rect 16761 40885 16773 40888
rect 16807 40885 16819 40919
rect 16761 40879 16819 40885
rect 18230 40876 18236 40928
rect 18288 40916 18294 40928
rect 18417 40919 18475 40925
rect 18417 40916 18429 40919
rect 18288 40888 18429 40916
rect 18288 40876 18294 40888
rect 18417 40885 18429 40888
rect 18463 40885 18475 40919
rect 18417 40879 18475 40885
rect 20165 40919 20223 40925
rect 20165 40885 20177 40919
rect 20211 40916 20223 40919
rect 20990 40916 20996 40928
rect 20211 40888 20996 40916
rect 20211 40885 20223 40888
rect 20165 40879 20223 40885
rect 20990 40876 20996 40888
rect 21048 40876 21054 40928
rect 22002 40876 22008 40928
rect 22060 40916 22066 40928
rect 23201 40919 23259 40925
rect 23201 40916 23213 40919
rect 22060 40888 23213 40916
rect 22060 40876 22066 40888
rect 23201 40885 23213 40888
rect 23247 40885 23259 40919
rect 23201 40879 23259 40885
rect 25866 40876 25872 40928
rect 25924 40876 25930 40928
rect 34149 40919 34207 40925
rect 34149 40885 34161 40919
rect 34195 40916 34207 40919
rect 34238 40916 34244 40928
rect 34195 40888 34244 40916
rect 34195 40885 34207 40888
rect 34149 40879 34207 40885
rect 34238 40876 34244 40888
rect 34296 40876 34302 40928
rect 34790 40876 34796 40928
rect 34848 40916 34854 40928
rect 35713 40919 35771 40925
rect 35713 40916 35725 40919
rect 34848 40888 35725 40916
rect 34848 40876 34854 40888
rect 35713 40885 35725 40888
rect 35759 40885 35771 40919
rect 35820 40916 35848 40956
rect 36173 40953 36185 40987
rect 36219 40984 36231 40987
rect 36262 40984 36268 40996
rect 36219 40956 36268 40984
rect 36219 40953 36231 40956
rect 36173 40947 36231 40953
rect 36262 40944 36268 40956
rect 36320 40944 36326 40996
rect 36538 40944 36544 40996
rect 36596 40984 36602 40996
rect 36648 40984 36676 41015
rect 36814 41012 36820 41024
rect 36872 41052 36878 41064
rect 37476 41052 37504 41228
rect 38933 41191 38991 41197
rect 36872 41024 37504 41052
rect 37568 41160 38148 41188
rect 36872 41012 36878 41024
rect 37568 40984 37596 41160
rect 37642 41080 37648 41132
rect 37700 41080 37706 41132
rect 38120 41129 38148 41160
rect 38933 41157 38945 41191
rect 38979 41188 38991 41191
rect 39390 41188 39396 41200
rect 38979 41160 39396 41188
rect 38979 41157 38991 41160
rect 38933 41151 38991 41157
rect 39390 41148 39396 41160
rect 39448 41148 39454 41200
rect 38105 41123 38163 41129
rect 38105 41089 38117 41123
rect 38151 41089 38163 41123
rect 38105 41083 38163 41089
rect 36596 40956 37596 40984
rect 37660 40984 37688 41080
rect 38120 41052 38148 41083
rect 38378 41080 38384 41132
rect 38436 41080 38442 41132
rect 38654 41080 38660 41132
rect 38712 41080 38718 41132
rect 38838 41080 38844 41132
rect 38896 41080 38902 41132
rect 38930 41052 38936 41064
rect 38120 41024 38936 41052
rect 38930 41012 38936 41024
rect 38988 41012 38994 41064
rect 39206 41012 39212 41064
rect 39264 41052 39270 41064
rect 39301 41055 39359 41061
rect 39301 41052 39313 41055
rect 39264 41024 39313 41052
rect 39264 41012 39270 41024
rect 39301 41021 39313 41024
rect 39347 41021 39359 41055
rect 39301 41015 39359 41021
rect 39393 41055 39451 41061
rect 39393 41021 39405 41055
rect 39439 41052 39451 41055
rect 39500 41052 39528 41228
rect 40126 41052 40132 41064
rect 39439 41024 40132 41052
rect 39439 41021 39451 41024
rect 39393 41015 39451 41021
rect 40126 41012 40132 41024
rect 40184 41012 40190 41064
rect 38470 40984 38476 40996
rect 37660 40956 38476 40984
rect 36596 40944 36602 40956
rect 38470 40944 38476 40956
rect 38528 40944 38534 40996
rect 38565 40987 38623 40993
rect 38565 40953 38577 40987
rect 38611 40984 38623 40987
rect 39577 40987 39635 40993
rect 39577 40984 39589 40987
rect 38611 40956 39589 40984
rect 38611 40953 38623 40956
rect 38565 40947 38623 40953
rect 39577 40953 39589 40956
rect 39623 40953 39635 40987
rect 39577 40947 39635 40953
rect 36354 40916 36360 40928
rect 35820 40888 36360 40916
rect 35713 40879 35771 40885
rect 36354 40876 36360 40888
rect 36412 40876 36418 40928
rect 37090 40876 37096 40928
rect 37148 40916 37154 40928
rect 38197 40919 38255 40925
rect 38197 40916 38209 40919
rect 37148 40888 38209 40916
rect 37148 40876 37154 40888
rect 38197 40885 38209 40888
rect 38243 40885 38255 40919
rect 38197 40879 38255 40885
rect 1104 40826 47104 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 47104 40826
rect 1104 40752 47104 40774
rect 3513 40715 3571 40721
rect 3513 40681 3525 40715
rect 3559 40712 3571 40715
rect 10226 40712 10232 40724
rect 3559 40684 10232 40712
rect 3559 40681 3571 40684
rect 3513 40675 3571 40681
rect 2038 40468 2044 40520
rect 2096 40468 2102 40520
rect 2133 40511 2191 40517
rect 2133 40477 2145 40511
rect 2179 40508 2191 40511
rect 3418 40508 3424 40520
rect 2179 40480 3424 40508
rect 2179 40477 2191 40480
rect 2133 40471 2191 40477
rect 3418 40468 3424 40480
rect 3476 40468 3482 40520
rect 2378 40443 2436 40449
rect 2378 40440 2390 40443
rect 1872 40412 2390 40440
rect 1872 40381 1900 40412
rect 2378 40409 2390 40412
rect 2424 40409 2436 40443
rect 2378 40403 2436 40409
rect 1857 40375 1915 40381
rect 1857 40341 1869 40375
rect 1903 40341 1915 40375
rect 1857 40335 1915 40341
rect 2590 40332 2596 40384
rect 2648 40372 2654 40384
rect 3528 40372 3556 40675
rect 10226 40672 10232 40684
rect 10284 40672 10290 40724
rect 12158 40672 12164 40724
rect 12216 40672 12222 40724
rect 12526 40672 12532 40724
rect 12584 40712 12590 40724
rect 13998 40712 14004 40724
rect 12584 40684 14004 40712
rect 12584 40672 12590 40684
rect 13998 40672 14004 40684
rect 14056 40672 14062 40724
rect 16666 40712 16672 40724
rect 16316 40684 16672 40712
rect 10778 40576 10784 40588
rect 9968 40548 10784 40576
rect 8938 40468 8944 40520
rect 8996 40508 9002 40520
rect 9968 40508 9996 40548
rect 10778 40536 10784 40548
rect 10836 40536 10842 40588
rect 12452 40548 12664 40576
rect 8996 40480 9996 40508
rect 8996 40468 9002 40480
rect 10686 40468 10692 40520
rect 10744 40468 10750 40520
rect 12452 40517 12480 40548
rect 12437 40511 12495 40517
rect 12437 40477 12449 40511
rect 12483 40477 12495 40511
rect 12437 40471 12495 40477
rect 12526 40468 12532 40520
rect 12584 40468 12590 40520
rect 12636 40508 12664 40548
rect 13998 40536 14004 40588
rect 14056 40576 14062 40588
rect 14553 40579 14611 40585
rect 14553 40576 14565 40579
rect 14056 40548 14565 40576
rect 14056 40536 14062 40548
rect 14553 40545 14565 40548
rect 14599 40545 14611 40579
rect 14553 40539 14611 40545
rect 15841 40579 15899 40585
rect 15841 40545 15853 40579
rect 15887 40576 15899 40579
rect 16316 40576 16344 40684
rect 16666 40672 16672 40684
rect 16724 40712 16730 40724
rect 20165 40715 20223 40721
rect 16724 40684 18920 40712
rect 16724 40672 16730 40684
rect 17773 40647 17831 40653
rect 17773 40613 17785 40647
rect 17819 40644 17831 40647
rect 18892 40644 18920 40684
rect 20165 40681 20177 40715
rect 20211 40712 20223 40715
rect 20898 40712 20904 40724
rect 20211 40684 20904 40712
rect 20211 40681 20223 40684
rect 20165 40675 20223 40681
rect 20898 40672 20904 40684
rect 20956 40672 20962 40724
rect 21818 40672 21824 40724
rect 21876 40672 21882 40724
rect 22554 40672 22560 40724
rect 22612 40712 22618 40724
rect 22612 40684 34836 40712
rect 22612 40672 22618 40684
rect 34808 40644 34836 40684
rect 36722 40672 36728 40724
rect 36780 40712 36786 40724
rect 36909 40715 36967 40721
rect 36909 40712 36921 40715
rect 36780 40684 36921 40712
rect 36780 40672 36786 40684
rect 36909 40681 36921 40684
rect 36955 40681 36967 40715
rect 36909 40675 36967 40681
rect 38470 40672 38476 40724
rect 38528 40712 38534 40724
rect 39945 40715 40003 40721
rect 39945 40712 39957 40715
rect 38528 40684 39957 40712
rect 38528 40672 38534 40684
rect 39945 40681 39957 40684
rect 39991 40681 40003 40715
rect 39945 40675 40003 40681
rect 37826 40644 37832 40656
rect 17819 40616 18828 40644
rect 18892 40616 22508 40644
rect 34808 40616 37832 40644
rect 17819 40613 17831 40616
rect 17773 40607 17831 40613
rect 15887 40548 16344 40576
rect 15887 40545 15899 40548
rect 15841 40539 15899 40545
rect 18230 40536 18236 40588
rect 18288 40536 18294 40588
rect 18417 40579 18475 40585
rect 18417 40545 18429 40579
rect 18463 40576 18475 40579
rect 18690 40576 18696 40588
rect 18463 40548 18696 40576
rect 18463 40545 18475 40548
rect 18417 40539 18475 40545
rect 18690 40536 18696 40548
rect 18748 40536 18754 40588
rect 13170 40508 13176 40520
rect 12636 40480 13176 40508
rect 13170 40468 13176 40480
rect 13228 40468 13234 40520
rect 14277 40511 14335 40517
rect 14277 40477 14289 40511
rect 14323 40508 14335 40511
rect 15102 40508 15108 40520
rect 14323 40480 15108 40508
rect 14323 40477 14335 40480
rect 14277 40471 14335 40477
rect 15102 40468 15108 40480
rect 15160 40508 15166 40520
rect 16574 40517 16580 40520
rect 16301 40511 16359 40517
rect 16301 40508 16313 40511
rect 15160 40480 16313 40508
rect 15160 40468 15166 40480
rect 16301 40477 16313 40480
rect 16347 40477 16359 40511
rect 16568 40508 16580 40517
rect 16535 40480 16580 40508
rect 16301 40471 16359 40477
rect 16568 40471 16580 40480
rect 8846 40400 8852 40452
rect 8904 40440 8910 40452
rect 9186 40443 9244 40449
rect 9186 40440 9198 40443
rect 8904 40412 9198 40440
rect 8904 40400 8910 40412
rect 9186 40409 9198 40412
rect 9232 40409 9244 40443
rect 11026 40443 11084 40449
rect 11026 40440 11038 40443
rect 9186 40403 9244 40409
rect 10520 40412 11038 40440
rect 2648 40344 3556 40372
rect 5813 40375 5871 40381
rect 2648 40332 2654 40344
rect 5813 40341 5825 40375
rect 5859 40372 5871 40375
rect 6181 40375 6239 40381
rect 6181 40372 6193 40375
rect 5859 40344 6193 40372
rect 5859 40341 5871 40344
rect 5813 40335 5871 40341
rect 6181 40341 6193 40344
rect 6227 40372 6239 40375
rect 6549 40375 6607 40381
rect 6549 40372 6561 40375
rect 6227 40344 6561 40372
rect 6227 40341 6239 40344
rect 6181 40335 6239 40341
rect 6549 40341 6561 40344
rect 6595 40372 6607 40375
rect 6914 40372 6920 40384
rect 6595 40344 6920 40372
rect 6595 40341 6607 40344
rect 6549 40335 6607 40341
rect 6914 40332 6920 40344
rect 6972 40372 6978 40384
rect 7193 40375 7251 40381
rect 7193 40372 7205 40375
rect 6972 40344 7205 40372
rect 6972 40332 6978 40344
rect 7193 40341 7205 40344
rect 7239 40372 7251 40375
rect 7561 40375 7619 40381
rect 7561 40372 7573 40375
rect 7239 40344 7573 40372
rect 7239 40341 7251 40344
rect 7193 40335 7251 40341
rect 7561 40341 7573 40344
rect 7607 40341 7619 40375
rect 7561 40335 7619 40341
rect 10321 40375 10379 40381
rect 10321 40341 10333 40375
rect 10367 40372 10379 40375
rect 10410 40372 10416 40384
rect 10367 40344 10416 40372
rect 10367 40341 10379 40344
rect 10321 40335 10379 40341
rect 10410 40332 10416 40344
rect 10468 40332 10474 40384
rect 10520 40381 10548 40412
rect 11026 40409 11038 40412
rect 11072 40409 11084 40443
rect 12774 40443 12832 40449
rect 12774 40440 12786 40443
rect 11026 40403 11084 40409
rect 12406 40412 12786 40440
rect 10505 40375 10563 40381
rect 10505 40341 10517 40375
rect 10551 40341 10563 40375
rect 10505 40335 10563 40341
rect 12253 40375 12311 40381
rect 12253 40341 12265 40375
rect 12299 40372 12311 40375
rect 12406 40372 12434 40412
rect 12774 40409 12786 40412
rect 12820 40409 12832 40443
rect 12774 40403 12832 40409
rect 15470 40400 15476 40452
rect 15528 40440 15534 40452
rect 15657 40443 15715 40449
rect 15657 40440 15669 40443
rect 15528 40412 15669 40440
rect 15528 40400 15534 40412
rect 15657 40409 15669 40412
rect 15703 40409 15715 40443
rect 16316 40440 16344 40471
rect 16574 40468 16580 40471
rect 16632 40468 16638 40520
rect 18800 40517 18828 40616
rect 22480 40588 22508 40616
rect 37826 40604 37832 40616
rect 37884 40604 37890 40656
rect 38838 40604 38844 40656
rect 38896 40604 38902 40656
rect 20438 40536 20444 40588
rect 20496 40576 20502 40588
rect 20717 40579 20775 40585
rect 20717 40576 20729 40579
rect 20496 40548 20729 40576
rect 20496 40536 20502 40548
rect 20717 40545 20729 40548
rect 20763 40576 20775 40579
rect 20763 40548 21772 40576
rect 20763 40545 20775 40548
rect 20717 40539 20775 40545
rect 18785 40511 18843 40517
rect 18785 40477 18797 40511
rect 18831 40477 18843 40511
rect 18785 40471 18843 40477
rect 20533 40511 20591 40517
rect 20533 40477 20545 40511
rect 20579 40508 20591 40511
rect 21634 40508 21640 40520
rect 20579 40480 21640 40508
rect 20579 40477 20591 40480
rect 20533 40471 20591 40477
rect 21634 40468 21640 40480
rect 21692 40468 21698 40520
rect 17034 40440 17040 40452
rect 16316 40412 17040 40440
rect 15657 40403 15715 40409
rect 17034 40400 17040 40412
rect 17092 40440 17098 40452
rect 19058 40440 19064 40452
rect 17092 40412 19064 40440
rect 17092 40400 17098 40412
rect 19058 40400 19064 40412
rect 19116 40400 19122 40452
rect 21744 40440 21772 40548
rect 22462 40536 22468 40588
rect 22520 40536 22526 40588
rect 24302 40536 24308 40588
rect 24360 40576 24366 40588
rect 24765 40579 24823 40585
rect 24765 40576 24777 40579
rect 24360 40548 24777 40576
rect 24360 40536 24366 40548
rect 24765 40545 24777 40548
rect 24811 40545 24823 40579
rect 35115 40579 35173 40585
rect 24765 40539 24823 40545
rect 27356 40548 27568 40576
rect 22002 40468 22008 40520
rect 22060 40508 22066 40520
rect 22189 40511 22247 40517
rect 22189 40508 22201 40511
rect 22060 40480 22201 40508
rect 22060 40468 22066 40480
rect 22189 40477 22201 40480
rect 22235 40477 22247 40511
rect 22189 40471 22247 40477
rect 22649 40511 22707 40517
rect 22649 40477 22661 40511
rect 22695 40477 22707 40511
rect 24489 40511 24547 40517
rect 24489 40508 24501 40511
rect 23759 40484 24501 40508
rect 22649 40471 22707 40477
rect 23676 40480 24501 40484
rect 22554 40440 22560 40452
rect 21744 40412 22560 40440
rect 22554 40400 22560 40412
rect 22612 40400 22618 40452
rect 12299 40344 12434 40372
rect 12299 40341 12311 40344
rect 12253 40335 12311 40341
rect 13538 40332 13544 40384
rect 13596 40372 13602 40384
rect 13909 40375 13967 40381
rect 13909 40372 13921 40375
rect 13596 40344 13921 40372
rect 13596 40332 13602 40344
rect 13909 40341 13921 40344
rect 13955 40341 13967 40375
rect 13909 40335 13967 40341
rect 15194 40332 15200 40384
rect 15252 40332 15258 40384
rect 15378 40332 15384 40384
rect 15436 40372 15442 40384
rect 15565 40375 15623 40381
rect 15565 40372 15577 40375
rect 15436 40344 15577 40372
rect 15436 40332 15442 40344
rect 15565 40341 15577 40344
rect 15611 40341 15623 40375
rect 15565 40335 15623 40341
rect 17678 40332 17684 40384
rect 17736 40332 17742 40384
rect 17770 40332 17776 40384
rect 17828 40372 17834 40384
rect 18141 40375 18199 40381
rect 18141 40372 18153 40375
rect 17828 40344 18153 40372
rect 17828 40332 17834 40344
rect 18141 40341 18153 40344
rect 18187 40341 18199 40375
rect 18141 40335 18199 40341
rect 18598 40332 18604 40384
rect 18656 40332 18662 40384
rect 20622 40332 20628 40384
rect 20680 40332 20686 40384
rect 22278 40332 22284 40384
rect 22336 40332 22342 40384
rect 22664 40372 22692 40471
rect 23676 40456 23787 40480
rect 24489 40477 24501 40480
rect 24535 40508 24547 40511
rect 25685 40511 25743 40517
rect 25685 40508 25697 40511
rect 24535 40480 25697 40508
rect 24535 40477 24547 40480
rect 24489 40471 24547 40477
rect 25685 40477 25697 40480
rect 25731 40508 25743 40511
rect 27246 40508 27252 40520
rect 25731 40480 27252 40508
rect 25731 40477 25743 40480
rect 25685 40471 25743 40477
rect 27246 40468 27252 40480
rect 27304 40468 27310 40520
rect 27356 40517 27384 40548
rect 27341 40511 27399 40517
rect 27341 40477 27353 40511
rect 27387 40477 27399 40511
rect 27341 40471 27399 40477
rect 27430 40468 27436 40520
rect 27488 40468 27494 40520
rect 27540 40508 27568 40548
rect 35115 40545 35127 40579
rect 35161 40576 35173 40579
rect 36354 40576 36360 40588
rect 35161 40548 36360 40576
rect 35161 40545 35173 40548
rect 35115 40539 35173 40545
rect 36354 40536 36360 40548
rect 36412 40536 36418 40588
rect 36538 40536 36544 40588
rect 36596 40536 36602 40588
rect 40126 40536 40132 40588
rect 40184 40536 40190 40588
rect 29089 40511 29147 40517
rect 27540 40480 27844 40508
rect 22916 40443 22974 40449
rect 22916 40409 22928 40443
rect 22962 40440 22974 40443
rect 23014 40440 23020 40452
rect 22962 40412 23020 40440
rect 22962 40409 22974 40412
rect 22916 40403 22974 40409
rect 23014 40400 23020 40412
rect 23072 40400 23078 40452
rect 23676 40440 23704 40456
rect 23115 40412 23704 40440
rect 25952 40443 26010 40449
rect 23115 40372 23143 40412
rect 25952 40409 25964 40443
rect 25998 40440 26010 40443
rect 26234 40440 26240 40452
rect 25998 40412 26240 40440
rect 25998 40409 26010 40412
rect 25952 40403 26010 40409
rect 26234 40400 26240 40412
rect 26292 40400 26298 40452
rect 27678 40443 27736 40449
rect 27678 40440 27690 40443
rect 27172 40412 27690 40440
rect 22664 40344 23143 40372
rect 23566 40332 23572 40384
rect 23624 40372 23630 40384
rect 24029 40375 24087 40381
rect 24029 40372 24041 40375
rect 23624 40344 24041 40372
rect 23624 40332 23630 40344
rect 24029 40341 24041 40344
rect 24075 40341 24087 40375
rect 24029 40335 24087 40341
rect 27062 40332 27068 40384
rect 27120 40332 27126 40384
rect 27172 40381 27200 40412
rect 27678 40409 27690 40412
rect 27724 40409 27736 40443
rect 27816 40440 27844 40480
rect 29089 40477 29101 40511
rect 29135 40508 29147 40511
rect 29362 40508 29368 40520
rect 29135 40480 29368 40508
rect 29135 40477 29147 40480
rect 29089 40471 29147 40477
rect 29362 40468 29368 40480
rect 29420 40468 29426 40520
rect 30193 40511 30251 40517
rect 30193 40477 30205 40511
rect 30239 40508 30251 40511
rect 30926 40508 30932 40520
rect 30239 40480 30932 40508
rect 30239 40477 30251 40480
rect 30193 40471 30251 40477
rect 30926 40468 30932 40480
rect 30984 40468 30990 40520
rect 32953 40511 33011 40517
rect 32953 40477 32965 40511
rect 32999 40508 33011 40511
rect 33042 40508 33048 40520
rect 32999 40480 33048 40508
rect 32999 40477 33011 40480
rect 32953 40471 33011 40477
rect 33042 40468 33048 40480
rect 33100 40468 33106 40520
rect 34882 40468 34888 40520
rect 34940 40508 34946 40520
rect 34977 40511 35035 40517
rect 34977 40508 34989 40511
rect 34940 40480 34989 40508
rect 34940 40468 34946 40480
rect 34977 40477 34989 40480
rect 35023 40477 35035 40511
rect 34977 40471 35035 40477
rect 35342 40468 35348 40520
rect 35400 40508 35406 40520
rect 35529 40511 35587 40517
rect 35529 40508 35541 40511
rect 35400 40480 35541 40508
rect 35400 40468 35406 40480
rect 35529 40477 35541 40480
rect 35575 40477 35587 40511
rect 35529 40471 35587 40477
rect 35802 40468 35808 40520
rect 35860 40508 35866 40520
rect 36722 40508 36728 40520
rect 35860 40480 36728 40508
rect 35860 40468 35866 40480
rect 36722 40468 36728 40480
rect 36780 40468 36786 40520
rect 36814 40468 36820 40520
rect 36872 40508 36878 40520
rect 36909 40511 36967 40517
rect 36909 40508 36921 40511
rect 36872 40480 36921 40508
rect 36872 40468 36878 40480
rect 36909 40477 36921 40480
rect 36955 40477 36967 40511
rect 36909 40471 36967 40477
rect 37182 40468 37188 40520
rect 37240 40508 37246 40520
rect 37645 40511 37703 40517
rect 37645 40508 37657 40511
rect 37240 40480 37657 40508
rect 37240 40468 37246 40480
rect 37645 40477 37657 40480
rect 37691 40477 37703 40511
rect 37645 40471 37703 40477
rect 37921 40511 37979 40517
rect 37921 40477 37933 40511
rect 37967 40508 37979 40511
rect 38010 40508 38016 40520
rect 37967 40480 38016 40508
rect 37967 40477 37979 40480
rect 37921 40471 37979 40477
rect 38010 40468 38016 40480
rect 38068 40468 38074 40520
rect 38105 40511 38163 40517
rect 38105 40477 38117 40511
rect 38151 40508 38163 40511
rect 38654 40508 38660 40520
rect 38151 40480 38660 40508
rect 38151 40477 38163 40480
rect 38105 40471 38163 40477
rect 38654 40468 38660 40480
rect 38712 40468 38718 40520
rect 39206 40508 39212 40520
rect 38780 40480 39212 40508
rect 27890 40440 27896 40452
rect 27816 40412 27896 40440
rect 27678 40403 27736 40409
rect 27890 40400 27896 40412
rect 27948 40400 27954 40452
rect 30460 40443 30518 40449
rect 30460 40409 30472 40443
rect 30506 40440 30518 40443
rect 30558 40440 30564 40452
rect 30506 40412 30564 40440
rect 30506 40409 30518 40412
rect 30460 40403 30518 40409
rect 30558 40400 30564 40412
rect 30616 40400 30622 40452
rect 33220 40443 33278 40449
rect 33220 40409 33232 40443
rect 33266 40440 33278 40443
rect 34054 40440 34060 40452
rect 33266 40412 34060 40440
rect 33266 40409 33278 40412
rect 33220 40403 33278 40409
rect 34054 40400 34060 40412
rect 34112 40400 34118 40452
rect 36262 40400 36268 40452
rect 36320 40440 36326 40452
rect 38780 40440 38808 40480
rect 39206 40468 39212 40480
rect 39264 40508 39270 40520
rect 39853 40511 39911 40517
rect 39853 40508 39865 40511
rect 39264 40480 39865 40508
rect 39264 40468 39270 40480
rect 39853 40477 39865 40480
rect 39899 40477 39911 40511
rect 39853 40471 39911 40477
rect 45554 40468 45560 40520
rect 45612 40508 45618 40520
rect 46477 40511 46535 40517
rect 46477 40508 46489 40511
rect 45612 40480 46489 40508
rect 45612 40468 45618 40480
rect 46477 40477 46489 40480
rect 46523 40477 46535 40511
rect 46477 40471 46535 40477
rect 36320 40412 38808 40440
rect 38841 40443 38899 40449
rect 36320 40400 36326 40412
rect 38841 40409 38853 40443
rect 38887 40440 38899 40443
rect 38930 40440 38936 40452
rect 38887 40412 38936 40440
rect 38887 40409 38899 40412
rect 38841 40403 38899 40409
rect 38930 40400 38936 40412
rect 38988 40400 38994 40452
rect 39301 40443 39359 40449
rect 39301 40409 39313 40443
rect 39347 40440 39359 40443
rect 39347 40412 39896 40440
rect 39347 40409 39359 40412
rect 39301 40403 39359 40409
rect 39868 40384 39896 40412
rect 27157 40375 27215 40381
rect 27157 40341 27169 40375
rect 27203 40341 27215 40375
rect 27157 40335 27215 40341
rect 28258 40332 28264 40384
rect 28316 40372 28322 40384
rect 28813 40375 28871 40381
rect 28813 40372 28825 40375
rect 28316 40344 28825 40372
rect 28316 40332 28322 40344
rect 28813 40341 28825 40344
rect 28859 40341 28871 40375
rect 28813 40335 28871 40341
rect 28902 40332 28908 40384
rect 28960 40332 28966 40384
rect 31573 40375 31631 40381
rect 31573 40341 31585 40375
rect 31619 40372 31631 40375
rect 31754 40372 31760 40384
rect 31619 40344 31760 40372
rect 31619 40341 31631 40344
rect 31573 40335 31631 40341
rect 31754 40332 31760 40344
rect 31812 40332 31818 40384
rect 33594 40332 33600 40384
rect 33652 40372 33658 40384
rect 34333 40375 34391 40381
rect 34333 40372 34345 40375
rect 33652 40344 34345 40372
rect 33652 40332 33658 40344
rect 34333 40341 34345 40344
rect 34379 40341 34391 40375
rect 34333 40335 34391 40341
rect 34790 40332 34796 40384
rect 34848 40372 34854 40384
rect 34977 40375 35035 40381
rect 34977 40372 34989 40375
rect 34848 40344 34989 40372
rect 34848 40332 34854 40344
rect 34977 40341 34989 40344
rect 35023 40341 35035 40375
rect 34977 40335 35035 40341
rect 36354 40332 36360 40384
rect 36412 40372 36418 40384
rect 36725 40375 36783 40381
rect 36725 40372 36737 40375
rect 36412 40344 36737 40372
rect 36412 40332 36418 40344
rect 36725 40341 36737 40344
rect 36771 40341 36783 40375
rect 36725 40335 36783 40341
rect 36906 40332 36912 40384
rect 36964 40372 36970 40384
rect 37090 40372 37096 40384
rect 36964 40344 37096 40372
rect 36964 40332 36970 40344
rect 37090 40332 37096 40344
rect 37148 40332 37154 40384
rect 37458 40332 37464 40384
rect 37516 40332 37522 40384
rect 39390 40332 39396 40384
rect 39448 40332 39454 40384
rect 39574 40332 39580 40384
rect 39632 40332 39638 40384
rect 39850 40332 39856 40384
rect 39908 40332 39914 40384
rect 40402 40332 40408 40384
rect 40460 40332 40466 40384
rect 46658 40332 46664 40384
rect 46716 40332 46722 40384
rect 1104 40282 47104 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 35594 40282
rect 35646 40230 35658 40282
rect 35710 40230 35722 40282
rect 35774 40230 35786 40282
rect 35838 40230 35850 40282
rect 35902 40230 47104 40282
rect 1104 40208 47104 40230
rect 2038 40128 2044 40180
rect 2096 40168 2102 40180
rect 2225 40171 2283 40177
rect 2225 40168 2237 40171
rect 2096 40140 2237 40168
rect 2096 40128 2102 40140
rect 2225 40137 2237 40140
rect 2271 40137 2283 40171
rect 2225 40131 2283 40137
rect 2590 40128 2596 40180
rect 2648 40128 2654 40180
rect 8846 40128 8852 40180
rect 8904 40128 8910 40180
rect 9677 40171 9735 40177
rect 9677 40137 9689 40171
rect 9723 40137 9735 40171
rect 9677 40131 9735 40137
rect 11149 40171 11207 40177
rect 11149 40137 11161 40171
rect 11195 40137 11207 40171
rect 11149 40131 11207 40137
rect 9692 40100 9720 40131
rect 9048 40072 9720 40100
rect 1397 40035 1455 40041
rect 1397 40001 1409 40035
rect 1443 40032 1455 40035
rect 2038 40032 2044 40044
rect 1443 40004 2044 40032
rect 1443 40001 1455 40004
rect 1397 39995 1455 40001
rect 2038 39992 2044 40004
rect 2096 39992 2102 40044
rect 9048 40041 9076 40072
rect 10042 40060 10048 40112
rect 10100 40060 10106 40112
rect 11164 40100 11192 40131
rect 12434 40128 12440 40180
rect 12492 40168 12498 40180
rect 12897 40171 12955 40177
rect 12897 40168 12909 40171
rect 12492 40140 12909 40168
rect 12492 40128 12498 40140
rect 12897 40137 12909 40140
rect 12943 40137 12955 40171
rect 12897 40131 12955 40137
rect 13170 40128 13176 40180
rect 13228 40128 13234 40180
rect 13538 40128 13544 40180
rect 13596 40128 13602 40180
rect 14458 40128 14464 40180
rect 14516 40168 14522 40180
rect 14645 40171 14703 40177
rect 14645 40168 14657 40171
rect 14516 40140 14657 40168
rect 14516 40128 14522 40140
rect 14645 40137 14657 40140
rect 14691 40137 14703 40171
rect 14645 40131 14703 40137
rect 16942 40128 16948 40180
rect 17000 40168 17006 40180
rect 17313 40171 17371 40177
rect 17313 40168 17325 40171
rect 17000 40140 17325 40168
rect 17000 40128 17006 40140
rect 17313 40137 17325 40140
rect 17359 40137 17371 40171
rect 17313 40131 17371 40137
rect 17678 40128 17684 40180
rect 17736 40128 17742 40180
rect 23014 40128 23020 40180
rect 23072 40128 23078 40180
rect 24026 40128 24032 40180
rect 24084 40128 24090 40180
rect 24394 40128 24400 40180
rect 24452 40168 24458 40180
rect 24857 40171 24915 40177
rect 24857 40168 24869 40171
rect 24452 40140 24869 40168
rect 24452 40128 24458 40140
rect 24857 40137 24869 40140
rect 24903 40137 24915 40171
rect 24857 40131 24915 40137
rect 24946 40128 24952 40180
rect 25004 40168 25010 40180
rect 25317 40171 25375 40177
rect 25317 40168 25329 40171
rect 25004 40140 25329 40168
rect 25004 40128 25010 40140
rect 25317 40137 25329 40140
rect 25363 40168 25375 40171
rect 25866 40168 25872 40180
rect 25363 40140 25872 40168
rect 25363 40137 25375 40140
rect 25317 40131 25375 40137
rect 25866 40128 25872 40140
rect 25924 40128 25930 40180
rect 26234 40128 26240 40180
rect 26292 40128 26298 40180
rect 26878 40168 26884 40180
rect 26344 40140 26884 40168
rect 11762 40103 11820 40109
rect 11762 40100 11774 40103
rect 11164 40072 11774 40100
rect 11762 40069 11774 40072
rect 11808 40069 11820 40103
rect 11762 40063 11820 40069
rect 11882 40060 11888 40112
rect 11940 40100 11946 40112
rect 13556 40100 13584 40128
rect 15194 40100 15200 40112
rect 11940 40072 13584 40100
rect 14844 40072 15200 40100
rect 11940 40060 11946 40072
rect 9033 40035 9091 40041
rect 9033 40001 9045 40035
rect 9079 40001 9091 40035
rect 9033 39995 9091 40001
rect 10137 40035 10195 40041
rect 10137 40001 10149 40035
rect 10183 40032 10195 40035
rect 10410 40032 10416 40044
rect 10183 40004 10416 40032
rect 10183 40001 10195 40004
rect 10137 39995 10195 40001
rect 10410 39992 10416 40004
rect 10468 40032 10474 40044
rect 10594 40032 10600 40044
rect 10468 40004 10600 40032
rect 10468 39992 10474 40004
rect 10594 39992 10600 40004
rect 10652 39992 10658 40044
rect 11330 39992 11336 40044
rect 11388 39992 11394 40044
rect 11514 39992 11520 40044
rect 11572 39992 11578 40044
rect 14844 40041 14872 40072
rect 15194 40060 15200 40072
rect 15252 40060 15258 40112
rect 22278 40060 22284 40112
rect 22336 40100 22342 40112
rect 24486 40100 24492 40112
rect 22336 40072 24348 40100
rect 22336 40060 22342 40072
rect 14829 40035 14887 40041
rect 11624 40004 14780 40032
rect 2682 39924 2688 39976
rect 2740 39924 2746 39976
rect 2869 39967 2927 39973
rect 2869 39933 2881 39967
rect 2915 39933 2927 39967
rect 2869 39927 2927 39933
rect 2884 39896 2912 39927
rect 10226 39924 10232 39976
rect 10284 39924 10290 39976
rect 11624 39964 11652 40004
rect 10336 39936 11652 39964
rect 3142 39896 3148 39908
rect 2884 39868 3148 39896
rect 3142 39856 3148 39868
rect 3200 39896 3206 39908
rect 10336 39896 10364 39936
rect 13630 39924 13636 39976
rect 13688 39924 13694 39976
rect 13817 39967 13875 39973
rect 13817 39933 13829 39967
rect 13863 39933 13875 39967
rect 14752 39964 14780 40004
rect 14829 40001 14841 40035
rect 14875 40001 14887 40035
rect 20438 40032 20444 40044
rect 14829 39995 14887 40001
rect 17696 40004 20444 40032
rect 17696 39964 17724 40004
rect 20438 39992 20444 40004
rect 20496 39992 20502 40044
rect 23198 39992 23204 40044
rect 23256 39992 23262 40044
rect 14752 39936 17724 39964
rect 13817 39927 13875 39933
rect 3200 39868 10364 39896
rect 13832 39896 13860 39927
rect 17770 39924 17776 39976
rect 17828 39924 17834 39976
rect 17865 39967 17923 39973
rect 17865 39933 17877 39967
rect 17911 39964 17923 39967
rect 24320 39964 24348 40072
rect 24412 40072 24492 40100
rect 24412 40041 24440 40072
rect 24486 40060 24492 40072
rect 24544 40060 24550 40112
rect 24670 40060 24676 40112
rect 24728 40100 24734 40112
rect 26344 40100 26372 40140
rect 26878 40128 26884 40140
rect 26936 40128 26942 40180
rect 26973 40171 27031 40177
rect 26973 40137 26985 40171
rect 27019 40137 27031 40171
rect 26973 40131 27031 40137
rect 26988 40100 27016 40131
rect 27062 40128 27068 40180
rect 27120 40168 27126 40180
rect 27341 40171 27399 40177
rect 27341 40168 27353 40171
rect 27120 40140 27353 40168
rect 27120 40128 27126 40140
rect 27341 40137 27353 40140
rect 27387 40137 27399 40171
rect 27341 40131 27399 40137
rect 29362 40128 29368 40180
rect 29420 40128 29426 40180
rect 30558 40128 30564 40180
rect 30616 40128 30622 40180
rect 30837 40171 30895 40177
rect 30837 40137 30849 40171
rect 30883 40137 30895 40171
rect 30837 40131 30895 40137
rect 31205 40171 31263 40177
rect 31205 40137 31217 40171
rect 31251 40168 31263 40171
rect 31754 40168 31760 40180
rect 31251 40140 31760 40168
rect 31251 40137 31263 40140
rect 31205 40131 31263 40137
rect 24728 40072 26372 40100
rect 26436 40072 27016 40100
rect 24728 40060 24734 40072
rect 26436 40041 26464 40072
rect 27430 40060 27436 40112
rect 27488 40100 27494 40112
rect 28160 40103 28218 40109
rect 27488 40072 27936 40100
rect 27488 40060 27494 40072
rect 27908 40041 27936 40072
rect 28160 40069 28172 40103
rect 28206 40100 28218 40103
rect 28902 40100 28908 40112
rect 28206 40072 28908 40100
rect 28206 40069 28218 40072
rect 28160 40063 28218 40069
rect 28902 40060 28908 40072
rect 28960 40060 28966 40112
rect 30852 40100 30880 40131
rect 31754 40128 31760 40140
rect 31812 40168 31818 40180
rect 32766 40168 32772 40180
rect 31812 40140 32772 40168
rect 31812 40128 31818 40140
rect 32766 40128 32772 40140
rect 32824 40128 32830 40180
rect 34054 40128 34060 40180
rect 34112 40128 34118 40180
rect 36909 40171 36967 40177
rect 36909 40137 36921 40171
rect 36955 40168 36967 40171
rect 37550 40168 37556 40180
rect 36955 40140 37556 40168
rect 36955 40137 36967 40140
rect 36909 40131 36967 40137
rect 37550 40128 37556 40140
rect 37608 40128 37614 40180
rect 38473 40171 38531 40177
rect 38473 40137 38485 40171
rect 38519 40168 38531 40171
rect 38654 40168 38660 40180
rect 38519 40140 38660 40168
rect 38519 40137 38531 40140
rect 38473 40131 38531 40137
rect 38654 40128 38660 40140
rect 38712 40128 38718 40180
rect 39390 40168 39396 40180
rect 38764 40140 39396 40168
rect 30760 40072 30880 40100
rect 24397 40035 24455 40041
rect 24397 40001 24409 40035
rect 24443 40001 24455 40035
rect 25225 40035 25283 40041
rect 25225 40032 25237 40035
rect 24397 39995 24455 40001
rect 24504 40004 25237 40032
rect 24504 39973 24532 40004
rect 25225 40001 25237 40004
rect 25271 40001 25283 40035
rect 25225 39995 25283 40001
rect 26421 40035 26479 40041
rect 26421 40001 26433 40035
rect 26467 40001 26479 40035
rect 26421 39995 26479 40001
rect 27893 40035 27951 40041
rect 27893 40001 27905 40035
rect 27939 40032 27951 40035
rect 28442 40032 28448 40044
rect 27939 40004 28448 40032
rect 27939 40001 27951 40004
rect 27893 39995 27951 40001
rect 24489 39967 24547 39973
rect 24489 39964 24501 39967
rect 17911 39936 22094 39964
rect 24320 39936 24501 39964
rect 17911 39933 17923 39936
rect 17865 39927 17923 39933
rect 15010 39896 15016 39908
rect 13832 39868 15016 39896
rect 3200 39856 3206 39868
rect 15010 39856 15016 39868
rect 15068 39856 15074 39908
rect 15470 39856 15476 39908
rect 15528 39896 15534 39908
rect 17788 39896 17816 39924
rect 15528 39868 17816 39896
rect 22066 39896 22094 39936
rect 24489 39933 24501 39936
rect 24535 39933 24547 39967
rect 24489 39927 24547 39933
rect 24673 39967 24731 39973
rect 24673 39933 24685 39967
rect 24719 39964 24731 39967
rect 24762 39964 24768 39976
rect 24719 39936 24768 39964
rect 24719 39933 24731 39936
rect 24673 39927 24731 39933
rect 24688 39896 24716 39927
rect 24762 39924 24768 39936
rect 24820 39924 24826 39976
rect 22066 39868 24716 39896
rect 15528 39856 15534 39868
rect 934 39788 940 39840
rect 992 39828 998 39840
rect 1581 39831 1639 39837
rect 1581 39828 1593 39831
rect 992 39800 1593 39828
rect 992 39788 998 39800
rect 1581 39797 1593 39800
rect 1627 39797 1639 39831
rect 1581 39791 1639 39797
rect 2038 39788 2044 39840
rect 2096 39788 2102 39840
rect 6914 39788 6920 39840
rect 6972 39828 6978 39840
rect 7285 39831 7343 39837
rect 7285 39828 7297 39831
rect 6972 39800 7297 39828
rect 6972 39788 6978 39800
rect 7285 39797 7297 39800
rect 7331 39828 7343 39831
rect 7653 39831 7711 39837
rect 7653 39828 7665 39831
rect 7331 39800 7665 39828
rect 7331 39797 7343 39800
rect 7285 39791 7343 39797
rect 7653 39797 7665 39800
rect 7699 39828 7711 39831
rect 8021 39831 8079 39837
rect 8021 39828 8033 39831
rect 7699 39800 8033 39828
rect 7699 39797 7711 39800
rect 7653 39791 7711 39797
rect 8021 39797 8033 39800
rect 8067 39828 8079 39831
rect 8389 39831 8447 39837
rect 8389 39828 8401 39831
rect 8067 39800 8401 39828
rect 8067 39797 8079 39800
rect 8021 39791 8079 39797
rect 8389 39797 8401 39800
rect 8435 39828 8447 39831
rect 8757 39831 8815 39837
rect 8757 39828 8769 39831
rect 8435 39800 8769 39828
rect 8435 39797 8447 39800
rect 8389 39791 8447 39797
rect 8757 39797 8769 39800
rect 8803 39828 8815 39831
rect 9030 39828 9036 39840
rect 8803 39800 9036 39828
rect 8803 39797 8815 39800
rect 8757 39791 8815 39797
rect 9030 39788 9036 39800
rect 9088 39828 9094 39840
rect 9309 39831 9367 39837
rect 9309 39828 9321 39831
rect 9088 39800 9321 39828
rect 9088 39788 9094 39800
rect 9309 39797 9321 39800
rect 9355 39828 9367 39831
rect 10042 39828 10048 39840
rect 9355 39800 10048 39828
rect 9355 39797 9367 39800
rect 9309 39791 9367 39797
rect 10042 39788 10048 39800
rect 10100 39788 10106 39840
rect 10226 39788 10232 39840
rect 10284 39828 10290 39840
rect 17770 39828 17776 39840
rect 10284 39800 17776 39828
rect 10284 39788 10290 39800
rect 17770 39788 17776 39800
rect 17828 39788 17834 39840
rect 25240 39828 25268 39995
rect 28442 39992 28448 40004
rect 28500 39992 28506 40044
rect 29730 39992 29736 40044
rect 29788 39992 29794 40044
rect 30760 40041 30788 40072
rect 33134 40060 33140 40112
rect 33192 40100 33198 40112
rect 33192 40072 33456 40100
rect 33192 40060 33198 40072
rect 33428 40044 33456 40072
rect 33686 40060 33692 40112
rect 33744 40060 33750 40112
rect 33778 40060 33784 40112
rect 33836 40100 33842 40112
rect 34422 40100 34428 40112
rect 33836 40072 34428 40100
rect 33836 40060 33842 40072
rect 34422 40060 34428 40072
rect 34480 40100 34486 40112
rect 34790 40100 34796 40112
rect 34480 40072 34796 40100
rect 34480 40060 34486 40072
rect 34790 40060 34796 40072
rect 34848 40060 34854 40112
rect 34882 40060 34888 40112
rect 34940 40100 34946 40112
rect 35529 40103 35587 40109
rect 35529 40100 35541 40103
rect 34940 40072 35541 40100
rect 34940 40060 34946 40072
rect 35529 40069 35541 40072
rect 35575 40069 35587 40103
rect 35529 40063 35587 40069
rect 35713 40103 35771 40109
rect 35713 40069 35725 40103
rect 35759 40100 35771 40103
rect 35986 40100 35992 40112
rect 35759 40072 35992 40100
rect 35759 40069 35771 40072
rect 35713 40063 35771 40069
rect 35986 40060 35992 40072
rect 36044 40060 36050 40112
rect 37369 40103 37427 40109
rect 36096 40072 36308 40100
rect 30745 40035 30803 40041
rect 30745 40001 30757 40035
rect 30791 40001 30803 40035
rect 30745 39995 30803 40001
rect 33410 39992 33416 40044
rect 33468 39992 33474 40044
rect 33594 40041 33600 40044
rect 33561 40035 33600 40041
rect 33561 40001 33573 40035
rect 33561 39995 33600 40001
rect 33594 39992 33600 39995
rect 33652 39992 33658 40044
rect 33919 40035 33977 40041
rect 33919 40001 33931 40035
rect 33965 40032 33977 40035
rect 33965 40004 34100 40032
rect 33965 40001 33977 40004
rect 33919 39995 33977 40001
rect 25501 39967 25559 39973
rect 25501 39933 25513 39967
rect 25547 39964 25559 39967
rect 26234 39964 26240 39976
rect 25547 39936 26240 39964
rect 25547 39933 25559 39936
rect 25501 39927 25559 39933
rect 26234 39924 26240 39936
rect 26292 39924 26298 39976
rect 27430 39924 27436 39976
rect 27488 39924 27494 39976
rect 27522 39924 27528 39976
rect 27580 39924 27586 39976
rect 29825 39967 29883 39973
rect 29825 39964 29837 39967
rect 29288 39936 29837 39964
rect 28994 39856 29000 39908
rect 29052 39896 29058 39908
rect 29288 39905 29316 39936
rect 29825 39933 29837 39936
rect 29871 39933 29883 39967
rect 29825 39927 29883 39933
rect 30006 39924 30012 39976
rect 30064 39924 30070 39976
rect 31297 39967 31355 39973
rect 31297 39933 31309 39967
rect 31343 39933 31355 39967
rect 31297 39927 31355 39933
rect 29273 39899 29331 39905
rect 29273 39896 29285 39899
rect 29052 39868 29285 39896
rect 29052 39856 29058 39868
rect 29273 39865 29285 39868
rect 29319 39865 29331 39899
rect 29273 39859 29331 39865
rect 31312 39840 31340 39927
rect 31386 39924 31392 39976
rect 31444 39924 31450 39976
rect 34072 39964 34100 40004
rect 35250 39992 35256 40044
rect 35308 40032 35314 40044
rect 36096 40032 36124 40072
rect 35308 40004 36124 40032
rect 36173 40035 36231 40041
rect 35308 39992 35314 40004
rect 36173 40001 36185 40035
rect 36219 40001 36231 40035
rect 36173 39995 36231 40001
rect 34146 39964 34152 39976
rect 34072 39936 34152 39964
rect 34146 39924 34152 39936
rect 34204 39964 34210 39976
rect 34422 39964 34428 39976
rect 34204 39936 34428 39964
rect 34204 39924 34210 39936
rect 34422 39924 34428 39936
rect 34480 39924 34486 39976
rect 34790 39924 34796 39976
rect 34848 39964 34854 39976
rect 35268 39964 35296 39992
rect 34848 39936 35296 39964
rect 34848 39924 34854 39936
rect 35434 39924 35440 39976
rect 35492 39964 35498 39976
rect 35897 39967 35955 39973
rect 35897 39964 35909 39967
rect 35492 39936 35909 39964
rect 35492 39924 35498 39936
rect 35897 39933 35909 39936
rect 35943 39964 35955 39967
rect 36188 39964 36216 39995
rect 35943 39936 36216 39964
rect 36280 39964 36308 40072
rect 37369 40069 37381 40103
rect 37415 40100 37427 40103
rect 37458 40100 37464 40112
rect 37415 40072 37464 40100
rect 37415 40069 37427 40072
rect 37369 40063 37427 40069
rect 37458 40060 37464 40072
rect 37516 40060 37522 40112
rect 36354 39992 36360 40044
rect 36412 40032 36418 40044
rect 36449 40035 36507 40041
rect 36449 40032 36461 40035
rect 36412 40004 36461 40032
rect 36412 39992 36418 40004
rect 36449 40001 36461 40004
rect 36495 40001 36507 40035
rect 36449 39995 36507 40001
rect 36722 39992 36728 40044
rect 36780 39992 36786 40044
rect 38764 40041 38792 40140
rect 39390 40128 39396 40140
rect 39448 40128 39454 40180
rect 38838 40060 38844 40112
rect 38896 40100 38902 40112
rect 40402 40100 40408 40112
rect 38896 40072 39068 40100
rect 38896 40060 38902 40072
rect 39040 40041 39068 40072
rect 39684 40072 40408 40100
rect 39684 40041 39712 40072
rect 40402 40060 40408 40072
rect 40460 40060 40466 40112
rect 38381 40035 38439 40041
rect 38381 40001 38393 40035
rect 38427 40001 38439 40035
rect 38381 39995 38439 40001
rect 38565 40035 38623 40041
rect 38565 40001 38577 40035
rect 38611 40001 38623 40035
rect 38565 39995 38623 40001
rect 38749 40035 38807 40041
rect 38749 40001 38761 40035
rect 38795 40001 38807 40035
rect 38749 39995 38807 40001
rect 39025 40035 39083 40041
rect 39025 40001 39037 40035
rect 39071 40001 39083 40035
rect 39025 39995 39083 40001
rect 39669 40035 39727 40041
rect 39669 40001 39681 40035
rect 39715 40001 39727 40035
rect 39669 39995 39727 40001
rect 36541 39967 36599 39973
rect 36541 39964 36553 39967
rect 36280 39936 36553 39964
rect 35943 39933 35955 39936
rect 35897 39927 35955 39933
rect 36541 39933 36553 39936
rect 36587 39964 36599 39967
rect 36906 39964 36912 39976
rect 36587 39936 36912 39964
rect 36587 39933 36599 39936
rect 36541 39927 36599 39933
rect 36906 39924 36912 39936
rect 36964 39924 36970 39976
rect 36265 39899 36323 39905
rect 36265 39865 36277 39899
rect 36311 39896 36323 39899
rect 37826 39896 37832 39908
rect 36311 39868 37832 39896
rect 36311 39865 36323 39868
rect 36265 39859 36323 39865
rect 37826 39856 37832 39868
rect 37884 39856 37890 39908
rect 38396 39896 38424 39995
rect 38580 39964 38608 39995
rect 39850 39992 39856 40044
rect 39908 40032 39914 40044
rect 40221 40035 40279 40041
rect 40221 40032 40233 40035
rect 39908 40004 40233 40032
rect 39908 39992 39914 40004
rect 40221 40001 40233 40004
rect 40267 40001 40279 40035
rect 40221 39995 40279 40001
rect 38930 39964 38936 39976
rect 38580 39936 38936 39964
rect 38930 39924 38936 39936
rect 38988 39964 38994 39976
rect 39574 39964 39580 39976
rect 38988 39936 39580 39964
rect 38988 39924 38994 39936
rect 39574 39924 39580 39936
rect 39632 39964 39638 39976
rect 39761 39967 39819 39973
rect 39761 39964 39773 39967
rect 39632 39936 39773 39964
rect 39632 39924 39638 39936
rect 39761 39933 39773 39936
rect 39807 39933 39819 39967
rect 39761 39927 39819 39933
rect 39850 39896 39856 39908
rect 38396 39868 39856 39896
rect 39850 39856 39856 39868
rect 39908 39856 39914 39908
rect 40129 39899 40187 39905
rect 40129 39865 40141 39899
rect 40175 39865 40187 39899
rect 40129 39859 40187 39865
rect 31294 39828 31300 39840
rect 25240 39800 31300 39828
rect 31294 39788 31300 39800
rect 31352 39788 31358 39840
rect 36725 39831 36783 39837
rect 36725 39797 36737 39831
rect 36771 39828 36783 39831
rect 37182 39828 37188 39840
rect 36771 39800 37188 39828
rect 36771 39797 36783 39800
rect 36725 39791 36783 39797
rect 37182 39788 37188 39800
rect 37240 39788 37246 39840
rect 37274 39788 37280 39840
rect 37332 39828 37338 39840
rect 37461 39831 37519 39837
rect 37461 39828 37473 39831
rect 37332 39800 37473 39828
rect 37332 39788 37338 39800
rect 37461 39797 37473 39800
rect 37507 39797 37519 39831
rect 37461 39791 37519 39797
rect 37642 39788 37648 39840
rect 37700 39828 37706 39840
rect 40144 39828 40172 39859
rect 37700 39800 40172 39828
rect 37700 39788 37706 39800
rect 1104 39738 47104 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 47104 39738
rect 1104 39664 47104 39686
rect 1486 39584 1492 39636
rect 1544 39624 1550 39636
rect 13078 39624 13084 39636
rect 1544 39596 13084 39624
rect 1544 39584 1550 39596
rect 13078 39584 13084 39596
rect 13136 39584 13142 39636
rect 13188 39596 19334 39624
rect 2038 39516 2044 39568
rect 2096 39556 2102 39568
rect 2409 39559 2467 39565
rect 2409 39556 2421 39559
rect 2096 39528 2421 39556
rect 2096 39516 2102 39528
rect 2409 39525 2421 39528
rect 2455 39556 2467 39559
rect 2455 39528 5764 39556
rect 2455 39525 2467 39528
rect 2409 39519 2467 39525
rect 2792 39497 2820 39528
rect 2777 39491 2835 39497
rect 2777 39457 2789 39491
rect 2823 39488 2835 39491
rect 5736 39488 5764 39528
rect 6914 39516 6920 39568
rect 6972 39516 6978 39568
rect 11330 39516 11336 39568
rect 11388 39556 11394 39568
rect 11793 39559 11851 39565
rect 11793 39556 11805 39559
rect 11388 39528 11805 39556
rect 11388 39516 11394 39528
rect 11793 39525 11805 39528
rect 11839 39525 11851 39559
rect 13188 39556 13216 39596
rect 11793 39519 11851 39525
rect 12268 39528 13216 39556
rect 19306 39556 19334 39596
rect 23198 39584 23204 39636
rect 23256 39584 23262 39636
rect 27890 39584 27896 39636
rect 27948 39584 27954 39636
rect 30006 39624 30012 39636
rect 28000 39596 30012 39624
rect 25682 39556 25688 39568
rect 19306 39528 25688 39556
rect 12268 39488 12296 39528
rect 25682 39516 25688 39528
rect 25740 39516 25746 39568
rect 26234 39516 26240 39568
rect 26292 39556 26298 39568
rect 28000 39556 28028 39596
rect 30006 39584 30012 39596
rect 30064 39584 30070 39636
rect 30834 39584 30840 39636
rect 30892 39624 30898 39636
rect 32401 39627 32459 39633
rect 32401 39624 32413 39627
rect 30892 39596 32413 39624
rect 30892 39584 30898 39596
rect 32401 39593 32413 39596
rect 32447 39593 32459 39627
rect 32401 39587 32459 39593
rect 36541 39627 36599 39633
rect 36541 39593 36553 39627
rect 36587 39624 36599 39627
rect 36587 39596 37412 39624
rect 36587 39593 36599 39596
rect 36541 39587 36599 39593
rect 29730 39556 29736 39568
rect 26292 39528 28028 39556
rect 28368 39528 29736 39556
rect 26292 39516 26298 39528
rect 2823 39460 2857 39488
rect 5736 39460 12296 39488
rect 12345 39491 12403 39497
rect 2823 39457 2835 39460
rect 2777 39451 2835 39457
rect 12345 39457 12357 39491
rect 12391 39457 12403 39491
rect 12345 39451 12403 39457
rect 12360 39420 12388 39451
rect 13078 39448 13084 39500
rect 13136 39488 13142 39500
rect 13136 39460 15516 39488
rect 13136 39448 13142 39460
rect 13170 39420 13176 39432
rect 12360 39392 13176 39420
rect 13170 39380 13176 39392
rect 13228 39380 13234 39432
rect 13998 39380 14004 39432
rect 14056 39420 14062 39432
rect 15381 39423 15439 39429
rect 15381 39420 15393 39423
rect 14056 39392 15393 39420
rect 14056 39380 14062 39392
rect 15381 39389 15393 39392
rect 15427 39389 15439 39423
rect 15488 39420 15516 39460
rect 17310 39448 17316 39500
rect 17368 39488 17374 39500
rect 23753 39491 23811 39497
rect 23753 39488 23765 39491
rect 17368 39460 23765 39488
rect 17368 39448 17374 39460
rect 23753 39457 23765 39460
rect 23799 39488 23811 39491
rect 26786 39488 26792 39500
rect 23799 39460 26792 39488
rect 23799 39457 23811 39460
rect 23753 39451 23811 39457
rect 26786 39448 26792 39460
rect 26844 39448 26850 39500
rect 27430 39448 27436 39500
rect 27488 39488 27494 39500
rect 28368 39497 28396 39528
rect 29730 39516 29736 39528
rect 29788 39516 29794 39568
rect 36446 39516 36452 39568
rect 36504 39556 36510 39568
rect 37093 39559 37151 39565
rect 37093 39556 37105 39559
rect 36504 39528 37105 39556
rect 36504 39516 36510 39528
rect 37093 39525 37105 39528
rect 37139 39556 37151 39559
rect 37182 39556 37188 39568
rect 37139 39528 37188 39556
rect 37139 39525 37151 39528
rect 37093 39519 37151 39525
rect 37182 39516 37188 39528
rect 37240 39516 37246 39568
rect 37384 39556 37412 39596
rect 37458 39584 37464 39636
rect 37516 39624 37522 39636
rect 38013 39627 38071 39633
rect 38013 39624 38025 39627
rect 37516 39596 38025 39624
rect 37516 39584 37522 39596
rect 38013 39593 38025 39596
rect 38059 39593 38071 39627
rect 38013 39587 38071 39593
rect 39669 39627 39727 39633
rect 39669 39593 39681 39627
rect 39715 39624 39727 39627
rect 39850 39624 39856 39636
rect 39715 39596 39856 39624
rect 39715 39593 39727 39596
rect 39669 39587 39727 39593
rect 39850 39584 39856 39596
rect 39908 39584 39914 39636
rect 37642 39556 37648 39568
rect 37384 39528 37648 39556
rect 37642 39516 37648 39528
rect 37700 39516 37706 39568
rect 28353 39491 28411 39497
rect 28353 39488 28365 39491
rect 27488 39460 28365 39488
rect 27488 39448 27494 39460
rect 28353 39457 28365 39460
rect 28399 39457 28411 39491
rect 28353 39451 28411 39457
rect 28537 39491 28595 39497
rect 28537 39457 28549 39491
rect 28583 39488 28595 39491
rect 29086 39488 29092 39500
rect 28583 39460 29092 39488
rect 28583 39457 28595 39460
rect 28537 39451 28595 39457
rect 29086 39448 29092 39460
rect 29144 39488 29150 39500
rect 30190 39488 30196 39500
rect 29144 39460 30196 39488
rect 29144 39448 29150 39460
rect 30190 39448 30196 39460
rect 30248 39448 30254 39500
rect 30926 39448 30932 39500
rect 30984 39448 30990 39500
rect 31938 39448 31944 39500
rect 31996 39488 32002 39500
rect 32953 39491 33011 39497
rect 32953 39488 32965 39491
rect 31996 39460 32965 39488
rect 31996 39448 32002 39460
rect 32953 39457 32965 39460
rect 32999 39457 33011 39491
rect 32953 39451 33011 39457
rect 36173 39491 36231 39497
rect 36173 39457 36185 39491
rect 36219 39488 36231 39491
rect 36219 39460 36584 39488
rect 36219 39457 36231 39460
rect 36173 39451 36231 39457
rect 36556 39432 36584 39460
rect 36906 39448 36912 39500
rect 36964 39488 36970 39500
rect 36964 39460 37044 39488
rect 36964 39448 36970 39460
rect 19702 39420 19708 39432
rect 15488 39392 19708 39420
rect 15381 39383 15439 39389
rect 19702 39380 19708 39392
rect 19760 39380 19766 39432
rect 23566 39380 23572 39432
rect 23624 39380 23630 39432
rect 27614 39380 27620 39432
rect 27672 39420 27678 39432
rect 28258 39420 28264 39432
rect 27672 39392 28264 39420
rect 27672 39380 27678 39392
rect 28258 39380 28264 39392
rect 28316 39380 28322 39432
rect 30742 39420 30748 39432
rect 28368 39392 30748 39420
rect 14734 39312 14740 39364
rect 14792 39312 14798 39364
rect 15648 39355 15706 39361
rect 15648 39321 15660 39355
rect 15694 39352 15706 39355
rect 17494 39352 17500 39364
rect 15694 39324 17500 39352
rect 15694 39321 15706 39324
rect 15648 39315 15706 39321
rect 17494 39312 17500 39324
rect 17552 39312 17558 39364
rect 27982 39312 27988 39364
rect 28040 39352 28046 39364
rect 28368 39352 28396 39392
rect 30742 39380 30748 39392
rect 30800 39380 30806 39432
rect 30834 39380 30840 39432
rect 30892 39380 30898 39432
rect 36354 39380 36360 39432
rect 36412 39380 36418 39432
rect 36538 39380 36544 39432
rect 36596 39380 36602 39432
rect 36630 39380 36636 39432
rect 36688 39420 36694 39432
rect 37016 39429 37044 39460
rect 38286 39448 38292 39500
rect 38344 39448 38350 39500
rect 36817 39423 36875 39429
rect 36817 39420 36829 39423
rect 36688 39392 36829 39420
rect 36688 39380 36694 39392
rect 36817 39389 36829 39392
rect 36863 39389 36875 39423
rect 36817 39383 36875 39389
rect 37001 39423 37059 39429
rect 37001 39389 37013 39423
rect 37047 39420 37059 39423
rect 37737 39423 37795 39429
rect 37737 39420 37749 39423
rect 37047 39392 37749 39420
rect 37047 39389 37059 39392
rect 37001 39383 37059 39389
rect 37737 39389 37749 39392
rect 37783 39420 37795 39423
rect 37918 39420 37924 39432
rect 37783 39392 37924 39420
rect 37783 39389 37795 39392
rect 37737 39383 37795 39389
rect 37918 39380 37924 39392
rect 37976 39380 37982 39432
rect 31174 39355 31232 39361
rect 31174 39352 31186 39355
rect 28040 39324 28396 39352
rect 30668 39324 31186 39352
rect 28040 39312 28046 39324
rect 9030 39244 9036 39296
rect 9088 39284 9094 39296
rect 9309 39287 9367 39293
rect 9309 39284 9321 39287
rect 9088 39256 9321 39284
rect 9088 39244 9094 39256
rect 9309 39253 9321 39256
rect 9355 39253 9367 39287
rect 9309 39247 9367 39253
rect 12158 39244 12164 39296
rect 12216 39244 12222 39296
rect 12253 39287 12311 39293
rect 12253 39253 12265 39287
rect 12299 39284 12311 39287
rect 13630 39284 13636 39296
rect 12299 39256 13636 39284
rect 12299 39253 12311 39256
rect 12253 39247 12311 39253
rect 13630 39244 13636 39256
rect 13688 39284 13694 39296
rect 14829 39287 14887 39293
rect 14829 39284 14841 39287
rect 13688 39256 14841 39284
rect 13688 39244 13694 39256
rect 14829 39253 14841 39256
rect 14875 39284 14887 39287
rect 15470 39284 15476 39296
rect 14875 39256 15476 39284
rect 14875 39253 14887 39256
rect 14829 39247 14887 39253
rect 15470 39244 15476 39256
rect 15528 39244 15534 39296
rect 16758 39244 16764 39296
rect 16816 39244 16822 39296
rect 17126 39244 17132 39296
rect 17184 39284 17190 39296
rect 20162 39284 20168 39296
rect 17184 39256 20168 39284
rect 17184 39244 17190 39256
rect 20162 39244 20168 39256
rect 20220 39244 20226 39296
rect 23658 39244 23664 39296
rect 23716 39244 23722 39296
rect 24762 39244 24768 39296
rect 24820 39284 24826 39296
rect 29086 39284 29092 39296
rect 24820 39256 29092 39284
rect 24820 39244 24826 39256
rect 29086 39244 29092 39256
rect 29144 39244 29150 39296
rect 30668 39293 30696 39324
rect 31174 39321 31186 39324
rect 31220 39321 31232 39355
rect 35434 39352 35440 39364
rect 31174 39315 31232 39321
rect 31312 39324 35440 39352
rect 30653 39287 30711 39293
rect 30653 39253 30665 39287
rect 30699 39253 30711 39287
rect 30653 39247 30711 39253
rect 30742 39244 30748 39296
rect 30800 39284 30806 39296
rect 31312 39284 31340 39324
rect 35434 39312 35440 39324
rect 35492 39312 35498 39364
rect 35986 39312 35992 39364
rect 36044 39312 36050 39364
rect 36372 39352 36400 39380
rect 36906 39352 36912 39364
rect 36372 39324 36912 39352
rect 36906 39312 36912 39324
rect 36964 39312 36970 39364
rect 37553 39355 37611 39361
rect 37553 39321 37565 39355
rect 37599 39352 37611 39355
rect 37599 39324 37780 39352
rect 37599 39321 37611 39324
rect 37553 39315 37611 39321
rect 30800 39256 31340 39284
rect 32309 39287 32367 39293
rect 30800 39244 30806 39256
rect 32309 39253 32321 39287
rect 32355 39284 32367 39287
rect 32674 39284 32680 39296
rect 32355 39256 32680 39284
rect 32355 39253 32367 39256
rect 32309 39247 32367 39253
rect 32674 39244 32680 39256
rect 32732 39284 32738 39296
rect 32769 39287 32827 39293
rect 32769 39284 32781 39287
rect 32732 39256 32781 39284
rect 32732 39244 32738 39256
rect 32769 39253 32781 39256
rect 32815 39253 32827 39287
rect 32769 39247 32827 39253
rect 32858 39244 32864 39296
rect 32916 39244 32922 39296
rect 34330 39244 34336 39296
rect 34388 39284 34394 39296
rect 35158 39284 35164 39296
rect 34388 39256 35164 39284
rect 34388 39244 34394 39256
rect 35158 39244 35164 39256
rect 35216 39244 35222 39296
rect 36004 39284 36032 39312
rect 37752 39296 37780 39324
rect 37826 39312 37832 39364
rect 37884 39352 37890 39364
rect 38534 39355 38592 39361
rect 38534 39352 38546 39355
rect 37884 39324 38546 39352
rect 37884 39312 37890 39324
rect 38534 39321 38546 39324
rect 38580 39321 38592 39355
rect 38534 39315 38592 39321
rect 36630 39284 36636 39296
rect 36004 39256 36636 39284
rect 36630 39244 36636 39256
rect 36688 39244 36694 39296
rect 36722 39244 36728 39296
rect 36780 39244 36786 39296
rect 37734 39244 37740 39296
rect 37792 39284 37798 39296
rect 38029 39287 38087 39293
rect 38029 39284 38041 39287
rect 37792 39256 38041 39284
rect 37792 39244 37798 39256
rect 38029 39253 38041 39256
rect 38075 39253 38087 39287
rect 38029 39247 38087 39253
rect 38194 39244 38200 39296
rect 38252 39244 38258 39296
rect 1104 39194 47104 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 35594 39194
rect 35646 39142 35658 39194
rect 35710 39142 35722 39194
rect 35774 39142 35786 39194
rect 35838 39142 35850 39194
rect 35902 39142 47104 39194
rect 1104 39120 47104 39142
rect 3510 39040 3516 39092
rect 3568 39080 3574 39092
rect 31478 39080 31484 39092
rect 3568 39052 31484 39080
rect 3568 39040 3574 39052
rect 31478 39040 31484 39052
rect 31536 39040 31542 39092
rect 34330 39040 34336 39092
rect 34388 39080 34394 39092
rect 34425 39083 34483 39089
rect 34425 39080 34437 39083
rect 34388 39052 34437 39080
rect 34388 39040 34394 39052
rect 34425 39049 34437 39052
rect 34471 39049 34483 39083
rect 34425 39043 34483 39049
rect 34514 39040 34520 39092
rect 34572 39080 34578 39092
rect 35529 39083 35587 39089
rect 35529 39080 35541 39083
rect 34572 39052 35541 39080
rect 34572 39040 34578 39052
rect 35529 39049 35541 39052
rect 35575 39049 35587 39083
rect 37274 39080 37280 39092
rect 35529 39043 35587 39049
rect 36648 39052 37280 39080
rect 16390 38972 16396 39024
rect 16448 39012 16454 39024
rect 16448 38984 17724 39012
rect 16448 38972 16454 38984
rect 7561 38947 7619 38953
rect 7561 38913 7573 38947
rect 7607 38944 7619 38947
rect 7650 38944 7656 38956
rect 7607 38916 7656 38944
rect 7607 38913 7619 38916
rect 7561 38907 7619 38913
rect 7650 38904 7656 38916
rect 7708 38904 7714 38956
rect 9493 38947 9551 38953
rect 9493 38913 9505 38947
rect 9539 38944 9551 38947
rect 10502 38944 10508 38956
rect 9539 38916 10508 38944
rect 9539 38913 9551 38916
rect 9493 38907 9551 38913
rect 10502 38904 10508 38916
rect 10560 38904 10566 38956
rect 15102 38904 15108 38956
rect 15160 38904 15166 38956
rect 15372 38947 15430 38953
rect 15372 38913 15384 38947
rect 15418 38944 15430 38947
rect 15930 38944 15936 38956
rect 15418 38916 15936 38944
rect 15418 38913 15430 38916
rect 15372 38907 15430 38913
rect 15930 38904 15936 38916
rect 15988 38904 15994 38956
rect 17696 38953 17724 38984
rect 17770 38972 17776 39024
rect 17828 39012 17834 39024
rect 27982 39012 27988 39024
rect 17828 38984 27988 39012
rect 17828 38972 17834 38984
rect 27982 38972 27988 38984
rect 28040 38972 28046 39024
rect 29730 38972 29736 39024
rect 29788 39012 29794 39024
rect 30282 39012 30288 39024
rect 29788 38984 30288 39012
rect 29788 38972 29794 38984
rect 30282 38972 30288 38984
rect 30340 38972 30346 39024
rect 31202 38972 31208 39024
rect 31260 38972 31266 39024
rect 31294 38972 31300 39024
rect 31352 39012 31358 39024
rect 31389 39015 31447 39021
rect 31389 39012 31401 39015
rect 31352 38984 31401 39012
rect 31352 38972 31358 38984
rect 31389 38981 31401 38984
rect 31435 39012 31447 39015
rect 32858 39012 32864 39024
rect 31435 38984 32864 39012
rect 31435 38981 31447 38984
rect 31389 38975 31447 38981
rect 32858 38972 32864 38984
rect 32916 38972 32922 39024
rect 34146 39012 34152 39024
rect 33060 38984 34152 39012
rect 17037 38947 17095 38953
rect 17037 38944 17049 38947
rect 16500 38916 17049 38944
rect 16500 38817 16528 38916
rect 17037 38913 17049 38916
rect 17083 38944 17095 38947
rect 17681 38947 17739 38953
rect 17083 38916 17632 38944
rect 17083 38913 17095 38916
rect 17037 38907 17095 38913
rect 16850 38836 16856 38888
rect 16908 38876 16914 38888
rect 17129 38879 17187 38885
rect 17129 38876 17141 38879
rect 16908 38848 17141 38876
rect 16908 38836 16914 38848
rect 17129 38845 17141 38848
rect 17175 38845 17187 38879
rect 17129 38839 17187 38845
rect 17310 38836 17316 38888
rect 17368 38836 17374 38888
rect 17604 38876 17632 38916
rect 17681 38913 17693 38947
rect 17727 38913 17739 38947
rect 17681 38907 17739 38913
rect 19518 38904 19524 38956
rect 19576 38904 19582 38956
rect 20073 38947 20131 38953
rect 20073 38913 20085 38947
rect 20119 38944 20131 38947
rect 20622 38944 20628 38956
rect 20119 38916 20628 38944
rect 20119 38913 20131 38916
rect 20073 38907 20131 38913
rect 20622 38904 20628 38916
rect 20680 38904 20686 38956
rect 21726 38904 21732 38956
rect 21784 38944 21790 38956
rect 22094 38953 22100 38956
rect 21821 38947 21879 38953
rect 21821 38944 21833 38947
rect 21784 38916 21833 38944
rect 21784 38904 21790 38916
rect 21821 38913 21833 38916
rect 21867 38913 21879 38947
rect 21821 38907 21879 38913
rect 22088 38907 22100 38953
rect 22094 38904 22100 38907
rect 22152 38904 22158 38956
rect 24489 38947 24547 38953
rect 24489 38913 24501 38947
rect 24535 38944 24547 38947
rect 25314 38944 25320 38956
rect 24535 38916 25320 38944
rect 24535 38913 24547 38916
rect 24489 38907 24547 38913
rect 25314 38904 25320 38916
rect 25372 38944 25378 38956
rect 25774 38944 25780 38956
rect 25372 38916 25780 38944
rect 25372 38904 25378 38916
rect 25774 38904 25780 38916
rect 25832 38904 25838 38956
rect 30193 38947 30251 38953
rect 30193 38913 30205 38947
rect 30239 38944 30251 38947
rect 30926 38944 30932 38956
rect 30239 38916 30932 38944
rect 30239 38913 30251 38916
rect 30193 38907 30251 38913
rect 30926 38904 30932 38916
rect 30984 38904 30990 38956
rect 31938 38944 31944 38956
rect 31036 38916 31944 38944
rect 17954 38876 17960 38888
rect 17604 38848 17960 38876
rect 17954 38836 17960 38848
rect 18012 38876 18018 38888
rect 18230 38876 18236 38888
rect 18012 38848 18236 38876
rect 18012 38836 18018 38848
rect 18230 38836 18236 38848
rect 18288 38836 18294 38888
rect 20162 38836 20168 38888
rect 20220 38836 20226 38888
rect 20257 38879 20315 38885
rect 20257 38845 20269 38879
rect 20303 38845 20315 38879
rect 20257 38839 20315 38845
rect 16485 38811 16543 38817
rect 16485 38777 16497 38811
rect 16531 38777 16543 38811
rect 16868 38808 16896 38836
rect 16485 38771 16543 38777
rect 16592 38780 16896 38808
rect 7374 38700 7380 38752
rect 7432 38700 7438 38752
rect 9306 38700 9312 38752
rect 9364 38700 9370 38752
rect 14090 38700 14096 38752
rect 14148 38740 14154 38752
rect 14734 38740 14740 38752
rect 14148 38712 14740 38740
rect 14148 38700 14154 38712
rect 14734 38700 14740 38712
rect 14792 38740 14798 38752
rect 16592 38740 16620 38780
rect 17494 38768 17500 38820
rect 17552 38768 17558 38820
rect 20272 38808 20300 38839
rect 23658 38836 23664 38888
rect 23716 38876 23722 38888
rect 24581 38879 24639 38885
rect 24581 38876 24593 38879
rect 23716 38848 24593 38876
rect 23716 38836 23722 38848
rect 24581 38845 24593 38848
rect 24627 38845 24639 38879
rect 24581 38839 24639 38845
rect 24765 38879 24823 38885
rect 24765 38845 24777 38879
rect 24811 38876 24823 38879
rect 27338 38876 27344 38888
rect 24811 38848 27344 38876
rect 24811 38845 24823 38848
rect 24765 38839 24823 38845
rect 17604 38780 20300 38808
rect 24596 38808 24624 38839
rect 27338 38836 27344 38848
rect 27396 38836 27402 38888
rect 30469 38879 30527 38885
rect 30469 38845 30481 38879
rect 30515 38876 30527 38879
rect 31036 38876 31064 38916
rect 31938 38904 31944 38916
rect 31996 38904 32002 38956
rect 33060 38944 33088 38984
rect 34146 38972 34152 38984
rect 34204 38972 34210 39024
rect 36538 39012 36544 39024
rect 34348 38984 35046 39012
rect 34348 38956 34376 38984
rect 32876 38916 33088 38944
rect 33312 38947 33370 38953
rect 30515 38848 31064 38876
rect 30515 38845 30527 38848
rect 30469 38839 30527 38845
rect 24596 38780 31248 38808
rect 14792 38712 16620 38740
rect 14792 38700 14798 38712
rect 16666 38700 16672 38752
rect 16724 38700 16730 38752
rect 17218 38700 17224 38752
rect 17276 38740 17282 38752
rect 17604 38740 17632 38780
rect 31220 38752 31248 38780
rect 17276 38712 17632 38740
rect 17276 38700 17282 38712
rect 19334 38700 19340 38752
rect 19392 38700 19398 38752
rect 19705 38743 19763 38749
rect 19705 38709 19717 38743
rect 19751 38740 19763 38743
rect 20898 38740 20904 38752
rect 19751 38712 20904 38740
rect 19751 38709 19763 38712
rect 19705 38703 19763 38709
rect 20898 38700 20904 38712
rect 20956 38700 20962 38752
rect 23198 38700 23204 38752
rect 23256 38700 23262 38752
rect 24118 38700 24124 38752
rect 24176 38700 24182 38752
rect 29825 38743 29883 38749
rect 29825 38709 29837 38743
rect 29871 38740 29883 38743
rect 29914 38740 29920 38752
rect 29871 38712 29920 38740
rect 29871 38709 29883 38712
rect 29825 38703 29883 38709
rect 29914 38700 29920 38712
rect 29972 38700 29978 38752
rect 31202 38700 31208 38752
rect 31260 38740 31266 38752
rect 32876 38740 32904 38916
rect 33312 38913 33324 38947
rect 33358 38944 33370 38947
rect 33358 38916 34100 38944
rect 33358 38913 33370 38916
rect 33312 38907 33370 38913
rect 33042 38836 33048 38888
rect 33100 38836 33106 38888
rect 31260 38712 32904 38740
rect 34072 38740 34100 38916
rect 34330 38904 34336 38956
rect 34388 38904 34394 38956
rect 34701 38947 34759 38953
rect 34701 38913 34713 38947
rect 34747 38913 34759 38947
rect 34701 38907 34759 38913
rect 34716 38876 34744 38907
rect 34790 38904 34796 38956
rect 34848 38904 34854 38956
rect 34882 38904 34888 38956
rect 34940 38904 34946 38956
rect 35018 38953 35046 38984
rect 35728 38984 36544 39012
rect 35003 38947 35061 38953
rect 35003 38913 35015 38947
rect 35049 38913 35061 38947
rect 35003 38907 35061 38913
rect 35018 38876 35046 38907
rect 35158 38904 35164 38956
rect 35216 38904 35222 38956
rect 35342 38904 35348 38956
rect 35400 38944 35406 38956
rect 35728 38953 35756 38984
rect 36538 38972 36544 38984
rect 36596 38972 36602 39024
rect 35713 38947 35771 38953
rect 35713 38944 35725 38947
rect 35400 38916 35725 38944
rect 35400 38904 35406 38916
rect 35713 38913 35725 38916
rect 35759 38913 35771 38947
rect 35713 38907 35771 38913
rect 36170 38904 36176 38956
rect 36228 38904 36234 38956
rect 36449 38947 36507 38953
rect 36449 38913 36461 38947
rect 36495 38944 36507 38947
rect 36648 38944 36676 39052
rect 37274 39040 37280 39052
rect 37332 39040 37338 39092
rect 37645 39083 37703 39089
rect 37645 39049 37657 39083
rect 37691 39080 37703 39083
rect 37734 39080 37740 39092
rect 37691 39052 37740 39080
rect 37691 39049 37703 39052
rect 37645 39043 37703 39049
rect 37734 39040 37740 39052
rect 37792 39040 37798 39092
rect 38286 38972 38292 39024
rect 38344 39012 38350 39024
rect 38381 39015 38439 39021
rect 38381 39012 38393 39015
rect 38344 38984 38393 39012
rect 38344 38972 38350 38984
rect 38381 38981 38393 38984
rect 38427 38981 38439 39015
rect 38381 38975 38439 38981
rect 36495 38916 36676 38944
rect 36817 38947 36875 38953
rect 36495 38913 36507 38916
rect 36449 38907 36507 38913
rect 36817 38913 36829 38947
rect 36863 38913 36875 38947
rect 36817 38907 36875 38913
rect 35526 38876 35532 38888
rect 34716 38848 34836 38876
rect 35018 38848 35532 38876
rect 34517 38743 34575 38749
rect 34517 38740 34529 38743
rect 34072 38712 34529 38740
rect 31260 38700 31266 38712
rect 34517 38709 34529 38712
rect 34563 38709 34575 38743
rect 34808 38740 34836 38848
rect 35526 38836 35532 38848
rect 35584 38836 35590 38888
rect 35802 38836 35808 38888
rect 35860 38876 35866 38888
rect 36464 38876 36492 38907
rect 35860 38848 36492 38876
rect 35860 38836 35866 38848
rect 36538 38836 36544 38888
rect 36596 38876 36602 38888
rect 36832 38876 36860 38907
rect 36906 38904 36912 38956
rect 36964 38944 36970 38956
rect 37277 38947 37335 38953
rect 37277 38944 37289 38947
rect 36964 38916 37289 38944
rect 36964 38904 36970 38916
rect 37277 38913 37289 38916
rect 37323 38913 37335 38947
rect 37277 38907 37335 38913
rect 37458 38904 37464 38956
rect 37516 38904 37522 38956
rect 37553 38947 37611 38953
rect 37553 38913 37565 38947
rect 37599 38944 37611 38947
rect 37642 38944 37648 38956
rect 37599 38916 37648 38944
rect 37599 38913 37611 38916
rect 37553 38907 37611 38913
rect 37568 38876 37596 38907
rect 37642 38904 37648 38916
rect 37700 38904 37706 38956
rect 37737 38947 37795 38953
rect 37737 38913 37749 38947
rect 37783 38944 37795 38947
rect 38010 38944 38016 38956
rect 37783 38916 38016 38944
rect 37783 38913 37795 38916
rect 37737 38907 37795 38913
rect 38010 38904 38016 38916
rect 38068 38944 38074 38956
rect 38562 38944 38568 38956
rect 38068 38916 38568 38944
rect 38068 38904 38074 38916
rect 38562 38904 38568 38916
rect 38620 38904 38626 38956
rect 36596 38848 37596 38876
rect 36596 38836 36602 38848
rect 36998 38740 37004 38752
rect 34808 38712 37004 38740
rect 34517 38703 34575 38709
rect 36998 38700 37004 38712
rect 37056 38700 37062 38752
rect 37277 38743 37335 38749
rect 37277 38709 37289 38743
rect 37323 38740 37335 38743
rect 37458 38740 37464 38752
rect 37323 38712 37464 38740
rect 37323 38709 37335 38712
rect 37277 38703 37335 38709
rect 37458 38700 37464 38712
rect 37516 38700 37522 38752
rect 38010 38700 38016 38752
rect 38068 38740 38074 38752
rect 38473 38743 38531 38749
rect 38473 38740 38485 38743
rect 38068 38712 38485 38740
rect 38068 38700 38074 38712
rect 38473 38709 38485 38712
rect 38519 38709 38531 38743
rect 38473 38703 38531 38709
rect 1104 38650 47104 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 47104 38650
rect 1104 38576 47104 38598
rect 5350 38496 5356 38548
rect 5408 38536 5414 38548
rect 5408 38508 8156 38536
rect 5408 38496 5414 38508
rect 8128 38400 8156 38508
rect 10962 38496 10968 38548
rect 11020 38536 11026 38548
rect 11020 38508 15884 38536
rect 11020 38496 11026 38508
rect 15856 38468 15884 38508
rect 15930 38496 15936 38548
rect 15988 38536 15994 38548
rect 16025 38539 16083 38545
rect 16025 38536 16037 38539
rect 15988 38508 16037 38536
rect 15988 38496 15994 38508
rect 16025 38505 16037 38508
rect 16071 38505 16083 38539
rect 16025 38499 16083 38505
rect 16390 38496 16396 38548
rect 16448 38496 16454 38548
rect 20162 38536 20168 38548
rect 17144 38508 20168 38536
rect 17144 38468 17172 38508
rect 20162 38496 20168 38508
rect 20220 38496 20226 38548
rect 20622 38496 20628 38548
rect 20680 38496 20686 38548
rect 21450 38496 21456 38548
rect 21508 38536 21514 38548
rect 21508 38508 22876 38536
rect 21508 38496 21514 38508
rect 17678 38468 17684 38480
rect 15856 38440 17172 38468
rect 17236 38440 17684 38468
rect 13998 38400 14004 38412
rect 8128 38372 9168 38400
rect 4341 38335 4399 38341
rect 4341 38301 4353 38335
rect 4387 38332 4399 38335
rect 5258 38332 5264 38344
rect 4387 38304 5264 38332
rect 4387 38301 4399 38304
rect 4341 38295 4399 38301
rect 5258 38292 5264 38304
rect 5316 38292 5322 38344
rect 5626 38292 5632 38344
rect 5684 38292 5690 38344
rect 7374 38341 7380 38344
rect 7101 38335 7159 38341
rect 7101 38301 7113 38335
rect 7147 38301 7159 38335
rect 7368 38332 7380 38341
rect 7335 38304 7380 38332
rect 7101 38295 7159 38301
rect 7368 38295 7380 38304
rect 5896 38267 5954 38273
rect 5896 38233 5908 38267
rect 5942 38264 5954 38267
rect 5994 38264 6000 38276
rect 5942 38236 6000 38264
rect 5942 38233 5954 38236
rect 5896 38227 5954 38233
rect 5994 38224 6000 38236
rect 6052 38224 6058 38276
rect 7116 38264 7144 38295
rect 7374 38292 7380 38295
rect 7432 38292 7438 38344
rect 9033 38335 9091 38341
rect 9033 38301 9045 38335
rect 9079 38301 9091 38335
rect 9033 38295 9091 38301
rect 8938 38264 8944 38276
rect 7116 38236 8944 38264
rect 8938 38224 8944 38236
rect 8996 38264 9002 38276
rect 9048 38264 9076 38295
rect 8996 38236 9076 38264
rect 9140 38264 9168 38372
rect 12406 38372 14004 38400
rect 9306 38341 9312 38344
rect 9300 38332 9312 38341
rect 9267 38304 9312 38332
rect 9300 38295 9312 38304
rect 9306 38292 9312 38295
rect 9364 38292 9370 38344
rect 11149 38335 11207 38341
rect 11149 38301 11161 38335
rect 11195 38332 11207 38335
rect 12406 38332 12434 38372
rect 13998 38360 14004 38372
rect 14056 38400 14062 38412
rect 14093 38403 14151 38409
rect 14093 38400 14105 38403
rect 14056 38372 14105 38400
rect 14056 38360 14062 38372
rect 14093 38369 14105 38372
rect 14139 38369 14151 38403
rect 14093 38363 14151 38369
rect 16942 38360 16948 38412
rect 17000 38360 17006 38412
rect 17034 38360 17040 38412
rect 17092 38400 17098 38412
rect 17236 38409 17264 38440
rect 17678 38428 17684 38440
rect 17736 38428 17742 38480
rect 20640 38468 20668 38496
rect 17788 38440 18000 38468
rect 20640 38440 21956 38468
rect 17788 38412 17816 38440
rect 17221 38403 17279 38409
rect 17221 38400 17233 38403
rect 17092 38372 17233 38400
rect 17092 38360 17098 38372
rect 17221 38369 17233 38372
rect 17267 38369 17279 38403
rect 17770 38400 17776 38412
rect 17221 38363 17279 38369
rect 17328 38372 17776 38400
rect 11195 38304 12434 38332
rect 12805 38335 12863 38341
rect 11195 38301 11207 38304
rect 11149 38295 11207 38301
rect 12805 38301 12817 38335
rect 12851 38332 12863 38335
rect 13354 38332 13360 38344
rect 12851 38304 13360 38332
rect 12851 38301 12863 38304
rect 12805 38295 12863 38301
rect 13354 38292 13360 38304
rect 13412 38292 13418 38344
rect 13630 38292 13636 38344
rect 13688 38292 13694 38344
rect 13906 38292 13912 38344
rect 13964 38292 13970 38344
rect 16209 38335 16267 38341
rect 16209 38301 16221 38335
rect 16255 38332 16267 38335
rect 16666 38332 16672 38344
rect 16255 38304 16672 38332
rect 16255 38301 16267 38304
rect 16209 38295 16267 38301
rect 16666 38292 16672 38304
rect 16724 38292 16730 38344
rect 16758 38292 16764 38344
rect 16816 38332 16822 38344
rect 17328 38332 17356 38372
rect 17770 38360 17776 38372
rect 17828 38360 17834 38412
rect 17862 38360 17868 38412
rect 17920 38360 17926 38412
rect 17972 38400 18000 38440
rect 18141 38403 18199 38409
rect 18141 38400 18153 38403
rect 17972 38372 18153 38400
rect 18141 38369 18153 38372
rect 18187 38369 18199 38403
rect 18141 38363 18199 38369
rect 18230 38360 18236 38412
rect 18288 38409 18294 38412
rect 18288 38403 18316 38409
rect 18304 38369 18316 38403
rect 18288 38363 18316 38369
rect 18288 38360 18294 38363
rect 21174 38360 21180 38412
rect 21232 38360 21238 38412
rect 21821 38403 21879 38409
rect 21821 38400 21833 38403
rect 21284 38372 21833 38400
rect 16816 38304 17356 38332
rect 17405 38335 17463 38341
rect 16816 38292 16822 38304
rect 17405 38301 17417 38335
rect 17451 38301 17463 38335
rect 17405 38295 17463 38301
rect 9214 38264 9220 38276
rect 9140 38236 9220 38264
rect 8996 38224 9002 38236
rect 9214 38224 9220 38236
rect 9272 38264 9278 38276
rect 10686 38264 10692 38276
rect 9272 38236 10692 38264
rect 9272 38224 9278 38236
rect 10686 38224 10692 38236
rect 10744 38224 10750 38276
rect 11416 38267 11474 38273
rect 11416 38233 11428 38267
rect 11462 38264 11474 38267
rect 14338 38267 14396 38273
rect 14338 38264 14350 38267
rect 11462 38236 12664 38264
rect 11462 38233 11474 38236
rect 11416 38227 11474 38233
rect 4154 38156 4160 38208
rect 4212 38156 4218 38208
rect 7006 38156 7012 38208
rect 7064 38156 7070 38208
rect 8478 38156 8484 38208
rect 8536 38156 8542 38208
rect 8754 38156 8760 38208
rect 8812 38196 8818 38208
rect 10413 38199 10471 38205
rect 10413 38196 10425 38199
rect 8812 38168 10425 38196
rect 8812 38156 8818 38168
rect 10413 38165 10425 38168
rect 10459 38196 10471 38199
rect 10870 38196 10876 38208
rect 10459 38168 10876 38196
rect 10459 38165 10471 38168
rect 10413 38159 10471 38165
rect 10870 38156 10876 38168
rect 10928 38156 10934 38208
rect 12526 38156 12532 38208
rect 12584 38156 12590 38208
rect 12636 38205 12664 38236
rect 13464 38236 14350 38264
rect 13464 38205 13492 38236
rect 14338 38233 14350 38236
rect 14384 38233 14396 38267
rect 14338 38227 14396 38233
rect 12621 38199 12679 38205
rect 12621 38165 12633 38199
rect 12667 38165 12679 38199
rect 12621 38159 12679 38165
rect 13449 38199 13507 38205
rect 13449 38165 13461 38199
rect 13495 38165 13507 38199
rect 13449 38159 13507 38165
rect 13725 38199 13783 38205
rect 13725 38165 13737 38199
rect 13771 38196 13783 38199
rect 13814 38196 13820 38208
rect 13771 38168 13820 38196
rect 13771 38165 13783 38168
rect 13725 38159 13783 38165
rect 13814 38156 13820 38168
rect 13872 38156 13878 38208
rect 15470 38156 15476 38208
rect 15528 38156 15534 38208
rect 16850 38156 16856 38208
rect 16908 38156 16914 38208
rect 17420 38196 17448 38295
rect 18414 38292 18420 38344
rect 18472 38292 18478 38344
rect 19058 38292 19064 38344
rect 19116 38332 19122 38344
rect 19245 38335 19303 38341
rect 19245 38332 19257 38335
rect 19116 38304 19257 38332
rect 19116 38292 19122 38304
rect 19245 38301 19257 38304
rect 19291 38301 19303 38335
rect 19245 38295 19303 38301
rect 19444 38304 20852 38332
rect 18966 38224 18972 38276
rect 19024 38264 19030 38276
rect 19444 38264 19472 38304
rect 19024 38236 19472 38264
rect 19512 38267 19570 38273
rect 19024 38224 19030 38236
rect 19512 38233 19524 38267
rect 19558 38264 19570 38267
rect 20824 38264 20852 38304
rect 20898 38292 20904 38344
rect 20956 38292 20962 38344
rect 21284 38264 21312 38372
rect 21821 38369 21833 38372
rect 21867 38369 21879 38403
rect 21928 38400 21956 38440
rect 22097 38403 22155 38409
rect 22097 38400 22109 38403
rect 21928 38372 22109 38400
rect 21821 38363 21879 38369
rect 22097 38369 22109 38372
rect 22143 38400 22155 38403
rect 22738 38400 22744 38412
rect 22143 38372 22744 38400
rect 22143 38369 22155 38372
rect 22097 38363 22155 38369
rect 22738 38360 22744 38372
rect 22796 38360 22802 38412
rect 22848 38400 22876 38508
rect 23768 38508 25360 38536
rect 22922 38428 22928 38480
rect 22980 38468 22986 38480
rect 23768 38468 23796 38508
rect 22980 38440 23796 38468
rect 25332 38468 25360 38508
rect 25774 38496 25780 38548
rect 25832 38496 25838 38548
rect 25976 38508 30512 38536
rect 25976 38468 26004 38508
rect 25332 38440 26004 38468
rect 30484 38468 30512 38508
rect 30926 38496 30932 38548
rect 30984 38496 30990 38548
rect 31036 38508 33548 38536
rect 31036 38468 31064 38508
rect 33520 38477 33548 38508
rect 35434 38496 35440 38548
rect 35492 38536 35498 38548
rect 35529 38539 35587 38545
rect 35529 38536 35541 38539
rect 35492 38508 35541 38536
rect 35492 38496 35498 38508
rect 35529 38505 35541 38508
rect 35575 38505 35587 38539
rect 38194 38536 38200 38548
rect 35529 38499 35587 38505
rect 37384 38508 38200 38536
rect 30484 38440 31064 38468
rect 33505 38471 33563 38477
rect 22980 38428 22986 38440
rect 33505 38437 33517 38471
rect 33551 38437 33563 38471
rect 35802 38468 35808 38480
rect 33505 38431 33563 38437
rect 34716 38440 35808 38468
rect 23569 38403 23627 38409
rect 23569 38400 23581 38403
rect 22848 38372 23581 38400
rect 23569 38369 23581 38372
rect 23615 38400 23627 38403
rect 23658 38400 23664 38412
rect 23615 38372 23664 38400
rect 23615 38369 23627 38372
rect 23569 38363 23627 38369
rect 23658 38360 23664 38372
rect 23716 38360 23722 38412
rect 23753 38403 23811 38409
rect 23753 38369 23765 38403
rect 23799 38400 23811 38403
rect 23842 38400 23848 38412
rect 23799 38372 23848 38400
rect 23799 38369 23811 38372
rect 23753 38363 23811 38369
rect 23842 38360 23848 38372
rect 23900 38360 23906 38412
rect 24302 38360 24308 38412
rect 24360 38400 24366 38412
rect 24397 38403 24455 38409
rect 24397 38400 24409 38403
rect 24360 38372 24409 38400
rect 24360 38360 24366 38372
rect 24397 38369 24409 38372
rect 24443 38369 24455 38403
rect 24397 38363 24455 38369
rect 27338 38360 27344 38412
rect 27396 38400 27402 38412
rect 28353 38403 28411 38409
rect 28353 38400 28365 38403
rect 27396 38372 28365 38400
rect 27396 38360 27402 38372
rect 28353 38369 28365 38372
rect 28399 38369 28411 38403
rect 28353 38363 28411 38369
rect 28442 38360 28448 38412
rect 28500 38400 28506 38412
rect 29549 38403 29607 38409
rect 29549 38400 29561 38403
rect 28500 38372 29561 38400
rect 28500 38360 28506 38372
rect 29549 38369 29561 38372
rect 29595 38369 29607 38403
rect 29549 38363 29607 38369
rect 31018 38360 31024 38412
rect 31076 38400 31082 38412
rect 31662 38400 31668 38412
rect 31076 38372 31668 38400
rect 31076 38360 31082 38372
rect 31662 38360 31668 38372
rect 31720 38360 31726 38412
rect 34422 38360 34428 38412
rect 34480 38360 34486 38412
rect 21361 38335 21419 38341
rect 21361 38301 21373 38335
rect 21407 38301 21419 38335
rect 21361 38295 21419 38301
rect 19558 38236 20760 38264
rect 20824 38236 21312 38264
rect 19558 38233 19570 38236
rect 19512 38227 19570 38233
rect 18138 38196 18144 38208
rect 17420 38168 18144 38196
rect 18138 38156 18144 38168
rect 18196 38156 18202 38208
rect 19061 38199 19119 38205
rect 19061 38165 19073 38199
rect 19107 38196 19119 38199
rect 19426 38196 19432 38208
rect 19107 38168 19432 38196
rect 19107 38165 19119 38168
rect 19061 38159 19119 38165
rect 19426 38156 19432 38168
rect 19484 38156 19490 38208
rect 20732 38205 20760 38236
rect 20717 38199 20775 38205
rect 20717 38165 20729 38199
rect 20763 38165 20775 38199
rect 21376 38196 21404 38295
rect 22186 38292 22192 38344
rect 22244 38341 22250 38344
rect 22244 38335 22272 38341
rect 22260 38301 22272 38335
rect 22244 38295 22272 38301
rect 22244 38292 22250 38295
rect 22370 38292 22376 38344
rect 22428 38292 22434 38344
rect 23198 38292 23204 38344
rect 23256 38332 23262 38344
rect 23477 38335 23535 38341
rect 23477 38332 23489 38335
rect 23256 38304 23489 38332
rect 23256 38292 23262 38304
rect 23477 38301 23489 38304
rect 23523 38301 23535 38335
rect 23477 38295 23535 38301
rect 24118 38292 24124 38344
rect 24176 38292 24182 38344
rect 26329 38335 26387 38341
rect 26329 38301 26341 38335
rect 26375 38332 26387 38335
rect 26970 38332 26976 38344
rect 26375 38304 26976 38332
rect 26375 38301 26387 38304
rect 26329 38295 26387 38301
rect 26970 38292 26976 38304
rect 27028 38332 27034 38344
rect 27798 38332 27804 38344
rect 27028 38304 27804 38332
rect 27028 38292 27034 38304
rect 27798 38292 27804 38304
rect 27856 38292 27862 38344
rect 31570 38292 31576 38344
rect 31628 38292 31634 38344
rect 33597 38335 33655 38341
rect 33597 38301 33609 38335
rect 33643 38301 33655 38335
rect 33597 38295 33655 38301
rect 23216 38264 23244 38292
rect 26602 38273 26608 38276
rect 22848 38236 23244 38264
rect 24642 38267 24700 38273
rect 21910 38196 21916 38208
rect 21376 38168 21916 38196
rect 20717 38159 20775 38165
rect 21910 38156 21916 38168
rect 21968 38196 21974 38208
rect 22848 38196 22876 38236
rect 24642 38233 24654 38267
rect 24688 38233 24700 38267
rect 24642 38227 24700 38233
rect 26596 38227 26608 38273
rect 21968 38168 22876 38196
rect 21968 38156 21974 38168
rect 23014 38156 23020 38208
rect 23072 38156 23078 38208
rect 23106 38156 23112 38208
rect 23164 38156 23170 38208
rect 23937 38199 23995 38205
rect 23937 38165 23949 38199
rect 23983 38196 23995 38199
rect 24657 38196 24685 38227
rect 26602 38224 26608 38227
rect 26660 38224 26666 38276
rect 28074 38224 28080 38276
rect 28132 38264 28138 38276
rect 29822 38273 29828 38276
rect 28261 38267 28319 38273
rect 28261 38264 28273 38267
rect 28132 38236 28273 38264
rect 28132 38224 28138 38236
rect 28261 38233 28273 38236
rect 28307 38233 28319 38267
rect 28261 38227 28319 38233
rect 29816 38227 29828 38273
rect 29822 38224 29828 38227
rect 29880 38224 29886 38276
rect 31910 38267 31968 38273
rect 31910 38264 31922 38267
rect 31726 38236 31922 38264
rect 23983 38168 24685 38196
rect 23983 38165 23995 38168
rect 23937 38159 23995 38165
rect 27706 38156 27712 38208
rect 27764 38156 27770 38208
rect 27798 38156 27804 38208
rect 27856 38156 27862 38208
rect 28166 38156 28172 38208
rect 28224 38156 28230 38208
rect 31389 38199 31447 38205
rect 31389 38165 31401 38199
rect 31435 38196 31447 38199
rect 31726 38196 31754 38236
rect 31910 38233 31922 38236
rect 31956 38233 31968 38267
rect 31910 38227 31968 38233
rect 33226 38224 33232 38276
rect 33284 38264 33290 38276
rect 33612 38264 33640 38295
rect 33778 38292 33784 38344
rect 33836 38332 33842 38344
rect 33965 38335 34023 38341
rect 33965 38332 33977 38335
rect 33836 38304 33977 38332
rect 33836 38292 33842 38304
rect 33965 38301 33977 38304
rect 34011 38301 34023 38335
rect 33965 38295 34023 38301
rect 34606 38292 34612 38344
rect 34664 38332 34670 38344
rect 34716 38332 34744 38440
rect 35802 38428 35808 38440
rect 35860 38428 35866 38480
rect 37384 38412 37412 38508
rect 38194 38496 38200 38508
rect 38252 38496 38258 38548
rect 39301 38539 39359 38545
rect 39301 38505 39313 38539
rect 39347 38536 39359 38539
rect 39390 38536 39396 38548
rect 39347 38508 39396 38536
rect 39347 38505 39359 38508
rect 39301 38499 39359 38505
rect 39390 38496 39396 38508
rect 39448 38496 39454 38548
rect 34790 38360 34796 38412
rect 34848 38400 34854 38412
rect 35161 38403 35219 38409
rect 35161 38400 35173 38403
rect 34848 38372 35173 38400
rect 34848 38360 34854 38372
rect 35161 38369 35173 38372
rect 35207 38400 35219 38403
rect 35207 38372 36860 38400
rect 35207 38369 35219 38372
rect 35161 38363 35219 38369
rect 35069 38335 35127 38341
rect 35069 38332 35081 38335
rect 34664 38304 35081 38332
rect 34664 38292 34670 38304
rect 35069 38301 35081 38304
rect 35115 38301 35127 38335
rect 35069 38295 35127 38301
rect 35253 38335 35311 38341
rect 35253 38301 35265 38335
rect 35299 38332 35311 38335
rect 35342 38332 35348 38344
rect 35299 38304 35348 38332
rect 35299 38301 35311 38304
rect 35253 38295 35311 38301
rect 35342 38292 35348 38304
rect 35400 38292 35406 38344
rect 35437 38335 35495 38341
rect 35437 38301 35449 38335
rect 35483 38332 35495 38335
rect 35897 38335 35955 38341
rect 35897 38332 35909 38335
rect 35483 38304 35909 38332
rect 35483 38301 35495 38304
rect 35437 38295 35495 38301
rect 35897 38301 35909 38304
rect 35943 38332 35955 38335
rect 36722 38332 36728 38344
rect 35943 38304 36728 38332
rect 35943 38301 35955 38304
rect 35897 38295 35955 38301
rect 36722 38292 36728 38304
rect 36780 38292 36786 38344
rect 36832 38276 36860 38372
rect 36998 38360 37004 38412
rect 37056 38400 37062 38412
rect 37093 38403 37151 38409
rect 37093 38400 37105 38403
rect 37056 38372 37105 38400
rect 37056 38360 37062 38372
rect 37093 38369 37105 38372
rect 37139 38369 37151 38403
rect 37093 38363 37151 38369
rect 37182 38360 37188 38412
rect 37240 38360 37246 38412
rect 37274 38360 37280 38412
rect 37332 38360 37338 38412
rect 37366 38360 37372 38412
rect 37424 38360 37430 38412
rect 37921 38335 37979 38341
rect 37921 38301 37933 38335
rect 37967 38332 37979 38335
rect 38010 38332 38016 38344
rect 37967 38304 38016 38332
rect 37967 38301 37979 38304
rect 37921 38295 37979 38301
rect 38010 38292 38016 38304
rect 38068 38292 38074 38344
rect 33284 38236 35664 38264
rect 33284 38224 33290 38236
rect 31435 38168 31754 38196
rect 31435 38165 31447 38168
rect 31389 38159 31447 38165
rect 32490 38156 32496 38208
rect 32548 38196 32554 38208
rect 33045 38199 33103 38205
rect 33045 38196 33057 38199
rect 32548 38168 33057 38196
rect 32548 38156 32554 38168
rect 33045 38165 33057 38168
rect 33091 38165 33103 38199
rect 33045 38159 33103 38165
rect 34330 38156 34336 38208
rect 34388 38196 34394 38208
rect 35526 38196 35532 38208
rect 34388 38168 35532 38196
rect 34388 38156 34394 38168
rect 35526 38156 35532 38168
rect 35584 38156 35590 38208
rect 35636 38196 35664 38236
rect 35986 38224 35992 38276
rect 36044 38264 36050 38276
rect 36633 38267 36691 38273
rect 36633 38264 36645 38267
rect 36044 38236 36645 38264
rect 36044 38224 36050 38236
rect 36633 38233 36645 38236
rect 36679 38233 36691 38267
rect 36633 38227 36691 38233
rect 36814 38224 36820 38276
rect 36872 38264 36878 38276
rect 38166 38267 38224 38273
rect 38166 38264 38178 38267
rect 36872 38236 38178 38264
rect 36872 38224 36878 38236
rect 38166 38233 38178 38236
rect 38212 38233 38224 38267
rect 38166 38227 38224 38233
rect 36906 38196 36912 38208
rect 35636 38168 36912 38196
rect 36906 38156 36912 38168
rect 36964 38156 36970 38208
rect 1104 38106 47104 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 35594 38106
rect 35646 38054 35658 38106
rect 35710 38054 35722 38106
rect 35774 38054 35786 38106
rect 35838 38054 35850 38106
rect 35902 38054 47104 38106
rect 1104 38032 47104 38054
rect 5994 37952 6000 38004
rect 6052 37952 6058 38004
rect 7006 37952 7012 38004
rect 7064 37992 7070 38004
rect 9582 37992 9588 38004
rect 7064 37964 9588 37992
rect 7064 37952 7070 37964
rect 9582 37952 9588 37964
rect 9640 37952 9646 38004
rect 10502 37952 10508 38004
rect 10560 37952 10566 38004
rect 10870 37952 10876 38004
rect 10928 37952 10934 38004
rect 10962 37952 10968 38004
rect 11020 37952 11026 38004
rect 12526 37992 12532 38004
rect 11716 37964 12532 37992
rect 3418 37884 3424 37936
rect 3476 37924 3482 37936
rect 4056 37927 4114 37933
rect 3476 37896 3832 37924
rect 3476 37884 3482 37896
rect 3804 37868 3832 37896
rect 4056 37893 4068 37927
rect 4102 37924 4114 37927
rect 4154 37924 4160 37936
rect 4102 37896 4160 37924
rect 4102 37893 4114 37896
rect 4056 37887 4114 37893
rect 4154 37884 4160 37896
rect 4212 37884 4218 37936
rect 6454 37924 6460 37936
rect 6196 37896 6460 37924
rect 3694 37816 3700 37868
rect 3752 37816 3758 37868
rect 3786 37816 3792 37868
rect 3844 37856 3850 37868
rect 6196 37865 6224 37896
rect 6454 37884 6460 37896
rect 6512 37884 6518 37936
rect 6181 37859 6239 37865
rect 3844 37828 5672 37856
rect 3844 37816 3850 37828
rect 5644 37800 5672 37828
rect 6181 37825 6193 37859
rect 6227 37825 6239 37859
rect 6181 37819 6239 37825
rect 6270 37816 6276 37868
rect 6328 37856 6334 37868
rect 6621 37859 6679 37865
rect 6621 37856 6633 37859
rect 6328 37828 6633 37856
rect 6328 37816 6334 37828
rect 6621 37825 6633 37828
rect 6667 37825 6679 37859
rect 6621 37819 6679 37825
rect 8478 37816 8484 37868
rect 8536 37856 8542 37868
rect 8573 37859 8631 37865
rect 8573 37856 8585 37859
rect 8536 37828 8585 37856
rect 8536 37816 8542 37828
rect 8573 37825 8585 37828
rect 8619 37825 8631 37859
rect 8573 37819 8631 37825
rect 8754 37816 8760 37868
rect 8812 37816 8818 37868
rect 9582 37816 9588 37868
rect 9640 37865 9646 37868
rect 11716 37865 11744 37964
rect 12526 37952 12532 37964
rect 12584 37952 12590 38004
rect 13630 37952 13636 38004
rect 13688 37992 13694 38004
rect 15013 37995 15071 38001
rect 15013 37992 15025 37995
rect 13688 37964 15025 37992
rect 13688 37952 13694 37964
rect 15013 37961 15025 37964
rect 15059 37961 15071 37995
rect 15013 37955 15071 37961
rect 15381 37995 15439 38001
rect 15381 37961 15393 37995
rect 15427 37992 15439 37995
rect 15470 37992 15476 38004
rect 15427 37964 15476 37992
rect 15427 37961 15439 37964
rect 15381 37955 15439 37961
rect 15470 37952 15476 37964
rect 15528 37952 15534 38004
rect 18138 37992 18144 38004
rect 17144 37964 18144 37992
rect 13998 37924 14004 37936
rect 13556 37896 14004 37924
rect 9640 37859 9668 37865
rect 9656 37825 9668 37859
rect 9640 37819 9668 37825
rect 11701 37859 11759 37865
rect 11701 37825 11713 37859
rect 11747 37825 11759 37859
rect 11701 37819 11759 37825
rect 9640 37816 9646 37819
rect 12434 37816 12440 37868
rect 12492 37816 12498 37868
rect 13556 37865 13584 37896
rect 13998 37884 14004 37896
rect 14056 37884 14062 37936
rect 13814 37865 13820 37868
rect 13541 37859 13599 37865
rect 13541 37825 13553 37859
rect 13587 37825 13599 37859
rect 13808 37856 13820 37865
rect 13775 37828 13820 37856
rect 13541 37819 13599 37825
rect 13808 37819 13820 37828
rect 13814 37816 13820 37819
rect 13872 37816 13878 37868
rect 16945 37859 17003 37865
rect 16945 37825 16957 37859
rect 16991 37856 17003 37859
rect 17034 37856 17040 37868
rect 16991 37828 17040 37856
rect 16991 37825 17003 37828
rect 16945 37819 17003 37825
rect 17034 37816 17040 37828
rect 17092 37816 17098 37868
rect 17144 37865 17172 37964
rect 18138 37952 18144 37964
rect 18196 37952 18202 38004
rect 18414 37952 18420 38004
rect 18472 37992 18478 38004
rect 19794 37992 19800 38004
rect 18472 37964 19800 37992
rect 18472 37952 18478 37964
rect 19794 37952 19800 37964
rect 19852 37952 19858 38004
rect 20162 37952 20168 38004
rect 20220 37992 20226 38004
rect 20993 37995 21051 38001
rect 20993 37992 21005 37995
rect 20220 37964 21005 37992
rect 20220 37952 20226 37964
rect 20993 37961 21005 37964
rect 21039 37961 21051 37995
rect 23106 37992 23112 38004
rect 20993 37955 21051 37961
rect 21652 37964 23112 37992
rect 19334 37933 19340 37936
rect 19328 37924 19340 37933
rect 19295 37896 19340 37924
rect 19328 37887 19340 37896
rect 19334 37884 19340 37887
rect 19392 37884 19398 37936
rect 20901 37927 20959 37933
rect 20901 37893 20913 37927
rect 20947 37924 20959 37927
rect 21450 37924 21456 37936
rect 20947 37896 21456 37924
rect 20947 37893 20959 37896
rect 20901 37887 20959 37893
rect 21450 37884 21456 37896
rect 21508 37884 21514 37936
rect 17129 37859 17187 37865
rect 17129 37825 17141 37859
rect 17175 37825 17187 37859
rect 17129 37819 17187 37825
rect 17862 37816 17868 37868
rect 17920 37816 17926 37868
rect 17954 37816 17960 37868
rect 18012 37865 18018 37868
rect 18012 37859 18040 37865
rect 18028 37825 18040 37859
rect 18012 37819 18040 37825
rect 18012 37816 18018 37819
rect 19058 37816 19064 37868
rect 19116 37816 19122 37868
rect 21652 37865 21680 37964
rect 23106 37952 23112 37964
rect 23164 37952 23170 38004
rect 26513 37995 26571 38001
rect 26513 37961 26525 37995
rect 26559 37992 26571 37995
rect 26602 37992 26608 38004
rect 26559 37964 26608 37992
rect 26559 37961 26571 37964
rect 26513 37955 26571 37961
rect 26602 37952 26608 37964
rect 26660 37952 26666 38004
rect 29733 37995 29791 38001
rect 27172 37964 29408 37992
rect 22002 37924 22008 37936
rect 21836 37896 22008 37924
rect 21836 37865 21864 37896
rect 22002 37884 22008 37896
rect 22060 37884 22066 37936
rect 26142 37884 26148 37936
rect 26200 37924 26206 37936
rect 27172 37924 27200 37964
rect 27798 37924 27804 37936
rect 26200 37896 27200 37924
rect 27264 37896 27804 37924
rect 26200 37884 26206 37896
rect 21637 37859 21695 37865
rect 19168 37828 20576 37856
rect 5626 37748 5632 37800
rect 5684 37788 5690 37800
rect 6365 37791 6423 37797
rect 6365 37788 6377 37791
rect 5684 37760 6377 37788
rect 5684 37748 5690 37760
rect 6365 37757 6377 37760
rect 6411 37757 6423 37791
rect 9490 37788 9496 37800
rect 6365 37751 6423 37757
rect 7760 37760 9496 37788
rect 3513 37655 3571 37661
rect 3513 37621 3525 37655
rect 3559 37652 3571 37655
rect 4062 37652 4068 37664
rect 3559 37624 4068 37652
rect 3559 37621 3571 37624
rect 3513 37615 3571 37621
rect 4062 37612 4068 37624
rect 4120 37612 4126 37664
rect 5166 37612 5172 37664
rect 5224 37612 5230 37664
rect 6380 37652 6408 37751
rect 7760 37732 7788 37760
rect 9490 37748 9496 37760
rect 9548 37748 9554 37800
rect 9769 37791 9827 37797
rect 9769 37757 9781 37791
rect 9815 37788 9827 37791
rect 10318 37788 10324 37800
rect 9815 37760 10324 37788
rect 9815 37757 9827 37760
rect 9769 37751 9827 37757
rect 10318 37748 10324 37760
rect 10376 37748 10382 37800
rect 10502 37748 10508 37800
rect 10560 37788 10566 37800
rect 11057 37791 11115 37797
rect 11057 37788 11069 37791
rect 10560 37760 11069 37788
rect 10560 37748 10566 37760
rect 11057 37757 11069 37760
rect 11103 37757 11115 37791
rect 11057 37751 11115 37757
rect 11238 37748 11244 37800
rect 11296 37788 11302 37800
rect 11517 37791 11575 37797
rect 11517 37788 11529 37791
rect 11296 37760 11529 37788
rect 11296 37748 11302 37760
rect 11517 37757 11529 37760
rect 11563 37788 11575 37791
rect 11882 37788 11888 37800
rect 11563 37760 11888 37788
rect 11563 37757 11575 37760
rect 11517 37751 11575 37757
rect 11882 37748 11888 37760
rect 11940 37748 11946 37800
rect 12066 37748 12072 37800
rect 12124 37788 12130 37800
rect 12554 37791 12612 37797
rect 12554 37788 12566 37791
rect 12124 37760 12566 37788
rect 12124 37748 12130 37760
rect 7742 37680 7748 37732
rect 7800 37680 7806 37732
rect 9214 37680 9220 37732
rect 9272 37680 9278 37732
rect 11422 37720 11428 37732
rect 10152 37692 11428 37720
rect 10152 37652 10180 37692
rect 11422 37680 11428 37692
rect 11480 37680 11486 37732
rect 12161 37723 12219 37729
rect 12161 37689 12173 37723
rect 12207 37689 12219 37723
rect 12161 37683 12219 37689
rect 6380 37624 10180 37652
rect 10413 37655 10471 37661
rect 10413 37621 10425 37655
rect 10459 37652 10471 37655
rect 10870 37652 10876 37664
rect 10459 37624 10876 37652
rect 10459 37621 10471 37624
rect 10413 37615 10471 37621
rect 10870 37612 10876 37624
rect 10928 37612 10934 37664
rect 11054 37612 11060 37664
rect 11112 37652 11118 37664
rect 12176 37652 12204 37683
rect 12268 37664 12296 37760
rect 12554 37757 12566 37760
rect 12600 37757 12612 37791
rect 12554 37751 12612 37757
rect 12713 37791 12771 37797
rect 12713 37757 12725 37791
rect 12759 37788 12771 37791
rect 13078 37788 13084 37800
rect 12759 37760 13084 37788
rect 12759 37757 12771 37760
rect 12713 37751 12771 37757
rect 13078 37748 13084 37760
rect 13136 37748 13142 37800
rect 14734 37748 14740 37800
rect 14792 37788 14798 37800
rect 15473 37791 15531 37797
rect 15473 37788 15485 37791
rect 14792 37760 15485 37788
rect 14792 37748 14798 37760
rect 15473 37757 15485 37760
rect 15519 37757 15531 37791
rect 15473 37751 15531 37757
rect 15657 37791 15715 37797
rect 15657 37757 15669 37791
rect 15703 37788 15715 37791
rect 17218 37788 17224 37800
rect 15703 37760 17224 37788
rect 15703 37757 15715 37760
rect 15657 37751 15715 37757
rect 17218 37748 17224 37760
rect 17276 37748 17282 37800
rect 17494 37748 17500 37800
rect 17552 37788 17558 37800
rect 17589 37791 17647 37797
rect 17589 37788 17601 37791
rect 17552 37760 17601 37788
rect 17552 37748 17558 37760
rect 17589 37757 17601 37760
rect 17635 37788 17647 37791
rect 17678 37788 17684 37800
rect 17635 37760 17684 37788
rect 17635 37757 17647 37760
rect 17589 37751 17647 37757
rect 17678 37748 17684 37760
rect 17736 37748 17742 37800
rect 18141 37791 18199 37797
rect 18141 37757 18153 37791
rect 18187 37788 18199 37791
rect 18322 37788 18328 37800
rect 18187 37760 18328 37788
rect 18187 37757 18199 37760
rect 18141 37751 18199 37757
rect 18322 37748 18328 37760
rect 18380 37788 18386 37800
rect 19168 37788 19196 37828
rect 18380 37760 19196 37788
rect 18380 37748 18386 37760
rect 14844 37692 17356 37720
rect 11112 37624 12204 37652
rect 11112 37612 11118 37624
rect 12250 37612 12256 37664
rect 12308 37612 12314 37664
rect 13357 37655 13415 37661
rect 13357 37621 13369 37655
rect 13403 37652 13415 37655
rect 14844 37652 14872 37692
rect 13403 37624 14872 37652
rect 13403 37621 13415 37624
rect 13357 37615 13415 37621
rect 14918 37612 14924 37664
rect 14976 37612 14982 37664
rect 17328 37652 17356 37692
rect 18598 37652 18604 37664
rect 17328 37624 18604 37652
rect 18598 37612 18604 37624
rect 18656 37612 18662 37664
rect 18690 37612 18696 37664
rect 18748 37652 18754 37664
rect 18785 37655 18843 37661
rect 18785 37652 18797 37655
rect 18748 37624 18797 37652
rect 18748 37612 18754 37624
rect 18785 37621 18797 37624
rect 18831 37621 18843 37655
rect 18785 37615 18843 37621
rect 20438 37612 20444 37664
rect 20496 37612 20502 37664
rect 20548 37652 20576 37828
rect 21637 37825 21649 37859
rect 21683 37825 21695 37859
rect 21637 37819 21695 37825
rect 21821 37859 21879 37865
rect 21821 37825 21833 37859
rect 21867 37825 21879 37859
rect 21821 37819 21879 37825
rect 21174 37748 21180 37800
rect 21232 37788 21238 37800
rect 21836 37788 21864 37819
rect 22738 37816 22744 37868
rect 22796 37816 22802 37868
rect 24397 37859 24455 37865
rect 24397 37825 24409 37859
rect 24443 37856 24455 37859
rect 24486 37856 24492 37868
rect 24443 37828 24492 37856
rect 24443 37825 24455 37828
rect 24397 37819 24455 37825
rect 24486 37816 24492 37828
rect 24544 37816 24550 37868
rect 25314 37816 25320 37868
rect 25372 37816 25378 37868
rect 26694 37816 26700 37868
rect 26752 37816 26758 37868
rect 27264 37865 27292 37896
rect 27798 37884 27804 37896
rect 27856 37884 27862 37936
rect 27249 37859 27307 37865
rect 27249 37825 27261 37859
rect 27295 37825 27307 37859
rect 27249 37819 27307 37825
rect 27614 37816 27620 37868
rect 27672 37816 27678 37868
rect 27724 37828 27936 37856
rect 21232 37760 21864 37788
rect 21232 37748 21238 37760
rect 21910 37748 21916 37800
rect 21968 37788 21974 37800
rect 22005 37791 22063 37797
rect 22005 37788 22017 37791
rect 21968 37760 22017 37788
rect 21968 37748 21974 37760
rect 22005 37757 22017 37760
rect 22051 37757 22063 37791
rect 22005 37751 22063 37757
rect 22830 37748 22836 37800
rect 22888 37797 22894 37800
rect 22888 37791 22916 37797
rect 22904 37757 22916 37791
rect 22888 37751 22916 37757
rect 23017 37791 23075 37797
rect 23017 37757 23029 37791
rect 23063 37788 23075 37791
rect 23198 37788 23204 37800
rect 23063 37760 23204 37788
rect 23063 37757 23075 37760
rect 23017 37751 23075 37757
rect 22888 37748 22894 37751
rect 23198 37748 23204 37760
rect 23256 37748 23262 37800
rect 24578 37748 24584 37800
rect 24636 37788 24642 37800
rect 24946 37788 24952 37800
rect 24636 37760 24952 37788
rect 24636 37748 24642 37760
rect 24946 37748 24952 37760
rect 25004 37748 25010 37800
rect 25406 37788 25412 37800
rect 25464 37797 25470 37800
rect 25464 37791 25492 37797
rect 25148 37760 25412 37788
rect 21453 37723 21511 37729
rect 21453 37689 21465 37723
rect 21499 37720 21511 37723
rect 22094 37720 22100 37732
rect 21499 37692 22100 37720
rect 21499 37689 21511 37692
rect 21453 37683 21511 37689
rect 22094 37680 22100 37692
rect 22152 37680 22158 37732
rect 22462 37680 22468 37732
rect 22520 37680 22526 37732
rect 23566 37680 23572 37732
rect 23624 37720 23630 37732
rect 23624 37692 24992 37720
rect 23624 37680 23630 37692
rect 22370 37652 22376 37664
rect 20548 37624 22376 37652
rect 22370 37612 22376 37624
rect 22428 37612 22434 37664
rect 23658 37612 23664 37664
rect 23716 37612 23722 37664
rect 24964 37652 24992 37692
rect 25038 37680 25044 37732
rect 25096 37680 25102 37732
rect 25148 37652 25176 37760
rect 25406 37748 25412 37760
rect 25480 37757 25492 37791
rect 25464 37751 25492 37757
rect 25593 37791 25651 37797
rect 25593 37757 25605 37791
rect 25639 37788 25651 37791
rect 25958 37788 25964 37800
rect 25639 37760 25964 37788
rect 25639 37757 25651 37760
rect 25593 37751 25651 37757
rect 25464 37748 25470 37751
rect 25958 37748 25964 37760
rect 26016 37748 26022 37800
rect 26142 37748 26148 37800
rect 26200 37788 26206 37800
rect 27724 37788 27752 37828
rect 26200 37760 27752 37788
rect 27801 37791 27859 37797
rect 26200 37748 26206 37760
rect 27801 37757 27813 37791
rect 27847 37757 27859 37791
rect 27801 37751 27859 37757
rect 24964 37624 25176 37652
rect 26237 37655 26295 37661
rect 26237 37621 26249 37655
rect 26283 37652 26295 37655
rect 26418 37652 26424 37664
rect 26283 37624 26424 37652
rect 26283 37621 26295 37624
rect 26237 37615 26295 37621
rect 26418 37612 26424 37624
rect 26476 37612 26482 37664
rect 27062 37612 27068 37664
rect 27120 37612 27126 37664
rect 27816 37652 27844 37751
rect 27908 37720 27936 37828
rect 28166 37748 28172 37800
rect 28224 37788 28230 37800
rect 28718 37797 28724 37800
rect 28537 37791 28595 37797
rect 28537 37788 28549 37791
rect 28224 37760 28549 37788
rect 28224 37748 28230 37760
rect 28537 37757 28549 37760
rect 28583 37757 28595 37791
rect 28537 37751 28595 37757
rect 28675 37791 28724 37797
rect 28675 37757 28687 37791
rect 28721 37757 28724 37791
rect 28675 37751 28724 37757
rect 28718 37748 28724 37751
rect 28776 37748 28782 37800
rect 28813 37791 28871 37797
rect 28813 37757 28825 37791
rect 28859 37788 28871 37791
rect 29380 37788 29408 37964
rect 29733 37961 29745 37995
rect 29779 37992 29791 37995
rect 29822 37992 29828 38004
rect 29779 37964 29828 37992
rect 29779 37961 29791 37964
rect 29733 37955 29791 37961
rect 29822 37952 29828 37964
rect 29880 37952 29886 38004
rect 30282 37952 30288 38004
rect 30340 37992 30346 38004
rect 30653 37995 30711 38001
rect 30653 37992 30665 37995
rect 30340 37964 30665 37992
rect 30340 37952 30346 37964
rect 30653 37961 30665 37964
rect 30699 37961 30711 37995
rect 30653 37955 30711 37961
rect 31570 37952 31576 38004
rect 31628 37992 31634 38004
rect 32125 37995 32183 38001
rect 32125 37992 32137 37995
rect 31628 37964 32137 37992
rect 31628 37952 31634 37964
rect 32125 37961 32137 37964
rect 32171 37961 32183 37995
rect 32125 37955 32183 37961
rect 32490 37952 32496 38004
rect 32548 37952 32554 38004
rect 32585 37995 32643 38001
rect 32585 37961 32597 37995
rect 32631 37992 32643 37995
rect 32858 37992 32864 38004
rect 32631 37964 32864 37992
rect 32631 37961 32643 37964
rect 32585 37955 32643 37961
rect 32858 37952 32864 37964
rect 32916 37952 32922 38004
rect 33318 37952 33324 38004
rect 33376 37952 33382 38004
rect 36170 37952 36176 38004
rect 36228 37992 36234 38004
rect 36228 37964 37136 37992
rect 36228 37952 36234 37964
rect 33226 37884 33232 37936
rect 33284 37884 33290 37936
rect 29914 37816 29920 37868
rect 29972 37816 29978 37868
rect 30561 37859 30619 37865
rect 30561 37825 30573 37859
rect 30607 37856 30619 37859
rect 30742 37856 30748 37868
rect 30607 37828 30748 37856
rect 30607 37825 30619 37828
rect 30561 37819 30619 37825
rect 30742 37816 30748 37828
rect 30800 37816 30806 37868
rect 36464 37865 36492 37964
rect 36722 37924 36728 37936
rect 36648 37896 36728 37924
rect 36449 37859 36507 37865
rect 36449 37825 36461 37859
rect 36495 37825 36507 37859
rect 36449 37819 36507 37825
rect 36538 37816 36544 37868
rect 36596 37816 36602 37868
rect 36648 37865 36676 37896
rect 36722 37884 36728 37896
rect 36780 37924 36786 37936
rect 36998 37924 37004 37936
rect 36780 37896 37004 37924
rect 36780 37884 36786 37896
rect 36998 37884 37004 37896
rect 37056 37884 37062 37936
rect 36633 37859 36691 37865
rect 36633 37825 36645 37859
rect 36679 37825 36691 37859
rect 36633 37819 36691 37825
rect 36814 37816 36820 37868
rect 36872 37816 36878 37868
rect 37108 37856 37136 37964
rect 37458 37952 37464 38004
rect 37516 38001 37522 38004
rect 37516 37995 37535 38001
rect 37523 37992 37535 37995
rect 37523 37964 37780 37992
rect 37523 37961 37535 37964
rect 37516 37955 37535 37961
rect 37516 37952 37522 37955
rect 37274 37884 37280 37936
rect 37332 37884 37338 37936
rect 37752 37924 37780 37964
rect 39574 37952 39580 38004
rect 39632 37952 39638 38004
rect 38442 37927 38500 37933
rect 38442 37924 38454 37927
rect 37752 37896 38454 37924
rect 38442 37893 38454 37896
rect 38488 37893 38500 37927
rect 38442 37887 38500 37893
rect 38746 37856 38752 37868
rect 37108 37828 38752 37856
rect 38746 37816 38752 37828
rect 38804 37816 38810 37868
rect 44174 37816 44180 37868
rect 44232 37856 44238 37868
rect 46477 37859 46535 37865
rect 46477 37856 46489 37859
rect 44232 37828 46489 37856
rect 44232 37816 44238 37828
rect 46477 37825 46489 37828
rect 46523 37825 46535 37859
rect 46477 37819 46535 37825
rect 28859 37760 29408 37788
rect 30837 37791 30895 37797
rect 28859 37757 28871 37760
rect 28813 37751 28871 37757
rect 30837 37757 30849 37791
rect 30883 37788 30895 37791
rect 32582 37788 32588 37800
rect 30883 37760 32588 37788
rect 30883 37757 30895 37760
rect 30837 37751 30895 37757
rect 32582 37748 32588 37760
rect 32640 37788 32646 37800
rect 32677 37791 32735 37797
rect 32677 37788 32689 37791
rect 32640 37760 32689 37788
rect 32640 37748 32646 37760
rect 32677 37757 32689 37760
rect 32723 37757 32735 37791
rect 32677 37751 32735 37757
rect 34422 37748 34428 37800
rect 34480 37788 34486 37800
rect 38010 37788 38016 37800
rect 34480 37760 38016 37788
rect 34480 37748 34486 37760
rect 38010 37748 38016 37760
rect 38068 37788 38074 37800
rect 38197 37791 38255 37797
rect 38197 37788 38209 37791
rect 38068 37760 38209 37788
rect 38068 37748 38074 37760
rect 38197 37757 38209 37760
rect 38243 37757 38255 37791
rect 38197 37751 38255 37757
rect 28261 37723 28319 37729
rect 28261 37720 28273 37723
rect 27908 37692 28273 37720
rect 28261 37689 28273 37692
rect 28307 37689 28319 37723
rect 37918 37720 37924 37732
rect 28261 37683 28319 37689
rect 37476 37692 37924 37720
rect 27890 37652 27896 37664
rect 27816 37624 27896 37652
rect 27890 37612 27896 37624
rect 27948 37652 27954 37664
rect 28902 37652 28908 37664
rect 27948 37624 28908 37652
rect 27948 37612 27954 37624
rect 28902 37612 28908 37624
rect 28960 37612 28966 37664
rect 28994 37612 29000 37664
rect 29052 37652 29058 37664
rect 29457 37655 29515 37661
rect 29457 37652 29469 37655
rect 29052 37624 29469 37652
rect 29052 37612 29058 37624
rect 29457 37621 29469 37624
rect 29503 37621 29515 37655
rect 29457 37615 29515 37621
rect 29914 37612 29920 37664
rect 29972 37652 29978 37664
rect 30193 37655 30251 37661
rect 30193 37652 30205 37655
rect 29972 37624 30205 37652
rect 29972 37612 29978 37624
rect 30193 37621 30205 37624
rect 30239 37621 30251 37655
rect 30193 37615 30251 37621
rect 36170 37612 36176 37664
rect 36228 37612 36234 37664
rect 37476 37661 37504 37692
rect 37918 37680 37924 37692
rect 37976 37680 37982 37732
rect 37461 37655 37519 37661
rect 37461 37621 37473 37655
rect 37507 37621 37519 37655
rect 37461 37615 37519 37621
rect 37642 37612 37648 37664
rect 37700 37612 37706 37664
rect 46658 37612 46664 37664
rect 46716 37612 46722 37664
rect 1104 37562 47104 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 47104 37562
rect 1104 37488 47104 37510
rect 5258 37408 5264 37460
rect 5316 37408 5322 37460
rect 10502 37448 10508 37460
rect 5920 37420 10508 37448
rect 3786 37272 3792 37324
rect 3844 37272 3850 37324
rect 5920 37321 5948 37420
rect 10502 37408 10508 37420
rect 10560 37408 10566 37460
rect 10781 37451 10839 37457
rect 10781 37417 10793 37451
rect 10827 37448 10839 37451
rect 13173 37451 13231 37457
rect 10827 37420 12848 37448
rect 10827 37417 10839 37420
rect 10781 37411 10839 37417
rect 6273 37383 6331 37389
rect 6273 37349 6285 37383
rect 6319 37349 6331 37383
rect 6273 37343 6331 37349
rect 5905 37315 5963 37321
rect 5905 37281 5917 37315
rect 5951 37281 5963 37315
rect 5905 37275 5963 37281
rect 6288 37256 6316 37343
rect 6454 37340 6460 37392
rect 6512 37380 6518 37392
rect 6641 37383 6699 37389
rect 6641 37380 6653 37383
rect 6512 37352 6653 37380
rect 6512 37340 6518 37352
rect 6641 37349 6653 37352
rect 6687 37349 6699 37383
rect 9214 37380 9220 37392
rect 6641 37343 6699 37349
rect 7116 37352 9220 37380
rect 7116 37312 7144 37352
rect 6748 37284 7144 37312
rect 934 37204 940 37256
rect 992 37244 998 37256
rect 4062 37253 4068 37256
rect 1581 37247 1639 37253
rect 1581 37244 1593 37247
rect 992 37216 1593 37244
rect 992 37204 998 37216
rect 1581 37213 1593 37216
rect 1627 37213 1639 37247
rect 4056 37244 4068 37253
rect 4023 37216 4068 37244
rect 1581 37207 1639 37213
rect 4056 37207 4068 37216
rect 4062 37204 4068 37207
rect 4120 37204 4126 37256
rect 5166 37204 5172 37256
rect 5224 37244 5230 37256
rect 5629 37247 5687 37253
rect 5629 37244 5641 37247
rect 5224 37216 5641 37244
rect 5224 37204 5230 37216
rect 5629 37213 5641 37216
rect 5675 37213 5687 37247
rect 5629 37207 5687 37213
rect 6270 37204 6276 37256
rect 6328 37204 6334 37256
rect 6457 37247 6515 37253
rect 6457 37213 6469 37247
rect 6503 37244 6515 37247
rect 6638 37244 6644 37256
rect 6503 37216 6644 37244
rect 6503 37213 6515 37216
rect 6457 37207 6515 37213
rect 6638 37204 6644 37216
rect 6696 37204 6702 37256
rect 4706 37136 4712 37188
rect 4764 37176 4770 37188
rect 5184 37176 5212 37204
rect 4764 37148 5212 37176
rect 4764 37136 4770 37148
rect 5442 37136 5448 37188
rect 5500 37176 5506 37188
rect 6748 37176 6776 37284
rect 7190 37272 7196 37324
rect 7248 37272 7254 37324
rect 8220 37321 8248 37352
rect 9214 37340 9220 37352
rect 9272 37340 9278 37392
rect 9490 37340 9496 37392
rect 9548 37380 9554 37392
rect 9548 37352 9720 37380
rect 9548 37340 9554 37352
rect 8205 37315 8263 37321
rect 8205 37281 8217 37315
rect 8251 37281 8263 37315
rect 8205 37275 8263 37281
rect 8478 37272 8484 37324
rect 8536 37312 8542 37324
rect 8941 37315 8999 37321
rect 8941 37312 8953 37315
rect 8536 37284 8953 37312
rect 8536 37272 8542 37284
rect 8941 37281 8953 37284
rect 8987 37281 8999 37315
rect 8941 37275 8999 37281
rect 9306 37272 9312 37324
rect 9364 37312 9370 37324
rect 9582 37312 9588 37324
rect 9364 37284 9588 37312
rect 9364 37272 9370 37284
rect 9582 37272 9588 37284
rect 9640 37272 9646 37324
rect 9692 37312 9720 37352
rect 10686 37340 10692 37392
rect 10744 37380 10750 37392
rect 11885 37383 11943 37389
rect 11885 37380 11897 37383
rect 10744 37352 11897 37380
rect 10744 37340 10750 37352
rect 11885 37349 11897 37352
rect 11931 37349 11943 37383
rect 12820 37380 12848 37420
rect 13173 37417 13185 37451
rect 13219 37448 13231 37451
rect 13354 37448 13360 37460
rect 13219 37420 13360 37448
rect 13219 37417 13231 37420
rect 13173 37411 13231 37417
rect 13354 37408 13360 37420
rect 13412 37408 13418 37460
rect 13906 37408 13912 37460
rect 13964 37448 13970 37460
rect 14277 37451 14335 37457
rect 14277 37448 14289 37451
rect 13964 37420 14289 37448
rect 13964 37408 13970 37420
rect 14277 37417 14289 37420
rect 14323 37417 14335 37451
rect 14277 37411 14335 37417
rect 14826 37408 14832 37460
rect 14884 37448 14890 37460
rect 16206 37448 16212 37460
rect 14884 37420 16212 37448
rect 14884 37408 14890 37420
rect 16206 37408 16212 37420
rect 16264 37408 16270 37460
rect 19794 37408 19800 37460
rect 19852 37448 19858 37460
rect 23198 37448 23204 37460
rect 19852 37420 23204 37448
rect 19852 37408 19858 37420
rect 23198 37408 23204 37420
rect 23256 37408 23262 37460
rect 25038 37408 25044 37460
rect 25096 37448 25102 37460
rect 26142 37448 26148 37460
rect 25096 37420 26148 37448
rect 25096 37408 25102 37420
rect 26142 37408 26148 37420
rect 26200 37408 26206 37460
rect 26513 37451 26571 37457
rect 26513 37417 26525 37451
rect 26559 37448 26571 37451
rect 26694 37448 26700 37460
rect 26559 37420 26700 37448
rect 26559 37417 26571 37420
rect 26513 37411 26571 37417
rect 26694 37408 26700 37420
rect 26752 37408 26758 37460
rect 30742 37408 30748 37460
rect 30800 37448 30806 37460
rect 31389 37451 31447 37457
rect 31389 37448 31401 37451
rect 30800 37420 31401 37448
rect 30800 37408 30806 37420
rect 31389 37417 31401 37420
rect 31435 37417 31447 37451
rect 31389 37411 31447 37417
rect 19242 37380 19248 37392
rect 12820 37352 19248 37380
rect 11885 37343 11943 37349
rect 19242 37340 19248 37352
rect 19300 37340 19306 37392
rect 28074 37380 28080 37392
rect 27264 37352 28080 37380
rect 9861 37315 9919 37321
rect 9861 37312 9873 37315
rect 9692 37284 9873 37312
rect 9861 37281 9873 37284
rect 9907 37281 9919 37315
rect 9861 37275 9919 37281
rect 9950 37272 9956 37324
rect 10008 37321 10014 37324
rect 10008 37315 10036 37321
rect 10024 37281 10036 37315
rect 10008 37275 10036 37281
rect 10008 37272 10014 37275
rect 11238 37272 11244 37324
rect 11296 37272 11302 37324
rect 12158 37272 12164 37324
rect 12216 37272 12222 37324
rect 12250 37272 12256 37324
rect 12308 37321 12314 37324
rect 12308 37315 12336 37321
rect 12324 37281 12336 37315
rect 12308 37275 12336 37281
rect 12308 37272 12314 37275
rect 13078 37272 13084 37324
rect 13136 37272 13142 37324
rect 13725 37315 13783 37321
rect 13725 37281 13737 37315
rect 13771 37281 13783 37315
rect 13725 37275 13783 37281
rect 14829 37315 14887 37321
rect 14829 37281 14841 37315
rect 14875 37312 14887 37315
rect 15930 37312 15936 37324
rect 14875 37284 15936 37312
rect 14875 37281 14887 37284
rect 14829 37275 14887 37281
rect 7006 37204 7012 37256
rect 7064 37204 7070 37256
rect 8021 37247 8079 37253
rect 8021 37213 8033 37247
rect 8067 37244 8079 37247
rect 8496 37244 8524 37272
rect 8067 37216 8524 37244
rect 8067 37213 8079 37216
rect 8021 37207 8079 37213
rect 8754 37204 8760 37256
rect 8812 37244 8818 37256
rect 9125 37247 9183 37253
rect 9125 37244 9137 37247
rect 8812 37216 9137 37244
rect 8812 37204 8818 37216
rect 9125 37213 9137 37216
rect 9171 37213 9183 37247
rect 9125 37207 9183 37213
rect 10134 37204 10140 37256
rect 10192 37204 10198 37256
rect 11425 37247 11483 37253
rect 11425 37213 11437 37247
rect 11471 37213 11483 37247
rect 11425 37207 11483 37213
rect 5500 37148 6776 37176
rect 5500 37136 5506 37148
rect 7098 37136 7104 37188
rect 7156 37176 7162 37188
rect 7156 37148 8156 37176
rect 7156 37136 7162 37148
rect 1397 37111 1455 37117
rect 1397 37077 1409 37111
rect 1443 37108 1455 37111
rect 2406 37108 2412 37120
rect 1443 37080 2412 37108
rect 1443 37077 1455 37080
rect 1397 37071 1455 37077
rect 2406 37068 2412 37080
rect 2464 37068 2470 37120
rect 4430 37068 4436 37120
rect 4488 37108 4494 37120
rect 5169 37111 5227 37117
rect 5169 37108 5181 37111
rect 4488 37080 5181 37108
rect 4488 37068 4494 37080
rect 5169 37077 5181 37080
rect 5215 37077 5227 37111
rect 5169 37071 5227 37077
rect 5258 37068 5264 37120
rect 5316 37108 5322 37120
rect 5721 37111 5779 37117
rect 5721 37108 5733 37111
rect 5316 37080 5733 37108
rect 5316 37068 5322 37080
rect 5721 37077 5733 37080
rect 5767 37108 5779 37111
rect 7282 37108 7288 37120
rect 5767 37080 7288 37108
rect 5767 37077 5779 37080
rect 5721 37071 5779 37077
rect 7282 37068 7288 37080
rect 7340 37068 7346 37120
rect 7650 37068 7656 37120
rect 7708 37068 7714 37120
rect 8128 37117 8156 37148
rect 8113 37111 8171 37117
rect 8113 37077 8125 37111
rect 8159 37108 8171 37111
rect 10962 37108 10968 37120
rect 8159 37080 10968 37108
rect 8159 37077 8171 37080
rect 8113 37071 8171 37077
rect 10962 37068 10968 37080
rect 11020 37068 11026 37120
rect 11440 37108 11468 37207
rect 12434 37204 12440 37256
rect 12492 37204 12498 37256
rect 13740 37244 13768 37275
rect 15930 37272 15936 37284
rect 15988 37272 15994 37324
rect 17218 37272 17224 37324
rect 17276 37312 17282 37324
rect 17770 37312 17776 37324
rect 17276 37284 17776 37312
rect 17276 37272 17282 37284
rect 17770 37272 17776 37284
rect 17828 37272 17834 37324
rect 20165 37315 20223 37321
rect 20165 37281 20177 37315
rect 20211 37312 20223 37315
rect 21450 37312 21456 37324
rect 20211 37284 21456 37312
rect 20211 37281 20223 37284
rect 20165 37275 20223 37281
rect 21450 37272 21456 37284
rect 21508 37272 21514 37324
rect 22830 37312 22836 37324
rect 22204 37284 22836 37312
rect 22204 37256 22232 37284
rect 22830 37272 22836 37284
rect 22888 37272 22894 37324
rect 24397 37315 24455 37321
rect 24397 37281 24409 37315
rect 24443 37312 24455 37315
rect 24486 37312 24492 37324
rect 24443 37284 24492 37312
rect 24443 37281 24455 37284
rect 24397 37275 24455 37281
rect 24486 37272 24492 37284
rect 24544 37272 24550 37324
rect 24578 37272 24584 37324
rect 24636 37272 24642 37324
rect 25041 37315 25099 37321
rect 25041 37281 25053 37315
rect 25087 37312 25099 37315
rect 25130 37312 25136 37324
rect 25087 37284 25136 37312
rect 25087 37281 25099 37284
rect 25041 37275 25099 37281
rect 25130 37272 25136 37284
rect 25188 37272 25194 37324
rect 25314 37272 25320 37324
rect 25372 37272 25378 37324
rect 25406 37272 25412 37324
rect 25464 37321 25470 37324
rect 25464 37315 25492 37321
rect 25480 37281 25492 37315
rect 25464 37275 25492 37281
rect 25464 37272 25470 37275
rect 26234 37272 26240 37324
rect 26292 37272 26298 37324
rect 26786 37272 26792 37324
rect 26844 37312 26850 37324
rect 27065 37315 27123 37321
rect 27065 37312 27077 37315
rect 26844 37284 27077 37312
rect 26844 37272 26850 37284
rect 27065 37281 27077 37284
rect 27111 37281 27123 37315
rect 27065 37275 27123 37281
rect 14645 37247 14703 37253
rect 13740 37216 13952 37244
rect 13924 37176 13952 37216
rect 14645 37213 14657 37247
rect 14691 37244 14703 37247
rect 14918 37244 14924 37256
rect 14691 37216 14924 37244
rect 14691 37213 14703 37216
rect 14645 37207 14703 37213
rect 14918 37204 14924 37216
rect 14976 37244 14982 37256
rect 15654 37244 15660 37256
rect 14976 37216 15660 37244
rect 14976 37204 14982 37216
rect 15654 37204 15660 37216
rect 15712 37204 15718 37256
rect 19889 37247 19947 37253
rect 19889 37213 19901 37247
rect 19935 37244 19947 37247
rect 20438 37244 20444 37256
rect 19935 37216 20444 37244
rect 19935 37213 19947 37216
rect 19889 37207 19947 37213
rect 20438 37204 20444 37216
rect 20496 37244 20502 37256
rect 22186 37244 22192 37256
rect 20496 37216 22192 37244
rect 20496 37204 20502 37216
rect 22186 37204 22192 37216
rect 22244 37204 22250 37256
rect 22462 37204 22468 37256
rect 22520 37244 22526 37256
rect 24118 37244 24124 37256
rect 22520 37216 24124 37244
rect 22520 37204 22526 37216
rect 24118 37204 24124 37216
rect 24176 37204 24182 37256
rect 25590 37204 25596 37256
rect 25648 37204 25654 37256
rect 27264 37244 27292 37352
rect 28074 37340 28080 37352
rect 28132 37340 28138 37392
rect 35802 37340 35808 37392
rect 35860 37380 35866 37392
rect 35860 37352 38976 37380
rect 35860 37340 35866 37352
rect 27614 37312 27620 37324
rect 27448 37284 27620 37312
rect 26804 37216 27292 37244
rect 27341 37247 27399 37253
rect 15286 37176 15292 37188
rect 13924 37148 15292 37176
rect 15286 37136 15292 37148
rect 15344 37136 15350 37188
rect 19981 37179 20039 37185
rect 19981 37145 19993 37179
rect 20027 37176 20039 37179
rect 20162 37176 20168 37188
rect 20027 37148 20168 37176
rect 20027 37145 20039 37148
rect 19981 37139 20039 37145
rect 20162 37136 20168 37148
rect 20220 37136 20226 37188
rect 12526 37108 12532 37120
rect 11440 37080 12532 37108
rect 12526 37068 12532 37080
rect 12584 37108 12590 37120
rect 13541 37111 13599 37117
rect 13541 37108 13553 37111
rect 12584 37080 13553 37108
rect 12584 37068 12590 37080
rect 13541 37077 13553 37080
rect 13587 37077 13599 37111
rect 13541 37071 13599 37077
rect 13633 37111 13691 37117
rect 13633 37077 13645 37111
rect 13679 37108 13691 37111
rect 14090 37108 14096 37120
rect 13679 37080 14096 37108
rect 13679 37077 13691 37080
rect 13633 37071 13691 37077
rect 14090 37068 14096 37080
rect 14148 37068 14154 37120
rect 14274 37068 14280 37120
rect 14332 37108 14338 37120
rect 14734 37108 14740 37120
rect 14332 37080 14740 37108
rect 14332 37068 14338 37080
rect 14734 37068 14740 37080
rect 14792 37068 14798 37120
rect 19518 37068 19524 37120
rect 19576 37068 19582 37120
rect 23750 37068 23756 37120
rect 23808 37108 23814 37120
rect 26804 37108 26832 37216
rect 27341 37213 27353 37247
rect 27387 37244 27399 37247
rect 27448 37244 27476 37284
rect 27614 37272 27620 37284
rect 27672 37272 27678 37324
rect 27890 37312 27896 37324
rect 27724 37284 27896 37312
rect 27387 37216 27476 37244
rect 27525 37247 27583 37253
rect 27387 37213 27399 37216
rect 27341 37207 27399 37213
rect 27525 37213 27537 37247
rect 27571 37244 27583 37247
rect 27724 37244 27752 37284
rect 27890 37272 27896 37284
rect 27948 37272 27954 37324
rect 27982 37272 27988 37324
rect 28040 37272 28046 37324
rect 28258 37272 28264 37324
rect 28316 37272 28322 37324
rect 28350 37272 28356 37324
rect 28408 37321 28414 37324
rect 28408 37315 28436 37321
rect 28424 37312 28436 37315
rect 28718 37312 28724 37324
rect 28424 37284 28724 37312
rect 28424 37281 28436 37284
rect 28408 37275 28436 37281
rect 28408 37272 28414 37275
rect 28718 37272 28724 37284
rect 28776 37272 28782 37324
rect 29178 37272 29184 37324
rect 29236 37272 29242 37324
rect 31662 37272 31668 37324
rect 31720 37312 31726 37324
rect 38948 37321 38976 37352
rect 33965 37315 34023 37321
rect 33965 37312 33977 37315
rect 31720 37284 33977 37312
rect 31720 37272 31726 37284
rect 33965 37281 33977 37284
rect 34011 37312 34023 37315
rect 38933 37315 38991 37321
rect 34011 37284 34744 37312
rect 34011 37281 34023 37284
rect 33965 37275 34023 37281
rect 27571 37216 27752 37244
rect 27571 37213 27583 37216
rect 27525 37207 27583 37213
rect 28534 37204 28540 37256
rect 28592 37204 28598 37256
rect 29914 37204 29920 37256
rect 29972 37204 29978 37256
rect 30009 37247 30067 37253
rect 30009 37213 30021 37247
rect 30055 37244 30067 37247
rect 31680 37244 31708 37272
rect 30055 37216 31708 37244
rect 30055 37213 30067 37216
rect 30009 37207 30067 37213
rect 33134 37204 33140 37256
rect 33192 37244 33198 37256
rect 33781 37247 33839 37253
rect 33781 37244 33793 37247
rect 33192 37216 33793 37244
rect 33192 37204 33198 37216
rect 33781 37213 33793 37216
rect 33827 37244 33839 37247
rect 34422 37244 34428 37256
rect 33827 37216 34428 37244
rect 33827 37213 33839 37216
rect 33781 37207 33839 37213
rect 34422 37204 34428 37216
rect 34480 37204 34486 37256
rect 34716 37253 34744 37284
rect 36648 37284 36860 37312
rect 34701 37247 34759 37253
rect 34701 37213 34713 37247
rect 34747 37213 34759 37247
rect 34701 37207 34759 37213
rect 36449 37247 36507 37253
rect 36449 37213 36461 37247
rect 36495 37244 36507 37247
rect 36648 37244 36676 37284
rect 36495 37216 36676 37244
rect 36495 37213 36507 37216
rect 36449 37207 36507 37213
rect 36722 37204 36728 37256
rect 36780 37204 36786 37256
rect 36832 37244 36860 37284
rect 38933 37281 38945 37315
rect 38979 37281 38991 37315
rect 38933 37275 38991 37281
rect 37366 37244 37372 37256
rect 36832 37216 37372 37244
rect 37366 37204 37372 37216
rect 37424 37204 37430 37256
rect 39393 37247 39451 37253
rect 39393 37244 39405 37247
rect 38396 37216 39405 37244
rect 26881 37179 26939 37185
rect 26881 37145 26893 37179
rect 26927 37176 26939 37179
rect 30254 37179 30312 37185
rect 30254 37176 30266 37179
rect 26927 37148 27568 37176
rect 26927 37145 26939 37148
rect 26881 37139 26939 37145
rect 26973 37111 27031 37117
rect 26973 37108 26985 37111
rect 23808 37080 26985 37108
rect 23808 37068 23814 37080
rect 26973 37077 26985 37080
rect 27019 37077 27031 37111
rect 27540 37108 27568 37148
rect 29748 37148 30266 37176
rect 27706 37108 27712 37120
rect 27540 37080 27712 37108
rect 26973 37071 27031 37077
rect 27706 37068 27712 37080
rect 27764 37108 27770 37120
rect 28350 37108 28356 37120
rect 27764 37080 28356 37108
rect 27764 37068 27770 37080
rect 28350 37068 28356 37080
rect 28408 37068 28414 37120
rect 29748 37117 29776 37148
rect 30254 37145 30266 37148
rect 30300 37145 30312 37179
rect 30254 37139 30312 37145
rect 34514 37136 34520 37188
rect 34572 37176 34578 37188
rect 34946 37179 35004 37185
rect 34946 37176 34958 37179
rect 34572 37148 34958 37176
rect 34572 37136 34578 37148
rect 34946 37145 34958 37148
rect 34992 37145 35004 37179
rect 34946 37139 35004 37145
rect 36633 37179 36691 37185
rect 36633 37145 36645 37179
rect 36679 37176 36691 37179
rect 37182 37176 37188 37188
rect 36679 37148 37188 37176
rect 36679 37145 36691 37148
rect 36633 37139 36691 37145
rect 37182 37136 37188 37148
rect 37240 37136 37246 37188
rect 29733 37111 29791 37117
rect 29733 37077 29745 37111
rect 29779 37077 29791 37111
rect 29733 37071 29791 37077
rect 36078 37068 36084 37120
rect 36136 37068 36142 37120
rect 36538 37068 36544 37120
rect 36596 37117 36602 37120
rect 38396 37117 38424 37216
rect 39393 37213 39405 37216
rect 39439 37213 39451 37247
rect 39393 37207 39451 37213
rect 36596 37071 36605 37117
rect 38381 37111 38439 37117
rect 38381 37077 38393 37111
rect 38427 37077 38439 37111
rect 38381 37071 38439 37077
rect 36596 37068 36602 37071
rect 38562 37068 38568 37120
rect 38620 37108 38626 37120
rect 38749 37111 38807 37117
rect 38749 37108 38761 37111
rect 38620 37080 38761 37108
rect 38620 37068 38626 37080
rect 38749 37077 38761 37080
rect 38795 37077 38807 37111
rect 38749 37071 38807 37077
rect 38838 37068 38844 37120
rect 38896 37068 38902 37120
rect 39206 37068 39212 37120
rect 39264 37068 39270 37120
rect 1104 37018 47104 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 47104 37018
rect 1104 36944 47104 36966
rect 3694 36864 3700 36916
rect 3752 36904 3758 36916
rect 4065 36907 4123 36913
rect 4065 36904 4077 36907
rect 3752 36876 4077 36904
rect 3752 36864 3758 36876
rect 4065 36873 4077 36876
rect 4111 36873 4123 36907
rect 4065 36867 4123 36873
rect 4430 36864 4436 36916
rect 4488 36864 4494 36916
rect 4525 36907 4583 36913
rect 4525 36873 4537 36907
rect 4571 36904 4583 36907
rect 5258 36904 5264 36916
rect 4571 36876 5264 36904
rect 4571 36873 4583 36876
rect 4525 36867 4583 36873
rect 5258 36864 5264 36876
rect 5316 36864 5322 36916
rect 6638 36864 6644 36916
rect 6696 36864 6702 36916
rect 7009 36907 7067 36913
rect 7009 36873 7021 36907
rect 7055 36904 7067 36907
rect 7742 36904 7748 36916
rect 7055 36876 7748 36904
rect 7055 36873 7067 36876
rect 7009 36867 7067 36873
rect 7742 36864 7748 36876
rect 7800 36864 7806 36916
rect 10318 36864 10324 36916
rect 10376 36904 10382 36916
rect 12434 36904 12440 36916
rect 10376 36876 12440 36904
rect 10376 36864 10382 36876
rect 12434 36864 12440 36876
rect 12492 36864 12498 36916
rect 16482 36864 16488 36916
rect 16540 36904 16546 36916
rect 16669 36907 16727 36913
rect 16669 36904 16681 36907
rect 16540 36876 16681 36904
rect 16540 36864 16546 36876
rect 16669 36873 16681 36876
rect 16715 36873 16727 36907
rect 16669 36867 16727 36873
rect 16850 36864 16856 36916
rect 16908 36904 16914 36916
rect 17129 36907 17187 36913
rect 17129 36904 17141 36907
rect 16908 36876 17141 36904
rect 16908 36864 16914 36876
rect 17129 36873 17141 36876
rect 17175 36904 17187 36907
rect 17175 36876 27384 36904
rect 17175 36873 17187 36876
rect 17129 36867 17187 36873
rect 7098 36796 7104 36848
rect 7156 36796 7162 36848
rect 7282 36796 7288 36848
rect 7340 36836 7346 36848
rect 14458 36836 14464 36848
rect 7340 36808 14464 36836
rect 7340 36796 7346 36808
rect 14458 36796 14464 36808
rect 14516 36796 14522 36848
rect 16758 36796 16764 36848
rect 16816 36836 16822 36848
rect 16816 36808 20484 36836
rect 16816 36796 16822 36808
rect 16493 36780 16551 36781
rect 6914 36728 6920 36780
rect 6972 36768 6978 36780
rect 10134 36768 10140 36780
rect 6972 36740 10140 36768
rect 6972 36728 6978 36740
rect 10134 36728 10140 36740
rect 10192 36768 10198 36780
rect 12986 36768 12992 36780
rect 10192 36740 12992 36768
rect 10192 36728 10198 36740
rect 12986 36728 12992 36740
rect 13044 36728 13050 36780
rect 16482 36728 16488 36780
rect 16540 36735 16551 36780
rect 17037 36771 17095 36777
rect 17037 36737 17049 36771
rect 17083 36768 17095 36771
rect 17954 36768 17960 36780
rect 17083 36740 17960 36768
rect 17083 36737 17095 36740
rect 16540 36728 16546 36735
rect 17037 36731 17095 36737
rect 4709 36703 4767 36709
rect 4709 36669 4721 36703
rect 4755 36700 4767 36703
rect 5442 36700 5448 36712
rect 4755 36672 5448 36700
rect 4755 36669 4767 36672
rect 4709 36663 4767 36669
rect 5442 36660 5448 36672
rect 5500 36660 5506 36712
rect 7285 36703 7343 36709
rect 7285 36669 7297 36703
rect 7331 36700 7343 36703
rect 8202 36700 8208 36712
rect 7331 36672 8208 36700
rect 7331 36669 7343 36672
rect 7285 36663 7343 36669
rect 8202 36660 8208 36672
rect 8260 36660 8266 36712
rect 15838 36660 15844 36712
rect 15896 36700 15902 36712
rect 17052 36700 17080 36731
rect 17954 36728 17960 36740
rect 18012 36728 18018 36780
rect 15896 36672 17080 36700
rect 17313 36703 17371 36709
rect 15896 36660 15902 36672
rect 17313 36669 17325 36703
rect 17359 36700 17371 36703
rect 19150 36700 19156 36712
rect 17359 36672 19156 36700
rect 17359 36669 17371 36672
rect 17313 36663 17371 36669
rect 19150 36660 19156 36672
rect 19208 36660 19214 36712
rect 19245 36703 19303 36709
rect 19245 36669 19257 36703
rect 19291 36700 19303 36703
rect 20346 36700 20352 36712
rect 19291 36672 20352 36700
rect 19291 36669 19303 36672
rect 19245 36663 19303 36669
rect 20346 36660 20352 36672
rect 20404 36660 20410 36712
rect 20456 36700 20484 36808
rect 27062 36796 27068 36848
rect 27120 36836 27126 36848
rect 27218 36839 27276 36845
rect 27218 36836 27230 36839
rect 27120 36808 27230 36836
rect 27120 36796 27126 36808
rect 27218 36805 27230 36808
rect 27264 36805 27276 36839
rect 27218 36799 27276 36805
rect 23109 36771 23167 36777
rect 23109 36737 23121 36771
rect 23155 36768 23167 36771
rect 23750 36768 23756 36780
rect 23155 36740 23756 36768
rect 23155 36737 23167 36740
rect 23109 36731 23167 36737
rect 23750 36728 23756 36740
rect 23808 36728 23814 36780
rect 26970 36728 26976 36780
rect 27028 36728 27034 36780
rect 27356 36768 27384 36876
rect 28258 36864 28264 36916
rect 28316 36904 28322 36916
rect 28353 36907 28411 36913
rect 28353 36904 28365 36907
rect 28316 36876 28365 36904
rect 28316 36864 28322 36876
rect 28353 36873 28365 36876
rect 28399 36873 28411 36907
rect 28353 36867 28411 36873
rect 30116 36876 31754 36904
rect 28074 36796 28080 36848
rect 28132 36836 28138 36848
rect 30116 36845 30144 36876
rect 30101 36839 30159 36845
rect 30101 36836 30113 36839
rect 28132 36808 30113 36836
rect 28132 36796 28138 36808
rect 30101 36805 30113 36808
rect 30147 36805 30159 36839
rect 30101 36799 30159 36805
rect 30282 36796 30288 36848
rect 30340 36796 30346 36848
rect 31726 36836 31754 36876
rect 32398 36864 32404 36916
rect 32456 36904 32462 36916
rect 32858 36904 32864 36916
rect 32456 36876 32864 36904
rect 32456 36864 32462 36876
rect 32858 36864 32864 36876
rect 32916 36864 32922 36916
rect 34514 36864 34520 36916
rect 34572 36864 34578 36916
rect 36078 36904 36084 36916
rect 35176 36876 36084 36904
rect 32030 36836 32036 36848
rect 31726 36808 32036 36836
rect 32030 36796 32036 36808
rect 32088 36796 32094 36848
rect 33502 36796 33508 36848
rect 33560 36836 33566 36848
rect 34238 36836 34244 36848
rect 33560 36808 34244 36836
rect 33560 36796 33566 36808
rect 34238 36796 34244 36808
rect 34296 36796 34302 36848
rect 35176 36845 35204 36876
rect 36078 36864 36084 36876
rect 36136 36864 36142 36916
rect 36446 36864 36452 36916
rect 36504 36904 36510 36916
rect 36541 36907 36599 36913
rect 36541 36904 36553 36907
rect 36504 36876 36553 36904
rect 36504 36864 36510 36876
rect 36541 36873 36553 36876
rect 36587 36873 36599 36907
rect 36541 36867 36599 36873
rect 38838 36864 38844 36916
rect 38896 36904 38902 36916
rect 40221 36907 40279 36913
rect 40221 36904 40233 36907
rect 38896 36876 40233 36904
rect 38896 36864 38902 36876
rect 40221 36873 40233 36876
rect 40267 36904 40279 36907
rect 44174 36904 44180 36916
rect 40267 36876 44180 36904
rect 40267 36873 40279 36876
rect 40221 36867 40279 36873
rect 44174 36864 44180 36876
rect 44232 36864 44238 36916
rect 35161 36839 35219 36845
rect 35161 36805 35173 36839
rect 35207 36805 35219 36839
rect 36906 36836 36912 36848
rect 35161 36799 35219 36805
rect 36096 36808 36912 36836
rect 31570 36768 31576 36780
rect 27356 36740 31576 36768
rect 31570 36728 31576 36740
rect 31628 36728 31634 36780
rect 31662 36728 31668 36780
rect 31720 36768 31726 36780
rect 32585 36771 32643 36777
rect 32585 36768 32597 36771
rect 31720 36740 32597 36768
rect 31720 36728 31726 36740
rect 32585 36737 32597 36740
rect 32631 36737 32643 36771
rect 32585 36731 32643 36737
rect 32852 36771 32910 36777
rect 32852 36737 32864 36771
rect 32898 36768 32910 36771
rect 34606 36768 34612 36780
rect 32898 36740 34612 36768
rect 32898 36737 32910 36740
rect 32852 36731 32910 36737
rect 34606 36728 34612 36740
rect 34664 36728 34670 36780
rect 34790 36728 34796 36780
rect 34848 36728 34854 36780
rect 35434 36768 35440 36780
rect 34900 36740 35440 36768
rect 22002 36700 22008 36712
rect 20456 36672 22008 36700
rect 22002 36660 22008 36672
rect 22060 36700 22066 36712
rect 23293 36703 23351 36709
rect 23293 36700 23305 36703
rect 22060 36672 23305 36700
rect 22060 36660 22066 36672
rect 23293 36669 23305 36672
rect 23339 36669 23351 36703
rect 23293 36663 23351 36669
rect 34701 36703 34759 36709
rect 34701 36669 34713 36703
rect 34747 36700 34759 36703
rect 34900 36700 34928 36740
rect 35434 36728 35440 36740
rect 35492 36728 35498 36780
rect 36096 36777 36124 36808
rect 36906 36796 36912 36808
rect 36964 36796 36970 36848
rect 39108 36839 39166 36845
rect 39108 36805 39120 36839
rect 39154 36836 39166 36839
rect 39206 36836 39212 36848
rect 39154 36808 39212 36836
rect 39154 36805 39166 36808
rect 39108 36799 39166 36805
rect 39206 36796 39212 36808
rect 39264 36796 39270 36848
rect 36081 36771 36139 36777
rect 36081 36737 36093 36771
rect 36127 36737 36139 36771
rect 36081 36731 36139 36737
rect 36170 36728 36176 36780
rect 36228 36768 36234 36780
rect 36357 36771 36415 36777
rect 36357 36768 36369 36771
rect 36228 36740 36369 36768
rect 36228 36728 36234 36740
rect 36357 36737 36369 36740
rect 36403 36737 36415 36771
rect 37642 36768 37648 36780
rect 36357 36731 36415 36737
rect 36464 36740 37648 36768
rect 34747 36672 34928 36700
rect 35069 36703 35127 36709
rect 34747 36669 34759 36672
rect 34701 36663 34759 36669
rect 35069 36669 35081 36703
rect 35115 36669 35127 36703
rect 35069 36663 35127 36669
rect 15654 36592 15660 36644
rect 15712 36632 15718 36644
rect 16482 36632 16488 36644
rect 15712 36604 16488 36632
rect 15712 36592 15718 36604
rect 16482 36592 16488 36604
rect 16540 36592 16546 36644
rect 19426 36592 19432 36644
rect 19484 36632 19490 36644
rect 19521 36635 19579 36641
rect 19521 36632 19533 36635
rect 19484 36604 19533 36632
rect 19484 36592 19490 36604
rect 19521 36601 19533 36604
rect 19567 36601 19579 36635
rect 19521 36595 19579 36601
rect 29270 36592 29276 36644
rect 29328 36632 29334 36644
rect 29328 36604 32628 36632
rect 29328 36592 29334 36604
rect 16301 36567 16359 36573
rect 16301 36533 16313 36567
rect 16347 36564 16359 36567
rect 16758 36564 16764 36576
rect 16347 36536 16764 36564
rect 16347 36533 16359 36536
rect 16301 36527 16359 36533
rect 16758 36524 16764 36536
rect 16816 36524 16822 36576
rect 19702 36524 19708 36576
rect 19760 36524 19766 36576
rect 32600 36564 32628 36604
rect 33520 36604 34468 36632
rect 33520 36564 33548 36604
rect 32600 36536 33548 36564
rect 33965 36567 34023 36573
rect 33965 36533 33977 36567
rect 34011 36564 34023 36567
rect 34054 36564 34060 36576
rect 34011 36536 34060 36564
rect 34011 36533 34023 36536
rect 33965 36527 34023 36533
rect 34054 36524 34060 36536
rect 34112 36524 34118 36576
rect 34440 36564 34468 36604
rect 34514 36592 34520 36644
rect 34572 36632 34578 36644
rect 35084 36632 35112 36663
rect 34572 36604 35112 36632
rect 34572 36592 34578 36604
rect 35986 36592 35992 36644
rect 36044 36632 36050 36644
rect 36173 36635 36231 36641
rect 36173 36632 36185 36635
rect 36044 36604 36185 36632
rect 36044 36592 36050 36604
rect 36173 36601 36185 36604
rect 36219 36632 36231 36635
rect 36464 36632 36492 36740
rect 37642 36728 37648 36740
rect 37700 36728 37706 36780
rect 38010 36728 38016 36780
rect 38068 36768 38074 36780
rect 38841 36771 38899 36777
rect 38841 36768 38853 36771
rect 38068 36740 38853 36768
rect 38068 36728 38074 36740
rect 38841 36737 38853 36740
rect 38887 36737 38899 36771
rect 38841 36731 38899 36737
rect 38654 36700 38660 36712
rect 36219 36604 36492 36632
rect 36556 36672 38660 36700
rect 36219 36601 36231 36604
rect 36173 36595 36231 36601
rect 36556 36564 36584 36672
rect 38654 36660 38660 36672
rect 38712 36660 38718 36712
rect 34440 36536 36584 36564
rect 36630 36524 36636 36576
rect 36688 36564 36694 36576
rect 46842 36564 46848 36576
rect 36688 36536 46848 36564
rect 36688 36524 36694 36536
rect 46842 36524 46848 36536
rect 46900 36524 46906 36576
rect 1104 36474 47104 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 47104 36474
rect 1104 36400 47104 36422
rect 17497 36363 17555 36369
rect 16224 36332 17448 36360
rect 2130 36184 2136 36236
rect 2188 36224 2194 36236
rect 2501 36227 2559 36233
rect 2501 36224 2513 36227
rect 2188 36196 2513 36224
rect 2188 36184 2194 36196
rect 2501 36193 2513 36196
rect 2547 36193 2559 36227
rect 2501 36187 2559 36193
rect 4433 36227 4491 36233
rect 4433 36193 4445 36227
rect 4479 36224 4491 36227
rect 7190 36224 7196 36236
rect 4479 36196 7196 36224
rect 4479 36193 4491 36196
rect 4433 36187 4491 36193
rect 7190 36184 7196 36196
rect 7248 36224 7254 36236
rect 7650 36224 7656 36236
rect 7248 36196 7656 36224
rect 7248 36184 7254 36196
rect 7650 36184 7656 36196
rect 7708 36184 7714 36236
rect 9674 36184 9680 36236
rect 9732 36224 9738 36236
rect 10045 36227 10103 36233
rect 10045 36224 10057 36227
rect 9732 36196 10057 36224
rect 9732 36184 9738 36196
rect 10045 36193 10057 36196
rect 10091 36193 10103 36227
rect 10045 36187 10103 36193
rect 10502 36184 10508 36236
rect 10560 36224 10566 36236
rect 11241 36227 11299 36233
rect 11241 36224 11253 36227
rect 10560 36196 11253 36224
rect 10560 36184 10566 36196
rect 11241 36193 11253 36196
rect 11287 36193 11299 36227
rect 11241 36187 11299 36193
rect 15194 36184 15200 36236
rect 15252 36224 15258 36236
rect 15749 36227 15807 36233
rect 15749 36224 15761 36227
rect 15252 36196 15761 36224
rect 15252 36184 15258 36196
rect 15749 36193 15761 36196
rect 15795 36224 15807 36227
rect 15838 36224 15844 36236
rect 15795 36196 15844 36224
rect 15795 36193 15807 36196
rect 15749 36187 15807 36193
rect 15838 36184 15844 36196
rect 15896 36184 15902 36236
rect 16224 36233 16252 36332
rect 17420 36292 17448 36332
rect 17497 36329 17509 36363
rect 17543 36360 17555 36363
rect 19426 36360 19432 36372
rect 17543 36332 19432 36360
rect 17543 36329 17555 36332
rect 17497 36323 17555 36329
rect 19426 36320 19432 36332
rect 19484 36320 19490 36372
rect 19518 36320 19524 36372
rect 19576 36360 19582 36372
rect 19576 36332 22784 36360
rect 19576 36320 19582 36332
rect 18506 36292 18512 36304
rect 17420 36264 18512 36292
rect 18506 36252 18512 36264
rect 18564 36252 18570 36304
rect 18690 36252 18696 36304
rect 18748 36252 18754 36304
rect 20257 36295 20315 36301
rect 20257 36261 20269 36295
rect 20303 36292 20315 36295
rect 20438 36292 20444 36304
rect 20303 36264 20444 36292
rect 20303 36261 20315 36264
rect 20257 36255 20315 36261
rect 20438 36252 20444 36264
rect 20496 36252 20502 36304
rect 21637 36295 21695 36301
rect 21637 36261 21649 36295
rect 21683 36292 21695 36295
rect 22094 36292 22100 36304
rect 21683 36264 22100 36292
rect 21683 36261 21695 36264
rect 21637 36255 21695 36261
rect 22094 36252 22100 36264
rect 22152 36252 22158 36304
rect 16209 36227 16267 36233
rect 16209 36193 16221 36227
rect 16255 36193 16267 36227
rect 16209 36187 16267 36193
rect 16574 36184 16580 36236
rect 16632 36233 16638 36236
rect 16632 36227 16660 36233
rect 16648 36193 16660 36227
rect 16632 36187 16660 36193
rect 16761 36227 16819 36233
rect 16761 36193 16773 36227
rect 16807 36224 16819 36227
rect 18141 36227 18199 36233
rect 16807 36196 18092 36224
rect 16807 36193 16819 36196
rect 16761 36187 16819 36193
rect 16632 36184 16638 36187
rect 2225 36159 2283 36165
rect 2225 36125 2237 36159
rect 2271 36156 2283 36159
rect 3970 36156 3976 36168
rect 2271 36128 3976 36156
rect 2271 36125 2283 36128
rect 2225 36119 2283 36125
rect 3970 36116 3976 36128
rect 4028 36116 4034 36168
rect 4249 36159 4307 36165
rect 4249 36125 4261 36159
rect 4295 36156 4307 36159
rect 5258 36156 5264 36168
rect 4295 36128 5264 36156
rect 4295 36125 4307 36128
rect 4249 36119 4307 36125
rect 5258 36116 5264 36128
rect 5316 36116 5322 36168
rect 9769 36159 9827 36165
rect 9769 36125 9781 36159
rect 9815 36156 9827 36159
rect 9950 36156 9956 36168
rect 9815 36128 9956 36156
rect 9815 36125 9827 36128
rect 9769 36119 9827 36125
rect 9950 36116 9956 36128
rect 10008 36116 10014 36168
rect 13722 36116 13728 36168
rect 13780 36156 13786 36168
rect 13780 36128 14412 36156
rect 13780 36116 13786 36128
rect 9306 36048 9312 36100
rect 9364 36088 9370 36100
rect 9364 36060 11192 36088
rect 9364 36048 9370 36060
rect 3326 35980 3332 36032
rect 3384 36020 3390 36032
rect 3789 36023 3847 36029
rect 3789 36020 3801 36023
rect 3384 35992 3801 36020
rect 3384 35980 3390 35992
rect 3789 35989 3801 35992
rect 3835 35989 3847 36023
rect 3789 35983 3847 35989
rect 4154 35980 4160 36032
rect 4212 35980 4218 36032
rect 4522 35980 4528 36032
rect 4580 36020 4586 36032
rect 5350 36020 5356 36032
rect 4580 35992 5356 36020
rect 4580 35980 4586 35992
rect 5350 35980 5356 35992
rect 5408 35980 5414 36032
rect 9582 35980 9588 36032
rect 9640 36020 9646 36032
rect 10689 36023 10747 36029
rect 10689 36020 10701 36023
rect 9640 35992 10701 36020
rect 9640 35980 9646 35992
rect 10689 35989 10701 35992
rect 10735 35989 10747 36023
rect 10689 35983 10747 35989
rect 11054 35980 11060 36032
rect 11112 35980 11118 36032
rect 11164 36029 11192 36060
rect 14090 36048 14096 36100
rect 14148 36088 14154 36100
rect 14185 36091 14243 36097
rect 14185 36088 14197 36091
rect 14148 36060 14197 36088
rect 14148 36048 14154 36060
rect 14185 36057 14197 36060
rect 14231 36057 14243 36091
rect 14185 36051 14243 36057
rect 11149 36023 11207 36029
rect 11149 35989 11161 36023
rect 11195 36020 11207 36023
rect 14274 36020 14280 36032
rect 11195 35992 14280 36020
rect 11195 35989 11207 35992
rect 11149 35983 11207 35989
rect 14274 35980 14280 35992
rect 14332 35980 14338 36032
rect 14384 36020 14412 36128
rect 15470 36116 15476 36168
rect 15528 36156 15534 36168
rect 15565 36159 15623 36165
rect 15565 36156 15577 36159
rect 15528 36128 15577 36156
rect 15528 36116 15534 36128
rect 15565 36125 15577 36128
rect 15611 36125 15623 36159
rect 15565 36119 15623 36125
rect 16482 36116 16488 36168
rect 16540 36116 16546 36168
rect 18064 36156 18092 36196
rect 18141 36193 18153 36227
rect 18187 36224 18199 36227
rect 19610 36224 19616 36236
rect 18187 36196 19616 36224
rect 18187 36193 18199 36196
rect 18141 36187 18199 36193
rect 19610 36184 19616 36196
rect 19668 36184 19674 36236
rect 19705 36227 19763 36233
rect 19705 36193 19717 36227
rect 19751 36224 19763 36227
rect 19751 36196 22508 36224
rect 19751 36193 19763 36196
rect 19705 36187 19763 36193
rect 18230 36156 18236 36168
rect 18064 36128 18236 36156
rect 18230 36116 18236 36128
rect 18288 36116 18294 36168
rect 18325 36159 18383 36165
rect 18325 36125 18337 36159
rect 18371 36156 18383 36159
rect 19334 36156 19340 36168
rect 18371 36128 19340 36156
rect 18371 36125 18383 36128
rect 18325 36119 18383 36125
rect 19334 36116 19340 36128
rect 19392 36156 19398 36168
rect 19518 36156 19524 36168
rect 19392 36128 19524 36156
rect 19392 36116 19398 36128
rect 19518 36116 19524 36128
rect 19576 36116 19582 36168
rect 19886 36116 19892 36168
rect 19944 36116 19950 36168
rect 20165 36159 20223 36165
rect 20165 36125 20177 36159
rect 20211 36125 20223 36159
rect 20165 36119 20223 36125
rect 17405 36091 17463 36097
rect 17405 36057 17417 36091
rect 17451 36088 17463 36091
rect 17865 36091 17923 36097
rect 17865 36088 17877 36091
rect 17451 36060 17877 36088
rect 17451 36057 17463 36060
rect 17405 36051 17463 36057
rect 17865 36057 17877 36060
rect 17911 36057 17923 36091
rect 17865 36051 17923 36057
rect 18598 36048 18604 36100
rect 18656 36088 18662 36100
rect 18656 36060 18920 36088
rect 18656 36048 18662 36060
rect 17957 36023 18015 36029
rect 17957 36020 17969 36023
rect 14384 35992 17969 36020
rect 17957 35989 17969 35992
rect 18003 35989 18015 36023
rect 17957 35983 18015 35989
rect 18782 35980 18788 36032
rect 18840 35980 18846 36032
rect 18892 36020 18920 36060
rect 19242 36048 19248 36100
rect 19300 36088 19306 36100
rect 20073 36091 20131 36097
rect 20073 36088 20085 36091
rect 19300 36060 20085 36088
rect 19300 36048 19306 36060
rect 20073 36057 20085 36060
rect 20119 36057 20131 36091
rect 20180 36088 20208 36119
rect 20254 36116 20260 36168
rect 20312 36156 20318 36168
rect 20441 36159 20499 36165
rect 20441 36156 20453 36159
rect 20312 36128 20453 36156
rect 20312 36116 20318 36128
rect 20441 36125 20453 36128
rect 20487 36125 20499 36159
rect 20441 36119 20499 36125
rect 20622 36116 20628 36168
rect 20680 36156 20686 36168
rect 20717 36159 20775 36165
rect 20717 36156 20729 36159
rect 20680 36128 20729 36156
rect 20680 36116 20686 36128
rect 20717 36125 20729 36128
rect 20763 36125 20775 36159
rect 20717 36119 20775 36125
rect 21821 36159 21879 36165
rect 21821 36125 21833 36159
rect 21867 36156 21879 36159
rect 21867 36128 21956 36156
rect 21867 36125 21879 36128
rect 21821 36119 21879 36125
rect 20640 36088 20668 36116
rect 20180 36060 20668 36088
rect 20073 36051 20131 36057
rect 21928 36029 21956 36128
rect 22002 36116 22008 36168
rect 22060 36156 22066 36168
rect 22373 36159 22431 36165
rect 22373 36156 22385 36159
rect 22060 36128 22385 36156
rect 22060 36116 22066 36128
rect 22373 36125 22385 36128
rect 22419 36125 22431 36159
rect 22480 36156 22508 36196
rect 22554 36184 22560 36236
rect 22612 36184 22618 36236
rect 22756 36233 22784 36332
rect 29086 36320 29092 36372
rect 29144 36360 29150 36372
rect 29733 36363 29791 36369
rect 29733 36360 29745 36363
rect 29144 36332 29745 36360
rect 29144 36320 29150 36332
rect 29733 36329 29745 36332
rect 29779 36329 29791 36363
rect 32306 36360 32312 36372
rect 29733 36323 29791 36329
rect 31956 36332 32312 36360
rect 23014 36252 23020 36304
rect 23072 36252 23078 36304
rect 23658 36252 23664 36304
rect 23716 36252 23722 36304
rect 22741 36227 22799 36233
rect 22741 36193 22753 36227
rect 22787 36193 22799 36227
rect 22741 36187 22799 36193
rect 23198 36184 23204 36236
rect 23256 36224 23262 36236
rect 25498 36224 25504 36236
rect 23256 36196 25504 36224
rect 23256 36184 23262 36196
rect 25498 36184 25504 36196
rect 25556 36184 25562 36236
rect 25682 36184 25688 36236
rect 25740 36224 25746 36236
rect 31956 36233 31984 36332
rect 32306 36320 32312 36332
rect 32364 36360 32370 36372
rect 34054 36360 34060 36372
rect 32364 36332 34060 36360
rect 32364 36320 32370 36332
rect 34054 36320 34060 36332
rect 34112 36320 34118 36372
rect 34606 36320 34612 36372
rect 34664 36360 34670 36372
rect 34701 36363 34759 36369
rect 34701 36360 34713 36363
rect 34664 36332 34713 36360
rect 34664 36320 34670 36332
rect 34701 36329 34713 36332
rect 34747 36329 34759 36363
rect 34701 36323 34759 36329
rect 36170 36320 36176 36372
rect 36228 36360 36234 36372
rect 36725 36363 36783 36369
rect 36725 36360 36737 36363
rect 36228 36332 36737 36360
rect 36228 36320 36234 36332
rect 36725 36329 36737 36332
rect 36771 36329 36783 36363
rect 36725 36323 36783 36329
rect 37277 36363 37335 36369
rect 37277 36329 37289 36363
rect 37323 36360 37335 36363
rect 37642 36360 37648 36372
rect 37323 36332 37648 36360
rect 37323 36329 37335 36332
rect 37277 36323 37335 36329
rect 37642 36320 37648 36332
rect 37700 36320 37706 36372
rect 38654 36320 38660 36372
rect 38712 36360 38718 36372
rect 39022 36360 39028 36372
rect 38712 36332 39028 36360
rect 38712 36320 38718 36332
rect 39022 36320 39028 36332
rect 39080 36320 39086 36372
rect 32490 36292 32496 36304
rect 32324 36264 32496 36292
rect 31941 36227 31999 36233
rect 25740 36196 29776 36224
rect 25740 36184 25746 36196
rect 26050 36156 26056 36168
rect 22480 36128 26056 36156
rect 22373 36119 22431 36125
rect 26050 36116 26056 36128
rect 26108 36116 26114 36168
rect 29270 36116 29276 36168
rect 29328 36116 29334 36168
rect 23293 36091 23351 36097
rect 23293 36057 23305 36091
rect 23339 36088 23351 36091
rect 23382 36088 23388 36100
rect 23339 36060 23388 36088
rect 23339 36057 23351 36060
rect 23293 36051 23351 36057
rect 23382 36048 23388 36060
rect 23440 36048 23446 36100
rect 29454 36088 29460 36100
rect 29104 36060 29460 36088
rect 20625 36023 20683 36029
rect 20625 36020 20637 36023
rect 18892 35992 20637 36020
rect 20625 35989 20637 35992
rect 20671 35989 20683 36023
rect 20625 35983 20683 35989
rect 21913 36023 21971 36029
rect 21913 35989 21925 36023
rect 21959 35989 21971 36023
rect 21913 35983 21971 35989
rect 22278 35980 22284 36032
rect 22336 35980 22342 36032
rect 23201 36023 23259 36029
rect 23201 35989 23213 36023
rect 23247 36020 23259 36023
rect 23474 36020 23480 36032
rect 23247 35992 23480 36020
rect 23247 35989 23259 35992
rect 23201 35983 23259 35989
rect 23474 35980 23480 35992
rect 23532 35980 23538 36032
rect 23753 36023 23811 36029
rect 23753 35989 23765 36023
rect 23799 36020 23811 36023
rect 26142 36020 26148 36032
rect 23799 35992 26148 36020
rect 23799 35989 23811 35992
rect 23753 35983 23811 35989
rect 26142 35980 26148 35992
rect 26200 35980 26206 36032
rect 29104 36029 29132 36060
rect 29454 36048 29460 36060
rect 29512 36088 29518 36100
rect 29641 36091 29699 36097
rect 29641 36088 29653 36091
rect 29512 36060 29653 36088
rect 29512 36048 29518 36060
rect 29641 36057 29653 36060
rect 29687 36057 29699 36091
rect 29748 36088 29776 36196
rect 31941 36193 31953 36227
rect 31987 36193 31999 36227
rect 32324 36224 32352 36264
rect 32490 36252 32496 36264
rect 32548 36252 32554 36304
rect 33410 36252 33416 36304
rect 33468 36292 33474 36304
rect 33468 36264 35848 36292
rect 33468 36252 33474 36264
rect 34624 36236 34652 36264
rect 31941 36187 31999 36193
rect 32140 36196 32352 36224
rect 32140 36168 32168 36196
rect 32398 36184 32404 36236
rect 32456 36184 32462 36236
rect 32674 36184 32680 36236
rect 32732 36184 32738 36236
rect 32766 36184 32772 36236
rect 32824 36233 32830 36236
rect 32824 36227 32873 36233
rect 32824 36193 32827 36227
rect 32861 36224 32873 36227
rect 33134 36224 33140 36236
rect 32861 36196 33140 36224
rect 32861 36193 32873 36196
rect 32824 36187 32873 36193
rect 32824 36184 32830 36187
rect 33134 36184 33140 36196
rect 33192 36184 33198 36236
rect 33502 36184 33508 36236
rect 33560 36224 33566 36236
rect 34241 36227 34299 36233
rect 34241 36224 34253 36227
rect 33560 36196 34253 36224
rect 33560 36184 33566 36196
rect 34241 36193 34253 36196
rect 34287 36193 34299 36227
rect 34241 36187 34299 36193
rect 34606 36184 34612 36236
rect 34664 36184 34670 36236
rect 31757 36159 31815 36165
rect 31757 36125 31769 36159
rect 31803 36156 31815 36159
rect 32122 36156 32128 36168
rect 31803 36128 32128 36156
rect 31803 36125 31815 36128
rect 31757 36119 31815 36125
rect 32122 36116 32128 36128
rect 32180 36116 32186 36168
rect 32950 36116 32956 36168
rect 33008 36116 33014 36168
rect 35820 36165 35848 36264
rect 36538 36252 36544 36304
rect 36596 36252 36602 36304
rect 36556 36224 36584 36252
rect 36556 36196 37136 36224
rect 34885 36159 34943 36165
rect 34885 36156 34897 36159
rect 33704 36128 34897 36156
rect 29748 36060 31754 36088
rect 29641 36051 29699 36057
rect 29089 36023 29147 36029
rect 29089 35989 29101 36023
rect 29135 35989 29147 36023
rect 31726 36020 31754 36060
rect 33704 36029 33732 36128
rect 34885 36125 34897 36128
rect 34931 36125 34943 36159
rect 34885 36119 34943 36125
rect 35805 36159 35863 36165
rect 35805 36125 35817 36159
rect 35851 36125 35863 36159
rect 35805 36119 35863 36125
rect 35986 36116 35992 36168
rect 36044 36116 36050 36168
rect 36262 36116 36268 36168
rect 36320 36116 36326 36168
rect 36541 36159 36599 36165
rect 36541 36125 36553 36159
rect 36587 36125 36599 36159
rect 36541 36119 36599 36125
rect 34054 36048 34060 36100
rect 34112 36048 34118 36100
rect 35897 36091 35955 36097
rect 35897 36057 35909 36091
rect 35943 36088 35955 36091
rect 36556 36088 36584 36119
rect 36814 36116 36820 36168
rect 36872 36116 36878 36168
rect 37108 36165 37136 36196
rect 37093 36159 37151 36165
rect 37093 36125 37105 36159
rect 37139 36125 37151 36159
rect 37093 36119 37151 36125
rect 37366 36116 37372 36168
rect 37424 36116 37430 36168
rect 35943 36060 36584 36088
rect 35943 36057 35955 36060
rect 35897 36051 35955 36057
rect 33597 36023 33655 36029
rect 33597 36020 33609 36023
rect 31726 35992 33609 36020
rect 29089 35983 29147 35989
rect 33597 35989 33609 35992
rect 33643 35989 33655 36023
rect 33597 35983 33655 35989
rect 33689 36023 33747 36029
rect 33689 35989 33701 36023
rect 33735 35989 33747 36023
rect 33689 35983 33747 35989
rect 34146 35980 34152 36032
rect 34204 35980 34210 36032
rect 35986 35980 35992 36032
rect 36044 36020 36050 36032
rect 36081 36023 36139 36029
rect 36081 36020 36093 36023
rect 36044 35992 36093 36020
rect 36044 35980 36050 35992
rect 36081 35989 36093 35992
rect 36127 35989 36139 36023
rect 36081 35983 36139 35989
rect 36354 35980 36360 36032
rect 36412 35980 36418 36032
rect 36538 35980 36544 36032
rect 36596 36020 36602 36032
rect 36909 36023 36967 36029
rect 36909 36020 36921 36023
rect 36596 35992 36921 36020
rect 36596 35980 36602 35992
rect 36909 35989 36921 35992
rect 36955 35989 36967 36023
rect 36909 35983 36967 35989
rect 1104 35930 47104 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 47104 35930
rect 1104 35856 47104 35878
rect 1857 35819 1915 35825
rect 1857 35785 1869 35819
rect 1903 35785 1915 35819
rect 1857 35779 1915 35785
rect 3513 35819 3571 35825
rect 3513 35785 3525 35819
rect 3559 35816 3571 35819
rect 4154 35816 4160 35828
rect 3559 35788 4160 35816
rect 3559 35785 3571 35788
rect 3513 35779 3571 35785
rect 1872 35748 1900 35779
rect 4154 35776 4160 35788
rect 4212 35816 4218 35828
rect 5258 35816 5264 35828
rect 4212 35788 5264 35816
rect 4212 35776 4218 35788
rect 5258 35776 5264 35788
rect 5316 35776 5322 35828
rect 7101 35819 7159 35825
rect 7101 35785 7113 35819
rect 7147 35785 7159 35819
rect 10318 35816 10324 35828
rect 7101 35779 7159 35785
rect 7392 35788 10324 35816
rect 2378 35751 2436 35757
rect 2378 35748 2390 35751
rect 1872 35720 2390 35748
rect 2378 35717 2390 35720
rect 2424 35717 2436 35751
rect 2378 35711 2436 35717
rect 2041 35683 2099 35689
rect 2041 35649 2053 35683
rect 2087 35680 2099 35683
rect 3326 35680 3332 35692
rect 2087 35652 3332 35680
rect 2087 35649 2099 35652
rect 2041 35643 2099 35649
rect 3326 35640 3332 35652
rect 3384 35640 3390 35692
rect 3786 35640 3792 35692
rect 3844 35640 3850 35692
rect 4249 35683 4307 35689
rect 4249 35649 4261 35683
rect 4295 35680 4307 35683
rect 4614 35680 4620 35692
rect 4295 35652 4620 35680
rect 4295 35649 4307 35652
rect 4249 35643 4307 35649
rect 4614 35640 4620 35652
rect 4672 35640 4678 35692
rect 5258 35640 5264 35692
rect 5316 35689 5322 35692
rect 5316 35683 5344 35689
rect 5332 35649 5344 35683
rect 5316 35643 5344 35649
rect 7009 35683 7067 35689
rect 7009 35649 7021 35683
rect 7055 35680 7067 35683
rect 7116 35680 7144 35779
rect 7055 35652 7144 35680
rect 7055 35649 7067 35652
rect 7009 35643 7067 35649
rect 5316 35640 5322 35643
rect 2130 35572 2136 35624
rect 2188 35572 2194 35624
rect 4433 35615 4491 35621
rect 4433 35581 4445 35615
rect 4479 35581 4491 35615
rect 4433 35575 4491 35581
rect 4448 35544 4476 35575
rect 4522 35572 4528 35624
rect 4580 35612 4586 35624
rect 4893 35615 4951 35621
rect 4893 35612 4905 35615
rect 4580 35584 4905 35612
rect 4580 35572 4586 35584
rect 4893 35581 4905 35584
rect 4939 35612 4951 35615
rect 4982 35612 4988 35624
rect 4939 35584 4988 35612
rect 4939 35581 4951 35584
rect 4893 35575 4951 35581
rect 4982 35572 4988 35584
rect 5040 35572 5046 35624
rect 5166 35572 5172 35624
rect 5224 35572 5230 35624
rect 5445 35615 5503 35621
rect 5445 35581 5457 35615
rect 5491 35612 5503 35615
rect 5626 35612 5632 35624
rect 5491 35584 5632 35612
rect 5491 35581 5503 35584
rect 5445 35575 5503 35581
rect 5626 35572 5632 35584
rect 5684 35612 5690 35624
rect 7392 35612 7420 35788
rect 10318 35776 10324 35788
rect 10376 35776 10382 35828
rect 13078 35776 13084 35828
rect 13136 35816 13142 35828
rect 13449 35819 13507 35825
rect 13449 35816 13461 35819
rect 13136 35788 13461 35816
rect 13136 35776 13142 35788
rect 13449 35785 13461 35788
rect 13495 35785 13507 35819
rect 15470 35816 15476 35828
rect 13449 35779 13507 35785
rect 14660 35788 15476 35816
rect 7561 35751 7619 35757
rect 7561 35717 7573 35751
rect 7607 35748 7619 35751
rect 9306 35748 9312 35760
rect 7607 35720 9312 35748
rect 7607 35717 7619 35720
rect 7561 35711 7619 35717
rect 9306 35708 9312 35720
rect 9364 35708 9370 35760
rect 9922 35751 9980 35757
rect 9922 35748 9934 35751
rect 9416 35720 9934 35748
rect 7469 35683 7527 35689
rect 7469 35649 7481 35683
rect 7515 35680 7527 35683
rect 7926 35680 7932 35692
rect 7515 35652 7932 35680
rect 7515 35649 7527 35652
rect 7469 35643 7527 35649
rect 7926 35640 7932 35652
rect 7984 35640 7990 35692
rect 8389 35683 8447 35689
rect 8389 35649 8401 35683
rect 8435 35680 8447 35683
rect 8938 35680 8944 35692
rect 8435 35652 8944 35680
rect 8435 35649 8447 35652
rect 8389 35643 8447 35649
rect 8938 35640 8944 35652
rect 8996 35640 9002 35692
rect 5684 35584 7420 35612
rect 5684 35572 5690 35584
rect 7650 35572 7656 35624
rect 7708 35572 7714 35624
rect 4706 35544 4712 35556
rect 4448 35516 4712 35544
rect 4706 35504 4712 35516
rect 4764 35504 4770 35556
rect 9122 35544 9128 35556
rect 5828 35516 9128 35544
rect 3602 35436 3608 35488
rect 3660 35436 3666 35488
rect 4890 35436 4896 35488
rect 4948 35476 4954 35488
rect 5828 35476 5856 35516
rect 9122 35504 9128 35516
rect 9180 35504 9186 35556
rect 4948 35448 5856 35476
rect 4948 35436 4954 35448
rect 6086 35436 6092 35488
rect 6144 35436 6150 35488
rect 6822 35436 6828 35488
rect 6880 35436 6886 35488
rect 8205 35479 8263 35485
rect 8205 35445 8217 35479
rect 8251 35476 8263 35479
rect 8294 35476 8300 35488
rect 8251 35448 8300 35476
rect 8251 35445 8263 35448
rect 8205 35439 8263 35445
rect 8294 35436 8300 35448
rect 8352 35436 8358 35488
rect 9416 35485 9444 35720
rect 9922 35717 9934 35720
rect 9968 35717 9980 35751
rect 13814 35748 13820 35760
rect 9922 35711 9980 35717
rect 13280 35720 13820 35748
rect 9582 35640 9588 35692
rect 9640 35640 9646 35692
rect 13280 35689 13308 35720
rect 13814 35708 13820 35720
rect 13872 35708 13878 35760
rect 14660 35689 14688 35788
rect 15470 35776 15476 35788
rect 15528 35776 15534 35828
rect 15562 35776 15568 35828
rect 15620 35816 15626 35828
rect 16482 35816 16488 35828
rect 15620 35788 16488 35816
rect 15620 35776 15626 35788
rect 16482 35776 16488 35788
rect 16540 35776 16546 35828
rect 17954 35776 17960 35828
rect 18012 35816 18018 35828
rect 18049 35819 18107 35825
rect 18049 35816 18061 35819
rect 18012 35788 18061 35816
rect 18012 35776 18018 35788
rect 18049 35785 18061 35788
rect 18095 35785 18107 35819
rect 18049 35779 18107 35785
rect 20901 35819 20959 35825
rect 20901 35785 20913 35819
rect 20947 35785 20959 35819
rect 20901 35779 20959 35785
rect 21361 35819 21419 35825
rect 21361 35785 21373 35819
rect 21407 35816 21419 35819
rect 22002 35816 22008 35828
rect 21407 35788 22008 35816
rect 21407 35785 21419 35788
rect 21361 35779 21419 35785
rect 17402 35748 17408 35760
rect 16684 35720 17408 35748
rect 13265 35683 13323 35689
rect 13265 35649 13277 35683
rect 13311 35649 13323 35683
rect 13265 35643 13323 35649
rect 13541 35683 13599 35689
rect 13541 35649 13553 35683
rect 13587 35649 13599 35683
rect 13541 35643 13599 35649
rect 14645 35683 14703 35689
rect 14645 35649 14657 35683
rect 14691 35649 14703 35683
rect 14645 35643 14703 35649
rect 9677 35615 9735 35621
rect 9677 35612 9689 35615
rect 9600 35584 9689 35612
rect 9600 35556 9628 35584
rect 9677 35581 9689 35584
rect 9723 35581 9735 35615
rect 9677 35575 9735 35581
rect 12434 35572 12440 35624
rect 12492 35612 12498 35624
rect 13556 35612 13584 35643
rect 15562 35640 15568 35692
rect 15620 35640 15626 35692
rect 15654 35640 15660 35692
rect 15712 35689 15718 35692
rect 16684 35689 16712 35720
rect 17402 35708 17408 35720
rect 17460 35708 17466 35760
rect 19352 35720 19932 35748
rect 15712 35683 15740 35689
rect 15728 35649 15740 35683
rect 15712 35643 15740 35649
rect 16669 35683 16727 35689
rect 16669 35649 16681 35683
rect 16715 35649 16727 35683
rect 16669 35643 16727 35649
rect 15712 35640 15718 35643
rect 16758 35640 16764 35692
rect 16816 35680 16822 35692
rect 16925 35683 16983 35689
rect 16925 35680 16937 35683
rect 16816 35652 16937 35680
rect 16816 35640 16822 35652
rect 16925 35649 16937 35652
rect 16971 35649 16983 35683
rect 16925 35643 16983 35649
rect 18046 35640 18052 35692
rect 18104 35680 18110 35692
rect 19352 35689 19380 35720
rect 19904 35692 19932 35720
rect 18233 35683 18291 35689
rect 18233 35680 18245 35683
rect 18104 35652 18245 35680
rect 18104 35640 18110 35652
rect 18233 35649 18245 35652
rect 18279 35649 18291 35683
rect 18233 35643 18291 35649
rect 19337 35683 19395 35689
rect 19337 35649 19349 35683
rect 19383 35649 19395 35683
rect 19337 35643 19395 35649
rect 19426 35640 19432 35692
rect 19484 35640 19490 35692
rect 19702 35640 19708 35692
rect 19760 35640 19766 35692
rect 19886 35640 19892 35692
rect 19944 35680 19950 35692
rect 19981 35683 20039 35689
rect 19981 35680 19993 35683
rect 19944 35652 19993 35680
rect 19944 35640 19950 35652
rect 19981 35649 19993 35652
rect 20027 35680 20039 35683
rect 20070 35680 20076 35692
rect 20027 35652 20076 35680
rect 20027 35649 20039 35652
rect 19981 35643 20039 35649
rect 20070 35640 20076 35652
rect 20128 35640 20134 35692
rect 20162 35640 20168 35692
rect 20220 35640 20226 35692
rect 20257 35683 20315 35689
rect 20257 35649 20269 35683
rect 20303 35649 20315 35683
rect 20257 35643 20315 35649
rect 20809 35683 20867 35689
rect 20809 35649 20821 35683
rect 20855 35680 20867 35683
rect 20916 35680 20944 35779
rect 22002 35776 22008 35788
rect 22060 35776 22066 35828
rect 22278 35776 22284 35828
rect 22336 35816 22342 35828
rect 23201 35819 23259 35825
rect 23201 35816 23213 35819
rect 22336 35788 23213 35816
rect 22336 35776 22342 35788
rect 23201 35785 23213 35788
rect 23247 35816 23259 35819
rect 25038 35816 25044 35828
rect 23247 35788 25044 35816
rect 23247 35785 23259 35788
rect 23201 35779 23259 35785
rect 25038 35776 25044 35788
rect 25096 35816 25102 35828
rect 25314 35816 25320 35828
rect 25096 35788 25320 35816
rect 25096 35776 25102 35788
rect 25314 35776 25320 35788
rect 25372 35776 25378 35828
rect 30377 35819 30435 35825
rect 25976 35788 27660 35816
rect 22094 35757 22100 35760
rect 22088 35711 22100 35757
rect 22094 35708 22100 35711
rect 22152 35708 22158 35760
rect 23750 35708 23756 35760
rect 23808 35708 23814 35760
rect 20855 35652 20944 35680
rect 21269 35683 21327 35689
rect 20855 35649 20867 35652
rect 20809 35643 20867 35649
rect 21269 35649 21281 35683
rect 21315 35680 21327 35683
rect 21910 35680 21916 35692
rect 21315 35652 21916 35680
rect 21315 35649 21327 35652
rect 21269 35643 21327 35649
rect 13725 35615 13783 35621
rect 13725 35612 13737 35615
rect 12492 35584 13737 35612
rect 12492 35572 12498 35584
rect 13725 35581 13737 35584
rect 13771 35581 13783 35615
rect 14734 35612 14740 35624
rect 13725 35575 13783 35581
rect 14016 35584 14740 35612
rect 9582 35504 9588 35556
rect 9640 35504 9646 35556
rect 14016 35544 14044 35584
rect 14734 35572 14740 35584
rect 14792 35572 14798 35624
rect 14829 35615 14887 35621
rect 14829 35581 14841 35615
rect 14875 35612 14887 35615
rect 15194 35612 15200 35624
rect 14875 35584 15200 35612
rect 14875 35581 14887 35584
rect 14829 35575 14887 35581
rect 15194 35572 15200 35584
rect 15252 35572 15258 35624
rect 15838 35572 15844 35624
rect 15896 35612 15902 35624
rect 15896 35584 16712 35612
rect 15896 35572 15902 35584
rect 10888 35516 14044 35544
rect 14093 35547 14151 35553
rect 9401 35479 9459 35485
rect 9401 35445 9413 35479
rect 9447 35445 9459 35479
rect 9401 35439 9459 35445
rect 9950 35436 9956 35488
rect 10008 35476 10014 35488
rect 10888 35476 10916 35516
rect 14093 35513 14105 35547
rect 14139 35544 14151 35547
rect 14139 35516 15240 35544
rect 14139 35513 14151 35516
rect 14093 35507 14151 35513
rect 10008 35448 10916 35476
rect 10008 35436 10014 35448
rect 11054 35436 11060 35488
rect 11112 35436 11118 35488
rect 13078 35436 13084 35488
rect 13136 35436 13142 35488
rect 14185 35479 14243 35485
rect 14185 35445 14197 35479
rect 14231 35476 14243 35479
rect 14366 35476 14372 35488
rect 14231 35448 14372 35476
rect 14231 35445 14243 35448
rect 14185 35439 14243 35445
rect 14366 35436 14372 35448
rect 14424 35436 14430 35488
rect 15212 35476 15240 35516
rect 15286 35504 15292 35556
rect 15344 35504 15350 35556
rect 16485 35479 16543 35485
rect 16485 35476 16497 35479
rect 15212 35448 16497 35476
rect 16485 35445 16497 35448
rect 16531 35445 16543 35479
rect 16684 35476 16712 35584
rect 18506 35572 18512 35624
rect 18564 35572 18570 35624
rect 19150 35572 19156 35624
rect 19208 35572 19214 35624
rect 20272 35612 20300 35643
rect 21910 35640 21916 35652
rect 21968 35640 21974 35692
rect 23661 35683 23719 35689
rect 23661 35649 23673 35683
rect 23707 35680 23719 35683
rect 23707 35652 24348 35680
rect 23707 35649 23719 35652
rect 23661 35643 23719 35649
rect 20622 35612 20628 35624
rect 20272 35584 20628 35612
rect 20622 35572 20628 35584
rect 20680 35612 20686 35624
rect 21082 35612 21088 35624
rect 20680 35584 21088 35612
rect 20680 35572 20686 35584
rect 21082 35572 21088 35584
rect 21140 35572 21146 35624
rect 21450 35572 21456 35624
rect 21508 35612 21514 35624
rect 21726 35612 21732 35624
rect 21508 35584 21732 35612
rect 21508 35572 21514 35584
rect 21726 35572 21732 35584
rect 21784 35572 21790 35624
rect 21821 35615 21879 35621
rect 21821 35581 21833 35615
rect 21867 35581 21879 35615
rect 21821 35575 21879 35581
rect 19613 35547 19671 35553
rect 19613 35513 19625 35547
rect 19659 35544 19671 35547
rect 20438 35544 20444 35556
rect 19659 35516 20444 35544
rect 19659 35513 19671 35516
rect 19613 35507 19671 35513
rect 20438 35504 20444 35516
rect 20496 35504 20502 35556
rect 20806 35504 20812 35556
rect 20864 35544 20870 35556
rect 21836 35544 21864 35575
rect 23842 35572 23848 35624
rect 23900 35572 23906 35624
rect 24121 35615 24179 35621
rect 24121 35581 24133 35615
rect 24167 35612 24179 35615
rect 24210 35612 24216 35624
rect 24167 35584 24216 35612
rect 24167 35581 24179 35584
rect 24121 35575 24179 35581
rect 24210 35572 24216 35584
rect 24268 35572 24274 35624
rect 24320 35621 24348 35652
rect 25038 35640 25044 35692
rect 25096 35640 25102 35692
rect 24305 35615 24363 35621
rect 24305 35581 24317 35615
rect 24351 35612 24363 35615
rect 24670 35612 24676 35624
rect 24351 35584 24676 35612
rect 24351 35581 24363 35584
rect 24305 35575 24363 35581
rect 24670 35572 24676 35584
rect 24728 35572 24734 35624
rect 25222 35621 25228 35624
rect 25179 35615 25228 35621
rect 25179 35581 25191 35615
rect 25225 35581 25228 35615
rect 25179 35575 25228 35581
rect 25222 35572 25228 35575
rect 25280 35572 25286 35624
rect 25317 35615 25375 35621
rect 25317 35581 25329 35615
rect 25363 35612 25375 35615
rect 25498 35612 25504 35624
rect 25363 35584 25504 35612
rect 25363 35581 25375 35584
rect 25317 35575 25375 35581
rect 25498 35572 25504 35584
rect 25556 35572 25562 35624
rect 25976 35612 26004 35788
rect 26142 35708 26148 35760
rect 26200 35748 26206 35760
rect 26200 35720 27568 35748
rect 26200 35708 26206 35720
rect 26050 35640 26056 35692
rect 26108 35680 26114 35692
rect 27157 35683 27215 35689
rect 27157 35680 27169 35683
rect 26108 35652 26556 35680
rect 26108 35640 26114 35652
rect 26142 35612 26148 35624
rect 25976 35584 26148 35612
rect 26142 35572 26148 35584
rect 26200 35572 26206 35624
rect 20864 35516 21864 35544
rect 20864 35504 20870 35516
rect 19518 35476 19524 35488
rect 16684 35448 19524 35476
rect 16485 35439 16543 35445
rect 19518 35436 19524 35448
rect 19576 35436 19582 35488
rect 19794 35436 19800 35488
rect 19852 35436 19858 35488
rect 20625 35479 20683 35485
rect 20625 35445 20637 35479
rect 20671 35476 20683 35479
rect 20898 35476 20904 35488
rect 20671 35448 20904 35476
rect 20671 35445 20683 35448
rect 20625 35439 20683 35445
rect 20898 35436 20904 35448
rect 20956 35436 20962 35488
rect 21836 35476 21864 35516
rect 24765 35547 24823 35553
rect 24765 35513 24777 35547
rect 24811 35513 24823 35547
rect 24765 35507 24823 35513
rect 22186 35476 22192 35488
rect 21836 35448 22192 35476
rect 22186 35436 22192 35448
rect 22244 35436 22250 35488
rect 23293 35479 23351 35485
rect 23293 35445 23305 35479
rect 23339 35476 23351 35479
rect 24026 35476 24032 35488
rect 23339 35448 24032 35476
rect 23339 35445 23351 35448
rect 23293 35439 23351 35445
rect 24026 35436 24032 35448
rect 24084 35436 24090 35488
rect 24118 35436 24124 35488
rect 24176 35476 24182 35488
rect 24780 35476 24808 35507
rect 26418 35504 26424 35556
rect 26476 35504 26482 35556
rect 26528 35544 26556 35652
rect 26620 35652 27169 35680
rect 26620 35621 26648 35652
rect 27157 35649 27169 35652
rect 27203 35649 27215 35683
rect 27157 35643 27215 35649
rect 27246 35640 27252 35692
rect 27304 35640 27310 35692
rect 27540 35689 27568 35720
rect 27525 35683 27583 35689
rect 27525 35649 27537 35683
rect 27571 35649 27583 35683
rect 27632 35680 27660 35788
rect 30377 35785 30389 35819
rect 30423 35816 30435 35819
rect 30837 35819 30895 35825
rect 30837 35816 30849 35819
rect 30423 35788 30849 35816
rect 30423 35785 30435 35788
rect 30377 35779 30435 35785
rect 30837 35785 30849 35788
rect 30883 35816 30895 35819
rect 30926 35816 30932 35828
rect 30883 35788 30932 35816
rect 30883 35785 30895 35788
rect 30837 35779 30895 35785
rect 30926 35776 30932 35788
rect 30984 35776 30990 35828
rect 33965 35819 34023 35825
rect 33965 35816 33977 35819
rect 31726 35788 33977 35816
rect 27890 35708 27896 35760
rect 27948 35748 27954 35760
rect 31726 35748 31754 35788
rect 33965 35785 33977 35788
rect 34011 35785 34023 35819
rect 33965 35779 34023 35785
rect 36262 35776 36268 35828
rect 36320 35816 36326 35828
rect 36630 35816 36636 35828
rect 36320 35788 36636 35816
rect 36320 35776 36326 35788
rect 36630 35776 36636 35788
rect 36688 35776 36694 35828
rect 36814 35776 36820 35828
rect 36872 35816 36878 35828
rect 37093 35819 37151 35825
rect 37093 35816 37105 35819
rect 36872 35788 37105 35816
rect 36872 35776 36878 35788
rect 37093 35785 37105 35788
rect 37139 35785 37151 35819
rect 37093 35779 37151 35785
rect 27948 35720 31754 35748
rect 35980 35751 36038 35757
rect 27948 35708 27954 35720
rect 35980 35717 35992 35751
rect 36026 35748 36038 35751
rect 36354 35748 36360 35760
rect 36026 35720 36360 35748
rect 36026 35717 36038 35720
rect 35980 35711 36038 35717
rect 36354 35708 36360 35720
rect 36412 35708 36418 35760
rect 28445 35683 28503 35689
rect 28445 35680 28457 35683
rect 27632 35652 28457 35680
rect 27525 35643 27583 35649
rect 28445 35649 28457 35652
rect 28491 35649 28503 35683
rect 28445 35643 28503 35649
rect 28997 35683 29055 35689
rect 28997 35649 29009 35683
rect 29043 35680 29055 35683
rect 29086 35680 29092 35692
rect 29043 35652 29092 35680
rect 29043 35649 29055 35652
rect 28997 35643 29055 35649
rect 29086 35640 29092 35652
rect 29144 35640 29150 35692
rect 29264 35683 29322 35689
rect 29264 35649 29276 35683
rect 29310 35680 29322 35683
rect 29546 35680 29552 35692
rect 29310 35652 29552 35680
rect 29310 35649 29322 35652
rect 29264 35643 29322 35649
rect 29546 35640 29552 35652
rect 29604 35640 29610 35692
rect 30282 35640 30288 35692
rect 30340 35680 30346 35692
rect 30929 35683 30987 35689
rect 30929 35680 30941 35683
rect 30340 35652 30941 35680
rect 30340 35640 30346 35652
rect 30929 35649 30941 35652
rect 30975 35649 30987 35683
rect 30929 35643 30987 35649
rect 32122 35640 32128 35692
rect 32180 35640 32186 35692
rect 32306 35640 32312 35692
rect 32364 35640 32370 35692
rect 33134 35640 33140 35692
rect 33192 35689 33198 35692
rect 33192 35683 33220 35689
rect 33208 35649 33220 35683
rect 33192 35643 33220 35649
rect 33192 35640 33198 35643
rect 40034 35640 40040 35692
rect 40092 35640 40098 35692
rect 46477 35683 46535 35689
rect 46477 35649 46489 35683
rect 46523 35680 46535 35683
rect 46842 35680 46848 35692
rect 46523 35652 46848 35680
rect 46523 35649 46535 35652
rect 46477 35643 46535 35649
rect 46842 35640 46848 35652
rect 46900 35640 46906 35692
rect 26605 35615 26663 35621
rect 26605 35581 26617 35615
rect 26651 35581 26663 35615
rect 26605 35575 26663 35581
rect 26970 35572 26976 35624
rect 27028 35572 27034 35624
rect 28902 35612 28908 35624
rect 28828 35584 28908 35612
rect 28828 35553 28856 35584
rect 28902 35572 28908 35584
rect 28960 35572 28966 35624
rect 31113 35615 31171 35621
rect 31113 35581 31125 35615
rect 31159 35612 31171 35615
rect 31386 35612 31392 35624
rect 31159 35584 31392 35612
rect 31159 35581 31171 35584
rect 31113 35575 31171 35581
rect 31386 35572 31392 35584
rect 31444 35572 31450 35624
rect 32674 35572 32680 35624
rect 32732 35612 32738 35624
rect 33045 35615 33103 35621
rect 33045 35612 33057 35615
rect 32732 35584 33057 35612
rect 32732 35572 32738 35584
rect 33045 35581 33057 35584
rect 33091 35581 33103 35615
rect 33045 35575 33103 35581
rect 33318 35572 33324 35624
rect 33376 35572 33382 35624
rect 35713 35615 35771 35621
rect 35713 35581 35725 35615
rect 35759 35581 35771 35615
rect 35713 35575 35771 35581
rect 27433 35547 27491 35553
rect 27433 35544 27445 35547
rect 26528 35516 27445 35544
rect 27433 35513 27445 35516
rect 27479 35513 27491 35547
rect 27433 35507 27491 35513
rect 28813 35547 28871 35553
rect 28813 35513 28825 35547
rect 28859 35513 28871 35547
rect 28813 35507 28871 35513
rect 30558 35504 30564 35556
rect 30616 35544 30622 35556
rect 32769 35547 32827 35553
rect 32769 35544 32781 35547
rect 30616 35516 32781 35544
rect 30616 35504 30622 35516
rect 32769 35513 32781 35516
rect 32815 35513 32827 35547
rect 32769 35507 32827 35513
rect 24176 35448 24808 35476
rect 25961 35479 26019 35485
rect 24176 35436 24182 35448
rect 25961 35445 25973 35479
rect 26007 35476 26019 35479
rect 26878 35476 26884 35488
rect 26007 35448 26884 35476
rect 26007 35445 26019 35448
rect 25961 35439 26019 35445
rect 26878 35436 26884 35448
rect 26936 35436 26942 35488
rect 28905 35479 28963 35485
rect 28905 35445 28917 35479
rect 28951 35476 28963 35479
rect 28994 35476 29000 35488
rect 28951 35448 29000 35476
rect 28951 35445 28963 35448
rect 28905 35439 28963 35445
rect 28994 35436 29000 35448
rect 29052 35436 29058 35488
rect 29730 35436 29736 35488
rect 29788 35476 29794 35488
rect 30469 35479 30527 35485
rect 30469 35476 30481 35479
rect 29788 35448 30481 35476
rect 29788 35436 29794 35448
rect 30469 35445 30481 35448
rect 30515 35445 30527 35479
rect 35728 35476 35756 35575
rect 39758 35572 39764 35624
rect 39816 35572 39822 35624
rect 35986 35476 35992 35488
rect 35728 35448 35992 35476
rect 30469 35439 30527 35445
rect 35986 35436 35992 35448
rect 36044 35436 36050 35488
rect 40773 35479 40831 35485
rect 40773 35445 40785 35479
rect 40819 35476 40831 35479
rect 41230 35476 41236 35488
rect 40819 35448 41236 35476
rect 40819 35445 40831 35448
rect 40773 35439 40831 35445
rect 41230 35436 41236 35448
rect 41288 35436 41294 35488
rect 46658 35436 46664 35488
rect 46716 35436 46722 35488
rect 1104 35386 47104 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 47104 35386
rect 1104 35312 47104 35334
rect 4522 35232 4528 35284
rect 4580 35272 4586 35284
rect 4982 35272 4988 35284
rect 4580 35244 4988 35272
rect 4580 35232 4586 35244
rect 4982 35232 4988 35244
rect 5040 35232 5046 35284
rect 6086 35232 6092 35284
rect 6144 35272 6150 35284
rect 6144 35244 8892 35272
rect 6144 35232 6150 35244
rect 3418 35164 3424 35216
rect 3476 35204 3482 35216
rect 3513 35207 3571 35213
rect 3513 35204 3525 35207
rect 3476 35176 3525 35204
rect 3476 35164 3482 35176
rect 3513 35173 3525 35176
rect 3559 35204 3571 35207
rect 3559 35176 5028 35204
rect 3559 35173 3571 35176
rect 3513 35167 3571 35173
rect 4249 35139 4307 35145
rect 4249 35105 4261 35139
rect 4295 35136 4307 35139
rect 4614 35136 4620 35148
rect 4295 35108 4620 35136
rect 4295 35105 4307 35108
rect 4249 35099 4307 35105
rect 4614 35096 4620 35108
rect 4672 35096 4678 35148
rect 4890 35096 4896 35148
rect 4948 35096 4954 35148
rect 5000 35136 5028 35176
rect 7926 35164 7932 35216
rect 7984 35164 7990 35216
rect 8864 35204 8892 35244
rect 8938 35232 8944 35284
rect 8996 35232 9002 35284
rect 11885 35275 11943 35281
rect 10612 35244 11652 35272
rect 10612 35204 10640 35244
rect 8864 35176 10640 35204
rect 10686 35164 10692 35216
rect 10744 35213 10750 35216
rect 10744 35167 10753 35213
rect 10744 35164 10750 35167
rect 5166 35136 5172 35148
rect 5000 35108 5172 35136
rect 5166 35096 5172 35108
rect 5224 35096 5230 35148
rect 5258 35096 5264 35148
rect 5316 35145 5322 35148
rect 5316 35139 5344 35145
rect 5332 35105 5344 35139
rect 5316 35099 5344 35105
rect 5445 35139 5503 35145
rect 5445 35105 5457 35139
rect 5491 35136 5503 35139
rect 5491 35108 6040 35136
rect 5491 35105 5503 35108
rect 5445 35099 5503 35105
rect 5316 35096 5322 35099
rect 1762 35028 1768 35080
rect 1820 35068 1826 35080
rect 2130 35068 2136 35080
rect 1820 35040 2136 35068
rect 1820 35028 1826 35040
rect 2130 35028 2136 35040
rect 2188 35028 2194 35080
rect 2400 35071 2458 35077
rect 2400 35037 2412 35071
rect 2446 35068 2458 35071
rect 3602 35068 3608 35080
rect 2446 35040 3608 35068
rect 2446 35037 2458 35040
rect 2400 35031 2458 35037
rect 3602 35028 3608 35040
rect 3660 35028 3666 35080
rect 4433 35071 4491 35077
rect 4433 35037 4445 35071
rect 4479 35037 4491 35071
rect 4433 35031 4491 35037
rect 4448 34932 4476 35031
rect 6012 35000 6040 35108
rect 6086 35096 6092 35148
rect 6144 35096 6150 35148
rect 8202 35096 8208 35148
rect 8260 35136 8266 35148
rect 8573 35139 8631 35145
rect 8573 35136 8585 35139
rect 8260 35108 8585 35136
rect 8260 35096 8266 35108
rect 8573 35105 8585 35108
rect 8619 35105 8631 35139
rect 8573 35099 8631 35105
rect 8662 35096 8668 35148
rect 8720 35136 8726 35148
rect 9214 35136 9220 35148
rect 8720 35108 9220 35136
rect 8720 35096 8726 35108
rect 9214 35096 9220 35108
rect 9272 35136 9278 35148
rect 9493 35139 9551 35145
rect 9493 35136 9505 35139
rect 9272 35108 9505 35136
rect 9272 35096 9278 35108
rect 9493 35105 9505 35108
rect 9539 35105 9551 35139
rect 9493 35099 9551 35105
rect 10318 35096 10324 35148
rect 10376 35136 10382 35148
rect 11082 35139 11140 35145
rect 11082 35136 11094 35139
rect 10376 35108 11094 35136
rect 10376 35096 10382 35108
rect 11082 35105 11094 35108
rect 11128 35105 11140 35139
rect 11624 35136 11652 35244
rect 11885 35241 11897 35275
rect 11931 35272 11943 35275
rect 13722 35272 13728 35284
rect 11931 35244 13728 35272
rect 11931 35241 11943 35244
rect 11885 35235 11943 35241
rect 13722 35232 13728 35244
rect 13780 35232 13786 35284
rect 14553 35275 14611 35281
rect 14553 35241 14565 35275
rect 14599 35272 14611 35275
rect 18782 35272 18788 35284
rect 14599 35244 18788 35272
rect 14599 35241 14611 35244
rect 14553 35235 14611 35241
rect 18782 35232 18788 35244
rect 18840 35232 18846 35284
rect 19794 35232 19800 35284
rect 19852 35272 19858 35284
rect 19852 35244 23428 35272
rect 19852 35232 19858 35244
rect 12621 35207 12679 35213
rect 12621 35173 12633 35207
rect 12667 35204 12679 35207
rect 17310 35204 17316 35216
rect 12667 35176 17316 35204
rect 12667 35173 12679 35176
rect 12621 35167 12679 35173
rect 17310 35164 17316 35176
rect 17368 35164 17374 35216
rect 19610 35164 19616 35216
rect 19668 35204 19674 35216
rect 19668 35176 20300 35204
rect 19668 35164 19674 35176
rect 12345 35139 12403 35145
rect 12345 35136 12357 35139
rect 11624 35108 12357 35136
rect 11082 35099 11140 35105
rect 12345 35105 12357 35108
rect 12391 35105 12403 35139
rect 12345 35099 12403 35105
rect 13078 35096 13084 35148
rect 13136 35136 13142 35148
rect 13136 35108 14504 35136
rect 13136 35096 13142 35108
rect 6457 35071 6515 35077
rect 6457 35037 6469 35071
rect 6503 35037 6515 35071
rect 6457 35031 6515 35037
rect 6472 35000 6500 35031
rect 6546 35028 6552 35080
rect 6604 35028 6610 35080
rect 6822 35077 6828 35080
rect 6816 35068 6828 35077
rect 6783 35040 6828 35068
rect 6816 35031 6828 35040
rect 6822 35028 6828 35031
rect 6880 35028 6886 35080
rect 9309 35071 9367 35077
rect 9309 35037 9321 35071
rect 9355 35068 9367 35071
rect 9398 35068 9404 35080
rect 9355 35040 9404 35068
rect 9355 35037 9367 35040
rect 9309 35031 9367 35037
rect 9398 35028 9404 35040
rect 9456 35068 9462 35080
rect 10045 35071 10103 35077
rect 10045 35068 10057 35071
rect 9456 35040 10057 35068
rect 9456 35028 9462 35040
rect 10045 35037 10057 35040
rect 10091 35037 10103 35071
rect 10045 35031 10103 35037
rect 10229 35071 10287 35077
rect 10229 35037 10241 35071
rect 10275 35037 10287 35071
rect 10229 35031 10287 35037
rect 6012 34972 6408 35000
rect 6472 34972 8064 35000
rect 4706 34932 4712 34944
rect 4448 34904 4712 34932
rect 4706 34892 4712 34904
rect 4764 34892 4770 34944
rect 5534 34892 5540 34944
rect 5592 34932 5598 34944
rect 6012 34932 6040 34972
rect 5592 34904 6040 34932
rect 5592 34892 5598 34904
rect 6270 34892 6276 34944
rect 6328 34892 6334 34944
rect 6380 34932 6408 34972
rect 6914 34932 6920 34944
rect 6380 34904 6920 34932
rect 6914 34892 6920 34904
rect 6972 34892 6978 34944
rect 8036 34941 8064 34972
rect 8386 34960 8392 35012
rect 8444 35000 8450 35012
rect 9490 35000 9496 35012
rect 8444 34972 9496 35000
rect 8444 34960 8450 34972
rect 9490 34960 9496 34972
rect 9548 34960 9554 35012
rect 9674 34960 9680 35012
rect 9732 35000 9738 35012
rect 10244 35000 10272 35031
rect 10962 35028 10968 35080
rect 11020 35028 11026 35080
rect 11238 35028 11244 35080
rect 11296 35028 11302 35080
rect 12434 35028 12440 35080
rect 12492 35028 12498 35080
rect 13541 35071 13599 35077
rect 13541 35037 13553 35071
rect 13587 35037 13599 35071
rect 13541 35031 13599 35037
rect 9732 34972 10272 35000
rect 9732 34960 9738 34972
rect 8021 34935 8079 34941
rect 8021 34901 8033 34935
rect 8067 34901 8079 34935
rect 8021 34895 8079 34901
rect 8481 34935 8539 34941
rect 8481 34901 8493 34935
rect 8527 34932 8539 34935
rect 9306 34932 9312 34944
rect 8527 34904 9312 34932
rect 8527 34901 8539 34904
rect 8481 34895 8539 34901
rect 9306 34892 9312 34904
rect 9364 34932 9370 34944
rect 9401 34935 9459 34941
rect 9401 34932 9413 34935
rect 9364 34904 9413 34932
rect 9364 34892 9370 34904
rect 9401 34901 9413 34904
rect 9447 34901 9459 34935
rect 10244 34932 10272 34972
rect 11790 34960 11796 35012
rect 11848 35000 11854 35012
rect 13556 35000 13584 35031
rect 13630 35028 13636 35080
rect 13688 35028 13694 35080
rect 13817 35071 13875 35077
rect 13817 35037 13829 35071
rect 13863 35068 13875 35071
rect 14277 35071 14335 35077
rect 14277 35068 14289 35071
rect 13863 35040 14289 35068
rect 13863 35037 13875 35040
rect 13817 35031 13875 35037
rect 14277 35037 14289 35040
rect 14323 35037 14335 35071
rect 14277 35031 14335 35037
rect 14366 35028 14372 35080
rect 14424 35028 14430 35080
rect 14476 35068 14504 35108
rect 14734 35096 14740 35148
rect 14792 35136 14798 35148
rect 19978 35136 19984 35148
rect 14792 35108 17816 35136
rect 14792 35096 14798 35108
rect 14645 35071 14703 35077
rect 14645 35068 14657 35071
rect 14476 35040 14657 35068
rect 14645 35037 14657 35040
rect 14691 35037 14703 35071
rect 14645 35031 14703 35037
rect 17678 35028 17684 35080
rect 17736 35028 17742 35080
rect 17788 35068 17816 35108
rect 19444 35108 19984 35136
rect 18506 35068 18512 35080
rect 17788 35040 18512 35068
rect 18506 35028 18512 35040
rect 18564 35028 18570 35080
rect 19444 35077 19472 35108
rect 19978 35096 19984 35108
rect 20036 35096 20042 35148
rect 20272 35136 20300 35176
rect 20346 35164 20352 35216
rect 20404 35164 20410 35216
rect 21910 35164 21916 35216
rect 21968 35204 21974 35216
rect 22189 35207 22247 35213
rect 22189 35204 22201 35207
rect 21968 35176 22201 35204
rect 21968 35164 21974 35176
rect 22189 35173 22201 35176
rect 22235 35173 22247 35207
rect 22189 35167 22247 35173
rect 20438 35136 20444 35148
rect 20272 35108 20444 35136
rect 20438 35096 20444 35108
rect 20496 35096 20502 35148
rect 20806 35096 20812 35148
rect 20864 35096 20870 35148
rect 23400 35136 23428 35244
rect 23474 35232 23480 35284
rect 23532 35232 23538 35284
rect 27246 35232 27252 35284
rect 27304 35272 27310 35284
rect 27525 35275 27583 35281
rect 27525 35272 27537 35275
rect 27304 35244 27537 35272
rect 27304 35232 27310 35244
rect 27525 35241 27537 35244
rect 27571 35241 27583 35275
rect 27525 35235 27583 35241
rect 29086 35232 29092 35284
rect 29144 35272 29150 35284
rect 29270 35272 29276 35284
rect 29144 35244 29276 35272
rect 29144 35232 29150 35244
rect 29270 35232 29276 35244
rect 29328 35232 29334 35284
rect 29546 35232 29552 35284
rect 29604 35232 29610 35284
rect 37366 35232 37372 35284
rect 37424 35232 37430 35284
rect 26237 35207 26295 35213
rect 24320 35176 25176 35204
rect 24320 35136 24348 35176
rect 23400 35108 24348 35136
rect 24394 35096 24400 35148
rect 24452 35096 24458 35148
rect 25038 35136 25044 35148
rect 24504 35108 25044 35136
rect 19429 35071 19487 35077
rect 19429 35037 19441 35071
rect 19475 35037 19487 35071
rect 19429 35031 19487 35037
rect 19527 35040 20300 35068
rect 11848 34972 13584 35000
rect 11848 34960 11854 34972
rect 14090 34960 14096 35012
rect 14148 34960 14154 35012
rect 17948 35003 18006 35009
rect 17948 34969 17960 35003
rect 17994 35000 18006 35003
rect 18322 35000 18328 35012
rect 17994 34972 18328 35000
rect 17994 34969 18006 34972
rect 17948 34963 18006 34969
rect 18322 34960 18328 34972
rect 18380 34960 18386 35012
rect 19527 35000 19555 35040
rect 18432 34972 19555 35000
rect 11054 34932 11060 34944
rect 10244 34904 11060 34932
rect 9401 34895 9459 34901
rect 11054 34892 11060 34904
rect 11112 34892 11118 34944
rect 11514 34892 11520 34944
rect 11572 34932 11578 34944
rect 11977 34935 12035 34941
rect 11977 34932 11989 34935
rect 11572 34904 11989 34932
rect 11572 34892 11578 34904
rect 11977 34901 11989 34904
rect 12023 34901 12035 34935
rect 11977 34895 12035 34901
rect 13173 34935 13231 34941
rect 13173 34901 13185 34935
rect 13219 34932 13231 34935
rect 13814 34932 13820 34944
rect 13219 34904 13820 34932
rect 13219 34901 13231 34904
rect 13173 34895 13231 34901
rect 13814 34892 13820 34904
rect 13872 34892 13878 34944
rect 16022 34892 16028 34944
rect 16080 34932 16086 34944
rect 18432 34932 18460 34972
rect 19978 34960 19984 35012
rect 20036 35000 20042 35012
rect 20165 35003 20223 35009
rect 20165 35000 20177 35003
rect 20036 34972 20177 35000
rect 20036 34960 20042 34972
rect 20165 34969 20177 34972
rect 20211 34969 20223 35003
rect 20272 35000 20300 35040
rect 20898 35028 20904 35080
rect 20956 35068 20962 35080
rect 21065 35071 21123 35077
rect 21065 35068 21077 35071
rect 20956 35040 21077 35068
rect 20956 35028 20962 35040
rect 21065 35037 21077 35040
rect 21111 35037 21123 35071
rect 21065 35031 21123 35037
rect 22738 35028 22744 35080
rect 22796 35068 22802 35080
rect 23201 35071 23259 35077
rect 23201 35068 23213 35071
rect 22796 35040 23213 35068
rect 22796 35028 22802 35040
rect 23201 35037 23213 35040
rect 23247 35037 23259 35071
rect 23201 35031 23259 35037
rect 23290 35028 23296 35080
rect 23348 35028 23354 35080
rect 23569 35071 23627 35077
rect 23569 35037 23581 35071
rect 23615 35037 23627 35071
rect 23569 35031 23627 35037
rect 23584 35000 23612 35031
rect 24026 35028 24032 35080
rect 24084 35028 24090 35080
rect 24210 35028 24216 35080
rect 24268 35068 24274 35080
rect 24504 35068 24532 35108
rect 25038 35096 25044 35108
rect 25096 35096 25102 35148
rect 25148 35136 25176 35176
rect 26237 35173 26249 35207
rect 26283 35204 26295 35207
rect 26605 35207 26663 35213
rect 26605 35204 26617 35207
rect 26283 35176 26617 35204
rect 26283 35173 26295 35176
rect 26237 35167 26295 35173
rect 26605 35173 26617 35176
rect 26651 35173 26663 35207
rect 26605 35167 26663 35173
rect 26878 35164 26884 35216
rect 26936 35204 26942 35216
rect 27157 35207 27215 35213
rect 27157 35204 27169 35207
rect 26936 35176 27169 35204
rect 26936 35164 26942 35176
rect 27157 35173 27169 35176
rect 27203 35173 27215 35207
rect 27157 35167 27215 35173
rect 27341 35207 27399 35213
rect 27341 35173 27353 35207
rect 27387 35204 27399 35207
rect 30650 35204 30656 35216
rect 27387 35176 29408 35204
rect 27387 35173 27399 35176
rect 27341 35167 27399 35173
rect 29273 35139 29331 35145
rect 29273 35136 29285 35139
rect 25148 35108 29285 35136
rect 29273 35105 29285 35108
rect 29319 35105 29331 35139
rect 29273 35099 29331 35105
rect 24268 35040 24532 35068
rect 24581 35071 24639 35077
rect 24268 35028 24274 35040
rect 24581 35037 24593 35071
rect 24627 35068 24639 35071
rect 24762 35068 24768 35080
rect 24627 35040 24768 35068
rect 24627 35037 24639 35040
rect 24581 35031 24639 35037
rect 24762 35028 24768 35040
rect 24820 35028 24826 35080
rect 25314 35028 25320 35080
rect 25372 35028 25378 35080
rect 25406 35028 25412 35080
rect 25464 35077 25470 35080
rect 25464 35071 25492 35077
rect 25480 35037 25492 35071
rect 25464 35031 25492 35037
rect 25464 35028 25470 35031
rect 25590 35028 25596 35080
rect 25648 35028 25654 35080
rect 26786 35028 26792 35080
rect 26844 35068 26850 35080
rect 26881 35071 26939 35077
rect 26881 35068 26893 35071
rect 26844 35040 26893 35068
rect 26844 35028 26850 35040
rect 26881 35037 26893 35040
rect 26927 35037 26939 35071
rect 26881 35031 26939 35037
rect 27706 35028 27712 35080
rect 27764 35028 27770 35080
rect 27890 35028 27896 35080
rect 27948 35028 27954 35080
rect 27985 35071 28043 35077
rect 27985 35037 27997 35071
rect 28031 35068 28043 35071
rect 28074 35068 28080 35080
rect 28031 35040 28080 35068
rect 28031 35037 28043 35040
rect 27985 35031 28043 35037
rect 28074 35028 28080 35040
rect 28132 35068 28138 35080
rect 28718 35068 28724 35080
rect 28132 35040 28724 35068
rect 28132 35028 28138 35040
rect 28718 35028 28724 35040
rect 28776 35028 28782 35080
rect 28813 35071 28871 35077
rect 28813 35037 28825 35071
rect 28859 35068 28871 35071
rect 28902 35068 28908 35080
rect 28859 35040 28908 35068
rect 28859 35037 28871 35040
rect 28813 35031 28871 35037
rect 28902 35028 28908 35040
rect 28960 35028 28966 35080
rect 28994 35028 29000 35080
rect 29052 35028 29058 35080
rect 29086 35028 29092 35080
rect 29144 35028 29150 35080
rect 29380 35077 29408 35176
rect 29932 35176 30656 35204
rect 29932 35080 29960 35176
rect 30650 35164 30656 35176
rect 30708 35164 30714 35216
rect 30558 35096 30564 35148
rect 30616 35096 30622 35148
rect 30834 35096 30840 35148
rect 30892 35096 30898 35148
rect 30926 35096 30932 35148
rect 30984 35145 30990 35148
rect 30984 35139 31012 35145
rect 31000 35105 31012 35139
rect 33318 35136 33324 35148
rect 30984 35099 31012 35105
rect 31128 35108 33324 35136
rect 30984 35096 30990 35099
rect 31128 35080 31156 35108
rect 33318 35096 33324 35108
rect 33376 35096 33382 35148
rect 29365 35071 29423 35077
rect 29365 35037 29377 35071
rect 29411 35037 29423 35071
rect 29365 35031 29423 35037
rect 29730 35028 29736 35080
rect 29788 35028 29794 35080
rect 29914 35028 29920 35080
rect 29972 35028 29978 35080
rect 30101 35071 30159 35077
rect 30101 35037 30113 35071
rect 30147 35068 30159 35071
rect 30282 35068 30288 35080
rect 30147 35040 30288 35068
rect 30147 35037 30159 35040
rect 30101 35031 30159 35037
rect 30282 35028 30288 35040
rect 30340 35028 30346 35080
rect 31110 35028 31116 35080
rect 31168 35028 31174 35080
rect 33594 35028 33600 35080
rect 33652 35068 33658 35080
rect 34238 35068 34244 35080
rect 33652 35040 34244 35068
rect 33652 35028 33658 35040
rect 34238 35028 34244 35040
rect 34296 35028 34302 35080
rect 34701 35071 34759 35077
rect 34701 35068 34713 35071
rect 34440 35040 34713 35068
rect 20272 34972 23612 35000
rect 26329 35003 26387 35009
rect 20165 34963 20223 34969
rect 26329 34969 26341 35003
rect 26375 34969 26387 35003
rect 27798 35000 27804 35012
rect 26329 34963 26387 34969
rect 27264 34972 27804 35000
rect 16080 34904 18460 34932
rect 16080 34892 16086 34904
rect 19058 34892 19064 34944
rect 19116 34892 19122 34944
rect 20180 34932 20208 34963
rect 20530 34932 20536 34944
rect 20180 34904 20536 34932
rect 20530 34892 20536 34904
rect 20588 34892 20594 34944
rect 23014 34892 23020 34944
rect 23072 34892 23078 34944
rect 23845 34935 23903 34941
rect 23845 34901 23857 34935
rect 23891 34932 23903 34935
rect 23934 34932 23940 34944
rect 23891 34904 23940 34932
rect 23891 34901 23903 34904
rect 23845 34895 23903 34901
rect 23934 34892 23940 34904
rect 23992 34892 23998 34944
rect 25866 34892 25872 34944
rect 25924 34932 25930 34944
rect 26344 34932 26372 34963
rect 25924 34904 26372 34932
rect 26789 34935 26847 34941
rect 25924 34892 25930 34904
rect 26789 34901 26801 34935
rect 26835 34932 26847 34935
rect 27264 34932 27292 34972
rect 27798 34960 27804 34972
rect 27856 34960 27862 35012
rect 34440 34944 34468 35040
rect 34701 35037 34713 35040
rect 34747 35037 34759 35071
rect 34701 35031 34759 35037
rect 34974 35028 34980 35080
rect 35032 35028 35038 35080
rect 35986 35028 35992 35080
rect 36044 35028 36050 35080
rect 36256 35071 36314 35077
rect 36256 35037 36268 35071
rect 36302 35068 36314 35071
rect 36538 35068 36544 35080
rect 36302 35040 36544 35068
rect 36302 35037 36314 35040
rect 36256 35031 36314 35037
rect 36538 35028 36544 35040
rect 36596 35028 36602 35080
rect 39022 35028 39028 35080
rect 39080 35068 39086 35080
rect 39209 35071 39267 35077
rect 39209 35068 39221 35071
rect 39080 35040 39221 35068
rect 39080 35028 39086 35040
rect 39209 35037 39221 35040
rect 39255 35037 39267 35071
rect 39209 35031 39267 35037
rect 39758 35028 39764 35080
rect 39816 35068 39822 35080
rect 39853 35071 39911 35077
rect 39853 35068 39865 35071
rect 39816 35040 39865 35068
rect 39816 35028 39822 35040
rect 39853 35037 39865 35040
rect 39899 35037 39911 35071
rect 39853 35031 39911 35037
rect 40126 35028 40132 35080
rect 40184 35028 40190 35080
rect 36630 34960 36636 35012
rect 36688 35000 36694 35012
rect 38289 35003 38347 35009
rect 38289 35000 38301 35003
rect 36688 34972 38301 35000
rect 36688 34960 36694 34972
rect 38289 34969 38301 34972
rect 38335 35000 38347 35003
rect 38335 34972 38516 35000
rect 38335 34969 38347 34972
rect 38289 34963 38347 34969
rect 26835 34904 27292 34932
rect 26835 34901 26847 34904
rect 26789 34895 26847 34901
rect 27706 34892 27712 34944
rect 27764 34932 27770 34944
rect 29546 34932 29552 34944
rect 27764 34904 29552 34932
rect 27764 34892 27770 34904
rect 29546 34892 29552 34904
rect 29604 34892 29610 34944
rect 29730 34892 29736 34944
rect 29788 34932 29794 34944
rect 31757 34935 31815 34941
rect 31757 34932 31769 34935
rect 29788 34904 31769 34932
rect 29788 34892 29794 34904
rect 31757 34901 31769 34904
rect 31803 34901 31815 34935
rect 31757 34895 31815 34901
rect 34422 34892 34428 34944
rect 34480 34892 34486 34944
rect 35713 34935 35771 34941
rect 35713 34901 35725 34935
rect 35759 34932 35771 34935
rect 37826 34932 37832 34944
rect 35759 34904 37832 34932
rect 35759 34901 35771 34904
rect 35713 34895 35771 34901
rect 37826 34892 37832 34904
rect 37884 34892 37890 34944
rect 38378 34892 38384 34944
rect 38436 34892 38442 34944
rect 38488 34932 38516 34972
rect 39301 34935 39359 34941
rect 39301 34932 39313 34935
rect 38488 34904 39313 34932
rect 39301 34901 39313 34904
rect 39347 34901 39359 34935
rect 39301 34895 39359 34901
rect 40865 34935 40923 34941
rect 40865 34901 40877 34935
rect 40911 34932 40923 34935
rect 41414 34932 41420 34944
rect 40911 34904 41420 34932
rect 40911 34901 40923 34904
rect 40865 34895 40923 34901
rect 41414 34892 41420 34904
rect 41472 34892 41478 34944
rect 1104 34842 47104 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 47104 34842
rect 1104 34768 47104 34790
rect 3053 34731 3111 34737
rect 3053 34697 3065 34731
rect 3099 34728 3111 34731
rect 3786 34728 3792 34740
rect 3099 34700 3792 34728
rect 3099 34697 3111 34700
rect 3053 34691 3111 34697
rect 3786 34688 3792 34700
rect 3844 34688 3850 34740
rect 7929 34731 7987 34737
rect 7929 34697 7941 34731
rect 7975 34728 7987 34731
rect 8386 34728 8392 34740
rect 7975 34700 8392 34728
rect 7975 34697 7987 34700
rect 7929 34691 7987 34697
rect 8386 34688 8392 34700
rect 8444 34688 8450 34740
rect 9398 34688 9404 34740
rect 9456 34688 9462 34740
rect 9490 34688 9496 34740
rect 9548 34728 9554 34740
rect 10410 34728 10416 34740
rect 9548 34700 10416 34728
rect 9548 34688 9554 34700
rect 10410 34688 10416 34700
rect 10468 34728 10474 34740
rect 10962 34728 10968 34740
rect 10468 34700 10968 34728
rect 10468 34688 10474 34700
rect 10962 34688 10968 34700
rect 11020 34688 11026 34740
rect 11333 34731 11391 34737
rect 11333 34697 11345 34731
rect 11379 34728 11391 34731
rect 11790 34728 11796 34740
rect 11379 34700 11796 34728
rect 11379 34697 11391 34700
rect 11333 34691 11391 34697
rect 11790 34688 11796 34700
rect 11848 34688 11854 34740
rect 14182 34688 14188 34740
rect 14240 34728 14246 34740
rect 14461 34731 14519 34737
rect 14461 34728 14473 34731
rect 14240 34700 14473 34728
rect 14240 34688 14246 34700
rect 14461 34697 14473 34700
rect 14507 34728 14519 34731
rect 14921 34731 14979 34737
rect 14921 34728 14933 34731
rect 14507 34700 14933 34728
rect 14507 34697 14519 34700
rect 14461 34691 14519 34697
rect 14921 34697 14933 34700
rect 14967 34697 14979 34731
rect 14921 34691 14979 34697
rect 16117 34731 16175 34737
rect 16117 34697 16129 34731
rect 16163 34697 16175 34731
rect 16117 34691 16175 34697
rect 1486 34620 1492 34672
rect 1544 34620 1550 34672
rect 3418 34620 3424 34672
rect 3476 34620 3482 34672
rect 3513 34663 3571 34669
rect 3513 34629 3525 34663
rect 3559 34660 3571 34663
rect 5350 34660 5356 34672
rect 3559 34632 5356 34660
rect 3559 34629 3571 34632
rect 3513 34623 3571 34629
rect 5350 34620 5356 34632
rect 5408 34620 5414 34672
rect 6270 34620 6276 34672
rect 6328 34660 6334 34672
rect 6794 34663 6852 34669
rect 6794 34660 6806 34663
rect 6328 34632 6806 34660
rect 6328 34620 6334 34632
rect 6794 34629 6806 34632
rect 6840 34629 6852 34663
rect 6794 34623 6852 34629
rect 8018 34620 8024 34672
rect 8076 34660 8082 34672
rect 8076 34632 9352 34660
rect 8076 34620 8082 34632
rect 6546 34552 6552 34604
rect 6604 34552 6610 34604
rect 8294 34601 8300 34604
rect 8288 34592 8300 34601
rect 8255 34564 8300 34592
rect 8288 34555 8300 34564
rect 8294 34552 8300 34555
rect 8352 34552 8358 34604
rect 3605 34527 3663 34533
rect 3605 34493 3617 34527
rect 3651 34493 3663 34527
rect 3605 34487 3663 34493
rect 8021 34527 8079 34533
rect 8021 34493 8033 34527
rect 8067 34493 8079 34527
rect 9324 34524 9352 34632
rect 9416 34592 9444 34688
rect 12345 34663 12403 34669
rect 12345 34629 12357 34663
rect 12391 34660 12403 34663
rect 16022 34660 16028 34672
rect 12391 34632 16028 34660
rect 12391 34629 12403 34632
rect 12345 34623 12403 34629
rect 16022 34620 16028 34632
rect 16080 34620 16086 34672
rect 16132 34660 16160 34691
rect 17310 34688 17316 34740
rect 17368 34728 17374 34740
rect 17368 34700 23244 34728
rect 17368 34688 17374 34700
rect 16914 34663 16972 34669
rect 16914 34660 16926 34663
rect 16132 34632 16926 34660
rect 16914 34629 16926 34632
rect 16960 34629 16972 34663
rect 16914 34623 16972 34629
rect 18233 34663 18291 34669
rect 18233 34629 18245 34663
rect 18279 34660 18291 34663
rect 18506 34660 18512 34672
rect 18279 34632 18512 34660
rect 18279 34629 18291 34632
rect 18233 34623 18291 34629
rect 18506 34620 18512 34632
rect 18564 34620 18570 34672
rect 19058 34620 19064 34672
rect 19116 34660 19122 34672
rect 19429 34663 19487 34669
rect 19429 34660 19441 34663
rect 19116 34632 19441 34660
rect 19116 34620 19122 34632
rect 19429 34629 19441 34632
rect 19475 34629 19487 34663
rect 23216 34660 23244 34700
rect 23290 34688 23296 34740
rect 23348 34728 23354 34740
rect 25225 34731 25283 34737
rect 25225 34728 25237 34731
rect 23348 34700 25237 34728
rect 23348 34688 23354 34700
rect 25225 34697 25237 34700
rect 25271 34697 25283 34731
rect 25225 34691 25283 34697
rect 25593 34731 25651 34737
rect 25593 34697 25605 34731
rect 25639 34728 25651 34731
rect 26234 34728 26240 34740
rect 25639 34700 26240 34728
rect 25639 34697 25651 34700
rect 25593 34691 25651 34697
rect 26234 34688 26240 34700
rect 26292 34688 26298 34740
rect 28537 34731 28595 34737
rect 28537 34697 28549 34731
rect 28583 34697 28595 34731
rect 28537 34691 28595 34697
rect 28552 34660 28580 34691
rect 29086 34688 29092 34740
rect 29144 34728 29150 34740
rect 29365 34731 29423 34737
rect 29365 34728 29377 34731
rect 29144 34700 29377 34728
rect 29144 34688 29150 34700
rect 29365 34697 29377 34700
rect 29411 34697 29423 34731
rect 29365 34691 29423 34697
rect 29730 34688 29736 34740
rect 29788 34688 29794 34740
rect 31757 34731 31815 34737
rect 31757 34728 31769 34731
rect 30116 34700 31769 34728
rect 23216 34632 25912 34660
rect 19429 34623 19487 34629
rect 9493 34595 9551 34601
rect 9493 34592 9505 34595
rect 9416 34564 9505 34592
rect 9493 34561 9505 34564
rect 9539 34561 9551 34595
rect 9493 34555 9551 34561
rect 9674 34552 9680 34604
rect 9732 34552 9738 34604
rect 10410 34552 10416 34604
rect 10468 34552 10474 34604
rect 13354 34601 13360 34604
rect 12069 34595 12127 34601
rect 12069 34592 12081 34595
rect 11256 34564 12081 34592
rect 9324 34496 10088 34524
rect 8021 34487 8079 34493
rect 3620 34456 3648 34487
rect 3694 34456 3700 34468
rect 3620 34428 3700 34456
rect 3694 34416 3700 34428
rect 3752 34416 3758 34468
rect 1578 34348 1584 34400
rect 1636 34348 1642 34400
rect 3970 34348 3976 34400
rect 4028 34388 4034 34400
rect 8036 34388 8064 34487
rect 10060 34456 10088 34496
rect 10134 34484 10140 34536
rect 10192 34484 10198 34536
rect 10226 34484 10232 34536
rect 10284 34524 10290 34536
rect 10530 34527 10588 34533
rect 10530 34524 10542 34527
rect 10284 34496 10542 34524
rect 10284 34484 10290 34496
rect 10530 34493 10542 34496
rect 10576 34493 10588 34527
rect 10530 34487 10588 34493
rect 10686 34484 10692 34536
rect 10744 34484 10750 34536
rect 10870 34484 10876 34536
rect 10928 34524 10934 34536
rect 11256 34524 11284 34564
rect 12069 34561 12081 34564
rect 12115 34561 12127 34595
rect 12069 34555 12127 34561
rect 13348 34555 13360 34601
rect 13354 34552 13360 34555
rect 13412 34552 13418 34604
rect 15010 34552 15016 34604
rect 15068 34552 15074 34604
rect 16298 34552 16304 34604
rect 16356 34552 16362 34604
rect 17678 34592 17684 34604
rect 16684 34564 17684 34592
rect 10928 34496 11284 34524
rect 10928 34484 10934 34496
rect 11514 34484 11520 34536
rect 11572 34524 11578 34536
rect 11701 34527 11759 34533
rect 11701 34524 11713 34527
rect 11572 34496 11713 34524
rect 11572 34484 11578 34496
rect 11701 34493 11713 34496
rect 11747 34493 11759 34527
rect 11701 34487 11759 34493
rect 12161 34527 12219 34533
rect 12161 34493 12173 34527
rect 12207 34524 12219 34527
rect 12434 34524 12440 34536
rect 12207 34496 12440 34524
rect 12207 34493 12219 34496
rect 12161 34487 12219 34493
rect 12434 34484 12440 34496
rect 12492 34484 12498 34536
rect 12618 34484 12624 34536
rect 12676 34524 12682 34536
rect 13081 34527 13139 34533
rect 13081 34524 13093 34527
rect 12676 34496 13093 34524
rect 12676 34484 12682 34496
rect 13081 34493 13093 34496
rect 13127 34493 13139 34527
rect 13081 34487 13139 34493
rect 14090 34484 14096 34536
rect 14148 34524 14154 34536
rect 14148 34496 15056 34524
rect 14148 34484 14154 34496
rect 10244 34456 10272 34484
rect 10060 34428 10272 34456
rect 15028 34456 15056 34496
rect 15102 34484 15108 34536
rect 15160 34484 15166 34536
rect 16684 34533 16712 34564
rect 17678 34552 17684 34564
rect 17736 34592 17742 34604
rect 18417 34595 18475 34601
rect 18417 34592 18429 34595
rect 17736 34564 18429 34592
rect 17736 34552 17742 34564
rect 18417 34561 18429 34564
rect 18463 34561 18475 34595
rect 18417 34555 18475 34561
rect 20346 34552 20352 34604
rect 20404 34592 20410 34604
rect 23290 34592 23296 34604
rect 20404 34564 23296 34592
rect 20404 34552 20410 34564
rect 23290 34552 23296 34564
rect 23348 34552 23354 34604
rect 23934 34601 23940 34604
rect 23928 34592 23940 34601
rect 23895 34564 23940 34592
rect 23928 34555 23940 34564
rect 23934 34552 23940 34555
rect 23992 34552 23998 34604
rect 25682 34552 25688 34604
rect 25740 34552 25746 34604
rect 16669 34527 16727 34533
rect 16669 34493 16681 34527
rect 16715 34493 16727 34527
rect 16669 34487 16727 34493
rect 16684 34456 16712 34487
rect 18690 34484 18696 34536
rect 18748 34524 18754 34536
rect 19521 34527 19579 34533
rect 19521 34524 19533 34527
rect 18748 34496 19533 34524
rect 18748 34484 18754 34496
rect 19521 34493 19533 34496
rect 19567 34493 19579 34527
rect 19521 34487 19579 34493
rect 19705 34527 19763 34533
rect 19705 34493 19717 34527
rect 19751 34493 19763 34527
rect 19705 34487 19763 34493
rect 15028 34428 16712 34456
rect 19720 34456 19748 34487
rect 23658 34484 23664 34536
rect 23716 34484 23722 34536
rect 24762 34484 24768 34536
rect 24820 34524 24826 34536
rect 24820 34496 25084 34524
rect 24820 34484 24826 34496
rect 23566 34456 23572 34468
rect 19720 34428 23572 34456
rect 23566 34416 23572 34428
rect 23624 34416 23630 34468
rect 25056 34465 25084 34496
rect 25774 34484 25780 34536
rect 25832 34484 25838 34536
rect 25884 34524 25912 34632
rect 27632 34632 28580 34660
rect 28997 34663 29055 34669
rect 27632 34601 27660 34632
rect 28997 34629 29009 34663
rect 29043 34660 29055 34663
rect 30116 34660 30144 34700
rect 31757 34697 31769 34700
rect 31803 34697 31815 34731
rect 31757 34691 31815 34697
rect 35437 34731 35495 34737
rect 35437 34697 35449 34731
rect 35483 34728 35495 34731
rect 37090 34728 37096 34740
rect 35483 34700 37096 34728
rect 35483 34697 35495 34700
rect 35437 34691 35495 34697
rect 37090 34688 37096 34700
rect 37148 34688 37154 34740
rect 37550 34688 37556 34740
rect 37608 34728 37614 34740
rect 37737 34731 37795 34737
rect 37737 34728 37749 34731
rect 37608 34700 37749 34728
rect 37608 34688 37614 34700
rect 37737 34697 37749 34700
rect 37783 34697 37795 34731
rect 37737 34691 37795 34697
rect 37826 34688 37832 34740
rect 37884 34728 37890 34740
rect 38010 34728 38016 34740
rect 37884 34700 38016 34728
rect 37884 34688 37890 34700
rect 38010 34688 38016 34700
rect 38068 34728 38074 34740
rect 39485 34731 39543 34737
rect 38068 34700 38516 34728
rect 38068 34688 38074 34700
rect 29043 34632 30144 34660
rect 37369 34663 37427 34669
rect 29043 34629 29055 34632
rect 28997 34623 29055 34629
rect 37369 34629 37381 34663
rect 37415 34660 37427 34663
rect 38350 34663 38408 34669
rect 38350 34660 38362 34663
rect 37415 34632 38362 34660
rect 37415 34629 37427 34632
rect 37369 34623 37427 34629
rect 38350 34629 38362 34632
rect 38396 34629 38408 34663
rect 38488 34660 38516 34700
rect 39485 34697 39497 34731
rect 39531 34728 39543 34731
rect 39574 34728 39580 34740
rect 39531 34700 39580 34728
rect 39531 34697 39543 34700
rect 39485 34691 39543 34697
rect 39574 34688 39580 34700
rect 39632 34688 39638 34740
rect 40589 34731 40647 34737
rect 40589 34697 40601 34731
rect 40635 34728 40647 34731
rect 44174 34728 44180 34740
rect 40635 34700 44180 34728
rect 40635 34697 40647 34700
rect 40589 34691 40647 34697
rect 44174 34688 44180 34700
rect 44232 34688 44238 34740
rect 38488 34632 42196 34660
rect 38350 34623 38408 34629
rect 42168 34604 42196 34632
rect 27617 34595 27675 34601
rect 27617 34561 27629 34595
rect 27663 34561 27675 34595
rect 27617 34555 27675 34561
rect 27709 34595 27767 34601
rect 27709 34561 27721 34595
rect 27755 34561 27767 34595
rect 27709 34555 27767 34561
rect 27433 34527 27491 34533
rect 25884 34496 27384 34524
rect 25041 34459 25099 34465
rect 25041 34425 25053 34459
rect 25087 34425 25099 34459
rect 25041 34419 25099 34425
rect 9398 34388 9404 34400
rect 4028 34360 9404 34388
rect 4028 34348 4034 34360
rect 9398 34348 9404 34360
rect 9456 34348 9462 34400
rect 14550 34348 14556 34400
rect 14608 34348 14614 34400
rect 16666 34348 16672 34400
rect 16724 34388 16730 34400
rect 18049 34391 18107 34397
rect 18049 34388 18061 34391
rect 16724 34360 18061 34388
rect 16724 34348 16730 34360
rect 18049 34357 18061 34360
rect 18095 34357 18107 34391
rect 18049 34351 18107 34357
rect 18506 34348 18512 34400
rect 18564 34388 18570 34400
rect 19061 34391 19119 34397
rect 19061 34388 19073 34391
rect 18564 34360 19073 34388
rect 18564 34348 18570 34360
rect 19061 34357 19073 34360
rect 19107 34357 19119 34391
rect 19061 34351 19119 34357
rect 22646 34348 22652 34400
rect 22704 34388 22710 34400
rect 26142 34388 26148 34400
rect 22704 34360 26148 34388
rect 22704 34348 22710 34360
rect 26142 34348 26148 34360
rect 26200 34348 26206 34400
rect 27356 34388 27384 34496
rect 27433 34493 27445 34527
rect 27479 34524 27491 34527
rect 27724 34524 27752 34555
rect 27798 34552 27804 34604
rect 27856 34592 27862 34604
rect 27985 34595 28043 34601
rect 27985 34592 27997 34595
rect 27856 34564 27997 34592
rect 27856 34552 27862 34564
rect 27985 34561 27997 34564
rect 28031 34561 28043 34595
rect 27985 34555 28043 34561
rect 28077 34595 28135 34601
rect 28077 34561 28089 34595
rect 28123 34592 28135 34595
rect 28350 34592 28356 34604
rect 28123 34564 28356 34592
rect 28123 34561 28135 34564
rect 28077 34555 28135 34561
rect 28350 34552 28356 34564
rect 28408 34552 28414 34604
rect 28534 34552 28540 34604
rect 28592 34592 28598 34604
rect 28813 34595 28871 34601
rect 28813 34592 28825 34595
rect 28592 34564 28825 34592
rect 28592 34552 28598 34564
rect 28813 34561 28825 34564
rect 28859 34561 28871 34595
rect 28813 34555 28871 34561
rect 29086 34552 29092 34604
rect 29144 34552 29150 34604
rect 29546 34552 29552 34604
rect 29604 34592 29610 34604
rect 29730 34592 29736 34604
rect 29604 34564 29736 34592
rect 29604 34552 29610 34564
rect 29730 34552 29736 34564
rect 29788 34552 29794 34604
rect 29825 34595 29883 34601
rect 29825 34561 29837 34595
rect 29871 34561 29883 34595
rect 29825 34555 29883 34561
rect 28629 34527 28687 34533
rect 28629 34524 28641 34527
rect 27479 34496 27660 34524
rect 27724 34496 28028 34524
rect 27479 34493 27491 34496
rect 27433 34487 27491 34493
rect 27632 34468 27660 34496
rect 27614 34416 27620 34468
rect 27672 34416 27678 34468
rect 28000 34456 28028 34496
rect 28184 34496 28641 34524
rect 28184 34456 28212 34496
rect 28629 34493 28641 34496
rect 28675 34493 28687 34527
rect 28629 34487 28687 34493
rect 28718 34484 28724 34536
rect 28776 34524 28782 34536
rect 29840 34524 29868 34555
rect 29914 34552 29920 34604
rect 29972 34552 29978 34604
rect 30834 34552 30840 34604
rect 30892 34552 30898 34604
rect 30926 34552 30932 34604
rect 30984 34601 30990 34604
rect 30984 34595 31012 34601
rect 31000 34561 31012 34595
rect 30984 34555 31012 34561
rect 30984 34552 30990 34555
rect 33042 34552 33048 34604
rect 33100 34592 33106 34604
rect 34701 34595 34759 34601
rect 34701 34592 34713 34595
rect 33100 34564 34713 34592
rect 33100 34552 33106 34564
rect 34701 34561 34713 34564
rect 34747 34561 34759 34595
rect 34701 34555 34759 34561
rect 35621 34595 35679 34601
rect 35621 34561 35633 34595
rect 35667 34592 35679 34595
rect 36078 34592 36084 34604
rect 35667 34564 36084 34592
rect 35667 34561 35679 34564
rect 35621 34555 35679 34561
rect 36078 34552 36084 34564
rect 36136 34552 36142 34604
rect 37458 34552 37464 34604
rect 37516 34592 37522 34604
rect 37553 34595 37611 34601
rect 37553 34592 37565 34595
rect 37516 34564 37565 34592
rect 37516 34552 37522 34564
rect 37553 34561 37565 34564
rect 37599 34561 37611 34595
rect 37553 34555 37611 34561
rect 37826 34552 37832 34604
rect 37884 34552 37890 34604
rect 37918 34552 37924 34604
rect 37976 34592 37982 34604
rect 39577 34595 39635 34601
rect 39577 34592 39589 34595
rect 37976 34564 39589 34592
rect 37976 34552 37982 34564
rect 39577 34561 39589 34564
rect 39623 34592 39635 34595
rect 39758 34592 39764 34604
rect 39623 34564 39764 34592
rect 39623 34561 39635 34564
rect 39577 34555 39635 34561
rect 39758 34552 39764 34564
rect 39816 34552 39822 34604
rect 39850 34552 39856 34604
rect 39908 34552 39914 34604
rect 41230 34552 41236 34604
rect 41288 34592 41294 34604
rect 41782 34592 41788 34604
rect 41288 34564 41788 34592
rect 41288 34552 41294 34564
rect 41782 34552 41788 34564
rect 41840 34552 41846 34604
rect 42150 34552 42156 34604
rect 42208 34592 42214 34604
rect 42521 34595 42579 34601
rect 42521 34592 42533 34595
rect 42208 34564 42533 34592
rect 42208 34552 42214 34564
rect 42521 34561 42533 34564
rect 42567 34561 42579 34595
rect 42521 34555 42579 34561
rect 43349 34595 43407 34601
rect 43349 34561 43361 34595
rect 43395 34561 43407 34595
rect 43349 34555 43407 34561
rect 28776 34496 29868 34524
rect 30101 34527 30159 34533
rect 28776 34484 28782 34496
rect 30101 34493 30113 34527
rect 30147 34524 30159 34527
rect 30466 34524 30472 34536
rect 30147 34496 30472 34524
rect 30147 34493 30159 34496
rect 30101 34487 30159 34493
rect 30466 34484 30472 34496
rect 30524 34484 30530 34536
rect 30561 34527 30619 34533
rect 30561 34493 30573 34527
rect 30607 34524 30619 34527
rect 31113 34527 31171 34533
rect 30607 34496 30696 34524
rect 30607 34493 30619 34496
rect 30561 34487 30619 34493
rect 28000 34428 28212 34456
rect 28445 34459 28503 34465
rect 28445 34425 28457 34459
rect 28491 34456 28503 34459
rect 29178 34456 29184 34468
rect 28491 34428 29184 34456
rect 28491 34425 28503 34428
rect 28445 34419 28503 34425
rect 29178 34416 29184 34428
rect 29236 34416 29242 34468
rect 27893 34391 27951 34397
rect 27893 34388 27905 34391
rect 27356 34360 27905 34388
rect 27893 34357 27905 34360
rect 27939 34357 27951 34391
rect 30668 34388 30696 34496
rect 31113 34493 31125 34527
rect 31159 34524 31171 34527
rect 33318 34524 33324 34536
rect 31159 34496 33324 34524
rect 31159 34493 31171 34496
rect 31113 34487 31171 34493
rect 33318 34484 33324 34496
rect 33376 34484 33382 34536
rect 34238 34484 34244 34536
rect 34296 34524 34302 34536
rect 34425 34527 34483 34533
rect 34425 34524 34437 34527
rect 34296 34496 34437 34524
rect 34296 34484 34302 34496
rect 34425 34493 34437 34496
rect 34471 34493 34483 34527
rect 34425 34487 34483 34493
rect 35802 34484 35808 34536
rect 35860 34484 35866 34536
rect 38105 34527 38163 34533
rect 38105 34493 38117 34527
rect 38151 34493 38163 34527
rect 38105 34487 38163 34493
rect 41509 34527 41567 34533
rect 41509 34493 41521 34527
rect 41555 34493 41567 34527
rect 41800 34524 41828 34552
rect 43364 34524 43392 34555
rect 41800 34496 43392 34524
rect 41509 34487 41567 34493
rect 31754 34388 31760 34400
rect 30668 34360 31760 34388
rect 27893 34351 27951 34357
rect 31754 34348 31760 34360
rect 31812 34348 31818 34400
rect 31846 34348 31852 34400
rect 31904 34388 31910 34400
rect 32306 34388 32312 34400
rect 31904 34360 32312 34388
rect 31904 34348 31910 34360
rect 32306 34348 32312 34360
rect 32364 34388 32370 34400
rect 38120 34388 38148 34487
rect 41524 34456 41552 34487
rect 41524 34428 42012 34456
rect 41984 34400 42012 34428
rect 42150 34416 42156 34468
rect 42208 34416 42214 34468
rect 42245 34459 42303 34465
rect 42245 34425 42257 34459
rect 42291 34456 42303 34459
rect 42702 34456 42708 34468
rect 42291 34428 42708 34456
rect 42291 34425 42303 34428
rect 42245 34419 42303 34425
rect 42702 34416 42708 34428
rect 42760 34416 42766 34468
rect 38378 34388 38384 34400
rect 32364 34360 38384 34388
rect 32364 34348 32370 34360
rect 38378 34348 38384 34360
rect 38436 34348 38442 34400
rect 41601 34391 41659 34397
rect 41601 34357 41613 34391
rect 41647 34388 41659 34391
rect 41690 34388 41696 34400
rect 41647 34360 41696 34388
rect 41647 34357 41659 34360
rect 41601 34351 41659 34357
rect 41690 34348 41696 34360
rect 41748 34348 41754 34400
rect 41966 34348 41972 34400
rect 42024 34388 42030 34400
rect 42613 34391 42671 34397
rect 42613 34388 42625 34391
rect 42024 34360 42625 34388
rect 42024 34348 42030 34360
rect 42613 34357 42625 34360
rect 42659 34388 42671 34391
rect 43441 34391 43499 34397
rect 43441 34388 43453 34391
rect 42659 34360 43453 34388
rect 42659 34357 42671 34360
rect 42613 34351 42671 34357
rect 43441 34357 43453 34360
rect 43487 34357 43499 34391
rect 43441 34351 43499 34357
rect 43806 34348 43812 34400
rect 43864 34348 43870 34400
rect 1104 34298 47104 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 47104 34298
rect 1104 34224 47104 34246
rect 9950 34144 9956 34196
rect 10008 34184 10014 34196
rect 10318 34184 10324 34196
rect 10008 34156 10324 34184
rect 10008 34144 10014 34156
rect 10318 34144 10324 34156
rect 10376 34144 10382 34196
rect 10502 34144 10508 34196
rect 10560 34184 10566 34196
rect 10870 34184 10876 34196
rect 10560 34156 10876 34184
rect 10560 34144 10566 34156
rect 10870 34144 10876 34156
rect 10928 34144 10934 34196
rect 13354 34144 13360 34196
rect 13412 34144 13418 34196
rect 16298 34144 16304 34196
rect 16356 34144 16362 34196
rect 18322 34144 18328 34196
rect 18380 34144 18386 34196
rect 24118 34144 24124 34196
rect 24176 34184 24182 34196
rect 34514 34184 34520 34196
rect 24176 34156 34520 34184
rect 24176 34144 24182 34156
rect 34514 34144 34520 34156
rect 34572 34144 34578 34196
rect 34606 34144 34612 34196
rect 34664 34184 34670 34196
rect 34664 34156 36032 34184
rect 34664 34144 34670 34156
rect 11238 34076 11244 34128
rect 11296 34116 11302 34128
rect 20993 34119 21051 34125
rect 20993 34116 21005 34119
rect 11296 34088 21005 34116
rect 11296 34076 11302 34088
rect 20993 34085 21005 34088
rect 21039 34116 21051 34119
rect 30926 34116 30932 34128
rect 21039 34088 30932 34116
rect 21039 34085 21051 34088
rect 20993 34079 21051 34085
rect 30926 34076 30932 34088
rect 30984 34076 30990 34128
rect 5077 34051 5135 34057
rect 5077 34017 5089 34051
rect 5123 34048 5135 34051
rect 5442 34048 5448 34060
rect 5123 34020 5448 34048
rect 5123 34017 5135 34020
rect 5077 34011 5135 34017
rect 5442 34008 5448 34020
rect 5500 34008 5506 34060
rect 11422 34008 11428 34060
rect 11480 34048 11486 34060
rect 15286 34048 15292 34060
rect 11480 34020 15292 34048
rect 11480 34008 11486 34020
rect 15286 34008 15292 34020
rect 15344 34008 15350 34060
rect 16758 34008 16764 34060
rect 16816 34048 16822 34060
rect 16853 34051 16911 34057
rect 16853 34048 16865 34051
rect 16816 34020 16865 34048
rect 16816 34008 16822 34020
rect 16853 34017 16865 34020
rect 16899 34048 16911 34051
rect 19702 34048 19708 34060
rect 16899 34020 19708 34048
rect 16899 34017 16911 34020
rect 16853 34011 16911 34017
rect 19702 34008 19708 34020
rect 19760 34008 19766 34060
rect 20070 34008 20076 34060
rect 20128 34048 20134 34060
rect 21174 34048 21180 34060
rect 20128 34020 21180 34048
rect 20128 34008 20134 34020
rect 21174 34008 21180 34020
rect 21232 34008 21238 34060
rect 23566 34008 23572 34060
rect 23624 34048 23630 34060
rect 30190 34048 30196 34060
rect 23624 34020 30196 34048
rect 23624 34008 23630 34020
rect 30190 34008 30196 34020
rect 30248 34048 30254 34060
rect 31018 34048 31024 34060
rect 30248 34020 31024 34048
rect 30248 34008 30254 34020
rect 31018 34008 31024 34020
rect 31076 34008 31082 34060
rect 34606 34048 34612 34060
rect 34256 34020 34612 34048
rect 3050 33940 3056 33992
rect 3108 33980 3114 33992
rect 3602 33980 3608 33992
rect 3108 33952 3608 33980
rect 3108 33940 3114 33952
rect 3602 33940 3608 33952
rect 3660 33980 3666 33992
rect 4893 33983 4951 33989
rect 4893 33980 4905 33983
rect 3660 33952 4905 33980
rect 3660 33940 3666 33952
rect 4893 33949 4905 33952
rect 4939 33949 4951 33983
rect 4893 33943 4951 33949
rect 13541 33983 13599 33989
rect 13541 33949 13553 33983
rect 13587 33980 13599 33983
rect 14550 33980 14556 33992
rect 13587 33952 14556 33980
rect 13587 33949 13599 33952
rect 13541 33943 13599 33949
rect 14550 33940 14556 33952
rect 14608 33940 14614 33992
rect 16666 33940 16672 33992
rect 16724 33940 16730 33992
rect 18506 33940 18512 33992
rect 18564 33940 18570 33992
rect 21266 33940 21272 33992
rect 21324 33940 21330 33992
rect 21910 33940 21916 33992
rect 21968 33940 21974 33992
rect 31662 33940 31668 33992
rect 31720 33940 31726 33992
rect 31757 33983 31815 33989
rect 31757 33949 31769 33983
rect 31803 33980 31815 33983
rect 31846 33980 31852 33992
rect 31803 33952 31852 33980
rect 31803 33949 31815 33952
rect 31757 33943 31815 33949
rect 31846 33940 31852 33952
rect 31904 33940 31910 33992
rect 34256 33989 34284 34020
rect 34606 34008 34612 34020
rect 34664 34008 34670 34060
rect 36004 34048 36032 34156
rect 36078 34144 36084 34196
rect 36136 34144 36142 34196
rect 41782 34076 41788 34128
rect 41840 34116 41846 34128
rect 42242 34116 42248 34128
rect 41840 34088 42248 34116
rect 41840 34076 41846 34088
rect 42242 34076 42248 34088
rect 42300 34076 42306 34128
rect 45005 34119 45063 34125
rect 45005 34116 45017 34119
rect 42352 34088 45017 34116
rect 36004 34020 37688 34048
rect 34241 33983 34299 33989
rect 34241 33949 34253 33983
rect 34287 33949 34299 33983
rect 34241 33943 34299 33949
rect 34514 33940 34520 33992
rect 34572 33940 34578 33992
rect 34701 33983 34759 33989
rect 34701 33949 34713 33983
rect 34747 33980 34759 33983
rect 35986 33980 35992 33992
rect 34747 33952 35992 33980
rect 34747 33949 34759 33952
rect 34701 33943 34759 33949
rect 35986 33940 35992 33952
rect 36044 33940 36050 33992
rect 37369 33983 37427 33989
rect 37369 33949 37381 33983
rect 37415 33980 37427 33983
rect 37458 33980 37464 33992
rect 37415 33952 37464 33980
rect 37415 33949 37427 33952
rect 37369 33943 37427 33949
rect 37458 33940 37464 33952
rect 37516 33940 37522 33992
rect 37660 33989 37688 34020
rect 42058 34008 42064 34060
rect 42116 34048 42122 34060
rect 42352 34048 42380 34088
rect 45005 34085 45017 34088
rect 45051 34085 45063 34119
rect 45005 34079 45063 34085
rect 43806 34048 43812 34060
rect 42116 34020 42380 34048
rect 43180 34020 43812 34048
rect 42116 34008 42122 34020
rect 37645 33983 37703 33989
rect 37645 33949 37657 33983
rect 37691 33949 37703 33983
rect 37645 33943 37703 33949
rect 37829 33983 37887 33989
rect 37829 33949 37841 33983
rect 37875 33980 37887 33983
rect 38654 33980 38660 33992
rect 37875 33952 38660 33980
rect 37875 33949 37887 33952
rect 37829 33943 37887 33949
rect 38654 33940 38660 33952
rect 38712 33940 38718 33992
rect 40957 33983 41015 33989
rect 40957 33949 40969 33983
rect 41003 33949 41015 33983
rect 40957 33943 41015 33949
rect 4614 33872 4620 33924
rect 4672 33912 4678 33924
rect 4801 33915 4859 33921
rect 4801 33912 4813 33915
rect 4672 33884 4813 33912
rect 4672 33872 4678 33884
rect 4801 33881 4813 33884
rect 4847 33912 4859 33915
rect 5350 33912 5356 33924
rect 4847 33884 5356 33912
rect 4847 33881 4859 33884
rect 4801 33875 4859 33881
rect 5350 33872 5356 33884
rect 5408 33872 5414 33924
rect 15102 33872 15108 33924
rect 15160 33912 15166 33924
rect 18322 33912 18328 33924
rect 15160 33884 18328 33912
rect 15160 33872 15166 33884
rect 18322 33872 18328 33884
rect 18380 33872 18386 33924
rect 20346 33872 20352 33924
rect 20404 33912 20410 33924
rect 20809 33915 20867 33921
rect 20809 33912 20821 33915
rect 20404 33884 20821 33912
rect 20404 33872 20410 33884
rect 20809 33881 20821 33884
rect 20855 33912 20867 33915
rect 20990 33912 20996 33924
rect 20855 33884 20996 33912
rect 20855 33881 20867 33884
rect 20809 33875 20867 33881
rect 20990 33872 20996 33884
rect 21048 33872 21054 33924
rect 21542 33872 21548 33924
rect 21600 33872 21606 33924
rect 32002 33915 32060 33921
rect 32002 33912 32014 33915
rect 31726 33884 32014 33912
rect 3878 33804 3884 33856
rect 3936 33844 3942 33856
rect 4433 33847 4491 33853
rect 4433 33844 4445 33847
rect 3936 33816 4445 33844
rect 3936 33804 3942 33816
rect 4433 33813 4445 33816
rect 4479 33813 4491 33847
rect 4433 33807 4491 33813
rect 15010 33804 15016 33856
rect 15068 33844 15074 33856
rect 16761 33847 16819 33853
rect 16761 33844 16773 33847
rect 15068 33816 16773 33844
rect 15068 33804 15074 33816
rect 16761 33813 16773 33816
rect 16807 33844 16819 33847
rect 16942 33844 16948 33856
rect 16807 33816 16948 33844
rect 16807 33813 16819 33816
rect 16761 33807 16819 33813
rect 16942 33804 16948 33816
rect 17000 33804 17006 33856
rect 22097 33847 22155 33853
rect 22097 33813 22109 33847
rect 22143 33844 22155 33847
rect 22738 33844 22744 33856
rect 22143 33816 22744 33844
rect 22143 33813 22155 33816
rect 22097 33807 22155 33813
rect 22738 33804 22744 33816
rect 22796 33804 22802 33856
rect 31481 33847 31539 33853
rect 31481 33813 31493 33847
rect 31527 33844 31539 33847
rect 31726 33844 31754 33884
rect 32002 33881 32014 33884
rect 32048 33881 32060 33915
rect 32002 33875 32060 33881
rect 34057 33915 34115 33921
rect 34057 33881 34069 33915
rect 34103 33912 34115 33915
rect 34946 33915 35004 33921
rect 34946 33912 34958 33915
rect 34103 33884 34958 33912
rect 34103 33881 34115 33884
rect 34057 33875 34115 33881
rect 34946 33881 34958 33884
rect 34992 33881 35004 33915
rect 37734 33912 37740 33924
rect 34946 33875 35004 33881
rect 35820 33884 37740 33912
rect 35820 33856 35848 33884
rect 37734 33872 37740 33884
rect 37792 33872 37798 33924
rect 40972 33912 41000 33943
rect 41046 33940 41052 33992
rect 41104 33940 41110 33992
rect 43180 33989 43208 34020
rect 43806 34008 43812 34020
rect 43864 34008 43870 34060
rect 44174 34008 44180 34060
rect 44232 34048 44238 34060
rect 45186 34048 45192 34060
rect 44232 34020 45192 34048
rect 44232 34008 44238 34020
rect 45186 34008 45192 34020
rect 45244 34048 45250 34060
rect 45738 34048 45744 34060
rect 45244 34020 45744 34048
rect 45244 34008 45250 34020
rect 45738 34008 45744 34020
rect 45796 34008 45802 34060
rect 43165 33983 43223 33989
rect 43165 33949 43177 33983
rect 43211 33949 43223 33983
rect 43165 33943 43223 33949
rect 43349 33983 43407 33989
rect 43349 33949 43361 33983
rect 43395 33980 43407 33983
rect 44450 33980 44456 33992
rect 43395 33952 44456 33980
rect 43395 33949 43407 33952
rect 43349 33943 43407 33949
rect 41138 33912 41144 33924
rect 40972 33884 41144 33912
rect 41138 33872 41144 33884
rect 41196 33872 41202 33924
rect 41598 33872 41604 33924
rect 41656 33912 41662 33924
rect 41966 33912 41972 33924
rect 41656 33884 41972 33912
rect 41656 33872 41662 33884
rect 41966 33872 41972 33884
rect 42024 33872 42030 33924
rect 43364 33912 43392 33943
rect 44450 33940 44456 33952
rect 44508 33940 44514 33992
rect 45281 33983 45339 33989
rect 45281 33949 45293 33983
rect 45327 33980 45339 33983
rect 45370 33980 45376 33992
rect 45327 33952 45376 33980
rect 45327 33949 45339 33952
rect 45281 33943 45339 33949
rect 45370 33940 45376 33952
rect 45428 33940 45434 33992
rect 42076 33884 43392 33912
rect 31527 33816 31754 33844
rect 31527 33813 31539 33816
rect 31481 33807 31539 33813
rect 32490 33804 32496 33856
rect 32548 33844 32554 33856
rect 33137 33847 33195 33853
rect 33137 33844 33149 33847
rect 32548 33816 33149 33844
rect 32548 33804 32554 33816
rect 33137 33813 33149 33816
rect 33183 33813 33195 33847
rect 33137 33807 33195 33813
rect 34425 33847 34483 33853
rect 34425 33813 34437 33847
rect 34471 33844 34483 33847
rect 35802 33844 35808 33856
rect 34471 33816 35808 33844
rect 34471 33813 34483 33816
rect 34425 33807 34483 33813
rect 35802 33804 35808 33816
rect 35860 33804 35866 33856
rect 37182 33804 37188 33856
rect 37240 33804 37246 33856
rect 40310 33804 40316 33856
rect 40368 33844 40374 33856
rect 41233 33847 41291 33853
rect 41233 33844 41245 33847
rect 40368 33816 41245 33844
rect 40368 33804 40374 33816
rect 41233 33813 41245 33816
rect 41279 33813 41291 33847
rect 41233 33807 41291 33813
rect 41690 33804 41696 33856
rect 41748 33844 41754 33856
rect 42076 33844 42104 33884
rect 45002 33872 45008 33924
rect 45060 33912 45066 33924
rect 46014 33912 46020 33924
rect 45060 33884 46020 33912
rect 45060 33872 45066 33884
rect 46014 33872 46020 33884
rect 46072 33872 46078 33924
rect 41748 33816 42104 33844
rect 41748 33804 41754 33816
rect 42426 33804 42432 33856
rect 42484 33804 42490 33856
rect 42518 33804 42524 33856
rect 42576 33844 42582 33856
rect 43257 33847 43315 33853
rect 43257 33844 43269 33847
rect 42576 33816 43269 33844
rect 42576 33804 42582 33816
rect 43257 33813 43269 33816
rect 43303 33813 43315 33847
rect 43257 33807 43315 33813
rect 45189 33847 45247 33853
rect 45189 33813 45201 33847
rect 45235 33844 45247 33847
rect 45370 33844 45376 33856
rect 45235 33816 45376 33844
rect 45235 33813 45247 33816
rect 45189 33807 45247 33813
rect 45370 33804 45376 33816
rect 45428 33804 45434 33856
rect 1104 33754 47104 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 47104 33754
rect 1104 33680 47104 33702
rect 2593 33643 2651 33649
rect 2593 33609 2605 33643
rect 2639 33609 2651 33643
rect 2593 33603 2651 33609
rect 2409 33507 2467 33513
rect 2409 33473 2421 33507
rect 2455 33504 2467 33507
rect 2608 33504 2636 33603
rect 3050 33600 3056 33652
rect 3108 33600 3114 33652
rect 3697 33643 3755 33649
rect 3697 33609 3709 33643
rect 3743 33609 3755 33643
rect 3697 33603 3755 33609
rect 3712 33572 3740 33603
rect 5350 33600 5356 33652
rect 5408 33600 5414 33652
rect 13814 33600 13820 33652
rect 13872 33640 13878 33652
rect 21910 33640 21916 33652
rect 13872 33612 21916 33640
rect 13872 33600 13878 33612
rect 21910 33600 21916 33612
rect 21968 33600 21974 33652
rect 23658 33600 23664 33652
rect 23716 33640 23722 33652
rect 24305 33643 24363 33649
rect 23716 33612 24256 33640
rect 23716 33600 23722 33612
rect 4218 33575 4276 33581
rect 4218 33572 4230 33575
rect 3712 33544 4230 33572
rect 4218 33541 4230 33544
rect 4264 33541 4276 33575
rect 4218 33535 4276 33541
rect 13081 33575 13139 33581
rect 13081 33541 13093 33575
rect 13127 33572 13139 33575
rect 13170 33572 13176 33584
rect 13127 33544 13176 33572
rect 13127 33541 13139 33544
rect 13081 33535 13139 33541
rect 13170 33532 13176 33544
rect 13228 33572 13234 33584
rect 15010 33572 15016 33584
rect 13228 33544 15016 33572
rect 13228 33532 13234 33544
rect 15010 33532 15016 33544
rect 15068 33532 15074 33584
rect 18598 33532 18604 33584
rect 18656 33572 18662 33584
rect 18969 33575 19027 33581
rect 18969 33572 18981 33575
rect 18656 33544 18981 33572
rect 18656 33532 18662 33544
rect 18969 33541 18981 33544
rect 19015 33541 19027 33575
rect 18969 33535 19027 33541
rect 20990 33532 20996 33584
rect 21048 33572 21054 33584
rect 23474 33572 23480 33584
rect 21048 33544 23480 33572
rect 21048 33532 21054 33544
rect 23474 33532 23480 33544
rect 23532 33572 23538 33584
rect 23532 33544 24164 33572
rect 23532 33532 23538 33544
rect 2455 33476 2636 33504
rect 2455 33473 2467 33476
rect 2409 33467 2467 33473
rect 2958 33464 2964 33516
rect 3016 33464 3022 33516
rect 3878 33464 3884 33516
rect 3936 33464 3942 33516
rect 3970 33464 3976 33516
rect 4028 33464 4034 33516
rect 9398 33464 9404 33516
rect 9456 33464 9462 33516
rect 12437 33507 12495 33513
rect 12437 33473 12449 33507
rect 12483 33504 12495 33507
rect 12483 33476 12664 33504
rect 12483 33473 12495 33476
rect 12437 33467 12495 33473
rect 3142 33396 3148 33448
rect 3200 33396 3206 33448
rect 9674 33396 9680 33448
rect 9732 33396 9738 33448
rect 10226 33328 10232 33380
rect 10284 33368 10290 33380
rect 12636 33377 12664 33476
rect 12986 33464 12992 33516
rect 13044 33464 13050 33516
rect 18785 33507 18843 33513
rect 18785 33473 18797 33507
rect 18831 33473 18843 33507
rect 18785 33467 18843 33473
rect 13078 33396 13084 33448
rect 13136 33436 13142 33448
rect 13173 33439 13231 33445
rect 13173 33436 13185 33439
rect 13136 33408 13185 33436
rect 13136 33396 13142 33408
rect 13173 33405 13185 33408
rect 13219 33436 13231 33439
rect 16574 33436 16580 33448
rect 13219 33408 16580 33436
rect 13219 33405 13231 33408
rect 13173 33399 13231 33405
rect 16574 33396 16580 33408
rect 16632 33396 16638 33448
rect 18800 33436 18828 33467
rect 22186 33464 22192 33516
rect 22244 33504 22250 33516
rect 22281 33507 22339 33513
rect 22281 33504 22293 33507
rect 22244 33476 22293 33504
rect 22244 33464 22250 33476
rect 22281 33473 22293 33476
rect 22327 33473 22339 33507
rect 22281 33467 22339 33473
rect 22548 33507 22606 33513
rect 22548 33473 22560 33507
rect 22594 33504 22606 33507
rect 23106 33504 23112 33516
rect 22594 33476 23112 33504
rect 22594 33473 22606 33476
rect 22548 33467 22606 33473
rect 23106 33464 23112 33476
rect 23164 33464 23170 33516
rect 24136 33513 24164 33544
rect 24121 33507 24179 33513
rect 24121 33473 24133 33507
rect 24167 33473 24179 33507
rect 24228 33504 24256 33612
rect 24305 33609 24317 33643
rect 24351 33640 24363 33643
rect 27706 33640 27712 33652
rect 24351 33612 27712 33640
rect 24351 33609 24363 33612
rect 24305 33603 24363 33609
rect 27706 33600 27712 33612
rect 27764 33600 27770 33652
rect 31662 33600 31668 33652
rect 31720 33640 31726 33652
rect 32125 33643 32183 33649
rect 32125 33640 32137 33643
rect 31720 33612 32137 33640
rect 31720 33600 31726 33612
rect 32125 33609 32137 33612
rect 32171 33609 32183 33643
rect 32490 33640 32496 33652
rect 32125 33603 32183 33609
rect 32324 33612 32496 33640
rect 29270 33572 29276 33584
rect 25424 33544 29276 33572
rect 25424 33513 25452 33544
rect 29270 33532 29276 33544
rect 29328 33532 29334 33584
rect 30466 33532 30472 33584
rect 30524 33572 30530 33584
rect 32324 33572 32352 33612
rect 32490 33600 32496 33612
rect 32548 33600 32554 33652
rect 41046 33600 41052 33652
rect 41104 33640 41110 33652
rect 41601 33643 41659 33649
rect 41601 33640 41613 33643
rect 41104 33612 41613 33640
rect 41104 33600 41110 33612
rect 41601 33609 41613 33612
rect 41647 33609 41659 33643
rect 41601 33603 41659 33609
rect 41785 33643 41843 33649
rect 41785 33609 41797 33643
rect 41831 33640 41843 33643
rect 41966 33640 41972 33652
rect 41831 33612 41972 33640
rect 41831 33609 41843 33612
rect 41785 33603 41843 33609
rect 41966 33600 41972 33612
rect 42024 33640 42030 33652
rect 46201 33643 46259 33649
rect 46201 33640 46213 33643
rect 42024 33612 43116 33640
rect 42024 33600 42030 33612
rect 30524 33544 32352 33572
rect 32416 33544 34744 33572
rect 30524 33532 30530 33544
rect 24489 33507 24547 33513
rect 24489 33504 24501 33507
rect 24228 33476 24501 33504
rect 24121 33467 24179 33473
rect 24489 33473 24501 33476
rect 24535 33504 24547 33507
rect 25409 33507 25467 33513
rect 25409 33504 25421 33507
rect 24535 33476 25421 33504
rect 24535 33473 24547 33476
rect 24489 33467 24547 33473
rect 25409 33473 25421 33476
rect 25455 33473 25467 33507
rect 25409 33467 25467 33473
rect 25676 33507 25734 33513
rect 25676 33473 25688 33507
rect 25722 33504 25734 33507
rect 26050 33504 26056 33516
rect 25722 33476 26056 33504
rect 25722 33473 25734 33476
rect 25676 33467 25734 33473
rect 26050 33464 26056 33476
rect 26108 33464 26114 33516
rect 27614 33464 27620 33516
rect 27672 33504 27678 33516
rect 32416 33504 32444 33544
rect 34716 33513 34744 33544
rect 37182 33532 37188 33584
rect 37240 33572 37246 33584
rect 37798 33575 37856 33581
rect 37798 33572 37810 33575
rect 37240 33544 37810 33572
rect 37240 33532 37246 33544
rect 37798 33541 37810 33544
rect 37844 33541 37856 33575
rect 37798 33535 37856 33541
rect 40788 33544 41736 33572
rect 27672 33476 32444 33504
rect 34701 33507 34759 33513
rect 27672 33464 27678 33476
rect 34701 33473 34713 33507
rect 34747 33473 34759 33507
rect 34701 33467 34759 33473
rect 35986 33464 35992 33516
rect 36044 33504 36050 33516
rect 37553 33507 37611 33513
rect 37553 33504 37565 33507
rect 36044 33476 37565 33504
rect 36044 33464 36050 33476
rect 37553 33473 37565 33476
rect 37599 33473 37611 33507
rect 37553 33467 37611 33473
rect 39298 33464 39304 33516
rect 39356 33464 39362 33516
rect 39393 33507 39451 33513
rect 39393 33473 39405 33507
rect 39439 33504 39451 33507
rect 39439 33476 40172 33504
rect 39439 33473 39451 33476
rect 39393 33467 39451 33473
rect 18800 33408 19012 33436
rect 12621 33371 12679 33377
rect 10284 33340 12434 33368
rect 10284 33328 10290 33340
rect 2038 33260 2044 33312
rect 2096 33300 2102 33312
rect 2225 33303 2283 33309
rect 2225 33300 2237 33303
rect 2096 33272 2237 33300
rect 2096 33260 2102 33272
rect 2225 33269 2237 33272
rect 2271 33269 2283 33303
rect 2225 33263 2283 33269
rect 12158 33260 12164 33312
rect 12216 33300 12222 33312
rect 12253 33303 12311 33309
rect 12253 33300 12265 33303
rect 12216 33272 12265 33300
rect 12216 33260 12222 33272
rect 12253 33269 12265 33272
rect 12299 33269 12311 33303
rect 12406 33300 12434 33340
rect 12621 33337 12633 33371
rect 12667 33337 12679 33371
rect 12621 33331 12679 33337
rect 18984 33312 19012 33408
rect 24578 33396 24584 33448
rect 24636 33436 24642 33448
rect 24765 33439 24823 33445
rect 24765 33436 24777 33439
rect 24636 33408 24777 33436
rect 24636 33396 24642 33408
rect 24765 33405 24777 33408
rect 24811 33405 24823 33439
rect 24765 33399 24823 33405
rect 32030 33396 32036 33448
rect 32088 33436 32094 33448
rect 32585 33439 32643 33445
rect 32585 33436 32597 33439
rect 32088 33408 32597 33436
rect 32088 33396 32094 33408
rect 32585 33405 32597 33408
rect 32631 33405 32643 33439
rect 32585 33399 32643 33405
rect 32769 33439 32827 33445
rect 32769 33405 32781 33439
rect 32815 33436 32827 33439
rect 33502 33436 33508 33448
rect 32815 33408 33508 33436
rect 32815 33405 32827 33408
rect 32769 33399 32827 33405
rect 31846 33328 31852 33380
rect 31904 33368 31910 33380
rect 32784 33368 32812 33399
rect 33502 33396 33508 33408
rect 33560 33396 33566 33448
rect 34422 33396 34428 33448
rect 34480 33396 34486 33448
rect 36170 33396 36176 33448
rect 36228 33436 36234 33448
rect 37182 33436 37188 33448
rect 36228 33408 37188 33436
rect 36228 33396 36234 33408
rect 37182 33396 37188 33408
rect 37240 33396 37246 33448
rect 39577 33439 39635 33445
rect 39577 33405 39589 33439
rect 39623 33405 39635 33439
rect 39577 33399 39635 33405
rect 31904 33340 32812 33368
rect 39117 33371 39175 33377
rect 31904 33328 31910 33340
rect 39117 33337 39129 33371
rect 39163 33368 39175 33371
rect 39592 33368 39620 33399
rect 40144 33377 40172 33476
rect 40310 33464 40316 33516
rect 40368 33464 40374 33516
rect 40788 33513 40816 33544
rect 41708 33516 41736 33544
rect 42426 33532 42432 33584
rect 42484 33572 42490 33584
rect 42484 33544 42840 33572
rect 42484 33532 42490 33544
rect 40773 33507 40831 33513
rect 40773 33473 40785 33507
rect 40819 33473 40831 33507
rect 40773 33467 40831 33473
rect 40865 33507 40923 33513
rect 40865 33473 40877 33507
rect 40911 33473 40923 33507
rect 40865 33467 40923 33473
rect 40880 33436 40908 33467
rect 41322 33464 41328 33516
rect 41380 33464 41386 33516
rect 41690 33464 41696 33516
rect 41748 33464 41754 33516
rect 42058 33464 42064 33516
rect 42116 33464 42122 33516
rect 42153 33507 42211 33513
rect 42153 33473 42165 33507
rect 42199 33504 42211 33507
rect 42518 33504 42524 33516
rect 42199 33476 42524 33504
rect 42199 33473 42211 33476
rect 42153 33467 42211 33473
rect 42518 33464 42524 33476
rect 42576 33464 42582 33516
rect 42702 33464 42708 33516
rect 42760 33464 42766 33516
rect 42812 33513 42840 33544
rect 43088 33513 43116 33612
rect 45526 33612 46213 33640
rect 43806 33532 43812 33584
rect 43864 33572 43870 33584
rect 43864 33544 45140 33572
rect 43864 33532 43870 33544
rect 42797 33507 42855 33513
rect 42797 33473 42809 33507
rect 42843 33473 42855 33507
rect 42797 33467 42855 33473
rect 42889 33507 42947 33513
rect 42889 33473 42901 33507
rect 42935 33473 42947 33507
rect 42889 33467 42947 33473
rect 43073 33507 43131 33513
rect 43073 33473 43085 33507
rect 43119 33473 43131 33507
rect 43073 33467 43131 33473
rect 40880 33408 41644 33436
rect 39163 33340 39620 33368
rect 40129 33371 40187 33377
rect 39163 33337 39175 33340
rect 39117 33331 39175 33337
rect 40129 33337 40141 33371
rect 40175 33337 40187 33371
rect 41616 33368 41644 33408
rect 41874 33396 41880 33448
rect 41932 33436 41938 33448
rect 42904 33436 42932 33467
rect 43898 33464 43904 33516
rect 43956 33464 43962 33516
rect 44192 33513 44220 33544
rect 44177 33507 44235 33513
rect 44177 33473 44189 33507
rect 44223 33473 44235 33507
rect 44177 33467 44235 33473
rect 44450 33464 44456 33516
rect 44508 33464 44514 33516
rect 44542 33464 44548 33516
rect 44600 33464 44606 33516
rect 44910 33464 44916 33516
rect 44968 33464 44974 33516
rect 45002 33464 45008 33516
rect 45060 33464 45066 33516
rect 45112 33513 45140 33544
rect 45370 33532 45376 33584
rect 45428 33572 45434 33584
rect 45526 33572 45554 33612
rect 46201 33609 46213 33612
rect 46247 33609 46259 33643
rect 46201 33603 46259 33609
rect 45428 33544 45554 33572
rect 45428 33532 45434 33544
rect 45098 33507 45156 33513
rect 45098 33473 45110 33507
rect 45144 33473 45156 33507
rect 45098 33467 45156 33473
rect 45281 33507 45339 33513
rect 45281 33473 45293 33507
rect 45327 33473 45339 33507
rect 45462 33504 45468 33516
rect 45520 33513 45526 33516
rect 45428 33476 45468 33504
rect 45281 33467 45339 33473
rect 41932 33408 42932 33436
rect 44468 33436 44496 33464
rect 45296 33436 45324 33467
rect 45462 33464 45468 33476
rect 45520 33467 45528 33513
rect 45520 33464 45526 33467
rect 45738 33464 45744 33516
rect 45796 33464 45802 33516
rect 46477 33507 46535 33513
rect 46477 33473 46489 33507
rect 46523 33473 46535 33507
rect 46477 33467 46535 33473
rect 46293 33439 46351 33445
rect 46293 33436 46305 33439
rect 44468 33408 45324 33436
rect 45526 33408 46305 33436
rect 41932 33396 41938 33408
rect 43993 33371 44051 33377
rect 43993 33368 44005 33371
rect 41616 33340 44005 33368
rect 40129 33331 40187 33337
rect 43993 33337 44005 33340
rect 44039 33368 44051 33371
rect 45526 33368 45554 33408
rect 46293 33405 46305 33408
rect 46339 33405 46351 33439
rect 46293 33399 46351 33405
rect 44039 33340 45554 33368
rect 45649 33371 45707 33377
rect 44039 33337 44051 33340
rect 43993 33331 44051 33337
rect 45649 33337 45661 33371
rect 45695 33368 45707 33371
rect 46492 33368 46520 33467
rect 45695 33340 46520 33368
rect 45695 33337 45707 33340
rect 45649 33331 45707 33337
rect 14826 33300 14832 33312
rect 12406 33272 14832 33300
rect 12253 33263 12311 33269
rect 14826 33260 14832 33272
rect 14884 33260 14890 33312
rect 16298 33260 16304 33312
rect 16356 33300 16362 33312
rect 18598 33300 18604 33312
rect 16356 33272 18604 33300
rect 16356 33260 16362 33272
rect 18598 33260 18604 33272
rect 18656 33260 18662 33312
rect 18966 33260 18972 33312
rect 19024 33300 19030 33312
rect 19061 33303 19119 33309
rect 19061 33300 19073 33303
rect 19024 33272 19073 33300
rect 19024 33260 19030 33272
rect 19061 33269 19073 33272
rect 19107 33269 19119 33303
rect 19061 33263 19119 33269
rect 23661 33303 23719 33309
rect 23661 33269 23673 33303
rect 23707 33300 23719 33303
rect 24394 33300 24400 33312
rect 23707 33272 24400 33300
rect 23707 33269 23719 33272
rect 23661 33263 23719 33269
rect 24394 33260 24400 33272
rect 24452 33260 24458 33312
rect 26510 33260 26516 33312
rect 26568 33300 26574 33312
rect 26789 33303 26847 33309
rect 26789 33300 26801 33303
rect 26568 33272 26801 33300
rect 26568 33260 26574 33272
rect 26789 33269 26801 33272
rect 26835 33269 26847 33303
rect 26789 33263 26847 33269
rect 35437 33303 35495 33309
rect 35437 33269 35449 33303
rect 35483 33300 35495 33303
rect 36998 33300 37004 33312
rect 35483 33272 37004 33300
rect 35483 33269 35495 33272
rect 35437 33263 35495 33269
rect 36998 33260 37004 33272
rect 37056 33260 37062 33312
rect 38933 33303 38991 33309
rect 38933 33269 38945 33303
rect 38979 33300 38991 33303
rect 39206 33300 39212 33312
rect 38979 33272 39212 33300
rect 38979 33269 38991 33272
rect 38933 33263 38991 33269
rect 39206 33260 39212 33272
rect 39264 33260 39270 33312
rect 40034 33260 40040 33312
rect 40092 33260 40098 33312
rect 41138 33260 41144 33312
rect 41196 33260 41202 33312
rect 41230 33260 41236 33312
rect 41288 33260 41294 33312
rect 41690 33260 41696 33312
rect 41748 33300 41754 33312
rect 42334 33300 42340 33312
rect 41748 33272 42340 33300
rect 41748 33260 41754 33272
rect 42334 33260 42340 33272
rect 42392 33260 42398 33312
rect 42429 33303 42487 33309
rect 42429 33269 42441 33303
rect 42475 33300 42487 33303
rect 43438 33300 43444 33312
rect 42475 33272 43444 33300
rect 42475 33269 42487 33272
rect 42429 33263 42487 33269
rect 43438 33260 43444 33272
rect 43496 33260 43502 33312
rect 44726 33260 44732 33312
rect 44784 33300 44790 33312
rect 45833 33303 45891 33309
rect 45833 33300 45845 33303
rect 44784 33272 45845 33300
rect 44784 33260 44790 33272
rect 45833 33269 45845 33272
rect 45879 33269 45891 33303
rect 45833 33263 45891 33269
rect 46106 33260 46112 33312
rect 46164 33300 46170 33312
rect 46661 33303 46719 33309
rect 46661 33300 46673 33303
rect 46164 33272 46673 33300
rect 46164 33260 46170 33272
rect 46661 33269 46673 33272
rect 46707 33269 46719 33303
rect 46661 33263 46719 33269
rect 1104 33210 47104 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 47104 33210
rect 1104 33136 47104 33158
rect 2958 33056 2964 33108
rect 3016 33096 3022 33108
rect 3145 33099 3203 33105
rect 3145 33096 3157 33099
rect 3016 33068 3157 33096
rect 3016 33056 3022 33068
rect 3145 33065 3157 33068
rect 3191 33096 3203 33099
rect 4062 33096 4068 33108
rect 3191 33068 4068 33096
rect 3191 33065 3203 33068
rect 3145 33059 3203 33065
rect 4062 33056 4068 33068
rect 4120 33096 4126 33108
rect 4120 33068 4844 33096
rect 4120 33056 4126 33068
rect 4706 32988 4712 33040
rect 4764 32988 4770 33040
rect 4065 32963 4123 32969
rect 4065 32929 4077 32963
rect 4111 32960 4123 32963
rect 4154 32960 4160 32972
rect 4111 32932 4160 32960
rect 4111 32929 4123 32932
rect 4065 32923 4123 32929
rect 4154 32920 4160 32932
rect 4212 32960 4218 32972
rect 4614 32960 4620 32972
rect 4212 32932 4620 32960
rect 4212 32920 4218 32932
rect 4614 32920 4620 32932
rect 4672 32920 4678 32972
rect 4816 32960 4844 33068
rect 6546 33056 6552 33108
rect 6604 33096 6610 33108
rect 9306 33096 9312 33108
rect 6604 33068 9312 33096
rect 6604 33056 6610 33068
rect 9306 33056 9312 33068
rect 9364 33096 9370 33108
rect 9674 33096 9680 33108
rect 9364 33068 9680 33096
rect 9364 33056 9370 33068
rect 9674 33056 9680 33068
rect 9732 33056 9738 33108
rect 10410 33056 10416 33108
rect 10468 33096 10474 33108
rect 10468 33068 12940 33096
rect 10468 33056 10474 33068
rect 7009 33031 7067 33037
rect 7009 32997 7021 33031
rect 7055 32997 7067 33031
rect 7009 32991 7067 32997
rect 5102 32963 5160 32969
rect 5102 32960 5114 32963
rect 4816 32932 5114 32960
rect 5102 32929 5114 32932
rect 5148 32929 5160 32963
rect 5102 32923 5160 32929
rect 5261 32963 5319 32969
rect 5261 32929 5273 32963
rect 5307 32960 5319 32963
rect 5626 32960 5632 32972
rect 5307 32932 5632 32960
rect 5307 32929 5319 32932
rect 5261 32923 5319 32929
rect 5626 32920 5632 32932
rect 5684 32920 5690 32972
rect 1670 32852 1676 32904
rect 1728 32852 1734 32904
rect 1762 32852 1768 32904
rect 1820 32852 1826 32904
rect 2038 32901 2044 32904
rect 2032 32892 2044 32901
rect 1999 32864 2044 32892
rect 2032 32855 2044 32864
rect 2038 32852 2044 32855
rect 2096 32852 2102 32904
rect 4246 32852 4252 32904
rect 4304 32852 4310 32904
rect 4982 32852 4988 32904
rect 5040 32852 5046 32904
rect 6917 32895 6975 32901
rect 6917 32861 6929 32895
rect 6963 32892 6975 32895
rect 7024 32892 7052 32991
rect 7098 32920 7104 32972
rect 7156 32960 7162 32972
rect 7650 32960 7656 32972
rect 7156 32932 7656 32960
rect 7156 32920 7162 32932
rect 7650 32920 7656 32932
rect 7708 32920 7714 32972
rect 8202 32960 8208 32972
rect 7760 32932 8208 32960
rect 6963 32864 7052 32892
rect 6963 32861 6975 32864
rect 6917 32855 6975 32861
rect 7558 32852 7564 32904
rect 7616 32892 7622 32904
rect 7760 32892 7788 32932
rect 8202 32920 8208 32932
rect 8260 32960 8266 32972
rect 8389 32963 8447 32969
rect 8389 32960 8401 32963
rect 8260 32932 8401 32960
rect 8260 32920 8266 32932
rect 8389 32929 8401 32932
rect 8435 32929 8447 32963
rect 12912 32960 12940 33068
rect 12986 33056 12992 33108
rect 13044 33096 13050 33108
rect 13265 33099 13323 33105
rect 13265 33096 13277 33099
rect 13044 33068 13277 33096
rect 13044 33056 13050 33068
rect 13265 33065 13277 33068
rect 13311 33096 13323 33099
rect 13311 33068 14228 33096
rect 13311 33065 13323 33068
rect 13265 33059 13323 33065
rect 14200 33028 14228 33068
rect 14274 33056 14280 33108
rect 14332 33096 14338 33108
rect 16025 33099 16083 33105
rect 14332 33068 15976 33096
rect 14332 33056 14338 33068
rect 14642 33028 14648 33040
rect 14200 33000 14648 33028
rect 14642 32988 14648 33000
rect 14700 33028 14706 33040
rect 15948 33028 15976 33068
rect 16025 33065 16037 33099
rect 16071 33096 16083 33099
rect 16071 33068 21220 33096
rect 16071 33065 16083 33068
rect 16025 33059 16083 33065
rect 18049 33031 18107 33037
rect 14700 33000 14964 33028
rect 15948 33000 18000 33028
rect 14700 32988 14706 33000
rect 13906 32960 13912 32972
rect 8389 32923 8447 32929
rect 9232 32932 9444 32960
rect 12912 32932 13912 32960
rect 9232 32901 9260 32932
rect 7616 32864 7788 32892
rect 9217 32895 9275 32901
rect 7616 32852 7622 32864
rect 9217 32861 9229 32895
rect 9263 32861 9275 32895
rect 9217 32855 9275 32861
rect 9306 32852 9312 32904
rect 9364 32852 9370 32904
rect 9416 32892 9444 32932
rect 13906 32920 13912 32932
rect 13964 32920 13970 32972
rect 14182 32920 14188 32972
rect 14240 32920 14246 32972
rect 14826 32920 14832 32972
rect 14884 32920 14890 32972
rect 14936 32960 14964 33000
rect 15105 32963 15163 32969
rect 15105 32960 15117 32963
rect 14936 32932 15117 32960
rect 15105 32929 15117 32932
rect 15151 32929 15163 32963
rect 15105 32923 15163 32929
rect 16942 32920 16948 32972
rect 17000 32920 17006 32972
rect 17034 32920 17040 32972
rect 17092 32960 17098 32972
rect 17773 32963 17831 32969
rect 17773 32960 17785 32963
rect 17092 32932 17785 32960
rect 17092 32920 17098 32932
rect 17773 32929 17785 32932
rect 17819 32960 17831 32963
rect 17862 32960 17868 32972
rect 17819 32932 17868 32960
rect 17819 32929 17831 32932
rect 17773 32923 17831 32929
rect 17862 32920 17868 32932
rect 17920 32920 17926 32972
rect 17972 32960 18000 33000
rect 18049 32997 18061 33031
rect 18095 33028 18107 33031
rect 18095 33000 19288 33028
rect 18095 32997 18107 33000
rect 18049 32991 18107 32997
rect 17972 32932 18552 32960
rect 12158 32901 12164 32904
rect 11885 32895 11943 32901
rect 9416 32864 9720 32892
rect 9692 32836 9720 32864
rect 11885 32861 11897 32895
rect 11931 32861 11943 32895
rect 12152 32892 12164 32901
rect 12119 32864 12164 32892
rect 11885 32855 11943 32861
rect 12152 32855 12164 32864
rect 5905 32827 5963 32833
rect 5905 32793 5917 32827
rect 5951 32824 5963 32827
rect 7469 32827 7527 32833
rect 5951 32796 6960 32824
rect 5951 32793 5963 32796
rect 5905 32787 5963 32793
rect 6932 32768 6960 32796
rect 7469 32793 7481 32827
rect 7515 32824 7527 32827
rect 9554 32827 9612 32833
rect 9554 32824 9566 32827
rect 7515 32796 8340 32824
rect 7515 32793 7527 32796
rect 7469 32787 7527 32793
rect 1486 32716 1492 32768
rect 1544 32716 1550 32768
rect 4522 32716 4528 32768
rect 4580 32756 4586 32768
rect 5350 32756 5356 32768
rect 4580 32728 5356 32756
rect 4580 32716 4586 32728
rect 5350 32716 5356 32728
rect 5408 32716 5414 32768
rect 6730 32716 6736 32768
rect 6788 32716 6794 32768
rect 6914 32716 6920 32768
rect 6972 32716 6978 32768
rect 7377 32759 7435 32765
rect 7377 32725 7389 32759
rect 7423 32756 7435 32759
rect 7742 32756 7748 32768
rect 7423 32728 7748 32756
rect 7423 32725 7435 32728
rect 7377 32719 7435 32725
rect 7742 32716 7748 32728
rect 7800 32716 7806 32768
rect 7834 32716 7840 32768
rect 7892 32716 7898 32768
rect 8202 32716 8208 32768
rect 8260 32716 8266 32768
rect 8312 32765 8340 32796
rect 9048 32796 9566 32824
rect 8297 32759 8355 32765
rect 8297 32725 8309 32759
rect 8343 32756 8355 32759
rect 8478 32756 8484 32768
rect 8343 32728 8484 32756
rect 8343 32725 8355 32728
rect 8297 32719 8355 32725
rect 8478 32716 8484 32728
rect 8536 32716 8542 32768
rect 9048 32765 9076 32796
rect 9554 32793 9566 32796
rect 9600 32793 9612 32827
rect 9554 32787 9612 32793
rect 9674 32784 9680 32836
rect 9732 32784 9738 32836
rect 9784 32796 10824 32824
rect 9033 32759 9091 32765
rect 9033 32725 9045 32759
rect 9079 32725 9091 32759
rect 9033 32719 9091 32725
rect 9122 32716 9128 32768
rect 9180 32756 9186 32768
rect 9784 32756 9812 32796
rect 9180 32728 9812 32756
rect 9180 32716 9186 32728
rect 9858 32716 9864 32768
rect 9916 32756 9922 32768
rect 10689 32759 10747 32765
rect 10689 32756 10701 32759
rect 9916 32728 10701 32756
rect 9916 32716 9922 32728
rect 10689 32725 10701 32728
rect 10735 32725 10747 32759
rect 10796 32756 10824 32796
rect 11790 32784 11796 32836
rect 11848 32824 11854 32836
rect 11900 32824 11928 32855
rect 12158 32852 12164 32855
rect 12216 32852 12222 32904
rect 14090 32852 14096 32904
rect 14148 32892 14154 32904
rect 14369 32895 14427 32901
rect 14369 32892 14381 32895
rect 14148 32864 14381 32892
rect 14148 32852 14154 32864
rect 14369 32861 14381 32864
rect 14415 32861 14427 32895
rect 14369 32855 14427 32861
rect 15194 32852 15200 32904
rect 15252 32901 15258 32904
rect 15252 32895 15280 32901
rect 15268 32861 15280 32895
rect 15252 32855 15280 32861
rect 15252 32852 15258 32855
rect 15378 32852 15384 32904
rect 15436 32852 15442 32904
rect 18233 32895 18291 32901
rect 18233 32888 18245 32895
rect 18156 32861 18245 32888
rect 18279 32861 18291 32895
rect 18156 32860 18291 32861
rect 12618 32824 12624 32836
rect 11848 32796 12624 32824
rect 11848 32784 11854 32796
rect 12618 32784 12624 32796
rect 12676 32784 12682 32836
rect 14274 32824 14280 32836
rect 13832 32796 14280 32824
rect 13832 32756 13860 32796
rect 14274 32784 14280 32796
rect 14332 32784 14338 32836
rect 15930 32784 15936 32836
rect 15988 32824 15994 32836
rect 16761 32827 16819 32833
rect 16761 32824 16773 32827
rect 15988 32796 16773 32824
rect 15988 32784 15994 32796
rect 16761 32793 16773 32796
rect 16807 32824 16819 32827
rect 17589 32827 17647 32833
rect 16807 32796 17540 32824
rect 16807 32793 16819 32796
rect 16761 32787 16819 32793
rect 10796 32728 13860 32756
rect 10689 32719 10747 32725
rect 13906 32716 13912 32768
rect 13964 32756 13970 32768
rect 15102 32756 15108 32768
rect 13964 32728 15108 32756
rect 13964 32716 13970 32728
rect 15102 32716 15108 32728
rect 15160 32716 15166 32768
rect 17218 32716 17224 32768
rect 17276 32716 17282 32768
rect 17512 32756 17540 32796
rect 17589 32793 17601 32827
rect 17635 32824 17647 32827
rect 18046 32824 18052 32836
rect 17635 32796 18052 32824
rect 17635 32793 17647 32796
rect 17589 32787 17647 32793
rect 18046 32784 18052 32796
rect 18104 32784 18110 32836
rect 17681 32759 17739 32765
rect 17681 32756 17693 32759
rect 17512 32728 17693 32756
rect 17681 32725 17693 32728
rect 17727 32756 17739 32759
rect 17954 32756 17960 32768
rect 17727 32728 17960 32756
rect 17727 32725 17739 32728
rect 17681 32719 17739 32725
rect 17954 32716 17960 32728
rect 18012 32716 18018 32768
rect 18156 32756 18184 32860
rect 18233 32855 18291 32860
rect 18524 32824 18552 32932
rect 18874 32920 18880 32972
rect 18932 32920 18938 32972
rect 19260 32960 19288 33000
rect 19260 32932 19380 32960
rect 18598 32852 18604 32904
rect 18656 32892 18662 32904
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 18656 32864 19257 32892
rect 18656 32852 18662 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 19352 32892 19380 32932
rect 20254 32920 20260 32972
rect 20312 32960 20318 32972
rect 20990 32960 20996 32972
rect 20312 32932 20996 32960
rect 20312 32920 20318 32932
rect 20990 32920 20996 32932
rect 21048 32920 21054 32972
rect 21192 32969 21220 33068
rect 23106 33056 23112 33108
rect 23164 33096 23170 33108
rect 23201 33099 23259 33105
rect 23201 33096 23213 33099
rect 23164 33068 23213 33096
rect 23164 33056 23170 33068
rect 23201 33065 23213 33068
rect 23247 33065 23259 33099
rect 25774 33096 25780 33108
rect 23201 33059 23259 33065
rect 24504 33068 25780 33096
rect 24504 33028 24532 33068
rect 25774 33056 25780 33068
rect 25832 33056 25838 33108
rect 26050 33056 26056 33108
rect 26108 33056 26114 33108
rect 30006 33096 30012 33108
rect 26160 33068 30012 33096
rect 22066 33000 24532 33028
rect 21177 32963 21235 32969
rect 21177 32929 21189 32963
rect 21223 32929 21235 32963
rect 21177 32923 21235 32929
rect 21361 32963 21419 32969
rect 21361 32929 21373 32963
rect 21407 32960 21419 32963
rect 22066 32960 22094 33000
rect 22370 32960 22376 32972
rect 21407 32932 22094 32960
rect 22296 32932 22376 32960
rect 21407 32929 21419 32932
rect 21361 32923 21419 32929
rect 19501 32895 19559 32901
rect 19501 32892 19513 32895
rect 19352 32864 19513 32892
rect 19245 32855 19303 32861
rect 19501 32861 19513 32864
rect 19547 32861 19559 32895
rect 19501 32855 19559 32861
rect 19794 32852 19800 32904
rect 19852 32892 19858 32904
rect 22296 32892 22324 32932
rect 22370 32920 22376 32932
rect 22428 32920 22434 32972
rect 22554 32920 22560 32972
rect 22612 32960 22618 32972
rect 22925 32963 22983 32969
rect 22925 32960 22937 32963
rect 22612 32932 22937 32960
rect 22612 32920 22618 32932
rect 22925 32929 22937 32932
rect 22971 32960 22983 32963
rect 23106 32960 23112 32972
rect 22971 32932 23112 32960
rect 22971 32929 22983 32932
rect 22925 32923 22983 32929
rect 23106 32920 23112 32932
rect 23164 32920 23170 32972
rect 23385 32895 23443 32901
rect 23385 32892 23397 32895
rect 19852 32864 22324 32892
rect 22388 32864 23397 32892
rect 19852 32852 19858 32864
rect 21634 32824 21640 32836
rect 18524 32796 21640 32824
rect 21634 32784 21640 32796
rect 21692 32784 21698 32836
rect 18325 32759 18383 32765
rect 18325 32756 18337 32759
rect 18156 32728 18337 32756
rect 18325 32725 18337 32728
rect 18371 32725 18383 32759
rect 18325 32719 18383 32725
rect 18506 32716 18512 32768
rect 18564 32756 18570 32768
rect 18693 32759 18751 32765
rect 18693 32756 18705 32759
rect 18564 32728 18705 32756
rect 18564 32716 18570 32728
rect 18693 32725 18705 32728
rect 18739 32725 18751 32759
rect 18693 32719 18751 32725
rect 18785 32759 18843 32765
rect 18785 32725 18797 32759
rect 18831 32756 18843 32759
rect 19150 32756 19156 32768
rect 18831 32728 19156 32756
rect 18831 32725 18843 32728
rect 18785 32719 18843 32725
rect 19150 32716 19156 32728
rect 19208 32756 19214 32768
rect 20625 32759 20683 32765
rect 20625 32756 20637 32759
rect 19208 32728 20637 32756
rect 19208 32716 19214 32728
rect 20625 32725 20637 32728
rect 20671 32725 20683 32759
rect 20625 32719 20683 32725
rect 20714 32716 20720 32768
rect 20772 32716 20778 32768
rect 20806 32716 20812 32768
rect 20864 32756 20870 32768
rect 22388 32765 22416 32864
rect 23385 32861 23397 32864
rect 23431 32861 23443 32895
rect 23385 32855 23443 32861
rect 24489 32895 24547 32901
rect 24489 32861 24501 32895
rect 24535 32892 24547 32895
rect 24578 32892 24584 32904
rect 24535 32864 24584 32892
rect 24535 32861 24547 32864
rect 24489 32855 24547 32861
rect 22462 32784 22468 32836
rect 22520 32824 22526 32836
rect 22833 32827 22891 32833
rect 22833 32824 22845 32827
rect 22520 32796 22845 32824
rect 22520 32784 22526 32796
rect 22833 32793 22845 32796
rect 22879 32793 22891 32827
rect 22833 32787 22891 32793
rect 22922 32784 22928 32836
rect 22980 32824 22986 32836
rect 24504 32824 24532 32855
rect 24578 32852 24584 32864
rect 24636 32852 24642 32904
rect 26160 32892 26188 33068
rect 30006 33056 30012 33068
rect 30064 33096 30070 33108
rect 30064 33068 30297 33096
rect 30064 33056 30070 33068
rect 26329 33031 26387 33037
rect 26329 32997 26341 33031
rect 26375 32997 26387 33031
rect 28994 33028 29000 33040
rect 26329 32991 26387 32997
rect 26804 33000 29000 33028
rect 24688 32864 26188 32892
rect 26237 32895 26295 32901
rect 24688 32824 24716 32864
rect 26237 32861 26249 32895
rect 26283 32892 26295 32895
rect 26344 32892 26372 32991
rect 26804 32972 26832 33000
rect 28994 32988 29000 33000
rect 29052 32988 29058 33040
rect 26786 32920 26792 32972
rect 26844 32920 26850 32972
rect 26878 32920 26884 32972
rect 26936 32960 26942 32972
rect 26973 32963 27031 32969
rect 26973 32960 26985 32963
rect 26936 32932 26985 32960
rect 26936 32920 26942 32932
rect 26973 32929 26985 32932
rect 27019 32960 27031 32963
rect 27154 32960 27160 32972
rect 27019 32932 27160 32960
rect 27019 32929 27031 32932
rect 26973 32923 27031 32929
rect 27154 32920 27160 32932
rect 27212 32920 27218 32972
rect 29638 32920 29644 32972
rect 29696 32960 29702 32972
rect 30009 32963 30067 32969
rect 30009 32960 30021 32963
rect 29696 32932 30021 32960
rect 29696 32920 29702 32932
rect 30009 32929 30021 32932
rect 30055 32929 30067 32963
rect 30009 32923 30067 32929
rect 30101 32963 30159 32969
rect 30101 32929 30113 32963
rect 30147 32960 30159 32963
rect 30269 32960 30297 33068
rect 32398 33056 32404 33108
rect 32456 33096 32462 33108
rect 33502 33096 33508 33108
rect 32456 33068 33508 33096
rect 32456 33056 32462 33068
rect 33502 33056 33508 33068
rect 33560 33056 33566 33108
rect 38654 33056 38660 33108
rect 38712 33056 38718 33108
rect 38933 33099 38991 33105
rect 38933 33065 38945 33099
rect 38979 33096 38991 33099
rect 39298 33096 39304 33108
rect 38979 33068 39304 33096
rect 38979 33065 38991 33068
rect 38933 33059 38991 33065
rect 39298 33056 39304 33068
rect 39356 33056 39362 33108
rect 41049 33099 41107 33105
rect 41049 33065 41061 33099
rect 41095 33096 41107 33099
rect 41874 33096 41880 33108
rect 41095 33068 41880 33096
rect 41095 33065 41107 33068
rect 41049 33059 41107 33065
rect 41874 33056 41880 33068
rect 41932 33056 41938 33108
rect 42334 33056 42340 33108
rect 42392 33096 42398 33108
rect 42392 33068 42472 33096
rect 42392 33056 42398 33068
rect 37185 33031 37243 33037
rect 37185 32997 37197 33031
rect 37231 33028 37243 33031
rect 37366 33028 37372 33040
rect 37231 33000 37372 33028
rect 37231 32997 37243 33000
rect 37185 32991 37243 32997
rect 37366 32988 37372 33000
rect 37424 32988 37430 33040
rect 41598 32988 41604 33040
rect 41656 32988 41662 33040
rect 30147 32932 30297 32960
rect 30147 32929 30159 32932
rect 30101 32923 30159 32929
rect 36814 32920 36820 32972
rect 36872 32920 36878 32972
rect 40865 32963 40923 32969
rect 40865 32929 40877 32963
rect 40911 32960 40923 32963
rect 41966 32960 41972 32972
rect 40911 32932 41972 32960
rect 40911 32929 40923 32932
rect 40865 32923 40923 32929
rect 41966 32920 41972 32932
rect 42024 32920 42030 32972
rect 26283 32864 26372 32892
rect 26283 32861 26295 32864
rect 26237 32855 26295 32861
rect 26510 32852 26516 32904
rect 26568 32892 26574 32904
rect 26697 32895 26755 32901
rect 26697 32892 26709 32895
rect 26568 32864 26709 32892
rect 26568 32852 26574 32864
rect 26697 32861 26709 32864
rect 26743 32892 26755 32895
rect 27522 32892 27528 32904
rect 26743 32864 27528 32892
rect 26743 32861 26755 32864
rect 26697 32855 26755 32861
rect 27522 32852 27528 32864
rect 27580 32852 27586 32904
rect 29365 32895 29423 32901
rect 29365 32861 29377 32895
rect 29411 32892 29423 32895
rect 30374 32892 30380 32904
rect 29411 32864 30380 32892
rect 29411 32861 29423 32864
rect 29365 32855 29423 32861
rect 30374 32852 30380 32864
rect 30432 32852 30438 32904
rect 32122 32852 32128 32904
rect 32180 32852 32186 32904
rect 32217 32895 32275 32901
rect 32217 32861 32229 32895
rect 32263 32892 32275 32895
rect 32306 32892 32312 32904
rect 32263 32864 32312 32892
rect 32263 32861 32275 32864
rect 32217 32855 32275 32861
rect 32306 32852 32312 32864
rect 32364 32892 32370 32904
rect 33410 32892 33416 32904
rect 32364 32864 33416 32892
rect 32364 32852 32370 32864
rect 33410 32852 33416 32864
rect 33468 32852 33474 32904
rect 34422 32852 34428 32904
rect 34480 32892 34486 32904
rect 35713 32895 35771 32901
rect 35713 32892 35725 32895
rect 34480 32864 35725 32892
rect 34480 32852 34486 32864
rect 35713 32861 35725 32864
rect 35759 32861 35771 32895
rect 35713 32855 35771 32861
rect 24762 32833 24768 32836
rect 22980 32796 24532 32824
rect 24596 32796 24716 32824
rect 22980 32784 22986 32796
rect 24596 32768 24624 32796
rect 24756 32787 24768 32833
rect 24762 32784 24768 32787
rect 24820 32784 24826 32836
rect 25332 32796 26556 32824
rect 21085 32759 21143 32765
rect 21085 32756 21097 32759
rect 20864 32728 21097 32756
rect 20864 32716 20870 32728
rect 21085 32725 21097 32728
rect 21131 32725 21143 32759
rect 21085 32719 21143 32725
rect 22373 32759 22431 32765
rect 22373 32725 22385 32759
rect 22419 32725 22431 32759
rect 22373 32719 22431 32725
rect 22741 32759 22799 32765
rect 22741 32725 22753 32759
rect 22787 32756 22799 32759
rect 24394 32756 24400 32768
rect 22787 32728 24400 32756
rect 22787 32725 22799 32728
rect 22741 32719 22799 32725
rect 24394 32716 24400 32728
rect 24452 32716 24458 32768
rect 24578 32716 24584 32768
rect 24636 32716 24642 32768
rect 24670 32716 24676 32768
rect 24728 32756 24734 32768
rect 25332 32756 25360 32796
rect 24728 32728 25360 32756
rect 24728 32716 24734 32728
rect 25406 32716 25412 32768
rect 25464 32756 25470 32768
rect 25869 32759 25927 32765
rect 25869 32756 25881 32759
rect 25464 32728 25881 32756
rect 25464 32716 25470 32728
rect 25869 32725 25881 32728
rect 25915 32725 25927 32759
rect 26528 32756 26556 32796
rect 26602 32784 26608 32836
rect 26660 32824 26666 32836
rect 30742 32824 30748 32836
rect 26660 32796 30748 32824
rect 26660 32784 26666 32796
rect 30742 32784 30748 32796
rect 30800 32784 30806 32836
rect 32473 32827 32531 32833
rect 32473 32824 32485 32827
rect 32416 32796 32485 32824
rect 28350 32756 28356 32768
rect 26528 32728 28356 32756
rect 25869 32719 25927 32725
rect 28350 32716 28356 32728
rect 28408 32716 28414 32768
rect 29181 32759 29239 32765
rect 29181 32725 29193 32759
rect 29227 32756 29239 32759
rect 29270 32756 29276 32768
rect 29227 32728 29276 32756
rect 29227 32725 29239 32728
rect 29181 32719 29239 32725
rect 29270 32716 29276 32728
rect 29328 32716 29334 32768
rect 29362 32716 29368 32768
rect 29420 32756 29426 32768
rect 29549 32759 29607 32765
rect 29549 32756 29561 32759
rect 29420 32728 29561 32756
rect 29420 32716 29426 32728
rect 29549 32725 29561 32728
rect 29595 32725 29607 32759
rect 29549 32719 29607 32725
rect 29917 32759 29975 32765
rect 29917 32725 29929 32759
rect 29963 32756 29975 32759
rect 30650 32756 30656 32768
rect 29963 32728 30656 32756
rect 29963 32725 29975 32728
rect 29917 32719 29975 32725
rect 30650 32716 30656 32728
rect 30708 32716 30714 32768
rect 31941 32759 31999 32765
rect 31941 32725 31953 32759
rect 31987 32756 31999 32759
rect 32416 32756 32444 32796
rect 32473 32793 32485 32796
rect 32519 32793 32531 32827
rect 35728 32824 35756 32855
rect 35986 32852 35992 32904
rect 36044 32852 36050 32904
rect 37090 32852 37096 32904
rect 37148 32892 37154 32904
rect 37148 32864 37780 32892
rect 37148 32852 37154 32864
rect 36078 32824 36084 32836
rect 35728 32796 36084 32824
rect 32473 32787 32531 32793
rect 36078 32784 36084 32796
rect 36136 32784 36142 32836
rect 37752 32824 37780 32864
rect 37826 32852 37832 32904
rect 37884 32892 37890 32904
rect 38194 32892 38200 32904
rect 37884 32864 38200 32892
rect 37884 32852 37890 32864
rect 38194 32852 38200 32864
rect 38252 32892 38258 32904
rect 38473 32895 38531 32901
rect 38473 32892 38485 32895
rect 38252 32864 38485 32892
rect 38252 32852 38258 32864
rect 38473 32861 38485 32864
rect 38519 32861 38531 32895
rect 40957 32895 41015 32901
rect 40957 32892 40969 32895
rect 38473 32855 38531 32861
rect 40512 32864 40969 32892
rect 40512 32836 40540 32864
rect 40957 32861 40969 32864
rect 41003 32861 41015 32895
rect 40957 32855 41015 32861
rect 41141 32895 41199 32901
rect 41141 32861 41153 32895
rect 41187 32861 41199 32895
rect 41141 32855 41199 32861
rect 38105 32827 38163 32833
rect 38105 32824 38117 32827
rect 36740 32796 37688 32824
rect 37752 32796 38117 32824
rect 31987 32728 32444 32756
rect 31987 32725 31999 32728
rect 31941 32719 31999 32725
rect 32674 32716 32680 32768
rect 32732 32756 32738 32768
rect 36740 32765 36768 32796
rect 37660 32768 37688 32796
rect 38105 32793 38117 32796
rect 38151 32793 38163 32827
rect 38105 32787 38163 32793
rect 38289 32827 38347 32833
rect 38289 32793 38301 32827
rect 38335 32824 38347 32827
rect 39022 32824 39028 32836
rect 38335 32796 39028 32824
rect 38335 32793 38347 32796
rect 38289 32787 38347 32793
rect 39022 32784 39028 32796
rect 39080 32784 39086 32836
rect 40494 32784 40500 32836
rect 40552 32784 40558 32836
rect 40681 32827 40739 32833
rect 40681 32793 40693 32827
rect 40727 32824 40739 32827
rect 40770 32824 40776 32836
rect 40727 32796 40776 32824
rect 40727 32793 40739 32796
rect 40681 32787 40739 32793
rect 40770 32784 40776 32796
rect 40828 32824 40834 32836
rect 41156 32824 41184 32855
rect 41782 32852 41788 32904
rect 41840 32852 41846 32904
rect 41878 32895 41936 32901
rect 41878 32861 41890 32895
rect 41924 32886 41936 32895
rect 41924 32861 42012 32886
rect 41878 32858 42012 32861
rect 41878 32855 41936 32858
rect 40828 32796 41184 32824
rect 41984 32824 42012 32858
rect 42058 32852 42064 32904
rect 42116 32852 42122 32904
rect 42242 32894 42248 32904
rect 42168 32866 42248 32894
rect 42168 32824 42196 32866
rect 42242 32852 42248 32866
rect 42300 32852 42306 32904
rect 42444 32901 42472 33068
rect 43806 33056 43812 33108
rect 43864 33096 43870 33108
rect 43864 33068 44312 33096
rect 43864 33056 43870 33068
rect 42518 32988 42524 33040
rect 42576 32988 42582 33040
rect 44284 32960 44312 33068
rect 44358 33056 44364 33108
rect 44416 33096 44422 33108
rect 44542 33096 44548 33108
rect 44416 33068 44548 33096
rect 44416 33056 44422 33068
rect 44542 33056 44548 33068
rect 44600 33056 44606 33108
rect 44634 33056 44640 33108
rect 44692 33096 44698 33108
rect 45097 33099 45155 33105
rect 45097 33096 45109 33099
rect 44692 33068 45109 33096
rect 44692 33056 44698 33068
rect 45097 33065 45109 33068
rect 45143 33065 45155 33099
rect 45097 33059 45155 33065
rect 45112 33028 45140 33059
rect 45462 33056 45468 33108
rect 45520 33056 45526 33108
rect 46014 33056 46020 33108
rect 46072 33056 46078 33108
rect 45830 33028 45836 33040
rect 45112 33000 45836 33028
rect 45830 32988 45836 33000
rect 45888 32988 45894 33040
rect 44284 32932 45554 32960
rect 42429 32895 42487 32901
rect 42429 32861 42441 32895
rect 42475 32861 42487 32895
rect 42429 32855 42487 32861
rect 42610 32852 42616 32904
rect 42668 32892 42674 32904
rect 42705 32895 42763 32901
rect 42705 32892 42717 32895
rect 42668 32864 42717 32892
rect 42668 32852 42674 32864
rect 42705 32861 42717 32864
rect 42751 32861 42763 32895
rect 42705 32855 42763 32861
rect 42797 32895 42855 32901
rect 42797 32861 42809 32895
rect 42843 32892 42855 32895
rect 42886 32892 42892 32904
rect 42843 32864 42892 32892
rect 42843 32861 42855 32864
rect 42797 32855 42855 32861
rect 42886 32852 42892 32864
rect 42944 32852 42950 32904
rect 44269 32895 44327 32901
rect 44269 32861 44281 32895
rect 44315 32892 44327 32895
rect 44315 32864 44956 32892
rect 44315 32861 44327 32864
rect 44269 32855 44327 32861
rect 41984 32796 42196 32824
rect 40828 32784 40834 32796
rect 42518 32784 42524 32836
rect 42576 32784 42582 32836
rect 44634 32824 44640 32836
rect 42812 32796 44640 32824
rect 42812 32768 42840 32796
rect 44634 32784 44640 32796
rect 44692 32784 44698 32836
rect 44928 32824 44956 32864
rect 45002 32852 45008 32904
rect 45060 32852 45066 32904
rect 45526 32892 45554 32932
rect 46477 32895 46535 32901
rect 46477 32892 46489 32895
rect 45526 32864 46489 32892
rect 46477 32861 46489 32864
rect 46523 32861 46535 32895
rect 46477 32855 46535 32861
rect 45094 32824 45100 32836
rect 44928 32796 45100 32824
rect 45094 32784 45100 32796
rect 45152 32824 45158 32836
rect 45557 32827 45615 32833
rect 45557 32824 45569 32827
rect 45152 32796 45569 32824
rect 45152 32784 45158 32796
rect 45557 32793 45569 32796
rect 45603 32793 45615 32827
rect 45557 32787 45615 32793
rect 33597 32759 33655 32765
rect 33597 32756 33609 32759
rect 32732 32728 33609 32756
rect 32732 32716 32738 32728
rect 33597 32725 33609 32728
rect 33643 32725 33655 32759
rect 33597 32719 33655 32725
rect 36725 32759 36783 32765
rect 36725 32725 36737 32759
rect 36771 32725 36783 32759
rect 36725 32719 36783 32725
rect 37274 32716 37280 32768
rect 37332 32716 37338 32768
rect 37642 32716 37648 32768
rect 37700 32756 37706 32768
rect 41690 32756 41696 32768
rect 37700 32728 41696 32756
rect 37700 32716 37706 32728
rect 41690 32716 41696 32728
rect 41748 32716 41754 32768
rect 42426 32716 42432 32768
rect 42484 32716 42490 32768
rect 42794 32716 42800 32768
rect 42852 32716 42858 32768
rect 44729 32759 44787 32765
rect 44729 32725 44741 32759
rect 44775 32756 44787 32759
rect 44910 32756 44916 32768
rect 44775 32728 44916 32756
rect 44775 32725 44787 32728
rect 44729 32719 44787 32725
rect 44910 32716 44916 32728
rect 44968 32716 44974 32768
rect 46658 32716 46664 32768
rect 46716 32716 46722 32768
rect 1104 32666 47104 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 47104 32666
rect 1104 32592 47104 32614
rect 1670 32512 1676 32564
rect 1728 32552 1734 32564
rect 3145 32555 3203 32561
rect 3145 32552 3157 32555
rect 1728 32524 3157 32552
rect 1728 32512 1734 32524
rect 3145 32521 3157 32524
rect 3191 32521 3203 32555
rect 3145 32515 3203 32521
rect 3513 32555 3571 32561
rect 3513 32521 3525 32555
rect 3559 32552 3571 32555
rect 4982 32552 4988 32564
rect 3559 32524 4988 32552
rect 3559 32521 3571 32524
rect 3513 32515 3571 32521
rect 1486 32444 1492 32496
rect 1544 32484 1550 32496
rect 1918 32487 1976 32493
rect 1918 32484 1930 32487
rect 1544 32456 1930 32484
rect 1544 32444 1550 32456
rect 1918 32453 1930 32456
rect 1964 32453 1976 32487
rect 1918 32447 1976 32453
rect 1673 32419 1731 32425
rect 1673 32385 1685 32419
rect 1719 32416 1731 32419
rect 1762 32416 1768 32428
rect 1719 32388 1768 32416
rect 1719 32385 1731 32388
rect 1673 32379 1731 32385
rect 1762 32376 1768 32388
rect 1820 32376 1826 32428
rect 3053 32283 3111 32289
rect 3053 32249 3065 32283
rect 3099 32280 3111 32283
rect 3528 32280 3556 32515
rect 4982 32512 4988 32524
rect 5040 32512 5046 32564
rect 5905 32555 5963 32561
rect 5905 32521 5917 32555
rect 5951 32552 5963 32555
rect 5951 32524 7696 32552
rect 5951 32521 5963 32524
rect 5905 32515 5963 32521
rect 3602 32444 3608 32496
rect 3660 32484 3666 32496
rect 3970 32484 3976 32496
rect 3660 32456 3976 32484
rect 3660 32444 3666 32456
rect 3970 32444 3976 32456
rect 4028 32444 4034 32496
rect 6632 32487 6690 32493
rect 6632 32453 6644 32487
rect 6678 32484 6690 32487
rect 6730 32484 6736 32496
rect 6678 32456 6736 32484
rect 6678 32453 6690 32456
rect 6632 32447 6690 32453
rect 6730 32444 6736 32456
rect 6788 32444 6794 32496
rect 7668 32484 7696 32524
rect 7742 32512 7748 32564
rect 7800 32552 7806 32564
rect 10502 32552 10508 32564
rect 7800 32524 10508 32552
rect 7800 32512 7806 32524
rect 10502 32512 10508 32524
rect 10560 32512 10566 32564
rect 11517 32555 11575 32561
rect 11517 32521 11529 32555
rect 11563 32552 11575 32555
rect 12066 32552 12072 32564
rect 11563 32524 12072 32552
rect 11563 32521 11575 32524
rect 11517 32515 11575 32521
rect 12066 32512 12072 32524
rect 12124 32512 12130 32564
rect 12618 32512 12624 32564
rect 12676 32512 12682 32564
rect 13173 32555 13231 32561
rect 13173 32521 13185 32555
rect 13219 32552 13231 32555
rect 13354 32552 13360 32564
rect 13219 32524 13360 32552
rect 13219 32521 13231 32524
rect 13173 32515 13231 32521
rect 13354 32512 13360 32524
rect 13412 32552 13418 32564
rect 14918 32552 14924 32564
rect 13412 32524 14924 32552
rect 13412 32512 13418 32524
rect 14918 32512 14924 32524
rect 14976 32552 14982 32564
rect 15194 32552 15200 32564
rect 14976 32524 15200 32552
rect 14976 32512 14982 32524
rect 15194 32512 15200 32524
rect 15252 32512 15258 32564
rect 15749 32555 15807 32561
rect 15749 32521 15761 32555
rect 15795 32552 15807 32555
rect 17954 32552 17960 32564
rect 15795 32524 17960 32552
rect 15795 32521 15807 32524
rect 15749 32515 15807 32521
rect 17954 32512 17960 32524
rect 18012 32512 18018 32564
rect 18046 32512 18052 32564
rect 18104 32512 18110 32564
rect 18138 32512 18144 32564
rect 18196 32552 18202 32564
rect 18601 32555 18659 32561
rect 18601 32552 18613 32555
rect 18196 32524 18613 32552
rect 18196 32512 18202 32524
rect 18601 32521 18613 32524
rect 18647 32552 18659 32555
rect 18782 32552 18788 32564
rect 18647 32524 18788 32552
rect 18647 32521 18659 32524
rect 18601 32515 18659 32521
rect 18782 32512 18788 32524
rect 18840 32512 18846 32564
rect 18892 32524 20668 32552
rect 9122 32484 9128 32496
rect 7668 32456 9128 32484
rect 9122 32444 9128 32456
rect 9180 32444 9186 32496
rect 12636 32484 12664 32512
rect 13998 32484 14004 32496
rect 12636 32456 14004 32484
rect 13998 32444 14004 32456
rect 14056 32444 14062 32496
rect 16914 32487 16972 32493
rect 16914 32484 16926 32487
rect 16132 32456 16926 32484
rect 4065 32419 4123 32425
rect 4065 32385 4077 32419
rect 4111 32416 4123 32419
rect 4154 32416 4160 32428
rect 4111 32388 4160 32416
rect 4111 32385 4123 32388
rect 4065 32379 4123 32385
rect 4154 32376 4160 32388
rect 4212 32376 4218 32428
rect 4982 32376 4988 32428
rect 5040 32376 5046 32428
rect 6181 32419 6239 32425
rect 6181 32385 6193 32419
rect 6227 32416 6239 32419
rect 7834 32416 7840 32428
rect 6227 32388 7840 32416
rect 6227 32385 6239 32388
rect 6181 32379 6239 32385
rect 7834 32376 7840 32388
rect 7892 32376 7898 32428
rect 8196 32419 8254 32425
rect 8196 32385 8208 32419
rect 8242 32416 8254 32419
rect 8938 32416 8944 32428
rect 8242 32388 8944 32416
rect 8242 32385 8254 32388
rect 8196 32379 8254 32385
rect 8938 32376 8944 32388
rect 8996 32376 9002 32428
rect 9677 32419 9735 32425
rect 9677 32385 9689 32419
rect 9723 32416 9735 32419
rect 9858 32416 9864 32428
rect 9723 32388 9864 32416
rect 9723 32385 9735 32388
rect 9677 32379 9735 32385
rect 9858 32376 9864 32388
rect 9916 32376 9922 32428
rect 10502 32376 10508 32428
rect 10560 32425 10566 32428
rect 10560 32419 10588 32425
rect 10576 32385 10588 32419
rect 10560 32379 10588 32385
rect 10560 32376 10566 32379
rect 10686 32376 10692 32428
rect 10744 32376 10750 32428
rect 11606 32376 11612 32428
rect 11664 32416 11670 32428
rect 12066 32425 12072 32428
rect 11701 32419 11759 32425
rect 11701 32416 11713 32419
rect 11664 32388 11713 32416
rect 11664 32376 11670 32388
rect 11701 32385 11713 32388
rect 11747 32385 11759 32419
rect 11701 32379 11759 32385
rect 12060 32379 12072 32425
rect 12124 32416 12130 32428
rect 12124 32388 12160 32416
rect 12066 32376 12072 32379
rect 12124 32376 12130 32388
rect 13814 32376 13820 32428
rect 13872 32376 13878 32428
rect 13909 32419 13967 32425
rect 13909 32385 13921 32419
rect 13955 32416 13967 32419
rect 13955 32388 14228 32416
rect 13955 32385 13967 32388
rect 13909 32379 13967 32385
rect 3694 32308 3700 32360
rect 3752 32308 3758 32360
rect 4246 32308 4252 32360
rect 4304 32348 4310 32360
rect 4614 32348 4620 32360
rect 4304 32320 4620 32348
rect 4304 32308 4310 32320
rect 4614 32308 4620 32320
rect 4672 32308 4678 32360
rect 5102 32351 5160 32357
rect 5102 32348 5114 32351
rect 4816 32320 5114 32348
rect 3099 32252 3556 32280
rect 3099 32249 3111 32252
rect 3053 32243 3111 32249
rect 4522 32240 4528 32292
rect 4580 32280 4586 32292
rect 4709 32283 4767 32289
rect 4709 32280 4721 32283
rect 4580 32252 4721 32280
rect 4580 32240 4586 32252
rect 4709 32249 4721 32252
rect 4755 32249 4767 32283
rect 4709 32243 4767 32249
rect 4062 32172 4068 32224
rect 4120 32212 4126 32224
rect 4816 32212 4844 32320
rect 5102 32317 5114 32320
rect 5148 32317 5160 32351
rect 5102 32311 5160 32317
rect 5261 32351 5319 32357
rect 5261 32317 5273 32351
rect 5307 32348 5319 32351
rect 5442 32348 5448 32360
rect 5307 32320 5448 32348
rect 5307 32317 5319 32320
rect 5261 32311 5319 32317
rect 5442 32308 5448 32320
rect 5500 32348 5506 32360
rect 5500 32320 5764 32348
rect 5500 32308 5506 32320
rect 5736 32292 5764 32320
rect 6362 32308 6368 32360
rect 6420 32308 6426 32360
rect 7929 32351 7987 32357
rect 7929 32317 7941 32351
rect 7975 32317 7987 32351
rect 9493 32351 9551 32357
rect 9493 32348 9505 32351
rect 7929 32311 7987 32317
rect 9324 32320 9505 32348
rect 5718 32240 5724 32292
rect 5776 32240 5782 32292
rect 4120 32184 4844 32212
rect 5997 32215 6055 32221
rect 4120 32172 4126 32184
rect 5997 32181 6009 32215
rect 6043 32212 6055 32215
rect 6638 32212 6644 32224
rect 6043 32184 6644 32212
rect 6043 32181 6055 32184
rect 5997 32175 6055 32181
rect 6638 32172 6644 32184
rect 6696 32172 6702 32224
rect 6730 32172 6736 32224
rect 6788 32212 6794 32224
rect 7944 32212 7972 32311
rect 9214 32240 9220 32292
rect 9272 32280 9278 32292
rect 9324 32289 9352 32320
rect 9493 32317 9505 32320
rect 9539 32317 9551 32351
rect 10413 32351 10471 32357
rect 10413 32348 10425 32351
rect 9493 32311 9551 32317
rect 9968 32320 10425 32348
rect 9309 32283 9367 32289
rect 9309 32280 9321 32283
rect 9272 32252 9321 32280
rect 9272 32240 9278 32252
rect 9309 32249 9321 32252
rect 9355 32249 9367 32283
rect 9309 32243 9367 32249
rect 9968 32224 9996 32320
rect 10413 32317 10425 32320
rect 10459 32317 10471 32351
rect 10704 32348 10732 32376
rect 14200 32360 14228 32388
rect 14918 32376 14924 32428
rect 14976 32425 14982 32428
rect 14976 32419 15004 32425
rect 14992 32385 15004 32419
rect 14976 32379 15004 32385
rect 14976 32376 14982 32379
rect 15102 32376 15108 32428
rect 15160 32376 15166 32428
rect 10704 32320 11744 32348
rect 10413 32311 10471 32317
rect 10134 32240 10140 32292
rect 10192 32240 10198 32292
rect 6788 32184 7972 32212
rect 6788 32172 6794 32184
rect 8202 32172 8208 32224
rect 8260 32212 8266 32224
rect 9950 32212 9956 32224
rect 8260 32184 9956 32212
rect 8260 32172 8266 32184
rect 9950 32172 9956 32184
rect 10008 32172 10014 32224
rect 10152 32212 10180 32240
rect 11146 32212 11152 32224
rect 10152 32184 11152 32212
rect 11146 32172 11152 32184
rect 11204 32172 11210 32224
rect 11330 32172 11336 32224
rect 11388 32172 11394 32224
rect 11716 32212 11744 32320
rect 11790 32308 11796 32360
rect 11848 32308 11854 32360
rect 14090 32308 14096 32360
rect 14148 32308 14154 32360
rect 14182 32308 14188 32360
rect 14240 32308 14246 32360
rect 14642 32308 14648 32360
rect 14700 32348 14706 32360
rect 14829 32351 14887 32357
rect 14829 32348 14841 32351
rect 14700 32320 14841 32348
rect 14700 32308 14706 32320
rect 14829 32317 14841 32320
rect 14875 32317 14887 32351
rect 14829 32311 14887 32317
rect 14553 32283 14611 32289
rect 14553 32280 14565 32283
rect 12728 32252 14565 32280
rect 11790 32212 11796 32224
rect 11716 32184 11796 32212
rect 11790 32172 11796 32184
rect 11848 32172 11854 32224
rect 12526 32172 12532 32224
rect 12584 32212 12590 32224
rect 12728 32212 12756 32252
rect 14553 32249 14565 32252
rect 14599 32249 14611 32283
rect 16132 32280 16160 32456
rect 16914 32453 16926 32456
rect 16960 32453 16972 32487
rect 18064 32484 18092 32512
rect 18064 32456 18736 32484
rect 16914 32447 16972 32453
rect 16209 32419 16267 32425
rect 16209 32385 16221 32419
rect 16255 32416 16267 32419
rect 16390 32416 16396 32428
rect 16255 32388 16396 32416
rect 16255 32385 16267 32388
rect 16209 32379 16267 32385
rect 16390 32376 16396 32388
rect 16448 32376 16454 32428
rect 16485 32419 16543 32425
rect 16485 32385 16497 32419
rect 16531 32416 16543 32419
rect 17218 32416 17224 32428
rect 16531 32388 17224 32416
rect 16531 32385 16543 32388
rect 16485 32379 16543 32385
rect 17218 32376 17224 32388
rect 17276 32376 17282 32428
rect 18506 32376 18512 32428
rect 18564 32376 18570 32428
rect 16669 32351 16727 32357
rect 16669 32348 16681 32351
rect 16592 32320 16681 32348
rect 16301 32283 16359 32289
rect 16301 32280 16313 32283
rect 16132 32252 16313 32280
rect 14553 32243 14611 32249
rect 16301 32249 16313 32252
rect 16347 32249 16359 32283
rect 16301 32243 16359 32249
rect 12584 32184 12756 32212
rect 13633 32215 13691 32221
rect 12584 32172 12590 32184
rect 13633 32181 13645 32215
rect 13679 32212 13691 32215
rect 14274 32212 14280 32224
rect 13679 32184 14280 32212
rect 13679 32181 13691 32184
rect 13633 32175 13691 32181
rect 14274 32172 14280 32184
rect 14332 32172 14338 32224
rect 16022 32172 16028 32224
rect 16080 32172 16086 32224
rect 16390 32172 16396 32224
rect 16448 32212 16454 32224
rect 16592 32212 16620 32320
rect 16669 32317 16681 32320
rect 16715 32317 16727 32351
rect 16669 32311 16727 32317
rect 18708 32280 18736 32456
rect 18785 32351 18843 32357
rect 18785 32317 18797 32351
rect 18831 32348 18843 32351
rect 18892 32348 18920 32524
rect 20640 32484 20668 32524
rect 20806 32512 20812 32564
rect 20864 32512 20870 32564
rect 21450 32552 21456 32564
rect 20916 32524 21456 32552
rect 20916 32484 20944 32524
rect 21450 32512 21456 32524
rect 21508 32512 21514 32564
rect 21542 32512 21548 32564
rect 21600 32552 21606 32564
rect 24578 32552 24584 32564
rect 21600 32524 24584 32552
rect 21600 32512 21606 32524
rect 24578 32512 24584 32524
rect 24636 32512 24642 32564
rect 24762 32512 24768 32564
rect 24820 32512 24826 32564
rect 25406 32512 25412 32564
rect 25464 32552 25470 32564
rect 27982 32552 27988 32564
rect 25464 32524 27988 32552
rect 25464 32512 25470 32524
rect 27982 32512 27988 32524
rect 28040 32512 28046 32564
rect 29178 32512 29184 32564
rect 29236 32512 29242 32564
rect 30374 32512 30380 32564
rect 30432 32512 30438 32564
rect 30742 32512 30748 32564
rect 30800 32512 30806 32564
rect 32122 32512 32128 32564
rect 32180 32512 32186 32564
rect 32490 32512 32496 32564
rect 32548 32552 32554 32564
rect 32674 32552 32680 32564
rect 32548 32524 32680 32552
rect 32548 32512 32554 32524
rect 32674 32512 32680 32524
rect 32732 32512 32738 32564
rect 32950 32512 32956 32564
rect 33008 32552 33014 32564
rect 34238 32552 34244 32564
rect 33008 32524 34244 32552
rect 33008 32512 33014 32524
rect 34238 32512 34244 32524
rect 34296 32512 34302 32564
rect 37366 32552 37372 32564
rect 36648 32524 37372 32552
rect 22738 32484 22744 32496
rect 20640 32456 20944 32484
rect 21080 32456 22744 32484
rect 18969 32419 19027 32425
rect 18969 32385 18981 32419
rect 19015 32416 19027 32419
rect 19058 32416 19064 32428
rect 19015 32388 19064 32416
rect 19015 32385 19027 32388
rect 18969 32379 19027 32385
rect 19058 32376 19064 32388
rect 19116 32376 19122 32428
rect 19150 32376 19156 32428
rect 19208 32376 19214 32428
rect 20898 32376 20904 32428
rect 20956 32376 20962 32428
rect 21080 32425 21108 32456
rect 22738 32444 22744 32456
rect 22796 32444 22802 32496
rect 25501 32487 25559 32493
rect 25501 32484 25513 32487
rect 24872 32456 25513 32484
rect 21080 32419 21143 32425
rect 21080 32392 21097 32419
rect 21085 32385 21097 32392
rect 21131 32385 21143 32419
rect 21085 32379 21143 32385
rect 21177 32419 21235 32425
rect 21177 32385 21189 32419
rect 21223 32385 21235 32419
rect 21453 32419 21511 32425
rect 21453 32416 21465 32419
rect 21177 32379 21235 32385
rect 21284 32388 21465 32416
rect 19886 32348 19892 32360
rect 18831 32320 18920 32348
rect 18984 32320 19892 32348
rect 18831 32317 18843 32320
rect 18785 32311 18843 32317
rect 18984 32280 19012 32320
rect 19886 32308 19892 32320
rect 19944 32308 19950 32360
rect 19978 32308 19984 32360
rect 20036 32357 20042 32360
rect 20036 32351 20064 32357
rect 20052 32317 20064 32351
rect 20036 32311 20064 32317
rect 20036 32308 20042 32311
rect 20162 32308 20168 32360
rect 20220 32308 20226 32360
rect 20714 32308 20720 32360
rect 20772 32348 20778 32360
rect 21192 32348 21220 32379
rect 20772 32320 21220 32348
rect 20772 32308 20778 32320
rect 18708 32252 19012 32280
rect 19613 32283 19671 32289
rect 19613 32249 19625 32283
rect 19659 32280 19671 32283
rect 19702 32280 19708 32292
rect 19659 32252 19708 32280
rect 19659 32249 19671 32252
rect 19613 32243 19671 32249
rect 19702 32240 19708 32252
rect 19760 32240 19766 32292
rect 20806 32240 20812 32292
rect 20864 32280 20870 32292
rect 21284 32280 21312 32388
rect 21453 32385 21465 32388
rect 21499 32385 21511 32419
rect 21453 32379 21511 32385
rect 22186 32376 22192 32428
rect 22244 32376 22250 32428
rect 23569 32419 23627 32425
rect 23569 32385 23581 32419
rect 23615 32416 23627 32419
rect 24872 32416 24900 32456
rect 25501 32453 25513 32456
rect 25547 32484 25559 32487
rect 26786 32484 26792 32496
rect 25547 32456 26792 32484
rect 25547 32453 25559 32456
rect 25501 32447 25559 32453
rect 26786 32444 26792 32456
rect 26844 32444 26850 32496
rect 29196 32484 29224 32512
rect 29546 32484 29552 32496
rect 28920 32456 29552 32484
rect 23615 32388 24900 32416
rect 23615 32385 23627 32388
rect 23569 32379 23627 32385
rect 24670 32308 24676 32360
rect 24728 32348 24734 32360
rect 24872 32348 24900 32388
rect 24949 32419 25007 32425
rect 24949 32385 24961 32419
rect 24995 32416 25007 32419
rect 26326 32416 26332 32428
rect 24995 32388 25084 32416
rect 24995 32385 25007 32388
rect 24949 32379 25007 32385
rect 24728 32320 24900 32348
rect 24728 32308 24734 32320
rect 20864 32252 21312 32280
rect 20864 32240 20870 32252
rect 21450 32240 21456 32292
rect 21508 32280 21514 32292
rect 25056 32289 25084 32388
rect 25700 32388 26332 32416
rect 25700 32357 25728 32388
rect 26326 32376 26332 32388
rect 26384 32416 26390 32428
rect 26694 32416 26700 32428
rect 26384 32388 26700 32416
rect 26384 32376 26390 32388
rect 26694 32376 26700 32388
rect 26752 32376 26758 32428
rect 27982 32376 27988 32428
rect 28040 32425 28046 32428
rect 28920 32425 28948 32456
rect 29546 32444 29552 32456
rect 29604 32444 29610 32496
rect 36648 32493 36676 32524
rect 37366 32512 37372 32524
rect 37424 32512 37430 32564
rect 42058 32552 42064 32564
rect 41800 32524 42064 32552
rect 32585 32487 32643 32493
rect 32585 32484 32597 32487
rect 30852 32456 32597 32484
rect 29178 32425 29184 32428
rect 28040 32419 28068 32425
rect 28056 32385 28068 32419
rect 28040 32379 28068 32385
rect 28905 32419 28963 32425
rect 28905 32385 28917 32419
rect 28951 32385 28963 32419
rect 28905 32379 28963 32385
rect 29172 32379 29184 32425
rect 28040 32376 28046 32379
rect 29178 32376 29184 32379
rect 29236 32376 29242 32428
rect 25685 32351 25743 32357
rect 25685 32317 25697 32351
rect 25731 32317 25743 32351
rect 25685 32311 25743 32317
rect 25041 32283 25099 32289
rect 21508 32252 24532 32280
rect 21508 32240 21514 32252
rect 16448 32184 16620 32212
rect 16448 32172 16454 32184
rect 18138 32172 18144 32224
rect 18196 32172 18202 32224
rect 18874 32172 18880 32224
rect 18932 32212 18938 32224
rect 19242 32212 19248 32224
rect 18932 32184 19248 32212
rect 18932 32172 18938 32184
rect 19242 32172 19248 32184
rect 19300 32172 19306 32224
rect 20346 32172 20352 32224
rect 20404 32212 20410 32224
rect 20898 32212 20904 32224
rect 20404 32184 20904 32212
rect 20404 32172 20410 32184
rect 20898 32172 20904 32184
rect 20956 32172 20962 32224
rect 21358 32172 21364 32224
rect 21416 32172 21422 32224
rect 22005 32215 22063 32221
rect 22005 32181 22017 32215
rect 22051 32212 22063 32215
rect 22094 32212 22100 32224
rect 22051 32184 22100 32212
rect 22051 32181 22063 32184
rect 22005 32175 22063 32181
rect 22094 32172 22100 32184
rect 22152 32172 22158 32224
rect 22462 32172 22468 32224
rect 22520 32212 22526 32224
rect 23661 32215 23719 32221
rect 23661 32212 23673 32215
rect 22520 32184 23673 32212
rect 22520 32172 22526 32184
rect 23661 32181 23673 32184
rect 23707 32181 23719 32215
rect 24504 32212 24532 32252
rect 25041 32249 25053 32283
rect 25087 32249 25099 32283
rect 25041 32243 25099 32249
rect 25700 32212 25728 32311
rect 26602 32308 26608 32360
rect 26660 32348 26666 32360
rect 26973 32351 27031 32357
rect 26973 32348 26985 32351
rect 26660 32320 26985 32348
rect 26660 32308 26666 32320
rect 26973 32317 26985 32320
rect 27019 32317 27031 32351
rect 26973 32311 27031 32317
rect 27154 32308 27160 32360
rect 27212 32308 27218 32360
rect 27522 32308 27528 32360
rect 27580 32348 27586 32360
rect 27893 32351 27951 32357
rect 27893 32348 27905 32351
rect 27580 32320 27905 32348
rect 27580 32308 27586 32320
rect 27893 32317 27905 32320
rect 27939 32317 27951 32351
rect 27893 32311 27951 32317
rect 28166 32308 28172 32360
rect 28224 32308 28230 32360
rect 30650 32308 30656 32360
rect 30708 32348 30714 32360
rect 30852 32357 30880 32456
rect 32585 32453 32597 32456
rect 32631 32453 32643 32487
rect 32585 32447 32643 32453
rect 36633 32487 36691 32493
rect 36633 32453 36645 32487
rect 36679 32453 36691 32487
rect 38010 32484 38016 32496
rect 36633 32447 36691 32453
rect 37384 32456 38016 32484
rect 37384 32425 37412 32456
rect 38010 32444 38016 32456
rect 38068 32444 38074 32496
rect 40773 32487 40831 32493
rect 40773 32453 40785 32487
rect 40819 32484 40831 32487
rect 40819 32456 41276 32484
rect 40819 32453 40831 32456
rect 40773 32447 40831 32453
rect 41248 32428 41276 32456
rect 37369 32419 37427 32425
rect 37369 32385 37381 32419
rect 37415 32385 37427 32419
rect 37645 32419 37703 32425
rect 37645 32416 37657 32419
rect 37369 32379 37427 32385
rect 37476 32388 37657 32416
rect 30837 32351 30895 32357
rect 30837 32348 30849 32351
rect 30708 32320 30849 32348
rect 30708 32308 30714 32320
rect 30837 32317 30849 32320
rect 30883 32317 30895 32351
rect 30837 32311 30895 32317
rect 31018 32308 31024 32360
rect 31076 32308 31082 32360
rect 32674 32308 32680 32360
rect 32732 32308 32738 32360
rect 35342 32308 35348 32360
rect 35400 32348 35406 32360
rect 35400 32320 37044 32348
rect 35400 32308 35406 32320
rect 27614 32240 27620 32292
rect 27672 32240 27678 32292
rect 28552 32252 28948 32280
rect 24504 32184 25728 32212
rect 23661 32175 23719 32181
rect 27154 32172 27160 32224
rect 27212 32212 27218 32224
rect 28552 32212 28580 32252
rect 27212 32184 28580 32212
rect 27212 32172 27218 32184
rect 28626 32172 28632 32224
rect 28684 32212 28690 32224
rect 28813 32215 28871 32221
rect 28813 32212 28825 32215
rect 28684 32184 28825 32212
rect 28684 32172 28690 32184
rect 28813 32181 28825 32184
rect 28859 32181 28871 32215
rect 28920 32212 28948 32252
rect 30190 32240 30196 32292
rect 30248 32280 30254 32292
rect 31036 32280 31064 32308
rect 30248 32252 31064 32280
rect 30248 32240 30254 32252
rect 36814 32240 36820 32292
rect 36872 32280 36878 32292
rect 36909 32283 36967 32289
rect 36909 32280 36921 32283
rect 36872 32252 36921 32280
rect 36872 32240 36878 32252
rect 36909 32249 36921 32252
rect 36955 32249 36967 32283
rect 37016 32280 37044 32320
rect 37090 32308 37096 32360
rect 37148 32348 37154 32360
rect 37476 32348 37504 32388
rect 37645 32385 37657 32388
rect 37691 32385 37703 32419
rect 37645 32379 37703 32385
rect 40405 32419 40463 32425
rect 40405 32385 40417 32419
rect 40451 32416 40463 32419
rect 40494 32416 40500 32428
rect 40451 32388 40500 32416
rect 40451 32385 40463 32388
rect 40405 32379 40463 32385
rect 40494 32376 40500 32388
rect 40552 32416 40558 32428
rect 40681 32419 40739 32425
rect 40681 32416 40693 32419
rect 40552 32388 40693 32416
rect 40552 32376 40558 32388
rect 40681 32385 40693 32388
rect 40727 32385 40739 32419
rect 40681 32379 40739 32385
rect 40865 32419 40923 32425
rect 40865 32385 40877 32419
rect 40911 32385 40923 32419
rect 40865 32379 40923 32385
rect 37148 32320 37504 32348
rect 37148 32308 37154 32320
rect 37550 32308 37556 32360
rect 37608 32308 37614 32360
rect 40218 32308 40224 32360
rect 40276 32348 40282 32360
rect 40770 32348 40776 32360
rect 40276 32320 40776 32348
rect 40276 32308 40282 32320
rect 40770 32308 40776 32320
rect 40828 32348 40834 32360
rect 40880 32348 40908 32379
rect 41230 32376 41236 32428
rect 41288 32376 41294 32428
rect 41429 32419 41487 32425
rect 41429 32385 41441 32419
rect 41475 32416 41487 32419
rect 41800 32416 41828 32524
rect 42058 32512 42064 32524
rect 42116 32512 42122 32564
rect 42426 32512 42432 32564
rect 42484 32512 42490 32564
rect 43898 32512 43904 32564
rect 43956 32552 43962 32564
rect 44821 32555 44879 32561
rect 44821 32552 44833 32555
rect 43956 32524 44833 32552
rect 43956 32512 43962 32524
rect 44821 32521 44833 32524
rect 44867 32521 44879 32555
rect 44821 32515 44879 32521
rect 45462 32512 45468 32564
rect 45520 32552 45526 32564
rect 45520 32524 46060 32552
rect 45520 32512 45526 32524
rect 42702 32484 42708 32496
rect 41892 32456 42708 32484
rect 41892 32425 41920 32456
rect 42702 32444 42708 32456
rect 42760 32444 42766 32496
rect 43162 32444 43168 32496
rect 43220 32444 43226 32496
rect 44174 32444 44180 32496
rect 44232 32484 44238 32496
rect 44453 32487 44511 32493
rect 44453 32484 44465 32487
rect 44232 32456 44465 32484
rect 44232 32444 44238 32456
rect 44453 32453 44465 32456
rect 44499 32453 44511 32487
rect 44453 32447 44511 32453
rect 44910 32444 44916 32496
rect 44968 32484 44974 32496
rect 44968 32456 45508 32484
rect 44968 32444 44974 32456
rect 41475 32388 41828 32416
rect 41877 32419 41935 32425
rect 41475 32385 41487 32388
rect 41429 32379 41487 32385
rect 41877 32385 41889 32419
rect 41923 32385 41935 32419
rect 41877 32379 41935 32385
rect 40828 32320 40908 32348
rect 40828 32308 40834 32320
rect 38562 32280 38568 32292
rect 37016 32252 38568 32280
rect 36909 32243 36967 32249
rect 38562 32240 38568 32252
rect 38620 32240 38626 32292
rect 40589 32283 40647 32289
rect 40589 32249 40601 32283
rect 40635 32280 40647 32283
rect 41322 32280 41328 32292
rect 40635 32252 41328 32280
rect 40635 32249 40647 32252
rect 40589 32243 40647 32249
rect 41322 32240 41328 32252
rect 41380 32280 41386 32292
rect 41432 32280 41460 32379
rect 42150 32376 42156 32428
rect 42208 32376 42214 32428
rect 42610 32376 42616 32428
rect 42668 32416 42674 32428
rect 42797 32419 42855 32425
rect 42797 32416 42809 32419
rect 42668 32388 42809 32416
rect 42668 32376 42674 32388
rect 42797 32385 42809 32388
rect 42843 32385 42855 32419
rect 42797 32379 42855 32385
rect 43349 32419 43407 32425
rect 43349 32385 43361 32419
rect 43395 32385 43407 32419
rect 43349 32379 43407 32385
rect 41969 32351 42027 32357
rect 41969 32317 41981 32351
rect 42015 32348 42027 32351
rect 42334 32348 42340 32360
rect 42015 32320 42340 32348
rect 42015 32317 42027 32320
rect 41969 32311 42027 32317
rect 42334 32308 42340 32320
rect 42392 32308 42398 32360
rect 42886 32308 42892 32360
rect 42944 32348 42950 32360
rect 43364 32348 43392 32379
rect 43438 32376 43444 32428
rect 43496 32376 43502 32428
rect 44085 32419 44143 32425
rect 44085 32385 44097 32419
rect 44131 32416 44143 32419
rect 44358 32416 44364 32428
rect 44131 32388 44364 32416
rect 44131 32385 44143 32388
rect 44085 32379 44143 32385
rect 44358 32376 44364 32388
rect 44416 32376 44422 32428
rect 44545 32419 44603 32425
rect 44545 32385 44557 32419
rect 44591 32416 44603 32419
rect 44591 32388 44956 32416
rect 44591 32385 44603 32388
rect 44545 32379 44603 32385
rect 44269 32351 44327 32357
rect 42944 32320 44128 32348
rect 42944 32308 42950 32320
rect 41380 32252 41460 32280
rect 42061 32283 42119 32289
rect 41380 32240 41386 32252
rect 42061 32249 42073 32283
rect 42107 32280 42119 32283
rect 42904 32280 42932 32308
rect 44100 32289 44128 32320
rect 44269 32317 44281 32351
rect 44315 32348 44327 32351
rect 44634 32348 44640 32360
rect 44315 32320 44640 32348
rect 44315 32317 44327 32320
rect 44269 32311 44327 32317
rect 44634 32308 44640 32320
rect 44692 32308 44698 32360
rect 44818 32308 44824 32360
rect 44876 32308 44882 32360
rect 44928 32348 44956 32388
rect 45002 32376 45008 32428
rect 45060 32376 45066 32428
rect 45480 32425 45508 32456
rect 46032 32425 46060 32524
rect 45465 32419 45523 32425
rect 45465 32385 45477 32419
rect 45511 32385 45523 32419
rect 45465 32379 45523 32385
rect 46017 32419 46075 32425
rect 46017 32385 46029 32419
rect 46063 32385 46075 32419
rect 46017 32379 46075 32385
rect 46201 32419 46259 32425
rect 46201 32385 46213 32419
rect 46247 32385 46259 32419
rect 46201 32379 46259 32385
rect 45925 32351 45983 32357
rect 44928 32320 45140 32348
rect 43165 32283 43223 32289
rect 43165 32280 43177 32283
rect 42107 32252 42932 32280
rect 42996 32252 43177 32280
rect 42107 32249 42119 32252
rect 42061 32243 42119 32249
rect 29638 32212 29644 32224
rect 28920 32184 29644 32212
rect 28813 32175 28871 32181
rect 29638 32172 29644 32184
rect 29696 32212 29702 32224
rect 30285 32215 30343 32221
rect 30285 32212 30297 32215
rect 29696 32184 30297 32212
rect 29696 32172 29702 32184
rect 30285 32181 30297 32184
rect 30331 32181 30343 32215
rect 30285 32175 30343 32181
rect 36538 32172 36544 32224
rect 36596 32212 36602 32224
rect 37093 32215 37151 32221
rect 37093 32212 37105 32215
rect 36596 32184 37105 32212
rect 36596 32172 36602 32184
rect 37093 32181 37105 32184
rect 37139 32181 37151 32215
rect 37093 32175 37151 32181
rect 37642 32172 37648 32224
rect 37700 32172 37706 32224
rect 37829 32215 37887 32221
rect 37829 32181 37841 32215
rect 37875 32212 37887 32215
rect 38470 32212 38476 32224
rect 37875 32184 38476 32212
rect 37875 32181 37887 32184
rect 37829 32175 37887 32181
rect 38470 32172 38476 32184
rect 38528 32172 38534 32224
rect 41233 32215 41291 32221
rect 41233 32181 41245 32215
rect 41279 32212 41291 32215
rect 41506 32212 41512 32224
rect 41279 32184 41512 32212
rect 41279 32181 41291 32184
rect 41233 32175 41291 32181
rect 41506 32172 41512 32184
rect 41564 32172 41570 32224
rect 41598 32172 41604 32224
rect 41656 32212 41662 32224
rect 41693 32215 41751 32221
rect 41693 32212 41705 32215
rect 41656 32184 41705 32212
rect 41656 32172 41662 32184
rect 41693 32181 41705 32184
rect 41739 32181 41751 32215
rect 41693 32175 41751 32181
rect 42518 32172 42524 32224
rect 42576 32212 42582 32224
rect 42996 32212 43024 32252
rect 43165 32249 43177 32252
rect 43211 32249 43223 32283
rect 43165 32243 43223 32249
rect 44085 32283 44143 32289
rect 44085 32249 44097 32283
rect 44131 32249 44143 32283
rect 44085 32243 44143 32249
rect 45112 32224 45140 32320
rect 45925 32317 45937 32351
rect 45971 32348 45983 32351
rect 46216 32348 46244 32379
rect 45971 32320 46244 32348
rect 45971 32317 45983 32320
rect 45925 32311 45983 32317
rect 45370 32240 45376 32292
rect 45428 32280 45434 32292
rect 46109 32283 46167 32289
rect 46109 32280 46121 32283
rect 45428 32252 46121 32280
rect 45428 32240 45434 32252
rect 46109 32249 46121 32252
rect 46155 32249 46167 32283
rect 46109 32243 46167 32249
rect 42576 32184 43024 32212
rect 42576 32172 42582 32184
rect 43070 32172 43076 32224
rect 43128 32172 43134 32224
rect 45094 32172 45100 32224
rect 45152 32212 45158 32224
rect 45557 32215 45615 32221
rect 45557 32212 45569 32215
rect 45152 32184 45569 32212
rect 45152 32172 45158 32184
rect 45557 32181 45569 32184
rect 45603 32181 45615 32215
rect 45557 32175 45615 32181
rect 1104 32122 47104 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 47104 32122
rect 1104 32048 47104 32070
rect 3694 31968 3700 32020
rect 3752 32008 3758 32020
rect 6270 32008 6276 32020
rect 3752 31980 6276 32008
rect 3752 31968 3758 31980
rect 6270 31968 6276 31980
rect 6328 32008 6334 32020
rect 7558 32008 7564 32020
rect 6328 31980 7564 32008
rect 6328 31968 6334 31980
rect 7558 31968 7564 31980
rect 7616 31968 7622 32020
rect 7745 32011 7803 32017
rect 7745 31977 7757 32011
rect 7791 32008 7803 32011
rect 8202 32008 8208 32020
rect 7791 31980 8208 32008
rect 7791 31977 7803 31980
rect 7745 31971 7803 31977
rect 8202 31968 8208 31980
rect 8260 31968 8266 32020
rect 8938 31968 8944 32020
rect 8996 31968 9002 32020
rect 12526 32008 12532 32020
rect 9876 31980 12532 32008
rect 4706 31900 4712 31952
rect 4764 31940 4770 31952
rect 5258 31940 5264 31952
rect 4764 31912 5264 31940
rect 4764 31900 4770 31912
rect 5258 31900 5264 31912
rect 5316 31900 5322 31952
rect 8021 31943 8079 31949
rect 8021 31909 8033 31943
rect 8067 31909 8079 31943
rect 8021 31903 8079 31909
rect 934 31832 940 31884
rect 992 31872 998 31884
rect 1397 31875 1455 31881
rect 1397 31872 1409 31875
rect 992 31844 1409 31872
rect 992 31832 998 31844
rect 1397 31841 1409 31844
rect 1443 31841 1455 31875
rect 1397 31835 1455 31841
rect 1670 31832 1676 31884
rect 1728 31832 1734 31884
rect 6362 31832 6368 31884
rect 6420 31832 6426 31884
rect 4706 31764 4712 31816
rect 4764 31804 4770 31816
rect 5350 31804 5356 31816
rect 4764 31776 5356 31804
rect 4764 31764 4770 31776
rect 5350 31764 5356 31776
rect 5408 31764 5414 31816
rect 6638 31813 6644 31816
rect 6632 31804 6644 31813
rect 6599 31776 6644 31804
rect 6632 31767 6644 31776
rect 6638 31764 6644 31767
rect 6696 31764 6702 31816
rect 8036 31804 8064 31903
rect 9582 31900 9588 31952
rect 9640 31940 9646 31952
rect 9876 31949 9904 31980
rect 12526 31968 12532 31980
rect 12584 31968 12590 32020
rect 12802 31968 12808 32020
rect 12860 32008 12866 32020
rect 13630 32008 13636 32020
rect 12860 31980 13636 32008
rect 12860 31968 12866 31980
rect 13630 31968 13636 31980
rect 13688 31968 13694 32020
rect 13906 31968 13912 32020
rect 13964 32008 13970 32020
rect 13964 31980 14136 32008
rect 13964 31968 13970 31980
rect 9861 31943 9919 31949
rect 9861 31940 9873 31943
rect 9640 31912 9873 31940
rect 9640 31900 9646 31912
rect 9861 31909 9873 31912
rect 9907 31909 9919 31943
rect 9861 31903 9919 31909
rect 11057 31943 11115 31949
rect 11057 31909 11069 31943
rect 11103 31940 11115 31943
rect 13998 31940 14004 31952
rect 11103 31912 14004 31940
rect 11103 31909 11115 31912
rect 11057 31903 11115 31909
rect 13998 31900 14004 31912
rect 14056 31900 14062 31952
rect 14108 31940 14136 31980
rect 14182 31968 14188 32020
rect 14240 32008 14246 32020
rect 17773 32011 17831 32017
rect 14240 31980 15332 32008
rect 14240 31968 14246 31980
rect 15304 31952 15332 31980
rect 17773 31977 17785 32011
rect 17819 32008 17831 32011
rect 18506 32008 18512 32020
rect 17819 31980 18512 32008
rect 17819 31977 17831 31980
rect 17773 31971 17831 31977
rect 18506 31968 18512 31980
rect 18564 32008 18570 32020
rect 19978 32008 19984 32020
rect 18564 31980 19984 32008
rect 18564 31968 18570 31980
rect 19978 31968 19984 31980
rect 20036 32008 20042 32020
rect 20254 32008 20260 32020
rect 20036 31980 20260 32008
rect 20036 31968 20042 31980
rect 20254 31968 20260 31980
rect 20312 31968 20318 32020
rect 20346 31968 20352 32020
rect 20404 32008 20410 32020
rect 21358 32008 21364 32020
rect 20404 31980 21364 32008
rect 20404 31968 20410 31980
rect 21358 31968 21364 31980
rect 21416 31968 21422 32020
rect 21726 31968 21732 32020
rect 21784 31968 21790 32020
rect 22002 32008 22008 32020
rect 21836 31980 22008 32008
rect 14108 31912 14228 31940
rect 8662 31832 8668 31884
rect 8720 31832 8726 31884
rect 9214 31832 9220 31884
rect 9272 31832 9278 31884
rect 9401 31875 9459 31881
rect 9401 31841 9413 31875
rect 9447 31872 9459 31875
rect 9766 31872 9772 31884
rect 9447 31844 9772 31872
rect 9447 31841 9459 31844
rect 9401 31835 9459 31841
rect 9766 31832 9772 31844
rect 9824 31832 9830 31884
rect 9950 31832 9956 31884
rect 10008 31872 10014 31884
rect 10137 31875 10195 31881
rect 10137 31872 10149 31875
rect 10008 31844 10149 31872
rect 10008 31832 10014 31844
rect 10137 31841 10149 31844
rect 10183 31841 10195 31875
rect 10137 31835 10195 31841
rect 10275 31875 10333 31881
rect 10275 31841 10287 31875
rect 10321 31872 10333 31875
rect 10594 31872 10600 31884
rect 10321 31844 10600 31872
rect 10321 31841 10333 31844
rect 10275 31835 10333 31841
rect 10594 31832 10600 31844
rect 10652 31832 10658 31884
rect 11330 31832 11336 31884
rect 11388 31872 11394 31884
rect 12253 31875 12311 31881
rect 12253 31872 12265 31875
rect 11388 31844 12265 31872
rect 11388 31832 11394 31844
rect 12253 31841 12265 31844
rect 12299 31841 12311 31875
rect 12253 31835 12311 31841
rect 12345 31875 12403 31881
rect 12345 31841 12357 31875
rect 12391 31872 12403 31875
rect 12391 31844 12480 31872
rect 12391 31841 12403 31844
rect 12345 31835 12403 31841
rect 9125 31807 9183 31813
rect 9125 31804 9137 31807
rect 8036 31776 9137 31804
rect 9125 31773 9137 31776
rect 9171 31773 9183 31807
rect 9125 31767 9183 31773
rect 8389 31739 8447 31745
rect 8389 31705 8401 31739
rect 8435 31736 8447 31739
rect 9232 31736 9260 31832
rect 10410 31764 10416 31816
rect 10468 31764 10474 31816
rect 12452 31804 12480 31844
rect 12526 31832 12532 31884
rect 12584 31832 12590 31884
rect 13081 31875 13139 31881
rect 13081 31841 13093 31875
rect 13127 31872 13139 31875
rect 13170 31872 13176 31884
rect 13127 31844 13176 31872
rect 13127 31841 13139 31844
rect 13081 31835 13139 31841
rect 13170 31832 13176 31844
rect 13228 31832 13234 31884
rect 13262 31832 13268 31884
rect 13320 31832 13326 31884
rect 14200 31881 14228 31912
rect 15286 31900 15292 31952
rect 15344 31940 15350 31952
rect 15565 31943 15623 31949
rect 15565 31940 15577 31943
rect 15344 31912 15577 31940
rect 15344 31900 15350 31912
rect 15565 31909 15577 31912
rect 15611 31909 15623 31943
rect 15565 31903 15623 31909
rect 19150 31900 19156 31952
rect 19208 31940 19214 31952
rect 19208 31912 19472 31940
rect 19208 31900 19214 31912
rect 14185 31875 14243 31881
rect 14185 31841 14197 31875
rect 14231 31841 14243 31875
rect 14185 31835 14243 31841
rect 16390 31832 16396 31884
rect 16448 31832 16454 31884
rect 19058 31832 19064 31884
rect 19116 31872 19122 31884
rect 19444 31881 19472 31912
rect 21082 31900 21088 31952
rect 21140 31940 21146 31952
rect 21450 31940 21456 31952
rect 21140 31912 21456 31940
rect 21140 31900 21146 31912
rect 21450 31900 21456 31912
rect 21508 31900 21514 31952
rect 19245 31875 19303 31881
rect 19245 31872 19257 31875
rect 19116 31844 19257 31872
rect 19116 31832 19122 31844
rect 19245 31841 19257 31844
rect 19291 31841 19303 31875
rect 19245 31835 19303 31841
rect 19429 31875 19487 31881
rect 19429 31841 19441 31875
rect 19475 31841 19487 31875
rect 19429 31835 19487 31841
rect 19518 31832 19524 31884
rect 19576 31872 19582 31884
rect 19889 31875 19947 31881
rect 19889 31872 19901 31875
rect 19576 31844 19901 31872
rect 19576 31832 19582 31844
rect 19889 31841 19901 31844
rect 19935 31841 19947 31875
rect 19889 31835 19947 31841
rect 20162 31832 20168 31884
rect 20220 31832 20226 31884
rect 20254 31832 20260 31884
rect 20312 31881 20318 31884
rect 20312 31875 20340 31881
rect 20328 31841 20340 31875
rect 20312 31835 20340 31841
rect 21008 31844 21496 31872
rect 20312 31832 20318 31835
rect 12802 31804 12808 31816
rect 12452 31776 12808 31804
rect 12802 31764 12808 31776
rect 12860 31764 12866 31816
rect 12989 31807 13047 31813
rect 12989 31773 13001 31807
rect 13035 31782 13047 31807
rect 13354 31804 13360 31816
rect 13096 31782 13360 31804
rect 13035 31776 13360 31782
rect 13035 31773 13124 31776
rect 12989 31767 13124 31773
rect 13004 31754 13124 31767
rect 13354 31764 13360 31776
rect 13412 31764 13418 31816
rect 14274 31764 14280 31816
rect 14332 31804 14338 31816
rect 14441 31807 14499 31813
rect 14441 31804 14453 31807
rect 14332 31776 14453 31804
rect 14332 31764 14338 31776
rect 14441 31773 14453 31776
rect 14487 31773 14499 31807
rect 14441 31767 14499 31773
rect 15930 31764 15936 31816
rect 15988 31764 15994 31816
rect 16022 31764 16028 31816
rect 16080 31804 16086 31816
rect 16649 31807 16707 31813
rect 16649 31804 16661 31807
rect 16080 31776 16661 31804
rect 16080 31764 16086 31776
rect 16649 31773 16661 31776
rect 16695 31773 16707 31807
rect 16649 31767 16707 31773
rect 20438 31764 20444 31816
rect 20496 31764 20502 31816
rect 8435 31708 9260 31736
rect 8435 31705 8447 31708
rect 8389 31699 8447 31705
rect 11514 31696 11520 31748
rect 11572 31736 11578 31748
rect 11885 31739 11943 31745
rect 11885 31736 11897 31739
rect 11572 31708 11897 31736
rect 11572 31696 11578 31708
rect 11885 31705 11897 31708
rect 11931 31705 11943 31739
rect 11885 31699 11943 31705
rect 15746 31696 15752 31748
rect 15804 31736 15810 31748
rect 21008 31736 21036 31844
rect 21174 31764 21180 31816
rect 21232 31804 21238 31816
rect 21361 31807 21419 31813
rect 21361 31804 21373 31807
rect 21232 31776 21373 31804
rect 21232 31764 21238 31776
rect 21361 31773 21373 31776
rect 21407 31773 21419 31807
rect 21361 31767 21419 31773
rect 15804 31708 16160 31736
rect 15804 31696 15810 31708
rect 8478 31628 8484 31680
rect 8536 31668 8542 31680
rect 10134 31668 10140 31680
rect 8536 31640 10140 31668
rect 8536 31628 8542 31640
rect 10134 31628 10140 31640
rect 10192 31628 10198 31680
rect 11606 31628 11612 31680
rect 11664 31668 11670 31680
rect 12621 31671 12679 31677
rect 12621 31668 12633 31671
rect 11664 31640 12633 31668
rect 11664 31628 11670 31640
rect 12621 31637 12633 31640
rect 12667 31637 12679 31671
rect 12621 31631 12679 31637
rect 16022 31628 16028 31680
rect 16080 31628 16086 31680
rect 16132 31668 16160 31708
rect 20916 31708 21036 31736
rect 20916 31668 20944 31708
rect 16132 31640 20944 31668
rect 20990 31628 20996 31680
rect 21048 31668 21054 31680
rect 21085 31671 21143 31677
rect 21085 31668 21097 31671
rect 21048 31640 21097 31668
rect 21048 31628 21054 31640
rect 21085 31637 21097 31640
rect 21131 31637 21143 31671
rect 21085 31631 21143 31637
rect 21174 31628 21180 31680
rect 21232 31628 21238 31680
rect 21376 31668 21404 31767
rect 21468 31736 21496 31844
rect 21744 31816 21772 31968
rect 21836 31881 21864 31980
rect 22002 31968 22008 31980
rect 22060 32008 22066 32020
rect 22060 31980 22784 32008
rect 22060 31968 22066 31980
rect 22756 31940 22784 31980
rect 23198 31968 23204 32020
rect 23256 32008 23262 32020
rect 28166 32008 28172 32020
rect 23256 31980 28172 32008
rect 23256 31968 23262 31980
rect 28166 31968 28172 31980
rect 28224 31968 28230 32020
rect 29178 31968 29184 32020
rect 29236 31968 29242 32020
rect 30650 32008 30656 32020
rect 29564 31980 30656 32008
rect 22830 31940 22836 31952
rect 22756 31912 22836 31940
rect 22830 31900 22836 31912
rect 22888 31900 22894 31952
rect 27249 31943 27307 31949
rect 27249 31909 27261 31943
rect 27295 31940 27307 31943
rect 27338 31940 27344 31952
rect 27295 31912 27344 31940
rect 27295 31909 27307 31912
rect 27249 31903 27307 31909
rect 27338 31900 27344 31912
rect 27396 31900 27402 31952
rect 28445 31943 28503 31949
rect 28445 31909 28457 31943
rect 28491 31940 28503 31943
rect 28813 31943 28871 31949
rect 28813 31940 28825 31943
rect 28491 31912 28825 31940
rect 28491 31909 28503 31912
rect 28445 31903 28503 31909
rect 28813 31909 28825 31912
rect 28859 31909 28871 31943
rect 28813 31903 28871 31909
rect 28902 31900 28908 31952
rect 28960 31940 28966 31952
rect 29564 31940 29592 31980
rect 30650 31968 30656 31980
rect 30708 31968 30714 32020
rect 30742 31968 30748 32020
rect 30800 32008 30806 32020
rect 30929 32011 30987 32017
rect 30929 32008 30941 32011
rect 30800 31980 30941 32008
rect 30800 31968 30806 31980
rect 30929 31977 30941 31980
rect 30975 31977 30987 32011
rect 30929 31971 30987 31977
rect 31018 31968 31024 32020
rect 31076 32008 31082 32020
rect 36817 32011 36875 32017
rect 31076 31980 36492 32008
rect 31076 31968 31082 31980
rect 28960 31912 29592 31940
rect 30668 31940 30696 31968
rect 31294 31949 31300 31952
rect 31251 31943 31300 31949
rect 31251 31940 31263 31943
rect 30668 31912 31263 31940
rect 28960 31900 28966 31912
rect 31251 31909 31263 31912
rect 31297 31909 31300 31943
rect 31251 31903 31300 31909
rect 31294 31900 31300 31903
rect 31352 31900 31358 31952
rect 32030 31900 32036 31952
rect 32088 31940 32094 31952
rect 35345 31943 35403 31949
rect 35345 31940 35357 31943
rect 32088 31912 35357 31940
rect 32088 31900 32094 31912
rect 35345 31909 35357 31912
rect 35391 31909 35403 31943
rect 36464 31940 36492 31980
rect 36817 31977 36829 32011
rect 36863 32008 36875 32011
rect 37550 32008 37556 32020
rect 36863 31980 37556 32008
rect 36863 31977 36875 31980
rect 36817 31971 36875 31977
rect 37550 31968 37556 31980
rect 37608 32008 37614 32020
rect 41966 32008 41972 32020
rect 37608 31980 41972 32008
rect 37608 31968 37614 31980
rect 38657 31943 38715 31949
rect 36464 31912 37596 31940
rect 35345 31903 35403 31909
rect 21821 31875 21879 31881
rect 21821 31841 21833 31875
rect 21867 31841 21879 31875
rect 21821 31835 21879 31841
rect 26602 31832 26608 31884
rect 26660 31832 26666 31884
rect 26789 31875 26847 31881
rect 26789 31841 26801 31875
rect 26835 31872 26847 31875
rect 27154 31872 27160 31884
rect 26835 31844 27160 31872
rect 26835 31841 26847 31844
rect 26789 31835 26847 31841
rect 27154 31832 27160 31844
rect 27212 31832 27218 31884
rect 27522 31832 27528 31884
rect 27580 31832 27586 31884
rect 27663 31875 27721 31881
rect 27663 31841 27675 31875
rect 27709 31872 27721 31875
rect 27982 31872 27988 31884
rect 27709 31844 27988 31872
rect 27709 31841 27721 31844
rect 27663 31835 27721 31841
rect 27982 31832 27988 31844
rect 28040 31832 28046 31884
rect 28350 31832 28356 31884
rect 28408 31872 28414 31884
rect 28537 31875 28595 31881
rect 28537 31872 28549 31875
rect 28408 31844 28549 31872
rect 28408 31832 28414 31844
rect 28537 31841 28549 31844
rect 28583 31841 28595 31875
rect 28537 31835 28595 31841
rect 29270 31832 29276 31884
rect 29328 31872 29334 31884
rect 29328 31844 29684 31872
rect 29328 31832 29334 31844
rect 21542 31764 21548 31816
rect 21600 31764 21606 31816
rect 21634 31764 21640 31816
rect 21692 31764 21698 31816
rect 21726 31764 21732 31816
rect 21784 31764 21790 31816
rect 22094 31813 22100 31816
rect 22088 31767 22100 31813
rect 22094 31764 22100 31767
rect 22152 31764 22158 31816
rect 22370 31764 22376 31816
rect 22428 31804 22434 31816
rect 26694 31804 26700 31816
rect 22428 31776 26700 31804
rect 22428 31764 22434 31776
rect 26694 31764 26700 31776
rect 26752 31764 26758 31816
rect 27798 31764 27804 31816
rect 27856 31764 27862 31816
rect 29362 31764 29368 31816
rect 29420 31764 29426 31816
rect 29546 31764 29552 31816
rect 29604 31764 29610 31816
rect 29656 31804 29684 31844
rect 30834 31832 30840 31884
rect 30892 31872 30898 31884
rect 30892 31844 31754 31872
rect 30892 31832 30898 31844
rect 29805 31807 29863 31813
rect 29805 31804 29817 31807
rect 29656 31776 29817 31804
rect 29805 31773 29817 31776
rect 29851 31773 29863 31807
rect 29805 31767 29863 31773
rect 30374 31764 30380 31816
rect 30432 31804 30438 31816
rect 31021 31807 31079 31813
rect 31021 31804 31033 31807
rect 30432 31776 31033 31804
rect 30432 31764 30438 31776
rect 31021 31773 31033 31776
rect 31067 31804 31079 31807
rect 31478 31804 31484 31816
rect 31067 31776 31484 31804
rect 31067 31773 31079 31776
rect 31021 31767 31079 31773
rect 31478 31764 31484 31776
rect 31536 31764 31542 31816
rect 31726 31804 31754 31844
rect 34716 31844 35664 31872
rect 31846 31804 31852 31816
rect 31726 31776 31852 31804
rect 31846 31764 31852 31776
rect 31904 31764 31910 31816
rect 34149 31807 34207 31813
rect 34149 31773 34161 31807
rect 34195 31804 34207 31807
rect 34606 31804 34612 31816
rect 34195 31776 34612 31804
rect 34195 31773 34207 31776
rect 34149 31767 34207 31773
rect 34606 31764 34612 31776
rect 34664 31764 34670 31816
rect 34716 31813 34744 31844
rect 34882 31813 34888 31816
rect 34701 31807 34759 31813
rect 34701 31773 34713 31807
rect 34747 31773 34759 31807
rect 34701 31767 34759 31773
rect 34849 31807 34888 31813
rect 34849 31773 34861 31807
rect 34849 31767 34888 31773
rect 34882 31764 34888 31767
rect 34940 31764 34946 31816
rect 35250 31813 35256 31816
rect 35069 31807 35127 31813
rect 35069 31773 35081 31807
rect 35115 31804 35127 31807
rect 35207 31807 35256 31813
rect 35115 31776 35149 31804
rect 35115 31773 35127 31776
rect 35069 31767 35127 31773
rect 35207 31773 35219 31807
rect 35253 31773 35256 31807
rect 35207 31767 35256 31773
rect 34514 31736 34520 31748
rect 21468 31708 24716 31736
rect 21818 31668 21824 31680
rect 21376 31640 21824 31668
rect 21818 31628 21824 31640
rect 21876 31628 21882 31680
rect 22370 31628 22376 31680
rect 22428 31668 22434 31680
rect 23201 31671 23259 31677
rect 23201 31668 23213 31671
rect 22428 31640 23213 31668
rect 22428 31628 22434 31640
rect 23201 31637 23213 31640
rect 23247 31668 23259 31671
rect 24578 31668 24584 31680
rect 23247 31640 24584 31668
rect 23247 31637 23259 31640
rect 23201 31631 23259 31637
rect 24578 31628 24584 31640
rect 24636 31628 24642 31680
rect 24688 31668 24716 31708
rect 28276 31708 34520 31736
rect 28276 31668 28304 31708
rect 34514 31696 34520 31708
rect 34572 31696 34578 31748
rect 34977 31739 35035 31745
rect 34977 31705 34989 31739
rect 35023 31705 35035 31739
rect 35084 31736 35112 31767
rect 35250 31764 35256 31767
rect 35308 31764 35314 31816
rect 35342 31764 35348 31816
rect 35400 31764 35406 31816
rect 35636 31804 35664 31844
rect 35805 31807 35863 31813
rect 35636 31776 35756 31804
rect 35360 31736 35388 31764
rect 35084 31708 35388 31736
rect 35728 31736 35756 31776
rect 35805 31773 35817 31807
rect 35851 31804 35863 31807
rect 35986 31804 35992 31816
rect 35851 31776 35992 31804
rect 35851 31773 35863 31776
rect 35805 31767 35863 31773
rect 35986 31764 35992 31776
rect 36044 31764 36050 31816
rect 36078 31764 36084 31816
rect 36136 31764 36142 31816
rect 37458 31804 37464 31816
rect 36188 31776 37464 31804
rect 36188 31736 36216 31776
rect 37458 31764 37464 31776
rect 37516 31764 37522 31816
rect 35728 31708 36216 31736
rect 37568 31736 37596 31912
rect 38657 31909 38669 31943
rect 38703 31909 38715 31943
rect 38657 31903 38715 31909
rect 37642 31832 37648 31884
rect 37700 31832 37706 31884
rect 37921 31807 37979 31813
rect 37921 31804 37933 31807
rect 37752 31776 37933 31804
rect 37752 31736 37780 31776
rect 37921 31773 37933 31776
rect 37967 31773 37979 31807
rect 38672 31804 38700 31903
rect 39868 31881 39896 31980
rect 41966 31968 41972 31980
rect 42024 31968 42030 32020
rect 42334 31968 42340 32020
rect 42392 32008 42398 32020
rect 42429 32011 42487 32017
rect 42429 32008 42441 32011
rect 42392 31980 42441 32008
rect 42392 31968 42398 31980
rect 42429 31977 42441 31980
rect 42475 31977 42487 32011
rect 42429 31971 42487 31977
rect 44634 31968 44640 32020
rect 44692 32008 44698 32020
rect 45097 32011 45155 32017
rect 45097 32008 45109 32011
rect 44692 31980 45109 32008
rect 44692 31968 44698 31980
rect 45097 31977 45109 31980
rect 45143 31977 45155 32011
rect 45097 31971 45155 31977
rect 45002 31940 45008 31952
rect 40052 31912 45008 31940
rect 39853 31875 39911 31881
rect 39853 31841 39865 31875
rect 39899 31841 39911 31875
rect 39853 31835 39911 31841
rect 40052 31804 40080 31912
rect 45002 31900 45008 31912
rect 45060 31900 45066 31952
rect 41506 31832 41512 31884
rect 41564 31872 41570 31884
rect 42613 31875 42671 31881
rect 42613 31872 42625 31875
rect 41564 31844 42625 31872
rect 41564 31832 41570 31844
rect 42613 31841 42625 31844
rect 42659 31841 42671 31875
rect 42613 31835 42671 31841
rect 38672 31776 40080 31804
rect 40129 31807 40187 31813
rect 37921 31767 37979 31773
rect 40129 31773 40141 31807
rect 40175 31804 40187 31807
rect 40218 31804 40224 31816
rect 40175 31776 40224 31804
rect 40175 31773 40187 31776
rect 40129 31767 40187 31773
rect 40218 31764 40224 31776
rect 40276 31764 40282 31816
rect 40586 31764 40592 31816
rect 40644 31804 40650 31816
rect 42242 31804 42248 31816
rect 40644 31776 42248 31804
rect 40644 31764 40650 31776
rect 42242 31764 42248 31776
rect 42300 31764 42306 31816
rect 42337 31807 42395 31813
rect 42337 31773 42349 31807
rect 42383 31804 42395 31807
rect 42702 31804 42708 31816
rect 42383 31776 42708 31804
rect 42383 31773 42395 31776
rect 42337 31767 42395 31773
rect 42702 31764 42708 31776
rect 42760 31764 42766 31816
rect 43714 31804 43720 31816
rect 42812 31776 43720 31804
rect 37568 31708 37780 31736
rect 42613 31739 42671 31745
rect 34977 31699 35035 31705
rect 42613 31705 42625 31739
rect 42659 31736 42671 31739
rect 42812 31736 42840 31776
rect 43714 31764 43720 31776
rect 43772 31764 43778 31816
rect 44910 31764 44916 31816
rect 44968 31804 44974 31816
rect 45005 31807 45063 31813
rect 45005 31804 45017 31807
rect 44968 31776 45017 31804
rect 44968 31764 44974 31776
rect 45005 31773 45017 31776
rect 45051 31773 45063 31807
rect 45005 31767 45063 31773
rect 42659 31708 42840 31736
rect 42659 31705 42671 31708
rect 42613 31699 42671 31705
rect 24688 31640 28304 31668
rect 28994 31628 29000 31680
rect 29052 31628 29058 31680
rect 33962 31628 33968 31680
rect 34020 31628 34026 31680
rect 34992 31668 35020 31699
rect 35158 31668 35164 31680
rect 34992 31640 35164 31668
rect 35158 31628 35164 31640
rect 35216 31628 35222 31680
rect 1104 31578 47104 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 47104 31578
rect 1104 31504 47104 31526
rect 9674 31424 9680 31476
rect 9732 31424 9738 31476
rect 9858 31424 9864 31476
rect 9916 31464 9922 31476
rect 10045 31467 10103 31473
rect 10045 31464 10057 31467
rect 9916 31436 10057 31464
rect 9916 31424 9922 31436
rect 10045 31433 10057 31436
rect 10091 31433 10103 31467
rect 10045 31427 10103 31433
rect 11514 31424 11520 31476
rect 11572 31464 11578 31476
rect 11793 31467 11851 31473
rect 11793 31464 11805 31467
rect 11572 31436 11805 31464
rect 11572 31424 11578 31436
rect 11793 31433 11805 31436
rect 11839 31433 11851 31467
rect 11793 31427 11851 31433
rect 13814 31424 13820 31476
rect 13872 31464 13878 31476
rect 14921 31467 14979 31473
rect 14921 31464 14933 31467
rect 13872 31436 14933 31464
rect 13872 31424 13878 31436
rect 14921 31433 14933 31436
rect 14967 31433 14979 31467
rect 14921 31427 14979 31433
rect 15286 31424 15292 31476
rect 15344 31424 15350 31476
rect 15381 31467 15439 31473
rect 15381 31433 15393 31467
rect 15427 31464 15439 31467
rect 15930 31464 15936 31476
rect 15427 31436 15936 31464
rect 15427 31433 15439 31436
rect 15381 31427 15439 31433
rect 15930 31424 15936 31436
rect 15988 31424 15994 31476
rect 17954 31424 17960 31476
rect 18012 31464 18018 31476
rect 21453 31467 21511 31473
rect 21453 31464 21465 31467
rect 18012 31436 21465 31464
rect 18012 31424 18018 31436
rect 21453 31433 21465 31436
rect 21499 31433 21511 31467
rect 21453 31427 21511 31433
rect 21542 31424 21548 31476
rect 21600 31464 21606 31476
rect 22278 31464 22284 31476
rect 21600 31436 22284 31464
rect 21600 31424 21606 31436
rect 22278 31424 22284 31436
rect 22336 31424 22342 31476
rect 22370 31424 22376 31476
rect 22428 31424 22434 31476
rect 22462 31424 22468 31476
rect 22520 31424 22526 31476
rect 30834 31464 30840 31476
rect 22572 31436 30840 31464
rect 20438 31356 20444 31408
rect 20496 31356 20502 31408
rect 22572 31396 22600 31436
rect 30834 31424 30840 31436
rect 30892 31424 30898 31476
rect 31294 31424 31300 31476
rect 31352 31464 31358 31476
rect 31573 31467 31631 31473
rect 31573 31464 31585 31467
rect 31352 31436 31585 31464
rect 31352 31424 31358 31436
rect 31573 31433 31585 31436
rect 31619 31464 31631 31467
rect 32585 31467 32643 31473
rect 32585 31464 32597 31467
rect 31619 31436 32597 31464
rect 31619 31433 31631 31436
rect 31573 31427 31631 31433
rect 32585 31433 32597 31436
rect 32631 31433 32643 31467
rect 32585 31427 32643 31433
rect 34606 31424 34612 31476
rect 34664 31464 34670 31476
rect 35161 31467 35219 31473
rect 35161 31464 35173 31467
rect 34664 31436 35173 31464
rect 34664 31424 34670 31436
rect 35161 31433 35173 31436
rect 35207 31433 35219 31467
rect 35161 31427 35219 31433
rect 35434 31424 35440 31476
rect 35492 31464 35498 31476
rect 35621 31467 35679 31473
rect 35621 31464 35633 31467
rect 35492 31436 35633 31464
rect 35492 31424 35498 31436
rect 35621 31433 35633 31436
rect 35667 31433 35679 31467
rect 35621 31427 35679 31433
rect 41506 31424 41512 31476
rect 41564 31424 41570 31476
rect 44818 31424 44824 31476
rect 44876 31464 44882 31476
rect 45189 31467 45247 31473
rect 45189 31464 45201 31467
rect 44876 31436 45201 31464
rect 44876 31424 44882 31436
rect 45189 31433 45201 31436
rect 45235 31464 45247 31467
rect 45462 31464 45468 31476
rect 45235 31436 45468 31464
rect 45235 31433 45247 31436
rect 45189 31427 45247 31433
rect 45462 31424 45468 31436
rect 45520 31424 45526 31476
rect 28537 31399 28595 31405
rect 21192 31368 22600 31396
rect 26160 31368 28120 31396
rect 2222 31288 2228 31340
rect 2280 31288 2286 31340
rect 6914 31288 6920 31340
rect 6972 31328 6978 31340
rect 12161 31331 12219 31337
rect 12161 31328 12173 31331
rect 6972 31300 12173 31328
rect 6972 31288 6978 31300
rect 12161 31297 12173 31300
rect 12207 31297 12219 31331
rect 12161 31291 12219 31297
rect 20162 31288 20168 31340
rect 20220 31328 20226 31340
rect 20625 31331 20683 31337
rect 20625 31328 20637 31331
rect 20220 31300 20637 31328
rect 20220 31288 20226 31300
rect 20625 31297 20637 31300
rect 20671 31297 20683 31331
rect 20625 31291 20683 31297
rect 20714 31288 20720 31340
rect 20772 31288 20778 31340
rect 20993 31331 21051 31337
rect 20993 31297 21005 31331
rect 21039 31328 21051 31331
rect 21085 31331 21143 31337
rect 21085 31328 21097 31331
rect 21039 31300 21097 31328
rect 21039 31297 21051 31300
rect 20993 31291 21051 31297
rect 21085 31297 21097 31300
rect 21131 31297 21143 31331
rect 21085 31291 21143 31297
rect 4982 31220 4988 31272
rect 5040 31260 5046 31272
rect 5442 31260 5448 31272
rect 5040 31232 5448 31260
rect 5040 31220 5046 31232
rect 5442 31220 5448 31232
rect 5500 31220 5506 31272
rect 10134 31220 10140 31272
rect 10192 31220 10198 31272
rect 10229 31263 10287 31269
rect 10229 31229 10241 31263
rect 10275 31260 10287 31263
rect 10870 31260 10876 31272
rect 10275 31232 10876 31260
rect 10275 31229 10287 31232
rect 10229 31223 10287 31229
rect 9766 31152 9772 31204
rect 9824 31192 9830 31204
rect 10244 31192 10272 31223
rect 10870 31220 10876 31232
rect 10928 31220 10934 31272
rect 12253 31263 12311 31269
rect 12253 31229 12265 31263
rect 12299 31229 12311 31263
rect 12253 31223 12311 31229
rect 9824 31164 10272 31192
rect 9824 31152 9830 31164
rect 12158 31152 12164 31204
rect 12216 31192 12222 31204
rect 12268 31192 12296 31223
rect 15470 31220 15476 31272
rect 15528 31260 15534 31272
rect 15565 31263 15623 31269
rect 15565 31260 15577 31263
rect 15528 31232 15577 31260
rect 15528 31220 15534 31232
rect 15565 31229 15577 31232
rect 15611 31260 15623 31263
rect 21192 31260 21220 31368
rect 21269 31331 21327 31337
rect 21269 31297 21281 31331
rect 21315 31297 21327 31331
rect 21269 31291 21327 31297
rect 21545 31331 21603 31337
rect 21545 31297 21557 31331
rect 21591 31328 21603 31331
rect 21634 31328 21640 31340
rect 21591 31300 21640 31328
rect 21591 31297 21603 31300
rect 21545 31291 21603 31297
rect 15611 31232 21220 31260
rect 15611 31229 15623 31232
rect 15565 31223 15623 31229
rect 21284 31204 21312 31291
rect 21634 31288 21640 31300
rect 21692 31288 21698 31340
rect 21726 31220 21732 31272
rect 21784 31260 21790 31272
rect 22370 31260 22376 31272
rect 21784 31232 22376 31260
rect 21784 31220 21790 31232
rect 22370 31220 22376 31232
rect 22428 31260 22434 31272
rect 22557 31263 22615 31269
rect 22557 31260 22569 31263
rect 22428 31232 22569 31260
rect 22428 31220 22434 31232
rect 22557 31229 22569 31232
rect 22603 31229 22615 31263
rect 22557 31223 22615 31229
rect 23566 31220 23572 31272
rect 23624 31220 23630 31272
rect 23750 31220 23756 31272
rect 23808 31220 23814 31272
rect 24210 31220 24216 31272
rect 24268 31220 24274 31272
rect 24486 31220 24492 31272
rect 24544 31220 24550 31272
rect 24578 31220 24584 31272
rect 24636 31269 24642 31272
rect 24636 31263 24664 31269
rect 24652 31229 24664 31263
rect 24636 31223 24664 31229
rect 24765 31263 24823 31269
rect 24765 31229 24777 31263
rect 24811 31260 24823 31263
rect 25590 31260 25596 31272
rect 24811 31232 25596 31260
rect 24811 31229 24823 31232
rect 24765 31223 24823 31229
rect 24636 31220 24642 31223
rect 25590 31220 25596 31232
rect 25648 31220 25654 31272
rect 25685 31263 25743 31269
rect 25685 31229 25697 31263
rect 25731 31260 25743 31263
rect 25774 31260 25780 31272
rect 25731 31232 25780 31260
rect 25731 31229 25743 31232
rect 25685 31223 25743 31229
rect 25774 31220 25780 31232
rect 25832 31220 25838 31272
rect 26160 31269 26188 31368
rect 28092 31337 28120 31368
rect 28537 31365 28549 31399
rect 28583 31396 28595 31399
rect 33778 31396 33784 31408
rect 28583 31368 33784 31396
rect 28583 31365 28595 31368
rect 28537 31359 28595 31365
rect 33778 31356 33784 31368
rect 33836 31356 33842 31408
rect 33962 31405 33968 31408
rect 33956 31359 33968 31405
rect 33962 31356 33968 31359
rect 34020 31356 34026 31408
rect 36078 31396 36084 31408
rect 34072 31368 36084 31396
rect 27709 31331 27767 31337
rect 27709 31297 27721 31331
rect 27755 31297 27767 31331
rect 27709 31291 27767 31297
rect 27801 31331 27859 31337
rect 27801 31297 27813 31331
rect 27847 31297 27859 31331
rect 27801 31291 27859 31297
rect 28077 31331 28135 31337
rect 28077 31297 28089 31331
rect 28123 31297 28135 31331
rect 28077 31291 28135 31297
rect 26145 31263 26203 31269
rect 26145 31229 26157 31263
rect 26191 31229 26203 31263
rect 26145 31223 26203 31229
rect 12216 31164 12296 31192
rect 12360 31164 21220 31192
rect 12216 31152 12222 31164
rect 2038 31084 2044 31136
rect 2096 31084 2102 31136
rect 7650 31084 7656 31136
rect 7708 31124 7714 31136
rect 12360 31124 12388 31164
rect 7708 31096 12388 31124
rect 12437 31127 12495 31133
rect 7708 31084 7714 31096
rect 12437 31093 12449 31127
rect 12483 31124 12495 31127
rect 20806 31124 20812 31136
rect 12483 31096 20812 31124
rect 12483 31093 12495 31096
rect 12437 31087 12495 31093
rect 20806 31084 20812 31096
rect 20864 31084 20870 31136
rect 20901 31127 20959 31133
rect 20901 31093 20913 31127
rect 20947 31124 20959 31127
rect 21082 31124 21088 31136
rect 20947 31096 21088 31124
rect 20947 31093 20959 31096
rect 20901 31087 20959 31093
rect 21082 31084 21088 31096
rect 21140 31084 21146 31136
rect 21192 31124 21220 31164
rect 21266 31152 21272 31204
rect 21324 31152 21330 31204
rect 22005 31195 22063 31201
rect 22005 31161 22017 31195
rect 22051 31192 22063 31195
rect 22186 31192 22192 31204
rect 22051 31164 22192 31192
rect 22051 31161 22063 31164
rect 22005 31155 22063 31161
rect 22186 31152 22192 31164
rect 22244 31152 22250 31204
rect 23658 31152 23664 31204
rect 23716 31192 23722 31204
rect 24228 31192 24256 31220
rect 23716 31164 24256 31192
rect 25409 31195 25467 31201
rect 23716 31152 23722 31164
rect 25409 31161 25421 31195
rect 25455 31192 25467 31195
rect 25961 31195 26019 31201
rect 25961 31192 25973 31195
rect 25455 31164 25973 31192
rect 25455 31161 25467 31164
rect 25409 31155 25467 31161
rect 25961 31161 25973 31164
rect 26007 31161 26019 31195
rect 27724 31192 27752 31291
rect 27816 31260 27844 31291
rect 28258 31288 28264 31340
rect 28316 31328 28322 31340
rect 28353 31331 28411 31337
rect 28353 31328 28365 31331
rect 28316 31300 28365 31328
rect 28316 31288 28322 31300
rect 28353 31297 28365 31300
rect 28399 31328 28411 31331
rect 28442 31328 28448 31340
rect 28399 31300 28448 31328
rect 28399 31297 28411 31300
rect 28353 31291 28411 31297
rect 28442 31288 28448 31300
rect 28500 31288 28506 31340
rect 28629 31331 28687 31337
rect 28629 31297 28641 31331
rect 28675 31328 28687 31331
rect 29086 31328 29092 31340
rect 28675 31300 29092 31328
rect 28675 31297 28687 31300
rect 28629 31291 28687 31297
rect 29086 31288 29092 31300
rect 29144 31288 29150 31340
rect 31021 31331 31079 31337
rect 31021 31297 31033 31331
rect 31067 31328 31079 31331
rect 31481 31331 31539 31337
rect 31067 31300 31156 31328
rect 31067 31297 31079 31300
rect 31021 31291 31079 31297
rect 28169 31263 28227 31269
rect 28169 31260 28181 31263
rect 27816 31232 28181 31260
rect 28169 31229 28181 31232
rect 28215 31229 28227 31263
rect 28169 31223 28227 31229
rect 28994 31192 29000 31204
rect 27724 31164 29000 31192
rect 25961 31155 26019 31161
rect 28994 31152 29000 31164
rect 29052 31152 29058 31204
rect 31128 31201 31156 31300
rect 31481 31297 31493 31331
rect 31527 31328 31539 31331
rect 31938 31328 31944 31340
rect 31527 31300 31944 31328
rect 31527 31297 31539 31300
rect 31481 31291 31539 31297
rect 31938 31288 31944 31300
rect 31996 31288 32002 31340
rect 32493 31331 32551 31337
rect 32493 31297 32505 31331
rect 32539 31328 32551 31331
rect 33042 31328 33048 31340
rect 32539 31300 33048 31328
rect 32539 31297 32551 31300
rect 32493 31291 32551 31297
rect 33042 31288 33048 31300
rect 33100 31288 33106 31340
rect 34072 31328 34100 31368
rect 36078 31356 36084 31368
rect 36136 31356 36142 31408
rect 41524 31396 41552 31424
rect 41524 31368 41736 31396
rect 33152 31300 34100 31328
rect 35529 31331 35587 31337
rect 31386 31220 31392 31272
rect 31444 31260 31450 31272
rect 31665 31263 31723 31269
rect 31665 31260 31677 31263
rect 31444 31232 31677 31260
rect 31444 31220 31450 31232
rect 31665 31229 31677 31232
rect 31711 31229 31723 31263
rect 31665 31223 31723 31229
rect 32030 31220 32036 31272
rect 32088 31260 32094 31272
rect 32582 31260 32588 31272
rect 32088 31232 32588 31260
rect 32088 31220 32094 31232
rect 32582 31220 32588 31232
rect 32640 31260 32646 31272
rect 32677 31263 32735 31269
rect 32677 31260 32689 31263
rect 32640 31232 32689 31260
rect 32640 31220 32646 31232
rect 32677 31229 32689 31232
rect 32723 31229 32735 31263
rect 32677 31223 32735 31229
rect 31113 31195 31171 31201
rect 31113 31161 31125 31195
rect 31159 31161 31171 31195
rect 31113 31155 31171 31161
rect 31202 31152 31208 31204
rect 31260 31192 31266 31204
rect 32125 31195 32183 31201
rect 32125 31192 32137 31195
rect 31260 31164 32137 31192
rect 31260 31152 31266 31164
rect 32125 31161 32137 31164
rect 32171 31161 32183 31195
rect 33152 31192 33180 31300
rect 35529 31297 35541 31331
rect 35575 31297 35587 31331
rect 35529 31291 35587 31297
rect 33410 31220 33416 31272
rect 33468 31260 33474 31272
rect 33689 31263 33747 31269
rect 33689 31260 33701 31263
rect 33468 31232 33701 31260
rect 33468 31220 33474 31232
rect 33689 31229 33701 31232
rect 33735 31229 33747 31263
rect 33689 31223 33747 31229
rect 32125 31155 32183 31161
rect 32232 31164 33180 31192
rect 35069 31195 35127 31201
rect 22922 31124 22928 31136
rect 21192 31096 22928 31124
rect 22922 31084 22928 31096
rect 22980 31084 22986 31136
rect 23842 31084 23848 31136
rect 23900 31124 23906 31136
rect 24762 31124 24768 31136
rect 23900 31096 24768 31124
rect 23900 31084 23906 31096
rect 24762 31084 24768 31096
rect 24820 31084 24826 31136
rect 27522 31084 27528 31136
rect 27580 31084 27586 31136
rect 27982 31084 27988 31136
rect 28040 31084 28046 31136
rect 30834 31084 30840 31136
rect 30892 31084 30898 31136
rect 31846 31084 31852 31136
rect 31904 31124 31910 31136
rect 32232 31124 32260 31164
rect 35069 31161 35081 31195
rect 35115 31192 35127 31195
rect 35544 31192 35572 31291
rect 36354 31288 36360 31340
rect 36412 31328 36418 31340
rect 36449 31331 36507 31337
rect 36449 31328 36461 31331
rect 36412 31300 36461 31328
rect 36412 31288 36418 31300
rect 36449 31297 36461 31300
rect 36495 31328 36507 31331
rect 36538 31328 36544 31340
rect 36495 31300 36544 31328
rect 36495 31297 36507 31300
rect 36449 31291 36507 31297
rect 36538 31288 36544 31300
rect 36596 31288 36602 31340
rect 36725 31331 36783 31337
rect 36725 31297 36737 31331
rect 36771 31328 36783 31331
rect 37274 31328 37280 31340
rect 36771 31300 37280 31328
rect 36771 31297 36783 31300
rect 36725 31291 36783 31297
rect 37274 31288 37280 31300
rect 37332 31288 37338 31340
rect 37550 31288 37556 31340
rect 37608 31288 37614 31340
rect 41708 31337 41736 31368
rect 41325 31331 41383 31337
rect 41325 31297 41337 31331
rect 41371 31297 41383 31331
rect 41325 31291 41383 31297
rect 41601 31331 41659 31337
rect 41601 31297 41613 31331
rect 41647 31297 41659 31331
rect 41601 31291 41659 31297
rect 41693 31331 41751 31337
rect 41693 31297 41705 31331
rect 41739 31297 41751 31331
rect 41693 31291 41751 31297
rect 41785 31331 41843 31337
rect 41785 31297 41797 31331
rect 41831 31328 41843 31331
rect 43070 31328 43076 31340
rect 41831 31300 43076 31328
rect 41831 31297 41843 31300
rect 41785 31291 41843 31297
rect 35710 31220 35716 31272
rect 35768 31220 35774 31272
rect 35115 31164 35572 31192
rect 35115 31161 35127 31164
rect 35069 31155 35127 31161
rect 31904 31096 32260 31124
rect 31904 31084 31910 31096
rect 32306 31084 32312 31136
rect 32364 31124 32370 31136
rect 35084 31124 35112 31155
rect 35618 31152 35624 31204
rect 35676 31192 35682 31204
rect 41340 31192 41368 31291
rect 41616 31260 41644 31291
rect 41800 31260 41828 31291
rect 43070 31288 43076 31300
rect 43128 31288 43134 31340
rect 41616 31232 41828 31260
rect 41969 31263 42027 31269
rect 41969 31229 41981 31263
rect 42015 31260 42027 31263
rect 42702 31260 42708 31272
rect 42015 31232 42708 31260
rect 42015 31229 42027 31232
rect 41969 31223 42027 31229
rect 42702 31220 42708 31232
rect 42760 31220 42766 31272
rect 44726 31220 44732 31272
rect 44784 31220 44790 31272
rect 41877 31195 41935 31201
rect 41877 31192 41889 31195
rect 35676 31164 36952 31192
rect 41340 31164 41889 31192
rect 35676 31152 35682 31164
rect 32364 31096 35112 31124
rect 32364 31084 32370 31096
rect 35158 31084 35164 31136
rect 35216 31124 35222 31136
rect 35636 31124 35664 31152
rect 36924 31136 36952 31164
rect 41877 31161 41889 31164
rect 41923 31161 41935 31195
rect 41877 31155 41935 31161
rect 45002 31152 45008 31204
rect 45060 31192 45066 31204
rect 45097 31195 45155 31201
rect 45097 31192 45109 31195
rect 45060 31164 45109 31192
rect 45060 31152 45066 31164
rect 45097 31161 45109 31164
rect 45143 31192 45155 31195
rect 45186 31192 45192 31204
rect 45143 31164 45192 31192
rect 45143 31161 45155 31164
rect 45097 31155 45155 31161
rect 45186 31152 45192 31164
rect 45244 31152 45250 31204
rect 35216 31096 35664 31124
rect 35216 31084 35222 31096
rect 36538 31084 36544 31136
rect 36596 31124 36602 31136
rect 36722 31124 36728 31136
rect 36596 31096 36728 31124
rect 36596 31084 36602 31096
rect 36722 31084 36728 31096
rect 36780 31084 36786 31136
rect 36906 31084 36912 31136
rect 36964 31084 36970 31136
rect 37366 31084 37372 31136
rect 37424 31124 37430 31136
rect 37645 31127 37703 31133
rect 37645 31124 37657 31127
rect 37424 31096 37657 31124
rect 37424 31084 37430 31096
rect 37645 31093 37657 31096
rect 37691 31124 37703 31127
rect 37918 31124 37924 31136
rect 37691 31096 37924 31124
rect 37691 31093 37703 31096
rect 37645 31087 37703 31093
rect 37918 31084 37924 31096
rect 37976 31084 37982 31136
rect 40402 31084 40408 31136
rect 40460 31124 40466 31136
rect 41325 31127 41383 31133
rect 41325 31124 41337 31127
rect 40460 31096 41337 31124
rect 40460 31084 40466 31096
rect 41325 31093 41337 31096
rect 41371 31093 41383 31127
rect 41325 31087 41383 31093
rect 1104 31034 47104 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 47104 31034
rect 1104 30960 47104 30982
rect 4982 30880 4988 30932
rect 5040 30880 5046 30932
rect 12894 30880 12900 30932
rect 12952 30920 12958 30932
rect 13081 30923 13139 30929
rect 13081 30920 13093 30923
rect 12952 30892 13093 30920
rect 12952 30880 12958 30892
rect 13081 30889 13093 30892
rect 13127 30889 13139 30923
rect 13081 30883 13139 30889
rect 13354 30880 13360 30932
rect 13412 30920 13418 30932
rect 17954 30920 17960 30932
rect 13412 30892 17960 30920
rect 13412 30880 13418 30892
rect 17954 30880 17960 30892
rect 18012 30880 18018 30932
rect 21082 30880 21088 30932
rect 21140 30880 21146 30932
rect 21634 30880 21640 30932
rect 21692 30920 21698 30932
rect 22189 30923 22247 30929
rect 22189 30920 22201 30923
rect 21692 30892 22201 30920
rect 21692 30880 21698 30892
rect 22189 30889 22201 30892
rect 22235 30889 22247 30923
rect 22189 30883 22247 30889
rect 23750 30880 23756 30932
rect 23808 30920 23814 30932
rect 24213 30923 24271 30929
rect 24213 30920 24225 30923
rect 23808 30892 24225 30920
rect 23808 30880 23814 30892
rect 24213 30889 24225 30892
rect 24259 30889 24271 30923
rect 24213 30883 24271 30889
rect 4065 30855 4123 30861
rect 4065 30821 4077 30855
rect 4111 30821 4123 30855
rect 4065 30815 4123 30821
rect 1762 30676 1768 30728
rect 1820 30676 1826 30728
rect 2038 30725 2044 30728
rect 2032 30716 2044 30725
rect 1999 30688 2044 30716
rect 2032 30679 2044 30688
rect 2038 30676 2044 30679
rect 2096 30676 2102 30728
rect 3973 30719 4031 30725
rect 3973 30685 3985 30719
rect 4019 30716 4031 30719
rect 4080 30716 4108 30815
rect 4709 30787 4767 30793
rect 4709 30753 4721 30787
rect 4755 30784 4767 30787
rect 5000 30784 5028 30880
rect 10134 30812 10140 30864
rect 10192 30852 10198 30864
rect 10192 30824 16804 30852
rect 10192 30812 10198 30824
rect 4755 30756 5028 30784
rect 4755 30753 4767 30756
rect 4709 30747 4767 30753
rect 10962 30744 10968 30796
rect 11020 30744 11026 30796
rect 13630 30744 13636 30796
rect 13688 30744 13694 30796
rect 16776 30784 16804 30824
rect 20990 30812 20996 30864
rect 21048 30812 21054 30864
rect 22462 30784 22468 30796
rect 16776 30756 22468 30784
rect 22462 30744 22468 30756
rect 22520 30744 22526 30796
rect 22830 30744 22836 30796
rect 22888 30744 22894 30796
rect 4019 30688 4108 30716
rect 4019 30685 4031 30688
rect 3973 30679 4031 30685
rect 4798 30676 4804 30728
rect 4856 30716 4862 30728
rect 4985 30719 5043 30725
rect 4985 30716 4997 30719
rect 4856 30688 4997 30716
rect 4856 30676 4862 30688
rect 4985 30685 4997 30688
rect 5031 30685 5043 30719
rect 16022 30716 16028 30728
rect 4985 30679 5043 30685
rect 5184 30688 16028 30716
rect 1780 30648 1808 30676
rect 2590 30648 2596 30660
rect 1780 30620 2596 30648
rect 2590 30608 2596 30620
rect 2648 30608 2654 30660
rect 4433 30651 4491 30657
rect 4433 30617 4445 30651
rect 4479 30648 4491 30651
rect 4614 30648 4620 30660
rect 4479 30620 4620 30648
rect 4479 30617 4491 30620
rect 4433 30611 4491 30617
rect 4614 30608 4620 30620
rect 4672 30608 4678 30660
rect 3142 30540 3148 30592
rect 3200 30540 3206 30592
rect 3786 30540 3792 30592
rect 3844 30540 3850 30592
rect 4154 30540 4160 30592
rect 4212 30580 4218 30592
rect 4525 30583 4583 30589
rect 4525 30580 4537 30583
rect 4212 30552 4537 30580
rect 4212 30540 4218 30552
rect 4525 30549 4537 30552
rect 4571 30580 4583 30583
rect 5184 30580 5212 30688
rect 16022 30676 16028 30688
rect 16080 30716 16086 30728
rect 16482 30716 16488 30728
rect 16080 30688 16488 30716
rect 16080 30676 16086 30688
rect 16482 30676 16488 30688
rect 16540 30676 16546 30728
rect 20625 30719 20683 30725
rect 20625 30685 20637 30719
rect 20671 30716 20683 30719
rect 21910 30716 21916 30728
rect 20671 30688 21916 30716
rect 20671 30685 20683 30688
rect 20625 30679 20683 30685
rect 21910 30676 21916 30688
rect 21968 30676 21974 30728
rect 24228 30716 24256 30883
rect 24486 30880 24492 30932
rect 24544 30920 24550 30932
rect 24854 30920 24860 30932
rect 24544 30892 24860 30920
rect 24544 30880 24550 30892
rect 24854 30880 24860 30892
rect 24912 30880 24918 30932
rect 27522 30880 27528 30932
rect 27580 30920 27586 30932
rect 31846 30920 31852 30932
rect 27580 30892 31852 30920
rect 27580 30880 27586 30892
rect 31846 30880 31852 30892
rect 31904 30880 31910 30932
rect 31938 30880 31944 30932
rect 31996 30920 32002 30932
rect 33134 30920 33140 30932
rect 31996 30892 33140 30920
rect 31996 30880 32002 30892
rect 33134 30880 33140 30892
rect 33192 30880 33198 30932
rect 33778 30880 33784 30932
rect 33836 30920 33842 30932
rect 33965 30923 34023 30929
rect 33965 30920 33977 30923
rect 33836 30892 33977 30920
rect 33836 30880 33842 30892
rect 33965 30889 33977 30892
rect 34011 30889 34023 30923
rect 33965 30883 34023 30889
rect 34330 30880 34336 30932
rect 34388 30920 34394 30932
rect 35066 30920 35072 30932
rect 34388 30892 35072 30920
rect 34388 30880 34394 30892
rect 35066 30880 35072 30892
rect 35124 30880 35130 30932
rect 35345 30923 35403 30929
rect 35345 30889 35357 30923
rect 35391 30920 35403 30923
rect 35434 30920 35440 30932
rect 35391 30892 35440 30920
rect 35391 30889 35403 30892
rect 35345 30883 35403 30889
rect 35434 30880 35440 30892
rect 35492 30880 35498 30932
rect 38381 30923 38439 30929
rect 36188 30892 38148 30920
rect 24397 30855 24455 30861
rect 24397 30821 24409 30855
rect 24443 30852 24455 30855
rect 24443 30824 25452 30852
rect 24443 30821 24455 30824
rect 24397 30815 24455 30821
rect 24670 30744 24676 30796
rect 24728 30784 24734 30796
rect 24857 30787 24915 30793
rect 24857 30784 24869 30787
rect 24728 30756 24869 30784
rect 24728 30744 24734 30756
rect 24857 30753 24869 30756
rect 24903 30753 24915 30787
rect 24857 30747 24915 30753
rect 24946 30744 24952 30796
rect 25004 30744 25010 30796
rect 25424 30725 25452 30824
rect 27338 30812 27344 30864
rect 27396 30852 27402 30864
rect 27982 30852 27988 30864
rect 27396 30824 27988 30852
rect 27396 30812 27402 30824
rect 27982 30812 27988 30824
rect 28040 30812 28046 30864
rect 31662 30812 31668 30864
rect 31720 30852 31726 30864
rect 31720 30824 32904 30852
rect 31720 30812 31726 30824
rect 27798 30744 27804 30796
rect 27856 30744 27862 30796
rect 30558 30744 30564 30796
rect 30616 30744 30622 30796
rect 32122 30744 32128 30796
rect 32180 30784 32186 30796
rect 32490 30784 32496 30796
rect 32180 30756 32496 30784
rect 32180 30744 32186 30756
rect 32490 30744 32496 30756
rect 32548 30744 32554 30796
rect 32766 30744 32772 30796
rect 32824 30744 32830 30796
rect 32876 30784 32904 30824
rect 34514 30812 34520 30864
rect 34572 30852 34578 30864
rect 36081 30855 36139 30861
rect 34572 30824 35664 30852
rect 34572 30812 34578 30824
rect 32876 30756 35572 30784
rect 24765 30719 24823 30725
rect 24765 30716 24777 30719
rect 24228 30688 24777 30716
rect 24765 30685 24777 30688
rect 24811 30685 24823 30719
rect 24765 30679 24823 30685
rect 25409 30719 25467 30725
rect 25409 30685 25421 30719
rect 25455 30685 25467 30719
rect 25409 30679 25467 30685
rect 27617 30719 27675 30725
rect 27617 30685 27629 30719
rect 27663 30716 27675 30719
rect 28626 30716 28632 30728
rect 27663 30688 28632 30716
rect 27663 30685 27675 30688
rect 27617 30679 27675 30685
rect 28626 30676 28632 30688
rect 28684 30676 28690 30728
rect 30834 30725 30840 30728
rect 30469 30719 30527 30725
rect 30469 30685 30481 30719
rect 30515 30685 30527 30719
rect 30828 30716 30840 30725
rect 30795 30688 30840 30716
rect 30469 30679 30527 30685
rect 30828 30679 30840 30688
rect 5252 30651 5310 30657
rect 5252 30617 5264 30651
rect 5298 30648 5310 30651
rect 5442 30648 5448 30660
rect 5298 30620 5448 30648
rect 5298 30617 5310 30620
rect 5252 30611 5310 30617
rect 5442 30608 5448 30620
rect 5500 30608 5506 30660
rect 8294 30608 8300 30660
rect 8352 30648 8358 30660
rect 10781 30651 10839 30657
rect 10781 30648 10793 30651
rect 8352 30620 10793 30648
rect 8352 30608 8358 30620
rect 10781 30617 10793 30620
rect 10827 30617 10839 30651
rect 10781 30611 10839 30617
rect 10873 30651 10931 30657
rect 10873 30617 10885 30651
rect 10919 30648 10931 30651
rect 13354 30648 13360 30660
rect 10919 30620 13360 30648
rect 10919 30617 10931 30620
rect 10873 30611 10931 30617
rect 13354 30608 13360 30620
rect 13412 30608 13418 30660
rect 13449 30651 13507 30657
rect 13449 30617 13461 30651
rect 13495 30648 13507 30651
rect 15746 30648 15752 30660
rect 13495 30620 15752 30648
rect 13495 30617 13507 30620
rect 13449 30611 13507 30617
rect 15746 30608 15752 30620
rect 15804 30608 15810 30660
rect 21726 30608 21732 30660
rect 21784 30648 21790 30660
rect 22097 30651 22155 30657
rect 22097 30648 22109 30651
rect 21784 30620 22109 30648
rect 21784 30608 21790 30620
rect 22097 30617 22109 30620
rect 22143 30617 22155 30651
rect 22097 30611 22155 30617
rect 23100 30651 23158 30657
rect 23100 30617 23112 30651
rect 23146 30648 23158 30651
rect 23146 30620 25268 30648
rect 23146 30617 23158 30620
rect 23100 30611 23158 30617
rect 4571 30552 5212 30580
rect 6365 30583 6423 30589
rect 4571 30549 4583 30552
rect 4525 30543 4583 30549
rect 6365 30549 6377 30583
rect 6411 30580 6423 30583
rect 6822 30580 6828 30592
rect 6411 30552 6828 30580
rect 6411 30549 6423 30552
rect 6365 30543 6423 30549
rect 6822 30540 6828 30552
rect 6880 30540 6886 30592
rect 10134 30540 10140 30592
rect 10192 30580 10198 30592
rect 10413 30583 10471 30589
rect 10413 30580 10425 30583
rect 10192 30552 10425 30580
rect 10192 30540 10198 30552
rect 10413 30549 10425 30552
rect 10459 30549 10471 30583
rect 10413 30543 10471 30549
rect 13538 30540 13544 30592
rect 13596 30540 13602 30592
rect 19334 30540 19340 30592
rect 19392 30580 19398 30592
rect 20806 30580 20812 30592
rect 19392 30552 20812 30580
rect 19392 30540 19398 30552
rect 20806 30540 20812 30552
rect 20864 30540 20870 30592
rect 21082 30540 21088 30592
rect 21140 30580 21146 30592
rect 21450 30580 21456 30592
rect 21140 30552 21456 30580
rect 21140 30540 21146 30552
rect 21450 30540 21456 30552
rect 21508 30540 21514 30592
rect 25240 30589 25268 30620
rect 26050 30608 26056 30660
rect 26108 30648 26114 30660
rect 29086 30648 29092 30660
rect 26108 30620 29092 30648
rect 26108 30608 26114 30620
rect 29086 30608 29092 30620
rect 29144 30608 29150 30660
rect 30484 30648 30512 30679
rect 30834 30676 30840 30679
rect 30892 30676 30898 30728
rect 32306 30676 32312 30728
rect 32364 30676 32370 30728
rect 33042 30676 33048 30728
rect 33100 30676 33106 30728
rect 33134 30676 33140 30728
rect 33192 30725 33198 30728
rect 33192 30719 33220 30725
rect 33208 30685 33220 30719
rect 33192 30679 33220 30685
rect 33192 30676 33198 30679
rect 33318 30676 33324 30728
rect 33376 30676 33382 30728
rect 34698 30676 34704 30728
rect 34756 30676 34762 30728
rect 34794 30719 34852 30725
rect 34794 30685 34806 30719
rect 34840 30685 34852 30719
rect 34794 30679 34852 30685
rect 31202 30648 31208 30660
rect 30484 30620 31208 30648
rect 31202 30608 31208 30620
rect 31260 30608 31266 30660
rect 25225 30583 25283 30589
rect 25225 30549 25237 30583
rect 25271 30549 25283 30583
rect 25225 30543 25283 30549
rect 25866 30540 25872 30592
rect 25924 30580 25930 30592
rect 27249 30583 27307 30589
rect 27249 30580 27261 30583
rect 25924 30552 27261 30580
rect 25924 30540 25930 30552
rect 27249 30549 27261 30552
rect 27295 30549 27307 30583
rect 27249 30543 27307 30549
rect 27709 30583 27767 30589
rect 27709 30549 27721 30583
rect 27755 30580 27767 30583
rect 29730 30580 29736 30592
rect 27755 30552 29736 30580
rect 27755 30549 27767 30552
rect 27709 30543 27767 30549
rect 29730 30540 29736 30552
rect 29788 30540 29794 30592
rect 30285 30583 30343 30589
rect 30285 30549 30297 30583
rect 30331 30580 30343 30583
rect 30834 30580 30840 30592
rect 30331 30552 30840 30580
rect 30331 30549 30343 30552
rect 30285 30543 30343 30549
rect 30834 30540 30840 30552
rect 30892 30540 30898 30592
rect 32214 30540 32220 30592
rect 32272 30580 32278 30592
rect 34808 30580 34836 30679
rect 35066 30676 35072 30728
rect 35124 30676 35130 30728
rect 35158 30676 35164 30728
rect 35216 30725 35222 30728
rect 35544 30725 35572 30756
rect 35216 30716 35224 30725
rect 35529 30719 35587 30725
rect 35216 30688 35261 30716
rect 35216 30679 35224 30688
rect 35529 30685 35541 30719
rect 35575 30685 35587 30719
rect 35636 30716 35664 30824
rect 36081 30821 36093 30855
rect 36127 30821 36139 30855
rect 36081 30815 36139 30821
rect 36096 30728 36124 30815
rect 35805 30719 35863 30725
rect 35805 30716 35817 30719
rect 35636 30688 35817 30716
rect 35529 30679 35587 30685
rect 35805 30685 35817 30688
rect 35851 30685 35863 30719
rect 35805 30679 35863 30685
rect 35897 30719 35955 30725
rect 35897 30685 35909 30719
rect 35943 30716 35955 30719
rect 35986 30716 35992 30728
rect 35943 30688 35992 30716
rect 35943 30685 35955 30688
rect 35897 30679 35955 30685
rect 35216 30676 35222 30679
rect 35986 30676 35992 30688
rect 36044 30676 36050 30728
rect 36078 30676 36084 30728
rect 36136 30676 36142 30728
rect 36188 30725 36216 30892
rect 38120 30852 38148 30892
rect 38381 30889 38393 30923
rect 38427 30920 38439 30923
rect 40494 30920 40500 30932
rect 38427 30892 40500 30920
rect 38427 30889 38439 30892
rect 38381 30883 38439 30889
rect 40494 30880 40500 30892
rect 40552 30920 40558 30932
rect 40589 30923 40647 30929
rect 40589 30920 40601 30923
rect 40552 30892 40601 30920
rect 40552 30880 40558 30892
rect 40589 30889 40601 30892
rect 40635 30889 40647 30923
rect 40589 30883 40647 30889
rect 46198 30852 46204 30864
rect 38120 30824 46204 30852
rect 46198 30812 46204 30824
rect 46256 30812 46262 30864
rect 36354 30784 36360 30796
rect 36280 30756 36360 30784
rect 36173 30719 36231 30725
rect 36173 30685 36185 30719
rect 36219 30685 36231 30719
rect 36173 30679 36231 30685
rect 34977 30651 35035 30657
rect 34977 30617 34989 30651
rect 35023 30617 35035 30651
rect 34977 30611 35035 30617
rect 35713 30651 35771 30657
rect 35713 30617 35725 30651
rect 35759 30617 35771 30651
rect 36004 30648 36032 30676
rect 36280 30648 36308 30756
rect 36354 30744 36360 30756
rect 36412 30784 36418 30796
rect 36412 30756 36584 30784
rect 36412 30744 36418 30756
rect 36446 30676 36452 30728
rect 36504 30676 36510 30728
rect 36556 30725 36584 30756
rect 39114 30744 39120 30796
rect 39172 30784 39178 30796
rect 40218 30784 40224 30796
rect 39172 30756 40224 30784
rect 39172 30744 39178 30756
rect 40218 30744 40224 30756
rect 40276 30784 40282 30796
rect 40276 30756 40540 30784
rect 40276 30744 40282 30756
rect 36541 30719 36599 30725
rect 36541 30685 36553 30719
rect 36587 30716 36599 30719
rect 36909 30719 36967 30725
rect 36909 30716 36921 30719
rect 36587 30688 36921 30716
rect 36587 30685 36599 30688
rect 36541 30679 36599 30685
rect 36909 30685 36921 30688
rect 36955 30685 36967 30719
rect 36909 30679 36967 30685
rect 37185 30719 37243 30725
rect 37185 30685 37197 30719
rect 37231 30716 37243 30719
rect 37274 30716 37280 30728
rect 37231 30688 37280 30716
rect 37231 30685 37243 30688
rect 37185 30679 37243 30685
rect 37274 30676 37280 30688
rect 37332 30676 37338 30728
rect 37366 30676 37372 30728
rect 37424 30676 37430 30728
rect 37642 30676 37648 30728
rect 37700 30676 37706 30728
rect 40034 30676 40040 30728
rect 40092 30676 40098 30728
rect 40129 30719 40187 30725
rect 40129 30685 40141 30719
rect 40175 30685 40187 30719
rect 40129 30679 40187 30685
rect 36004 30620 36308 30648
rect 35713 30611 35771 30617
rect 32272 30552 34836 30580
rect 34992 30580 35020 30611
rect 35618 30580 35624 30592
rect 34992 30552 35624 30580
rect 32272 30540 32278 30552
rect 35618 30540 35624 30552
rect 35676 30540 35682 30592
rect 35728 30580 35756 30611
rect 36354 30608 36360 30660
rect 36412 30608 36418 30660
rect 40144 30648 40172 30679
rect 40310 30676 40316 30728
rect 40368 30676 40374 30728
rect 40402 30676 40408 30728
rect 40460 30676 40466 30728
rect 40512 30725 40540 30756
rect 45370 30744 45376 30796
rect 45428 30744 45434 30796
rect 45738 30744 45744 30796
rect 45796 30784 45802 30796
rect 45833 30787 45891 30793
rect 45833 30784 45845 30787
rect 45796 30756 45845 30784
rect 45796 30744 45802 30756
rect 45833 30753 45845 30756
rect 45879 30753 45891 30787
rect 45833 30747 45891 30753
rect 40497 30719 40555 30725
rect 40497 30685 40509 30719
rect 40543 30685 40555 30719
rect 40497 30679 40555 30685
rect 45462 30676 45468 30728
rect 45520 30676 45526 30728
rect 46106 30676 46112 30728
rect 46164 30676 46170 30728
rect 40144 30620 40448 30648
rect 36372 30580 36400 30608
rect 40420 30592 40448 30620
rect 35728 30552 36400 30580
rect 36446 30540 36452 30592
rect 36504 30580 36510 30592
rect 36725 30583 36783 30589
rect 36725 30580 36737 30583
rect 36504 30552 36737 30580
rect 36504 30540 36510 30552
rect 36725 30549 36737 30552
rect 36771 30549 36783 30583
rect 36725 30543 36783 30549
rect 37185 30583 37243 30589
rect 37185 30549 37197 30583
rect 37231 30580 37243 30583
rect 37734 30580 37740 30592
rect 37231 30552 37740 30580
rect 37231 30549 37243 30552
rect 37185 30543 37243 30549
rect 37734 30540 37740 30552
rect 37792 30540 37798 30592
rect 39390 30540 39396 30592
rect 39448 30580 39454 30592
rect 39853 30583 39911 30589
rect 39853 30580 39865 30583
rect 39448 30552 39865 30580
rect 39448 30540 39454 30552
rect 39853 30549 39865 30552
rect 39899 30549 39911 30583
rect 39853 30543 39911 30549
rect 40402 30540 40408 30592
rect 40460 30540 40466 30592
rect 40954 30540 40960 30592
rect 41012 30540 41018 30592
rect 45922 30540 45928 30592
rect 45980 30540 45986 30592
rect 1104 30490 47104 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 47104 30490
rect 1104 30416 47104 30438
rect 1949 30379 2007 30385
rect 1949 30345 1961 30379
rect 1995 30376 2007 30379
rect 2222 30376 2228 30388
rect 1995 30348 2228 30376
rect 1995 30345 2007 30348
rect 1949 30339 2007 30345
rect 2222 30336 2228 30348
rect 2280 30336 2286 30388
rect 3142 30376 3148 30388
rect 2746 30348 3148 30376
rect 2406 30268 2412 30320
rect 2464 30268 2470 30320
rect 2317 30243 2375 30249
rect 2317 30209 2329 30243
rect 2363 30240 2375 30243
rect 2746 30240 2774 30348
rect 3142 30336 3148 30348
rect 3200 30376 3206 30388
rect 3200 30348 3924 30376
rect 3200 30336 3206 30348
rect 3596 30311 3654 30317
rect 3596 30277 3608 30311
rect 3642 30308 3654 30311
rect 3786 30308 3792 30320
rect 3642 30280 3792 30308
rect 3642 30277 3654 30280
rect 3596 30271 3654 30277
rect 3786 30268 3792 30280
rect 3844 30268 3850 30320
rect 3896 30308 3924 30348
rect 4614 30336 4620 30388
rect 4672 30376 4678 30388
rect 4709 30379 4767 30385
rect 4709 30376 4721 30379
rect 4672 30348 4721 30376
rect 4672 30336 4678 30348
rect 4709 30345 4721 30348
rect 4755 30345 4767 30379
rect 4709 30339 4767 30345
rect 5442 30336 5448 30388
rect 5500 30336 5506 30388
rect 6822 30336 6828 30388
rect 6880 30336 6886 30388
rect 18322 30336 18328 30388
rect 18380 30376 18386 30388
rect 18690 30376 18696 30388
rect 18380 30348 18696 30376
rect 18380 30336 18386 30348
rect 18690 30336 18696 30348
rect 18748 30336 18754 30388
rect 18782 30336 18788 30388
rect 18840 30376 18846 30388
rect 19334 30376 19340 30388
rect 18840 30348 19340 30376
rect 18840 30336 18846 30348
rect 19334 30336 19340 30348
rect 19392 30336 19398 30388
rect 19797 30379 19855 30385
rect 19797 30345 19809 30379
rect 19843 30376 19855 30379
rect 20346 30376 20352 30388
rect 19843 30348 20352 30376
rect 19843 30345 19855 30348
rect 19797 30339 19855 30345
rect 20346 30336 20352 30348
rect 20404 30336 20410 30388
rect 20530 30336 20536 30388
rect 20588 30376 20594 30388
rect 20588 30348 21864 30376
rect 20588 30336 20594 30348
rect 6733 30311 6791 30317
rect 6733 30308 6745 30311
rect 3896 30280 6745 30308
rect 6733 30277 6745 30280
rect 6779 30308 6791 30311
rect 8294 30308 8300 30320
rect 6779 30280 8300 30308
rect 6779 30277 6791 30280
rect 6733 30271 6791 30277
rect 8294 30268 8300 30280
rect 8352 30268 8358 30320
rect 16022 30268 16028 30320
rect 16080 30268 16086 30320
rect 16114 30268 16120 30320
rect 16172 30308 16178 30320
rect 16172 30280 16252 30308
rect 16172 30268 16178 30280
rect 2363 30212 2774 30240
rect 2961 30243 3019 30249
rect 2363 30209 2375 30212
rect 2317 30203 2375 30209
rect 2961 30209 2973 30243
rect 3007 30240 3019 30243
rect 3050 30240 3056 30252
rect 3007 30212 3056 30240
rect 3007 30209 3019 30212
rect 2961 30203 3019 30209
rect 3050 30200 3056 30212
rect 3108 30200 3114 30252
rect 5629 30243 5687 30249
rect 5629 30209 5641 30243
rect 5675 30240 5687 30243
rect 8196 30243 8254 30249
rect 5675 30212 6408 30240
rect 5675 30209 5687 30212
rect 5629 30203 5687 30209
rect 2406 30132 2412 30184
rect 2464 30172 2470 30184
rect 2501 30175 2559 30181
rect 2501 30172 2513 30175
rect 2464 30144 2513 30172
rect 2464 30132 2470 30144
rect 2501 30141 2513 30144
rect 2547 30141 2559 30175
rect 2501 30135 2559 30141
rect 2516 30104 2544 30135
rect 2590 30132 2596 30184
rect 2648 30172 2654 30184
rect 3329 30175 3387 30181
rect 3329 30172 3341 30175
rect 2648 30144 3341 30172
rect 2648 30132 2654 30144
rect 3329 30141 3341 30144
rect 3375 30141 3387 30175
rect 3329 30135 3387 30141
rect 6380 30113 6408 30212
rect 8196 30209 8208 30243
rect 8242 30240 8254 30243
rect 8570 30240 8576 30252
rect 8242 30212 8576 30240
rect 8242 30209 8254 30212
rect 8196 30203 8254 30209
rect 8570 30200 8576 30212
rect 8628 30200 8634 30252
rect 9950 30200 9956 30252
rect 10008 30240 10014 30252
rect 10321 30243 10379 30249
rect 10321 30240 10333 30243
rect 10008 30212 10333 30240
rect 10008 30200 10014 30212
rect 10321 30209 10333 30212
rect 10367 30209 10379 30243
rect 10321 30203 10379 30209
rect 11974 30200 11980 30252
rect 12032 30200 12038 30252
rect 13633 30243 13691 30249
rect 13633 30240 13645 30243
rect 12406 30212 13645 30240
rect 7009 30175 7067 30181
rect 7009 30141 7021 30175
rect 7055 30172 7067 30175
rect 7650 30172 7656 30184
rect 7055 30144 7656 30172
rect 7055 30141 7067 30144
rect 7009 30135 7067 30141
rect 7650 30132 7656 30144
rect 7708 30132 7714 30184
rect 7929 30175 7987 30181
rect 7929 30172 7941 30175
rect 7760 30144 7941 30172
rect 3145 30107 3203 30113
rect 3145 30104 3157 30107
rect 2516 30076 3157 30104
rect 3145 30073 3157 30076
rect 3191 30073 3203 30107
rect 3145 30067 3203 30073
rect 6365 30107 6423 30113
rect 6365 30073 6377 30107
rect 6411 30073 6423 30107
rect 6365 30067 6423 30073
rect 4798 29996 4804 30048
rect 4856 30036 4862 30048
rect 7760 30036 7788 30144
rect 7929 30141 7941 30144
rect 7975 30141 7987 30175
rect 10045 30175 10103 30181
rect 10045 30172 10057 30175
rect 7929 30135 7987 30141
rect 8956 30144 10057 30172
rect 8956 30036 8984 30144
rect 10045 30141 10057 30144
rect 10091 30141 10103 30175
rect 10045 30135 10103 30141
rect 10060 30104 10088 30135
rect 10502 30132 10508 30184
rect 10560 30172 10566 30184
rect 12406 30172 12434 30212
rect 13633 30209 13645 30212
rect 13679 30240 13691 30243
rect 13679 30212 15884 30240
rect 13679 30209 13691 30212
rect 13633 30203 13691 30209
rect 10560 30144 12434 30172
rect 10560 30132 10566 30144
rect 13722 30132 13728 30184
rect 13780 30132 13786 30184
rect 13817 30175 13875 30181
rect 13817 30141 13829 30175
rect 13863 30141 13875 30175
rect 15856 30172 15884 30212
rect 15930 30200 15936 30252
rect 15988 30200 15994 30252
rect 16224 30240 16252 30280
rect 16482 30268 16488 30320
rect 16540 30308 16546 30320
rect 17129 30311 17187 30317
rect 17129 30308 17141 30311
rect 16540 30280 17141 30308
rect 16540 30268 16546 30280
rect 17129 30277 17141 30280
rect 17175 30277 17187 30311
rect 17129 30271 17187 30277
rect 18049 30311 18107 30317
rect 18049 30277 18061 30311
rect 18095 30308 18107 30311
rect 18800 30308 18828 30336
rect 19978 30308 19984 30320
rect 18095 30280 18828 30308
rect 19444 30280 19984 30308
rect 18095 30277 18107 30280
rect 18049 30271 18107 30277
rect 16298 30240 16304 30252
rect 16224 30212 16304 30240
rect 16114 30172 16120 30184
rect 15856 30144 16120 30172
rect 13817 30135 13875 30141
rect 10686 30104 10692 30116
rect 10060 30076 10692 30104
rect 10686 30064 10692 30076
rect 10744 30064 10750 30116
rect 12710 30064 12716 30116
rect 12768 30104 12774 30116
rect 13265 30107 13323 30113
rect 13265 30104 13277 30107
rect 12768 30076 13277 30104
rect 12768 30064 12774 30076
rect 13265 30073 13277 30076
rect 13311 30073 13323 30107
rect 13832 30104 13860 30135
rect 16114 30132 16120 30144
rect 16172 30132 16178 30184
rect 16224 30181 16252 30212
rect 16298 30200 16304 30212
rect 16356 30200 16362 30252
rect 17034 30200 17040 30252
rect 17092 30200 17098 30252
rect 18693 30243 18751 30249
rect 17144 30212 18644 30240
rect 16209 30175 16267 30181
rect 16209 30141 16221 30175
rect 16255 30141 16267 30175
rect 16209 30135 16267 30141
rect 16390 30132 16396 30184
rect 16448 30172 16454 30184
rect 17144 30172 17172 30212
rect 16448 30144 17172 30172
rect 17313 30175 17371 30181
rect 16448 30132 16454 30144
rect 17313 30141 17325 30175
rect 17359 30172 17371 30175
rect 17678 30172 17684 30184
rect 17359 30144 17684 30172
rect 17359 30141 17371 30144
rect 17313 30135 17371 30141
rect 17678 30132 17684 30144
rect 17736 30132 17742 30184
rect 17954 30132 17960 30184
rect 18012 30172 18018 30184
rect 18506 30172 18512 30184
rect 18012 30144 18512 30172
rect 18012 30132 18018 30144
rect 18506 30132 18512 30144
rect 18564 30132 18570 30184
rect 18616 30172 18644 30212
rect 18693 30209 18705 30243
rect 18739 30240 18751 30243
rect 19444 30240 19472 30280
rect 19978 30268 19984 30280
rect 20036 30268 20042 30320
rect 21726 30308 21732 30320
rect 20916 30280 21732 30308
rect 20916 30252 20944 30280
rect 21726 30268 21732 30280
rect 21784 30268 21790 30320
rect 18739 30212 19472 30240
rect 18739 30209 18751 30212
rect 18693 30203 18751 30209
rect 20898 30200 20904 30252
rect 20956 30200 20962 30252
rect 21358 30200 21364 30252
rect 21416 30200 21422 30252
rect 21545 30243 21603 30249
rect 21545 30209 21557 30243
rect 21591 30209 21603 30243
rect 21545 30203 21603 30209
rect 18874 30172 18880 30184
rect 18616 30144 18880 30172
rect 18874 30132 18880 30144
rect 18932 30132 18938 30184
rect 18966 30132 18972 30184
rect 19024 30132 19030 30184
rect 19334 30132 19340 30184
rect 19392 30132 19398 30184
rect 19886 30132 19892 30184
rect 19944 30172 19950 30184
rect 21560 30172 21588 30203
rect 21634 30200 21640 30252
rect 21692 30200 21698 30252
rect 19944 30144 21588 30172
rect 21744 30172 21772 30268
rect 21836 30249 21864 30348
rect 21910 30336 21916 30388
rect 21968 30376 21974 30388
rect 24946 30376 24952 30388
rect 21968 30348 24952 30376
rect 21968 30336 21974 30348
rect 24946 30336 24952 30348
rect 25004 30336 25010 30388
rect 25130 30336 25136 30388
rect 25188 30376 25194 30388
rect 31662 30376 31668 30388
rect 25188 30348 31668 30376
rect 25188 30336 25194 30348
rect 31662 30336 31668 30348
rect 31720 30336 31726 30388
rect 31941 30379 31999 30385
rect 31941 30345 31953 30379
rect 31987 30345 31999 30379
rect 31941 30339 31999 30345
rect 30834 30317 30840 30320
rect 30828 30308 30840 30317
rect 25240 30280 27384 30308
rect 30795 30280 30840 30308
rect 21821 30243 21879 30249
rect 21821 30209 21833 30243
rect 21867 30240 21879 30243
rect 21910 30240 21916 30252
rect 21867 30212 21916 30240
rect 21867 30209 21879 30212
rect 21821 30203 21879 30209
rect 21910 30200 21916 30212
rect 21968 30200 21974 30252
rect 23017 30243 23075 30249
rect 23017 30240 23029 30243
rect 22480 30212 23029 30240
rect 22480 30184 22508 30212
rect 23017 30209 23029 30212
rect 23063 30209 23075 30243
rect 23017 30203 23075 30209
rect 23477 30243 23535 30249
rect 23477 30209 23489 30243
rect 23523 30240 23535 30243
rect 23566 30240 23572 30252
rect 23523 30212 23572 30240
rect 23523 30209 23535 30212
rect 23477 30203 23535 30209
rect 23566 30200 23572 30212
rect 23624 30240 23630 30252
rect 23624 30212 23888 30240
rect 23624 30200 23630 30212
rect 22097 30175 22155 30181
rect 22097 30172 22109 30175
rect 21744 30144 22109 30172
rect 19944 30132 19950 30144
rect 22097 30141 22109 30144
rect 22143 30172 22155 30175
rect 22462 30172 22468 30184
rect 22143 30144 22468 30172
rect 22143 30141 22155 30144
rect 22097 30135 22155 30141
rect 22462 30132 22468 30144
rect 22520 30132 22526 30184
rect 23661 30175 23719 30181
rect 23661 30141 23673 30175
rect 23707 30172 23719 30175
rect 23750 30172 23756 30184
rect 23707 30144 23756 30172
rect 23707 30141 23719 30144
rect 23661 30135 23719 30141
rect 23750 30132 23756 30144
rect 23808 30132 23814 30184
rect 23860 30172 23888 30212
rect 24394 30200 24400 30252
rect 24452 30200 24458 30252
rect 24578 30249 24584 30252
rect 24535 30243 24584 30249
rect 24535 30209 24547 30243
rect 24581 30209 24584 30243
rect 24535 30203 24584 30209
rect 24578 30200 24584 30203
rect 24636 30200 24642 30252
rect 24210 30172 24216 30184
rect 23860 30144 24216 30172
rect 24210 30132 24216 30144
rect 24268 30132 24274 30184
rect 24670 30132 24676 30184
rect 24728 30132 24734 30184
rect 13265 30067 13323 30073
rect 13740 30076 13860 30104
rect 4856 30008 8984 30036
rect 4856 29996 4862 30008
rect 9306 29996 9312 30048
rect 9364 29996 9370 30048
rect 11606 29996 11612 30048
rect 11664 30036 11670 30048
rect 11793 30039 11851 30045
rect 11793 30036 11805 30039
rect 11664 30008 11805 30036
rect 11664 29996 11670 30008
rect 11793 30005 11805 30008
rect 11839 30005 11851 30039
rect 11793 29999 11851 30005
rect 13170 29996 13176 30048
rect 13228 30036 13234 30048
rect 13630 30036 13636 30048
rect 13228 30008 13636 30036
rect 13228 29996 13234 30008
rect 13630 29996 13636 30008
rect 13688 30036 13694 30048
rect 13740 30036 13768 30076
rect 13998 30064 14004 30116
rect 14056 30104 14062 30116
rect 14056 30076 19196 30104
rect 14056 30064 14062 30076
rect 13688 30008 13768 30036
rect 13688 29996 13694 30008
rect 15378 29996 15384 30048
rect 15436 30036 15442 30048
rect 15565 30039 15623 30045
rect 15565 30036 15577 30039
rect 15436 30008 15577 30036
rect 15436 29996 15442 30008
rect 15565 30005 15577 30008
rect 15611 30005 15623 30039
rect 15565 29999 15623 30005
rect 15654 29996 15660 30048
rect 15712 30036 15718 30048
rect 16669 30039 16727 30045
rect 16669 30036 16681 30039
rect 15712 30008 16681 30036
rect 15712 29996 15718 30008
rect 16669 30005 16681 30008
rect 16715 30005 16727 30039
rect 16669 29999 16727 30005
rect 17034 29996 17040 30048
rect 17092 30036 17098 30048
rect 18138 30036 18144 30048
rect 17092 30008 18144 30036
rect 17092 29996 17098 30008
rect 18138 29996 18144 30008
rect 18196 29996 18202 30048
rect 18325 30039 18383 30045
rect 18325 30005 18337 30039
rect 18371 30036 18383 30039
rect 18414 30036 18420 30048
rect 18371 30008 18420 30036
rect 18371 30005 18383 30008
rect 18325 29999 18383 30005
rect 18414 29996 18420 30008
rect 18472 29996 18478 30048
rect 18506 29996 18512 30048
rect 18564 30036 18570 30048
rect 18782 30036 18788 30048
rect 18564 30008 18788 30036
rect 18564 29996 18570 30008
rect 18782 29996 18788 30008
rect 18840 30036 18846 30048
rect 19058 30036 19064 30048
rect 18840 30008 19064 30036
rect 18840 29996 18846 30008
rect 19058 29996 19064 30008
rect 19116 29996 19122 30048
rect 19168 30036 19196 30076
rect 19242 30064 19248 30116
rect 19300 30104 19306 30116
rect 19613 30107 19671 30113
rect 19300 30076 19472 30104
rect 19300 30064 19306 30076
rect 19334 30036 19340 30048
rect 19168 30008 19340 30036
rect 19334 29996 19340 30008
rect 19392 29996 19398 30048
rect 19444 30036 19472 30076
rect 19613 30073 19625 30107
rect 19659 30073 19671 30107
rect 19613 30067 19671 30073
rect 19628 30036 19656 30067
rect 23842 30064 23848 30116
rect 23900 30104 23906 30116
rect 24121 30107 24179 30113
rect 24121 30104 24133 30107
rect 23900 30076 24133 30104
rect 23900 30064 23906 30076
rect 24121 30073 24133 30076
rect 24167 30073 24179 30107
rect 24121 30067 24179 30073
rect 19444 30008 19656 30036
rect 20993 30039 21051 30045
rect 20993 30005 21005 30039
rect 21039 30036 21051 30039
rect 21082 30036 21088 30048
rect 21039 30008 21088 30036
rect 21039 30005 21051 30008
rect 20993 29999 21051 30005
rect 21082 29996 21088 30008
rect 21140 29996 21146 30048
rect 21174 29996 21180 30048
rect 21232 29996 21238 30048
rect 23201 30039 23259 30045
rect 23201 30005 23213 30039
rect 23247 30036 23259 30039
rect 25240 30036 25268 30280
rect 25314 30200 25320 30252
rect 25372 30240 25378 30252
rect 25777 30243 25835 30249
rect 25777 30240 25789 30243
rect 25372 30212 25789 30240
rect 25372 30200 25378 30212
rect 25777 30209 25789 30212
rect 25823 30209 25835 30243
rect 25777 30203 25835 30209
rect 25866 30200 25872 30252
rect 25924 30200 25930 30252
rect 26145 30243 26203 30249
rect 26145 30209 26157 30243
rect 26191 30209 26203 30243
rect 26145 30203 26203 30209
rect 25406 30132 25412 30184
rect 25464 30172 25470 30184
rect 26160 30172 26188 30203
rect 26786 30200 26792 30252
rect 26844 30200 26850 30252
rect 26973 30243 27031 30249
rect 27240 30244 27298 30249
rect 26973 30240 26985 30243
rect 26896 30212 26985 30240
rect 25464 30144 26188 30172
rect 25464 30132 25470 30144
rect 26234 30132 26240 30184
rect 26292 30172 26298 30184
rect 26896 30172 26924 30212
rect 26973 30209 26985 30212
rect 27019 30209 27031 30243
rect 27172 30243 27298 30244
rect 27172 30240 27252 30243
rect 26973 30203 27031 30209
rect 27080 30216 27252 30240
rect 27080 30212 27200 30216
rect 27080 30172 27108 30212
rect 27240 30209 27252 30216
rect 27286 30209 27298 30243
rect 27356 30240 27384 30280
rect 30828 30271 30840 30280
rect 30834 30268 30840 30271
rect 30892 30268 30898 30320
rect 31956 30308 31984 30339
rect 32030 30336 32036 30388
rect 32088 30376 32094 30388
rect 32766 30376 32772 30388
rect 32088 30348 32772 30376
rect 32088 30336 32094 30348
rect 32766 30336 32772 30348
rect 32824 30336 32830 30388
rect 33318 30336 33324 30388
rect 33376 30376 33382 30388
rect 34422 30376 34428 30388
rect 33376 30348 34428 30376
rect 33376 30336 33382 30348
rect 34422 30336 34428 30348
rect 34480 30336 34486 30388
rect 34698 30336 34704 30388
rect 34756 30376 34762 30388
rect 38749 30379 38807 30385
rect 38749 30376 38761 30379
rect 34756 30348 38761 30376
rect 34756 30336 34762 30348
rect 38749 30345 38761 30348
rect 38795 30345 38807 30379
rect 40773 30379 40831 30385
rect 40773 30376 40785 30379
rect 38749 30339 38807 30345
rect 38856 30348 40785 30376
rect 31956 30280 32352 30308
rect 28074 30240 28080 30252
rect 27356 30212 28080 30240
rect 27240 30203 27298 30209
rect 28074 30200 28080 30212
rect 28132 30200 28138 30252
rect 29730 30200 29736 30252
rect 29788 30240 29794 30252
rect 29788 30212 31754 30240
rect 29788 30200 29794 30212
rect 26292 30144 26924 30172
rect 26988 30144 27108 30172
rect 28092 30172 28120 30200
rect 30374 30172 30380 30184
rect 28092 30144 30380 30172
rect 26292 30132 26298 30144
rect 25593 30107 25651 30113
rect 25593 30073 25605 30107
rect 25639 30104 25651 30107
rect 26605 30107 26663 30113
rect 25639 30076 26556 30104
rect 25639 30073 25651 30076
rect 25593 30067 25651 30073
rect 23247 30008 25268 30036
rect 25317 30039 25375 30045
rect 23247 30005 23259 30008
rect 23201 29999 23259 30005
rect 25317 30005 25329 30039
rect 25363 30036 25375 30039
rect 25498 30036 25504 30048
rect 25363 30008 25504 30036
rect 25363 30005 25375 30008
rect 25317 29999 25375 30005
rect 25498 29996 25504 30008
rect 25556 29996 25562 30048
rect 25682 29996 25688 30048
rect 25740 30036 25746 30048
rect 26053 30039 26111 30045
rect 26053 30036 26065 30039
rect 25740 30008 26065 30036
rect 25740 29996 25746 30008
rect 26053 30005 26065 30008
rect 26099 30005 26111 30039
rect 26528 30036 26556 30076
rect 26605 30073 26617 30107
rect 26651 30104 26663 30107
rect 26988 30104 27016 30144
rect 30374 30132 30380 30144
rect 30432 30132 30438 30184
rect 30558 30132 30564 30184
rect 30616 30132 30622 30184
rect 26651 30076 27016 30104
rect 31726 30104 31754 30212
rect 32122 30200 32128 30252
rect 32180 30200 32186 30252
rect 32324 30240 32352 30280
rect 37274 30268 37280 30320
rect 37332 30308 37338 30320
rect 37369 30311 37427 30317
rect 37369 30308 37381 30311
rect 37332 30280 37381 30308
rect 37332 30268 37338 30280
rect 37369 30277 37381 30280
rect 37415 30277 37427 30311
rect 37369 30271 37427 30277
rect 37458 30268 37464 30320
rect 37516 30308 37522 30320
rect 38197 30311 38255 30317
rect 38197 30308 38209 30311
rect 37516 30280 38209 30308
rect 37516 30268 37522 30280
rect 38197 30277 38209 30280
rect 38243 30277 38255 30311
rect 38197 30271 38255 30277
rect 32324 30212 32536 30240
rect 32306 30132 32312 30184
rect 32364 30132 32370 30184
rect 32508 30172 32536 30212
rect 33134 30200 33140 30252
rect 33192 30249 33198 30252
rect 33192 30243 33220 30249
rect 33208 30209 33220 30243
rect 33192 30203 33220 30209
rect 33192 30200 33198 30203
rect 34698 30200 34704 30252
rect 34756 30240 34762 30252
rect 35066 30240 35072 30252
rect 34756 30212 35072 30240
rect 34756 30200 34762 30212
rect 35066 30200 35072 30212
rect 35124 30200 35130 30252
rect 36357 30243 36415 30249
rect 36357 30209 36369 30243
rect 36403 30240 36415 30243
rect 36446 30240 36452 30252
rect 36403 30212 36452 30240
rect 36403 30209 36415 30212
rect 36357 30203 36415 30209
rect 36446 30200 36452 30212
rect 36504 30200 36510 30252
rect 36541 30243 36599 30249
rect 36541 30209 36553 30243
rect 36587 30209 36599 30243
rect 36541 30203 36599 30209
rect 36633 30243 36691 30249
rect 36633 30209 36645 30243
rect 36679 30240 36691 30243
rect 36998 30240 37004 30252
rect 36679 30212 37004 30240
rect 36679 30209 36691 30212
rect 36633 30203 36691 30209
rect 33042 30172 33048 30184
rect 32508 30144 33048 30172
rect 33042 30132 33048 30144
rect 33100 30132 33106 30184
rect 33318 30132 33324 30184
rect 33376 30132 33382 30184
rect 36556 30172 36584 30203
rect 36998 30200 37004 30212
rect 37056 30200 37062 30252
rect 38378 30200 38384 30252
rect 38436 30200 38442 30252
rect 38657 30243 38715 30249
rect 38657 30209 38669 30243
rect 38703 30240 38715 30243
rect 38856 30240 38884 30348
rect 40773 30345 40785 30348
rect 40819 30345 40831 30379
rect 40773 30339 40831 30345
rect 42245 30379 42303 30385
rect 42245 30345 42257 30379
rect 42291 30345 42303 30379
rect 42245 30339 42303 30345
rect 44913 30379 44971 30385
rect 44913 30345 44925 30379
rect 44959 30376 44971 30379
rect 45370 30376 45376 30388
rect 44959 30348 45376 30376
rect 44959 30345 44971 30348
rect 44913 30339 44971 30345
rect 42260 30308 42288 30339
rect 45370 30336 45376 30348
rect 45428 30336 45434 30388
rect 40880 30280 42288 30308
rect 38703 30212 38884 30240
rect 38933 30243 38991 30249
rect 38703 30209 38715 30212
rect 38657 30203 38715 30209
rect 38933 30209 38945 30243
rect 38979 30240 38991 30243
rect 39114 30240 39120 30252
rect 38979 30212 39120 30240
rect 38979 30209 38991 30212
rect 38933 30203 38991 30209
rect 39114 30200 39120 30212
rect 39172 30200 39178 30252
rect 39209 30243 39267 30249
rect 39209 30209 39221 30243
rect 39255 30240 39267 30243
rect 39298 30240 39304 30252
rect 39255 30212 39304 30240
rect 39255 30209 39267 30212
rect 39209 30203 39267 30209
rect 39298 30200 39304 30212
rect 39356 30200 39362 30252
rect 39390 30200 39396 30252
rect 39448 30200 39454 30252
rect 40034 30200 40040 30252
rect 40092 30240 40098 30252
rect 40221 30243 40279 30249
rect 40221 30240 40233 30243
rect 40092 30212 40233 30240
rect 40092 30200 40098 30212
rect 40221 30209 40233 30212
rect 40267 30209 40279 30243
rect 40221 30203 40279 30209
rect 40310 30200 40316 30252
rect 40368 30240 40374 30252
rect 40405 30243 40463 30249
rect 40405 30240 40417 30243
rect 40368 30212 40417 30240
rect 40368 30200 40374 30212
rect 40405 30209 40417 30212
rect 40451 30209 40463 30243
rect 40405 30203 40463 30209
rect 40494 30200 40500 30252
rect 40552 30200 40558 30252
rect 40589 30243 40647 30249
rect 40589 30209 40601 30243
rect 40635 30209 40647 30243
rect 40589 30203 40647 30209
rect 36556 30144 39436 30172
rect 32769 30107 32827 30113
rect 31726 30076 32076 30104
rect 26651 30073 26663 30076
rect 26605 30067 26663 30073
rect 28258 30036 28264 30048
rect 26528 30008 28264 30036
rect 26053 29999 26111 30005
rect 28258 29996 28264 30008
rect 28316 29996 28322 30048
rect 28350 29996 28356 30048
rect 28408 29996 28414 30048
rect 32048 30036 32076 30076
rect 32769 30073 32781 30107
rect 32815 30104 32827 30107
rect 32858 30104 32864 30116
rect 32815 30076 32864 30104
rect 32815 30073 32827 30076
rect 32769 30067 32827 30073
rect 32858 30064 32864 30076
rect 32916 30064 32922 30116
rect 35618 30064 35624 30116
rect 35676 30104 35682 30116
rect 36354 30104 36360 30116
rect 35676 30076 36360 30104
rect 35676 30064 35682 30076
rect 36354 30064 36360 30076
rect 36412 30104 36418 30116
rect 38565 30107 38623 30113
rect 36412 30076 37320 30104
rect 36412 30064 36418 30076
rect 37292 30048 37320 30076
rect 38565 30073 38577 30107
rect 38611 30073 38623 30107
rect 38565 30067 38623 30073
rect 33965 30039 34023 30045
rect 33965 30036 33977 30039
rect 32048 30008 33977 30036
rect 33965 30005 33977 30008
rect 34011 30005 34023 30039
rect 33965 29999 34023 30005
rect 34054 29996 34060 30048
rect 34112 30036 34118 30048
rect 36173 30039 36231 30045
rect 36173 30036 36185 30039
rect 34112 30008 36185 30036
rect 34112 29996 34118 30008
rect 36173 30005 36185 30008
rect 36219 30005 36231 30039
rect 36173 29999 36231 30005
rect 36446 29996 36452 30048
rect 36504 30036 36510 30048
rect 36906 30036 36912 30048
rect 36504 30008 36912 30036
rect 36504 29996 36510 30008
rect 36906 29996 36912 30008
rect 36964 29996 36970 30048
rect 37274 29996 37280 30048
rect 37332 30036 37338 30048
rect 37461 30039 37519 30045
rect 37461 30036 37473 30039
rect 37332 30008 37473 30036
rect 37332 29996 37338 30008
rect 37461 30005 37473 30008
rect 37507 30036 37519 30039
rect 38010 30036 38016 30048
rect 37507 30008 38016 30036
rect 37507 30005 37519 30008
rect 37461 29999 37519 30005
rect 38010 29996 38016 30008
rect 38068 29996 38074 30048
rect 38580 30036 38608 30067
rect 38930 30064 38936 30116
rect 38988 30104 38994 30116
rect 39025 30107 39083 30113
rect 39025 30104 39037 30107
rect 38988 30076 39037 30104
rect 38988 30064 38994 30076
rect 39025 30073 39037 30076
rect 39071 30073 39083 30107
rect 39025 30067 39083 30073
rect 39114 30064 39120 30116
rect 39172 30064 39178 30116
rect 39408 30104 39436 30144
rect 39482 30132 39488 30184
rect 39540 30132 39546 30184
rect 39666 30132 39672 30184
rect 39724 30132 39730 30184
rect 40129 30175 40187 30181
rect 40129 30141 40141 30175
rect 40175 30172 40187 30175
rect 40604 30172 40632 30203
rect 40175 30144 40632 30172
rect 40175 30141 40187 30144
rect 40129 30135 40187 30141
rect 40880 30104 40908 30280
rect 42334 30268 42340 30320
rect 42392 30308 42398 30320
rect 43349 30311 43407 30317
rect 43349 30308 43361 30311
rect 42392 30280 43361 30308
rect 42392 30268 42398 30280
rect 43349 30277 43361 30280
rect 43395 30277 43407 30311
rect 43349 30271 43407 30277
rect 43640 30280 44772 30308
rect 41598 30200 41604 30252
rect 41656 30200 41662 30252
rect 41782 30249 41788 30252
rect 41749 30243 41788 30249
rect 41749 30209 41761 30243
rect 41749 30203 41788 30209
rect 41782 30200 41788 30203
rect 41840 30200 41846 30252
rect 41877 30243 41935 30249
rect 41877 30209 41889 30243
rect 41923 30209 41935 30243
rect 41877 30203 41935 30209
rect 41969 30243 42027 30249
rect 41969 30209 41981 30243
rect 42015 30209 42027 30243
rect 41969 30203 42027 30209
rect 42107 30243 42165 30249
rect 42107 30209 42119 30243
rect 42153 30240 42165 30243
rect 43073 30243 43131 30249
rect 42153 30212 43024 30240
rect 42153 30209 42165 30212
rect 42107 30203 42165 30209
rect 41230 30132 41236 30184
rect 41288 30172 41294 30184
rect 41892 30172 41920 30203
rect 41288 30144 41920 30172
rect 41288 30132 41294 30144
rect 39408 30076 40908 30104
rect 41046 30064 41052 30116
rect 41104 30104 41110 30116
rect 41984 30104 42012 30203
rect 41104 30076 42012 30104
rect 42996 30104 43024 30212
rect 43073 30209 43085 30243
rect 43119 30240 43131 30243
rect 43162 30240 43168 30252
rect 43119 30212 43168 30240
rect 43119 30209 43131 30212
rect 43073 30203 43131 30209
rect 43162 30200 43168 30212
rect 43220 30200 43226 30252
rect 43640 30249 43668 30280
rect 43625 30243 43683 30249
rect 43625 30209 43637 30243
rect 43671 30209 43683 30243
rect 43625 30203 43683 30209
rect 43714 30200 43720 30252
rect 43772 30240 43778 30252
rect 43901 30243 43959 30249
rect 43901 30240 43913 30243
rect 43772 30212 43913 30240
rect 43772 30200 43778 30212
rect 43901 30209 43913 30212
rect 43947 30209 43959 30243
rect 43901 30203 43959 30209
rect 44082 30200 44088 30252
rect 44140 30200 44146 30252
rect 44177 30243 44235 30249
rect 44177 30209 44189 30243
rect 44223 30209 44235 30243
rect 44177 30203 44235 30209
rect 44192 30172 44220 30203
rect 44266 30200 44272 30252
rect 44324 30200 44330 30252
rect 44450 30200 44456 30252
rect 44508 30240 44514 30252
rect 44744 30249 44772 30280
rect 44729 30243 44787 30249
rect 44508 30212 44680 30240
rect 44508 30200 44514 30212
rect 44361 30175 44419 30181
rect 44361 30172 44373 30175
rect 44192 30144 44373 30172
rect 44361 30141 44373 30144
rect 44407 30172 44419 30175
rect 44545 30175 44603 30181
rect 44545 30172 44557 30175
rect 44407 30144 44557 30172
rect 44407 30141 44419 30144
rect 44361 30135 44419 30141
rect 44545 30141 44557 30144
rect 44591 30141 44603 30175
rect 44652 30172 44680 30212
rect 44729 30209 44741 30243
rect 44775 30209 44787 30243
rect 44729 30203 44787 30209
rect 45005 30243 45063 30249
rect 45005 30209 45017 30243
rect 45051 30240 45063 30243
rect 45370 30240 45376 30252
rect 45051 30212 45376 30240
rect 45051 30209 45063 30212
rect 45005 30203 45063 30209
rect 45370 30200 45376 30212
rect 45428 30200 45434 30252
rect 45649 30243 45707 30249
rect 45649 30209 45661 30243
rect 45695 30240 45707 30243
rect 45922 30240 45928 30252
rect 45695 30212 45928 30240
rect 45695 30209 45707 30212
rect 45649 30203 45707 30209
rect 45922 30200 45928 30212
rect 45980 30200 45986 30252
rect 44910 30172 44916 30184
rect 44652 30144 44916 30172
rect 44545 30135 44603 30141
rect 44910 30132 44916 30144
rect 44968 30172 44974 30184
rect 45097 30175 45155 30181
rect 45097 30172 45109 30175
rect 44968 30144 45109 30172
rect 44968 30132 44974 30144
rect 45097 30141 45109 30144
rect 45143 30141 45155 30175
rect 45833 30175 45891 30181
rect 45097 30135 45155 30141
rect 45204 30144 45508 30172
rect 45204 30104 45232 30144
rect 42996 30076 45232 30104
rect 41104 30064 41110 30076
rect 45278 30064 45284 30116
rect 45336 30104 45342 30116
rect 45373 30107 45431 30113
rect 45373 30104 45385 30107
rect 45336 30076 45385 30104
rect 45336 30064 45342 30076
rect 45373 30073 45385 30076
rect 45419 30073 45431 30107
rect 45480 30104 45508 30144
rect 45833 30141 45845 30175
rect 45879 30172 45891 30175
rect 46198 30172 46204 30184
rect 45879 30144 46204 30172
rect 45879 30141 45891 30144
rect 45833 30135 45891 30141
rect 46198 30132 46204 30144
rect 46256 30132 46262 30184
rect 46017 30107 46075 30113
rect 46017 30104 46029 30107
rect 45480 30076 46029 30104
rect 45373 30067 45431 30073
rect 46017 30073 46029 30076
rect 46063 30073 46075 30107
rect 46017 30067 46075 30073
rect 39942 30036 39948 30048
rect 38580 30008 39948 30036
rect 39942 29996 39948 30008
rect 40000 29996 40006 30048
rect 40862 29996 40868 30048
rect 40920 30036 40926 30048
rect 42150 30036 42156 30048
rect 40920 30008 42156 30036
rect 40920 29996 40926 30008
rect 42150 29996 42156 30008
rect 42208 29996 42214 30048
rect 43898 29996 43904 30048
rect 43956 29996 43962 30048
rect 45462 29996 45468 30048
rect 45520 30036 45526 30048
rect 45557 30039 45615 30045
rect 45557 30036 45569 30039
rect 45520 30008 45569 30036
rect 45520 29996 45526 30008
rect 45557 30005 45569 30008
rect 45603 30005 45615 30039
rect 45557 29999 45615 30005
rect 1104 29946 47104 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 47104 29946
rect 1104 29872 47104 29894
rect 8570 29792 8576 29844
rect 8628 29792 8634 29844
rect 17034 29792 17040 29844
rect 17092 29832 17098 29844
rect 17129 29835 17187 29841
rect 17129 29832 17141 29835
rect 17092 29804 17141 29832
rect 17092 29792 17098 29804
rect 17129 29801 17141 29804
rect 17175 29801 17187 29835
rect 19702 29832 19708 29844
rect 17129 29795 17187 29801
rect 17997 29804 19708 29832
rect 5258 29724 5264 29776
rect 5316 29764 5322 29776
rect 9306 29764 9312 29776
rect 5316 29736 9312 29764
rect 5316 29724 5322 29736
rect 9306 29724 9312 29736
rect 9364 29764 9370 29776
rect 17871 29767 17929 29773
rect 9364 29736 9904 29764
rect 9364 29724 9370 29736
rect 1670 29656 1676 29708
rect 1728 29656 1734 29708
rect 6822 29656 6828 29708
rect 6880 29696 6886 29708
rect 7101 29699 7159 29705
rect 7101 29696 7113 29699
rect 6880 29668 7113 29696
rect 6880 29656 6886 29668
rect 7101 29665 7113 29668
rect 7147 29665 7159 29699
rect 7101 29659 7159 29665
rect 7285 29699 7343 29705
rect 7285 29665 7297 29699
rect 7331 29696 7343 29699
rect 7466 29696 7472 29708
rect 7331 29668 7472 29696
rect 7331 29665 7343 29668
rect 7285 29659 7343 29665
rect 7466 29656 7472 29668
rect 7524 29696 7530 29708
rect 9876 29705 9904 29736
rect 17871 29733 17883 29767
rect 17917 29764 17929 29767
rect 17997 29764 18025 29804
rect 19702 29792 19708 29804
rect 19760 29792 19766 29844
rect 20714 29792 20720 29844
rect 20772 29792 20778 29844
rect 21174 29792 21180 29844
rect 21232 29832 21238 29844
rect 25406 29832 25412 29844
rect 21232 29804 25412 29832
rect 21232 29792 21238 29804
rect 25406 29792 25412 29804
rect 25464 29792 25470 29844
rect 25682 29792 25688 29844
rect 25740 29792 25746 29844
rect 26786 29792 26792 29844
rect 26844 29832 26850 29844
rect 27157 29835 27215 29841
rect 27157 29832 27169 29835
rect 26844 29804 27169 29832
rect 26844 29792 26850 29804
rect 27157 29801 27169 29804
rect 27203 29801 27215 29835
rect 27157 29795 27215 29801
rect 27338 29792 27344 29844
rect 27396 29832 27402 29844
rect 27798 29832 27804 29844
rect 27396 29804 27804 29832
rect 27396 29792 27402 29804
rect 27798 29792 27804 29804
rect 27856 29792 27862 29844
rect 28258 29792 28264 29844
rect 28316 29832 28322 29844
rect 31478 29832 31484 29844
rect 28316 29804 31484 29832
rect 28316 29792 28322 29804
rect 31478 29792 31484 29804
rect 31536 29792 31542 29844
rect 38562 29792 38568 29844
rect 38620 29792 38626 29844
rect 39025 29835 39083 29841
rect 39025 29801 39037 29835
rect 39071 29832 39083 29835
rect 39666 29832 39672 29844
rect 39071 29804 39672 29832
rect 39071 29801 39083 29804
rect 39025 29795 39083 29801
rect 39666 29792 39672 29804
rect 39724 29792 39730 29844
rect 39942 29792 39948 29844
rect 40000 29832 40006 29844
rect 40678 29832 40684 29844
rect 40000 29804 40684 29832
rect 40000 29792 40006 29804
rect 40678 29792 40684 29804
rect 40736 29792 40742 29844
rect 40773 29835 40831 29841
rect 40773 29801 40785 29835
rect 40819 29832 40831 29835
rect 40819 29804 41414 29832
rect 40819 29801 40831 29804
rect 40773 29795 40831 29801
rect 17917 29736 18025 29764
rect 19061 29767 19119 29773
rect 17917 29733 17929 29736
rect 17871 29727 17929 29733
rect 19061 29733 19073 29767
rect 19107 29764 19119 29767
rect 20533 29767 20591 29773
rect 20533 29764 20545 29767
rect 19107 29736 20545 29764
rect 19107 29733 19119 29736
rect 19061 29727 19119 29733
rect 20533 29733 20545 29736
rect 20579 29733 20591 29767
rect 20533 29727 20591 29733
rect 23753 29767 23811 29773
rect 23753 29733 23765 29767
rect 23799 29764 23811 29767
rect 25314 29764 25320 29776
rect 23799 29736 25320 29764
rect 23799 29733 23811 29736
rect 23753 29727 23811 29733
rect 25314 29724 25320 29736
rect 25372 29724 25378 29776
rect 25498 29724 25504 29776
rect 25556 29724 25562 29776
rect 26142 29724 26148 29776
rect 26200 29764 26206 29776
rect 29365 29767 29423 29773
rect 29365 29764 29377 29767
rect 26200 29736 29377 29764
rect 26200 29724 26206 29736
rect 29365 29733 29377 29736
rect 29411 29764 29423 29767
rect 29411 29736 29592 29764
rect 29411 29733 29423 29736
rect 29365 29727 29423 29733
rect 7837 29699 7895 29705
rect 7837 29696 7849 29699
rect 7524 29668 7849 29696
rect 7524 29656 7530 29668
rect 7837 29665 7849 29668
rect 7883 29665 7895 29699
rect 7837 29659 7895 29665
rect 9861 29699 9919 29705
rect 9861 29665 9873 29699
rect 9907 29665 9919 29699
rect 9861 29659 9919 29665
rect 10045 29699 10103 29705
rect 10045 29665 10057 29699
rect 10091 29696 10103 29699
rect 10226 29696 10232 29708
rect 10091 29668 10232 29696
rect 10091 29665 10103 29668
rect 10045 29659 10103 29665
rect 10226 29656 10232 29668
rect 10284 29656 10290 29708
rect 10318 29656 10324 29708
rect 10376 29696 10382 29708
rect 10413 29699 10471 29705
rect 10413 29696 10425 29699
rect 10376 29668 10425 29696
rect 10376 29656 10382 29668
rect 10413 29665 10425 29668
rect 10459 29665 10471 29699
rect 10413 29659 10471 29665
rect 10686 29656 10692 29708
rect 10744 29656 10750 29708
rect 15102 29656 15108 29708
rect 15160 29696 15166 29708
rect 15160 29668 15792 29696
rect 15160 29656 15166 29668
rect 934 29588 940 29640
rect 992 29628 998 29640
rect 1397 29631 1455 29637
rect 1397 29628 1409 29631
rect 992 29600 1409 29628
rect 992 29588 998 29600
rect 1397 29597 1409 29600
rect 1443 29597 1455 29631
rect 1397 29591 1455 29597
rect 5629 29631 5687 29637
rect 5629 29597 5641 29631
rect 5675 29628 5687 29631
rect 6362 29628 6368 29640
rect 5675 29600 6368 29628
rect 5675 29597 5687 29600
rect 5629 29591 5687 29597
rect 6362 29588 6368 29600
rect 6420 29588 6426 29640
rect 7009 29631 7067 29637
rect 7009 29597 7021 29631
rect 7055 29628 7067 29631
rect 8294 29628 8300 29640
rect 7055 29600 8300 29628
rect 7055 29597 7067 29600
rect 7009 29591 7067 29597
rect 8294 29588 8300 29600
rect 8352 29588 8358 29640
rect 8757 29631 8815 29637
rect 8757 29597 8769 29631
rect 8803 29628 8815 29631
rect 9769 29631 9827 29637
rect 8803 29600 9444 29628
rect 8803 29597 8815 29600
rect 8757 29591 8815 29597
rect 7650 29520 7656 29572
rect 7708 29520 7714 29572
rect 5442 29452 5448 29504
rect 5500 29452 5506 29504
rect 6641 29495 6699 29501
rect 6641 29461 6653 29495
rect 6687 29492 6699 29495
rect 6914 29492 6920 29504
rect 6687 29464 6920 29492
rect 6687 29461 6699 29464
rect 6641 29455 6699 29461
rect 6914 29452 6920 29464
rect 6972 29452 6978 29504
rect 9416 29501 9444 29600
rect 9769 29597 9781 29631
rect 9815 29628 9827 29631
rect 10502 29628 10508 29640
rect 9815 29600 10508 29628
rect 9815 29597 9827 29600
rect 9769 29591 9827 29597
rect 10502 29588 10508 29600
rect 10560 29588 10566 29640
rect 11606 29637 11612 29640
rect 11333 29631 11391 29637
rect 11333 29597 11345 29631
rect 11379 29597 11391 29631
rect 11600 29628 11612 29637
rect 11567 29600 11612 29628
rect 11333 29591 11391 29597
rect 11600 29591 11612 29600
rect 11348 29560 11376 29591
rect 11606 29588 11612 29591
rect 11664 29588 11670 29640
rect 15378 29588 15384 29640
rect 15436 29588 15442 29640
rect 15654 29588 15660 29640
rect 15712 29588 15718 29640
rect 15764 29637 15792 29668
rect 16758 29656 16764 29708
rect 16816 29696 16822 29708
rect 17218 29696 17224 29708
rect 16816 29668 17224 29696
rect 16816 29656 16822 29668
rect 17218 29656 17224 29668
rect 17276 29656 17282 29708
rect 17770 29696 17776 29708
rect 17328 29668 17776 29696
rect 15749 29631 15807 29637
rect 15749 29597 15761 29631
rect 15795 29628 15807 29631
rect 17328 29628 17356 29668
rect 17770 29656 17776 29668
rect 17828 29656 17834 29708
rect 17954 29656 17960 29708
rect 18012 29696 18018 29708
rect 18138 29696 18144 29708
rect 18012 29668 18144 29696
rect 18012 29656 18018 29668
rect 18138 29656 18144 29668
rect 18196 29656 18202 29708
rect 18417 29699 18475 29705
rect 18417 29665 18429 29699
rect 18463 29696 18475 29699
rect 19886 29696 19892 29708
rect 18463 29668 19892 29696
rect 18463 29665 18475 29668
rect 18417 29659 18475 29665
rect 19886 29656 19892 29668
rect 19944 29656 19950 29708
rect 20438 29656 20444 29708
rect 20496 29696 20502 29708
rect 21082 29696 21088 29708
rect 20496 29668 21088 29696
rect 20496 29656 20502 29668
rect 21082 29656 21088 29668
rect 21140 29656 21146 29708
rect 21450 29656 21456 29708
rect 21508 29656 21514 29708
rect 22189 29699 22247 29705
rect 22189 29665 22201 29699
rect 22235 29696 22247 29699
rect 27338 29696 27344 29708
rect 22235 29668 27344 29696
rect 22235 29665 22247 29668
rect 22189 29659 22247 29665
rect 27338 29656 27344 29668
rect 27396 29656 27402 29708
rect 27522 29656 27528 29708
rect 27580 29696 27586 29708
rect 29564 29705 29592 29736
rect 37734 29724 37740 29776
rect 37792 29764 37798 29776
rect 39298 29764 39304 29776
rect 37792 29736 39304 29764
rect 37792 29724 37798 29736
rect 39298 29724 39304 29736
rect 39356 29724 39362 29776
rect 39577 29767 39635 29773
rect 39577 29733 39589 29767
rect 39623 29764 39635 29767
rect 40034 29764 40040 29776
rect 39623 29736 40040 29764
rect 39623 29733 39635 29736
rect 39577 29727 39635 29733
rect 40034 29724 40040 29736
rect 40092 29724 40098 29776
rect 41138 29764 41144 29776
rect 40604 29736 41144 29764
rect 27709 29699 27767 29705
rect 27709 29696 27721 29699
rect 27580 29668 27721 29696
rect 27580 29656 27586 29668
rect 27709 29665 27721 29668
rect 27755 29665 27767 29699
rect 27709 29659 27767 29665
rect 29549 29699 29607 29705
rect 29549 29665 29561 29699
rect 29595 29665 29607 29699
rect 38749 29699 38807 29705
rect 29549 29659 29607 29665
rect 30576 29668 35756 29696
rect 15795 29600 17356 29628
rect 15795 29597 15807 29600
rect 15749 29591 15807 29597
rect 17402 29588 17408 29640
rect 17460 29588 17466 29640
rect 18322 29637 18328 29640
rect 18279 29631 18328 29637
rect 18279 29597 18291 29631
rect 18325 29597 18328 29631
rect 18279 29591 18328 29597
rect 18322 29588 18328 29591
rect 18380 29588 18386 29640
rect 18984 29600 20392 29628
rect 15102 29560 15108 29572
rect 11348 29532 15108 29560
rect 15102 29520 15108 29532
rect 15160 29520 15166 29572
rect 15994 29563 16052 29569
rect 15994 29560 16006 29563
rect 15488 29532 16006 29560
rect 9401 29495 9459 29501
rect 9401 29461 9413 29495
rect 9447 29461 9459 29495
rect 9401 29455 9459 29461
rect 12618 29452 12624 29504
rect 12676 29492 12682 29504
rect 12713 29495 12771 29501
rect 12713 29492 12725 29495
rect 12676 29464 12725 29492
rect 12676 29452 12682 29464
rect 12713 29461 12725 29464
rect 12759 29461 12771 29495
rect 12713 29455 12771 29461
rect 15194 29452 15200 29504
rect 15252 29452 15258 29504
rect 15488 29501 15516 29532
rect 15994 29529 16006 29532
rect 16040 29529 16052 29563
rect 15994 29523 16052 29529
rect 15473 29495 15531 29501
rect 15473 29461 15485 29495
rect 15519 29461 15531 29495
rect 15473 29455 15531 29461
rect 16114 29452 16120 29504
rect 16172 29492 16178 29504
rect 18322 29492 18328 29504
rect 16172 29464 18328 29492
rect 16172 29452 16178 29464
rect 18322 29452 18328 29464
rect 18380 29492 18386 29504
rect 18506 29492 18512 29504
rect 18380 29464 18512 29492
rect 18380 29452 18386 29464
rect 18506 29452 18512 29464
rect 18564 29452 18570 29504
rect 18874 29452 18880 29504
rect 18932 29492 18938 29504
rect 18984 29492 19012 29600
rect 20257 29563 20315 29569
rect 20257 29529 20269 29563
rect 20303 29529 20315 29563
rect 20364 29560 20392 29600
rect 20898 29588 20904 29640
rect 20956 29588 20962 29640
rect 21174 29588 21180 29640
rect 21232 29628 21238 29640
rect 21468 29628 21496 29656
rect 21232 29600 21496 29628
rect 21232 29588 21238 29600
rect 21910 29588 21916 29640
rect 21968 29588 21974 29640
rect 22462 29588 22468 29640
rect 22520 29588 22526 29640
rect 22646 29588 22652 29640
rect 22704 29628 22710 29640
rect 23474 29628 23480 29640
rect 22704 29600 23480 29628
rect 22704 29588 22710 29600
rect 23474 29588 23480 29600
rect 23532 29628 23538 29640
rect 23569 29631 23627 29637
rect 23569 29628 23581 29631
rect 23532 29600 23581 29628
rect 23532 29588 23538 29600
rect 23569 29597 23581 29600
rect 23615 29597 23627 29631
rect 27617 29631 27675 29637
rect 23569 29591 23627 29597
rect 23676 29600 25360 29628
rect 20364 29532 21128 29560
rect 20257 29523 20315 29529
rect 18932 29464 19012 29492
rect 20272 29492 20300 29523
rect 20898 29492 20904 29504
rect 20272 29464 20904 29492
rect 18932 29452 18938 29464
rect 20898 29452 20904 29464
rect 20956 29492 20962 29504
rect 20993 29495 21051 29501
rect 20993 29492 21005 29495
rect 20956 29464 21005 29492
rect 20956 29452 20962 29464
rect 20993 29461 21005 29464
rect 21039 29461 21051 29495
rect 21100 29492 21128 29532
rect 21450 29520 21456 29572
rect 21508 29520 21514 29572
rect 23676 29560 23704 29600
rect 22066 29532 23704 29560
rect 22066 29492 22094 29532
rect 24946 29520 24952 29572
rect 25004 29560 25010 29572
rect 25222 29560 25228 29572
rect 25004 29532 25228 29560
rect 25004 29520 25010 29532
rect 25222 29520 25228 29532
rect 25280 29520 25286 29572
rect 25332 29560 25360 29600
rect 27617 29597 27629 29631
rect 27663 29628 27675 29631
rect 28902 29628 28908 29640
rect 27663 29600 28908 29628
rect 27663 29597 27675 29600
rect 27617 29591 27675 29597
rect 28902 29588 28908 29600
rect 28960 29588 28966 29640
rect 29086 29588 29092 29640
rect 29144 29628 29150 29640
rect 29181 29631 29239 29637
rect 29181 29628 29193 29631
rect 29144 29600 29193 29628
rect 29144 29588 29150 29600
rect 29181 29597 29193 29600
rect 29227 29628 29239 29631
rect 29454 29628 29460 29640
rect 29227 29600 29460 29628
rect 29227 29597 29239 29600
rect 29181 29591 29239 29597
rect 29454 29588 29460 29600
rect 29512 29588 29518 29640
rect 30576 29628 30604 29668
rect 29748 29600 30604 29628
rect 29748 29560 29776 29600
rect 35434 29588 35440 29640
rect 35492 29588 35498 29640
rect 35618 29588 35624 29640
rect 35676 29588 35682 29640
rect 35728 29637 35756 29668
rect 38749 29665 38761 29699
rect 38795 29696 38807 29699
rect 38795 29668 39252 29696
rect 38795 29665 38807 29668
rect 38749 29659 38807 29665
rect 35713 29631 35771 29637
rect 35713 29597 35725 29631
rect 35759 29597 35771 29631
rect 35713 29591 35771 29597
rect 35805 29631 35863 29637
rect 35805 29597 35817 29631
rect 35851 29628 35863 29631
rect 35986 29628 35992 29640
rect 35851 29600 35992 29628
rect 35851 29597 35863 29600
rect 35805 29591 35863 29597
rect 35986 29588 35992 29600
rect 36044 29588 36050 29640
rect 37090 29588 37096 29640
rect 37148 29628 37154 29640
rect 37148 29600 38148 29628
rect 37148 29588 37154 29600
rect 25332 29532 29776 29560
rect 29816 29563 29874 29569
rect 29816 29529 29828 29563
rect 29862 29560 29874 29563
rect 30006 29560 30012 29572
rect 29862 29532 30012 29560
rect 29862 29529 29874 29532
rect 29816 29523 29874 29529
rect 30006 29520 30012 29532
rect 30064 29520 30070 29572
rect 31570 29520 31576 29572
rect 31628 29560 31634 29572
rect 34054 29560 34060 29572
rect 31628 29532 34060 29560
rect 31628 29520 31634 29532
rect 34054 29520 34060 29532
rect 34112 29520 34118 29572
rect 36630 29560 36636 29572
rect 34164 29532 36636 29560
rect 21100 29464 22094 29492
rect 20993 29455 21051 29461
rect 22278 29452 22284 29504
rect 22336 29492 22342 29504
rect 22554 29492 22560 29504
rect 22336 29464 22560 29492
rect 22336 29452 22342 29464
rect 22554 29452 22560 29464
rect 22612 29492 22618 29504
rect 22649 29495 22707 29501
rect 22649 29492 22661 29495
rect 22612 29464 22661 29492
rect 22612 29452 22618 29464
rect 22649 29461 22661 29464
rect 22695 29461 22707 29495
rect 22649 29455 22707 29461
rect 24210 29452 24216 29504
rect 24268 29492 24274 29504
rect 27525 29495 27583 29501
rect 27525 29492 27537 29495
rect 24268 29464 27537 29492
rect 24268 29452 24274 29464
rect 27525 29461 27537 29464
rect 27571 29492 27583 29495
rect 28350 29492 28356 29504
rect 27571 29464 28356 29492
rect 27571 29461 27583 29464
rect 27525 29455 27583 29461
rect 28350 29452 28356 29464
rect 28408 29452 28414 29504
rect 29546 29452 29552 29504
rect 29604 29492 29610 29504
rect 30929 29495 30987 29501
rect 30929 29492 30941 29495
rect 29604 29464 30941 29492
rect 29604 29452 29610 29464
rect 30929 29461 30941 29464
rect 30975 29461 30987 29495
rect 30929 29455 30987 29461
rect 33594 29452 33600 29504
rect 33652 29492 33658 29504
rect 34164 29492 34192 29532
rect 36630 29520 36636 29532
rect 36688 29520 36694 29572
rect 37734 29520 37740 29572
rect 37792 29520 37798 29572
rect 38120 29560 38148 29600
rect 38194 29588 38200 29640
rect 38252 29628 38258 29640
rect 39224 29637 39252 29668
rect 38289 29631 38347 29637
rect 38289 29628 38301 29631
rect 38252 29600 38301 29628
rect 38252 29588 38258 29600
rect 38289 29597 38301 29600
rect 38335 29597 38347 29631
rect 38289 29591 38347 29597
rect 39209 29631 39267 29637
rect 39209 29597 39221 29631
rect 39255 29597 39267 29631
rect 39209 29591 39267 29597
rect 39853 29631 39911 29637
rect 39853 29597 39865 29631
rect 39899 29628 39911 29631
rect 40218 29628 40224 29640
rect 39899 29600 40224 29628
rect 39899 29597 39911 29600
rect 39853 29591 39911 29597
rect 40218 29588 40224 29600
rect 40276 29588 40282 29640
rect 40604 29569 40632 29736
rect 41138 29724 41144 29736
rect 41196 29724 41202 29776
rect 41386 29764 41414 29804
rect 42150 29792 42156 29844
rect 42208 29792 42214 29844
rect 44266 29792 44272 29844
rect 44324 29832 44330 29844
rect 45094 29832 45100 29844
rect 44324 29804 45100 29832
rect 44324 29792 44330 29804
rect 45094 29792 45100 29804
rect 45152 29792 45158 29844
rect 45649 29835 45707 29841
rect 45649 29801 45661 29835
rect 45695 29832 45707 29835
rect 46014 29832 46020 29844
rect 45695 29804 46020 29832
rect 45695 29801 45707 29804
rect 45649 29795 45707 29801
rect 46014 29792 46020 29804
rect 46072 29792 46078 29844
rect 42610 29764 42616 29776
rect 41386 29736 42616 29764
rect 42610 29724 42616 29736
rect 42668 29764 42674 29776
rect 43073 29767 43131 29773
rect 42668 29736 42932 29764
rect 42668 29724 42674 29736
rect 40954 29656 40960 29708
rect 41012 29696 41018 29708
rect 41049 29699 41107 29705
rect 41049 29696 41061 29699
rect 41012 29668 41061 29696
rect 41012 29656 41018 29668
rect 41049 29665 41061 29668
rect 41095 29665 41107 29699
rect 42429 29699 42487 29705
rect 42429 29696 42441 29699
rect 41049 29659 41107 29665
rect 42076 29668 42441 29696
rect 42076 29640 42104 29668
rect 42429 29665 42441 29668
rect 42475 29665 42487 29699
rect 42429 29659 42487 29665
rect 42518 29656 42524 29708
rect 42576 29696 42582 29708
rect 42702 29696 42708 29708
rect 42576 29668 42708 29696
rect 42576 29656 42582 29668
rect 42702 29656 42708 29668
rect 42760 29656 42766 29708
rect 40696 29600 41092 29628
rect 39393 29563 39451 29569
rect 39393 29560 39405 29563
rect 38120 29532 39405 29560
rect 39393 29529 39405 29532
rect 39439 29560 39451 29563
rect 40589 29563 40647 29569
rect 39439 29532 40540 29560
rect 39439 29529 39451 29532
rect 39393 29523 39451 29529
rect 33652 29464 34192 29492
rect 35989 29495 36047 29501
rect 33652 29452 33658 29464
rect 35989 29461 36001 29495
rect 36035 29492 36047 29495
rect 36538 29492 36544 29504
rect 36035 29464 36544 29492
rect 36035 29461 36047 29464
rect 35989 29455 36047 29461
rect 36538 29452 36544 29464
rect 36596 29452 36602 29504
rect 37458 29452 37464 29504
rect 37516 29492 37522 29504
rect 37829 29495 37887 29501
rect 37829 29492 37841 29495
rect 37516 29464 37841 29492
rect 37516 29452 37522 29464
rect 37829 29461 37841 29464
rect 37875 29492 37887 29495
rect 38378 29492 38384 29504
rect 37875 29464 38384 29492
rect 37875 29461 37887 29464
rect 37829 29455 37887 29461
rect 38378 29452 38384 29464
rect 38436 29452 38442 29504
rect 38838 29452 38844 29504
rect 38896 29492 38902 29504
rect 39022 29492 39028 29504
rect 38896 29464 39028 29492
rect 38896 29452 38902 29464
rect 39022 29452 39028 29464
rect 39080 29452 39086 29504
rect 40037 29495 40095 29501
rect 40037 29461 40049 29495
rect 40083 29492 40095 29495
rect 40126 29492 40132 29504
rect 40083 29464 40132 29492
rect 40083 29461 40095 29464
rect 40037 29455 40095 29461
rect 40126 29452 40132 29464
rect 40184 29452 40190 29504
rect 40512 29492 40540 29532
rect 40589 29529 40601 29563
rect 40635 29529 40647 29563
rect 40589 29523 40647 29529
rect 40696 29492 40724 29600
rect 40862 29569 40868 29572
rect 40805 29563 40868 29569
rect 40805 29529 40817 29563
rect 40851 29529 40868 29563
rect 40805 29523 40868 29529
rect 40862 29520 40868 29523
rect 40920 29520 40926 29572
rect 41064 29560 41092 29600
rect 41138 29588 41144 29640
rect 41196 29628 41202 29640
rect 41233 29631 41291 29637
rect 41233 29628 41245 29631
rect 41196 29600 41245 29628
rect 41196 29588 41202 29600
rect 41233 29597 41245 29600
rect 41279 29597 41291 29631
rect 41233 29591 41291 29597
rect 41785 29631 41843 29637
rect 41785 29597 41797 29631
rect 41831 29597 41843 29631
rect 41785 29591 41843 29597
rect 41690 29560 41696 29572
rect 41064 29532 41696 29560
rect 41690 29520 41696 29532
rect 41748 29520 41754 29572
rect 41800 29560 41828 29591
rect 42058 29588 42064 29640
rect 42116 29588 42122 29640
rect 42337 29631 42395 29637
rect 42337 29597 42349 29631
rect 42383 29597 42395 29631
rect 42337 29591 42395 29597
rect 42613 29631 42671 29637
rect 42613 29597 42625 29631
rect 42659 29628 42671 29631
rect 42797 29631 42855 29637
rect 42797 29628 42809 29631
rect 42659 29600 42809 29628
rect 42659 29597 42671 29600
rect 42613 29591 42671 29597
rect 42797 29597 42809 29600
rect 42843 29597 42855 29631
rect 42904 29628 42932 29736
rect 43073 29733 43085 29767
rect 43119 29764 43131 29767
rect 43162 29764 43168 29776
rect 43119 29736 43168 29764
rect 43119 29733 43131 29736
rect 43073 29727 43131 29733
rect 43162 29724 43168 29736
rect 43220 29724 43226 29776
rect 44174 29724 44180 29776
rect 44232 29764 44238 29776
rect 46293 29767 46351 29773
rect 46293 29764 46305 29767
rect 44232 29736 46305 29764
rect 44232 29724 44238 29736
rect 46293 29733 46305 29736
rect 46339 29733 46351 29767
rect 46293 29727 46351 29733
rect 43898 29696 43904 29708
rect 43180 29668 43904 29696
rect 42981 29631 43039 29637
rect 42981 29628 42993 29631
rect 42904 29600 42993 29628
rect 42797 29591 42855 29597
rect 42981 29597 42993 29600
rect 43027 29597 43039 29631
rect 42981 29591 43039 29597
rect 41874 29560 41880 29572
rect 41800 29532 41880 29560
rect 41874 29520 41880 29532
rect 41932 29560 41938 29572
rect 42352 29560 42380 29591
rect 43070 29588 43076 29640
rect 43128 29628 43134 29640
rect 43180 29637 43208 29668
rect 43898 29656 43904 29668
rect 43956 29656 43962 29708
rect 45002 29656 45008 29708
rect 45060 29656 45066 29708
rect 45480 29668 46336 29696
rect 45480 29640 45508 29668
rect 43165 29631 43223 29637
rect 43165 29628 43177 29631
rect 43128 29600 43177 29628
rect 43128 29588 43134 29600
rect 43165 29597 43177 29600
rect 43211 29597 43223 29631
rect 43165 29591 43223 29597
rect 43257 29631 43315 29637
rect 43257 29597 43269 29631
rect 43303 29597 43315 29631
rect 43257 29591 43315 29597
rect 41932 29532 42380 29560
rect 41932 29520 41938 29532
rect 42886 29520 42892 29572
rect 42944 29560 42950 29572
rect 43272 29560 43300 29591
rect 44726 29588 44732 29640
rect 44784 29628 44790 29640
rect 45189 29631 45247 29637
rect 45189 29628 45201 29631
rect 44784 29600 45201 29628
rect 44784 29588 44790 29600
rect 45189 29597 45201 29600
rect 45235 29597 45247 29631
rect 45189 29591 45247 29597
rect 45462 29588 45468 29640
rect 45520 29588 45526 29640
rect 45649 29631 45707 29637
rect 45649 29597 45661 29631
rect 45695 29597 45707 29631
rect 45649 29591 45707 29597
rect 42944 29532 43300 29560
rect 42944 29520 42950 29532
rect 45370 29520 45376 29572
rect 45428 29560 45434 29572
rect 45664 29560 45692 29591
rect 46014 29588 46020 29640
rect 46072 29628 46078 29640
rect 46308 29637 46336 29668
rect 46109 29631 46167 29637
rect 46109 29628 46121 29631
rect 46072 29600 46121 29628
rect 46072 29588 46078 29600
rect 46109 29597 46121 29600
rect 46155 29597 46167 29631
rect 46109 29591 46167 29597
rect 46293 29631 46351 29637
rect 46293 29597 46305 29631
rect 46339 29597 46351 29631
rect 46661 29631 46719 29637
rect 46661 29628 46673 29631
rect 46293 29591 46351 29597
rect 46400 29600 46673 29628
rect 46400 29560 46428 29600
rect 46661 29597 46673 29600
rect 46707 29597 46719 29631
rect 46661 29591 46719 29597
rect 45428 29532 46428 29560
rect 45428 29520 45434 29532
rect 40512 29464 40724 29492
rect 40954 29452 40960 29504
rect 41012 29452 41018 29504
rect 41138 29452 41144 29504
rect 41196 29492 41202 29504
rect 41509 29495 41567 29501
rect 41509 29492 41521 29495
rect 41196 29464 41521 29492
rect 41196 29452 41202 29464
rect 41509 29461 41521 29464
rect 41555 29461 41567 29495
rect 41509 29455 41567 29461
rect 45462 29452 45468 29504
rect 45520 29492 45526 29504
rect 45833 29495 45891 29501
rect 45833 29492 45845 29495
rect 45520 29464 45845 29492
rect 45520 29452 45526 29464
rect 45833 29461 45845 29464
rect 45879 29461 45891 29495
rect 45833 29455 45891 29461
rect 1104 29402 47104 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 47104 29402
rect 1104 29328 47104 29350
rect 2406 29248 2412 29300
rect 2464 29288 2470 29300
rect 2464 29260 6316 29288
rect 2464 29248 2470 29260
rect 5068 29223 5126 29229
rect 5068 29189 5080 29223
rect 5114 29220 5126 29223
rect 5442 29220 5448 29232
rect 5114 29192 5448 29220
rect 5114 29189 5126 29192
rect 5068 29183 5126 29189
rect 5442 29180 5448 29192
rect 5500 29180 5506 29232
rect 6288 29220 6316 29260
rect 6362 29248 6368 29300
rect 6420 29248 6426 29300
rect 9030 29248 9036 29300
rect 9088 29288 9094 29300
rect 9585 29291 9643 29297
rect 9585 29288 9597 29291
rect 9088 29260 9597 29288
rect 9088 29248 9094 29260
rect 9585 29257 9597 29260
rect 9631 29257 9643 29291
rect 9585 29251 9643 29257
rect 11517 29291 11575 29297
rect 11517 29257 11529 29291
rect 11563 29257 11575 29291
rect 11517 29251 11575 29257
rect 12437 29291 12495 29297
rect 12437 29257 12449 29291
rect 12483 29288 12495 29291
rect 13173 29291 13231 29297
rect 13173 29288 13185 29291
rect 12483 29260 13185 29288
rect 12483 29257 12495 29260
rect 12437 29251 12495 29257
rect 13173 29257 13185 29260
rect 13219 29288 13231 29291
rect 15470 29288 15476 29300
rect 13219 29260 15476 29288
rect 13219 29257 13231 29260
rect 13173 29251 13231 29257
rect 9398 29220 9404 29232
rect 6288 29192 9404 29220
rect 9398 29180 9404 29192
rect 9456 29180 9462 29232
rect 9950 29220 9956 29232
rect 9600 29192 9956 29220
rect 6730 29112 6736 29164
rect 6788 29112 6794 29164
rect 7650 29152 7656 29164
rect 7024 29124 7656 29152
rect 4614 29044 4620 29096
rect 4672 29084 4678 29096
rect 4798 29084 4804 29096
rect 4672 29056 4804 29084
rect 4672 29044 4678 29056
rect 4798 29044 4804 29056
rect 4856 29044 4862 29096
rect 7024 29093 7052 29124
rect 7650 29112 7656 29124
rect 7708 29112 7714 29164
rect 7834 29161 7840 29164
rect 7828 29115 7840 29161
rect 7834 29112 7840 29115
rect 7892 29112 7898 29164
rect 9306 29112 9312 29164
rect 9364 29152 9370 29164
rect 9493 29155 9551 29161
rect 9493 29152 9505 29155
rect 9364 29124 9505 29152
rect 9364 29112 9370 29124
rect 9493 29121 9505 29124
rect 9539 29121 9551 29155
rect 9493 29115 9551 29121
rect 6825 29087 6883 29093
rect 6825 29053 6837 29087
rect 6871 29053 6883 29087
rect 6825 29047 6883 29053
rect 7009 29087 7067 29093
rect 7009 29053 7021 29087
rect 7055 29053 7067 29087
rect 7009 29047 7067 29053
rect 7561 29087 7619 29093
rect 7561 29053 7573 29087
rect 7607 29053 7619 29087
rect 9600 29084 9628 29192
rect 9950 29180 9956 29192
rect 10008 29180 10014 29232
rect 10220 29223 10278 29229
rect 10220 29189 10232 29223
rect 10266 29220 10278 29223
rect 11532 29220 11560 29251
rect 15470 29248 15476 29260
rect 15528 29248 15534 29300
rect 15930 29248 15936 29300
rect 15988 29288 15994 29300
rect 16485 29291 16543 29297
rect 16485 29288 16497 29291
rect 15988 29260 16497 29288
rect 15988 29248 15994 29260
rect 16485 29257 16497 29260
rect 16531 29257 16543 29291
rect 16485 29251 16543 29257
rect 17402 29248 17408 29300
rect 17460 29288 17466 29300
rect 17460 29260 19104 29288
rect 17460 29248 17466 29260
rect 10266 29192 11560 29220
rect 13464 29192 14228 29220
rect 10266 29189 10278 29192
rect 10220 29183 10278 29189
rect 9784 29124 11008 29152
rect 9784 29093 9812 29124
rect 10980 29096 11008 29124
rect 11054 29112 11060 29164
rect 11112 29152 11118 29164
rect 11701 29155 11759 29161
rect 11701 29152 11713 29155
rect 11112 29124 11713 29152
rect 11112 29112 11118 29124
rect 11701 29121 11713 29124
rect 11747 29121 11759 29155
rect 11701 29115 11759 29121
rect 13078 29112 13084 29164
rect 13136 29112 13142 29164
rect 7561 29047 7619 29053
rect 8588 29056 9628 29084
rect 9769 29087 9827 29093
rect 6181 29019 6239 29025
rect 6181 28985 6193 29019
rect 6227 29016 6239 29019
rect 6840 29016 6868 29047
rect 7282 29016 7288 29028
rect 6227 28988 7288 29016
rect 6227 28985 6239 28988
rect 6181 28979 6239 28985
rect 7282 28976 7288 28988
rect 7340 28976 7346 29028
rect 7576 28948 7604 29047
rect 8588 29016 8616 29056
rect 9769 29053 9781 29087
rect 9815 29053 9827 29087
rect 9769 29047 9827 29053
rect 9950 29044 9956 29096
rect 10008 29044 10014 29096
rect 10962 29044 10968 29096
rect 11020 29084 11026 29096
rect 13357 29087 13415 29093
rect 13357 29084 13369 29087
rect 11020 29056 13369 29084
rect 11020 29044 11026 29056
rect 13357 29053 13369 29056
rect 13403 29084 13415 29087
rect 13464 29084 13492 29192
rect 13808 29155 13866 29161
rect 13808 29121 13820 29155
rect 13854 29152 13866 29155
rect 14090 29152 14096 29164
rect 13854 29124 14096 29152
rect 13854 29121 13866 29124
rect 13808 29115 13866 29121
rect 14090 29112 14096 29124
rect 14148 29112 14154 29164
rect 14200 29152 14228 29192
rect 15194 29180 15200 29232
rect 15252 29220 15258 29232
rect 15350 29223 15408 29229
rect 15350 29220 15362 29223
rect 15252 29192 15362 29220
rect 15252 29180 15258 29192
rect 15350 29189 15362 29192
rect 15396 29189 15408 29223
rect 17494 29220 17500 29232
rect 15350 29183 15408 29189
rect 15488 29192 17500 29220
rect 15488 29152 15516 29192
rect 17494 29180 17500 29192
rect 17552 29180 17558 29232
rect 14200 29124 15516 29152
rect 17218 29112 17224 29164
rect 17276 29152 17282 29164
rect 17604 29161 17632 29260
rect 19076 29220 19104 29260
rect 19242 29248 19248 29300
rect 19300 29248 19306 29300
rect 20717 29291 20775 29297
rect 20717 29257 20729 29291
rect 20763 29257 20775 29291
rect 20717 29251 20775 29257
rect 29181 29291 29239 29297
rect 29181 29257 29193 29291
rect 29227 29257 29239 29291
rect 36725 29291 36783 29297
rect 36725 29288 36737 29291
rect 29181 29251 29239 29257
rect 35912 29260 36737 29288
rect 19978 29220 19984 29232
rect 19076 29192 19984 29220
rect 19978 29180 19984 29192
rect 20036 29220 20042 29232
rect 20732 29220 20760 29251
rect 20036 29192 20760 29220
rect 29196 29220 29224 29251
rect 29196 29192 30236 29220
rect 20036 29180 20042 29192
rect 18506 29161 18512 29164
rect 17405 29155 17463 29161
rect 17405 29152 17417 29155
rect 17276 29124 17417 29152
rect 17276 29112 17282 29124
rect 17405 29121 17417 29124
rect 17451 29121 17463 29155
rect 17405 29115 17463 29121
rect 17589 29155 17647 29161
rect 17589 29121 17601 29155
rect 17635 29121 17647 29155
rect 17589 29115 17647 29121
rect 18463 29155 18512 29161
rect 18463 29121 18475 29155
rect 18509 29121 18512 29155
rect 18463 29115 18512 29121
rect 18506 29112 18512 29115
rect 18564 29112 18570 29164
rect 19242 29112 19248 29164
rect 19300 29152 19306 29164
rect 19593 29155 19651 29161
rect 19593 29152 19605 29155
rect 19300 29124 19605 29152
rect 19300 29112 19306 29124
rect 19593 29121 19605 29124
rect 19639 29121 19651 29155
rect 19593 29115 19651 29121
rect 20806 29112 20812 29164
rect 20864 29152 20870 29164
rect 29362 29152 29368 29164
rect 20864 29124 29368 29152
rect 20864 29112 20870 29124
rect 29362 29112 29368 29124
rect 29420 29112 29426 29164
rect 29546 29112 29552 29164
rect 29604 29112 29610 29164
rect 29638 29112 29644 29164
rect 29696 29112 29702 29164
rect 30208 29161 30236 29192
rect 34146 29180 34152 29232
rect 34204 29220 34210 29232
rect 35912 29220 35940 29260
rect 36725 29257 36737 29260
rect 36771 29257 36783 29291
rect 36725 29251 36783 29257
rect 37274 29248 37280 29300
rect 37332 29288 37338 29300
rect 38102 29288 38108 29300
rect 37332 29260 37504 29288
rect 37332 29248 37338 29260
rect 36814 29220 36820 29232
rect 34204 29192 35940 29220
rect 36096 29192 36820 29220
rect 34204 29180 34210 29192
rect 30193 29155 30251 29161
rect 30193 29121 30205 29155
rect 30239 29121 30251 29155
rect 30193 29115 30251 29121
rect 32122 29112 32128 29164
rect 32180 29152 32186 29164
rect 33594 29152 33600 29164
rect 32180 29124 33600 29152
rect 32180 29112 32186 29124
rect 33594 29112 33600 29124
rect 33652 29112 33658 29164
rect 33870 29161 33876 29164
rect 33864 29115 33876 29161
rect 33870 29112 33876 29115
rect 33928 29112 33934 29164
rect 36096 29161 36124 29192
rect 36814 29180 36820 29192
rect 36872 29180 36878 29232
rect 36081 29155 36139 29161
rect 36081 29121 36093 29155
rect 36127 29121 36139 29155
rect 36081 29115 36139 29121
rect 36174 29155 36232 29161
rect 36174 29121 36186 29155
rect 36220 29121 36232 29155
rect 36174 29115 36232 29121
rect 13403 29056 13492 29084
rect 13541 29087 13599 29093
rect 13403 29053 13415 29056
rect 13357 29047 13415 29053
rect 13541 29053 13553 29087
rect 13587 29053 13599 29087
rect 13541 29047 13599 29053
rect 8496 28988 8616 29016
rect 9125 29019 9183 29025
rect 8496 28948 8524 28988
rect 9125 28985 9137 29019
rect 9171 29016 9183 29019
rect 9858 29016 9864 29028
rect 9171 28988 9864 29016
rect 9171 28985 9183 28988
rect 9125 28979 9183 28985
rect 9858 28976 9864 28988
rect 9916 28976 9922 29028
rect 13170 29016 13176 29028
rect 11256 28988 11468 29016
rect 7576 28920 8524 28948
rect 8941 28951 8999 28957
rect 8941 28917 8953 28951
rect 8987 28948 8999 28951
rect 9306 28948 9312 28960
rect 8987 28920 9312 28948
rect 8987 28917 8999 28920
rect 8941 28911 8999 28917
rect 9306 28908 9312 28920
rect 9364 28908 9370 28960
rect 9398 28908 9404 28960
rect 9456 28948 9462 28960
rect 11256 28948 11284 28988
rect 9456 28920 11284 28948
rect 9456 28908 9462 28920
rect 11330 28908 11336 28960
rect 11388 28908 11394 28960
rect 11440 28948 11468 28988
rect 12636 28988 13176 29016
rect 12636 28948 12664 28988
rect 13170 28976 13176 28988
rect 13228 28976 13234 29028
rect 11440 28920 12664 28948
rect 12710 28908 12716 28960
rect 12768 28908 12774 28960
rect 13556 28948 13584 29047
rect 15102 29044 15108 29096
rect 15160 29044 15166 29096
rect 17310 29044 17316 29096
rect 17368 29084 17374 29096
rect 17368 29056 17908 29084
rect 17368 29044 17374 29056
rect 15120 29016 15148 29044
rect 14476 28988 15148 29016
rect 14476 28948 14504 28988
rect 16758 28976 16764 29028
rect 16816 29016 16822 29028
rect 17678 29016 17684 29028
rect 16816 28988 17684 29016
rect 16816 28976 16822 28988
rect 17678 28976 17684 28988
rect 17736 28976 17742 29028
rect 17880 29016 17908 29056
rect 17954 29044 17960 29096
rect 18012 29084 18018 29096
rect 18325 29087 18383 29093
rect 18325 29084 18337 29087
rect 18012 29056 18337 29084
rect 18012 29044 18018 29056
rect 18325 29053 18337 29056
rect 18371 29053 18383 29087
rect 18325 29047 18383 29053
rect 18598 29044 18604 29096
rect 18656 29044 18662 29096
rect 18782 29044 18788 29096
rect 18840 29084 18846 29096
rect 19337 29087 19395 29093
rect 19337 29084 19349 29087
rect 18840 29056 19349 29084
rect 18840 29044 18846 29056
rect 19337 29053 19349 29056
rect 19383 29053 19395 29087
rect 19337 29047 19395 29053
rect 29454 29044 29460 29096
rect 29512 29084 29518 29096
rect 29733 29087 29791 29093
rect 29733 29084 29745 29087
rect 29512 29056 29745 29084
rect 29512 29044 29518 29056
rect 29733 29053 29745 29056
rect 29779 29053 29791 29087
rect 32858 29084 32864 29096
rect 29733 29047 29791 29053
rect 29932 29056 32864 29084
rect 18049 29019 18107 29025
rect 18049 29016 18061 29019
rect 17880 28988 18061 29016
rect 18049 28985 18061 28988
rect 18095 29016 18107 29019
rect 18138 29016 18144 29028
rect 18095 28988 18144 29016
rect 18095 28985 18107 28988
rect 18049 28979 18107 28985
rect 18138 28976 18144 28988
rect 18196 28976 18202 29028
rect 21450 28976 21456 29028
rect 21508 29016 21514 29028
rect 29932 29016 29960 29056
rect 32858 29044 32864 29056
rect 32916 29084 32922 29096
rect 33226 29084 33232 29096
rect 32916 29056 33232 29084
rect 32916 29044 32922 29056
rect 33226 29044 33232 29056
rect 33284 29044 33290 29096
rect 34606 29044 34612 29096
rect 34664 29084 34670 29096
rect 34664 29056 35112 29084
rect 34664 29044 34670 29056
rect 21508 28988 29960 29016
rect 21508 28976 21514 28988
rect 30006 28976 30012 29028
rect 30064 28976 30070 29028
rect 34977 29019 35035 29025
rect 34977 29016 34989 29019
rect 34532 28988 34989 29016
rect 13556 28920 14504 28948
rect 14921 28951 14979 28957
rect 14921 28917 14933 28951
rect 14967 28948 14979 28951
rect 15102 28948 15108 28960
rect 14967 28920 15108 28948
rect 14967 28917 14979 28920
rect 14921 28911 14979 28917
rect 15102 28908 15108 28920
rect 15160 28908 15166 28960
rect 18690 28908 18696 28960
rect 18748 28948 18754 28960
rect 32674 28948 32680 28960
rect 18748 28920 32680 28948
rect 18748 28908 18754 28920
rect 32674 28908 32680 28920
rect 32732 28908 32738 28960
rect 33410 28908 33416 28960
rect 33468 28948 33474 28960
rect 34532 28948 34560 28988
rect 34977 28985 34989 28988
rect 35023 28985 35035 29019
rect 35084 29016 35112 29056
rect 35986 29044 35992 29096
rect 36044 29084 36050 29096
rect 36188 29084 36216 29115
rect 36354 29112 36360 29164
rect 36412 29112 36418 29164
rect 36449 29155 36507 29161
rect 36449 29121 36461 29155
rect 36495 29121 36507 29155
rect 36449 29115 36507 29121
rect 36587 29155 36645 29161
rect 36587 29121 36599 29155
rect 36633 29152 36645 29155
rect 36722 29152 36728 29164
rect 36633 29124 36728 29152
rect 36633 29121 36645 29124
rect 36587 29115 36645 29121
rect 36044 29056 36216 29084
rect 36044 29044 36050 29056
rect 36464 29016 36492 29115
rect 36722 29112 36728 29124
rect 36780 29112 36786 29164
rect 37274 29112 37280 29164
rect 37332 29112 37338 29164
rect 37476 29161 37504 29260
rect 37568 29260 38108 29288
rect 37568 29229 37596 29260
rect 38102 29248 38108 29260
rect 38160 29248 38166 29300
rect 38286 29248 38292 29300
rect 38344 29288 38350 29300
rect 38473 29291 38531 29297
rect 38473 29288 38485 29291
rect 38344 29260 38485 29288
rect 38344 29248 38350 29260
rect 38473 29257 38485 29260
rect 38519 29257 38531 29291
rect 38473 29251 38531 29257
rect 38838 29248 38844 29300
rect 38896 29248 38902 29300
rect 39482 29248 39488 29300
rect 39540 29288 39546 29300
rect 40957 29291 41015 29297
rect 40957 29288 40969 29291
rect 39540 29260 40969 29288
rect 39540 29248 39546 29260
rect 40957 29257 40969 29260
rect 41003 29257 41015 29291
rect 40957 29251 41015 29257
rect 41322 29248 41328 29300
rect 41380 29288 41386 29300
rect 41380 29260 41644 29288
rect 41380 29248 41386 29260
rect 37553 29223 37611 29229
rect 37553 29189 37565 29223
rect 37599 29189 37611 29223
rect 38856 29220 38884 29248
rect 39298 29220 39304 29232
rect 37553 29183 37611 29189
rect 38672 29192 38884 29220
rect 38948 29192 39304 29220
rect 37461 29155 37519 29161
rect 37461 29121 37473 29155
rect 37507 29121 37519 29155
rect 37645 29155 37703 29161
rect 37645 29152 37657 29155
rect 37461 29115 37519 29121
rect 37568 29124 37657 29152
rect 35084 28988 36492 29016
rect 36740 29016 36768 29112
rect 37568 29016 37596 29124
rect 37645 29121 37657 29124
rect 37691 29121 37703 29155
rect 37645 29115 37703 29121
rect 38102 29112 38108 29164
rect 38160 29112 38166 29164
rect 38672 29161 38700 29192
rect 38657 29155 38715 29161
rect 38657 29121 38669 29155
rect 38703 29121 38715 29155
rect 38657 29115 38715 29121
rect 38749 29155 38807 29161
rect 38749 29121 38761 29155
rect 38795 29152 38807 29155
rect 38838 29152 38844 29164
rect 38795 29124 38844 29152
rect 38795 29121 38807 29124
rect 38749 29115 38807 29121
rect 38672 29084 38700 29115
rect 38838 29112 38844 29124
rect 38896 29112 38902 29164
rect 38948 29161 38976 29192
rect 39298 29180 39304 29192
rect 39356 29180 39362 29232
rect 40126 29180 40132 29232
rect 40184 29220 40190 29232
rect 41230 29220 41236 29232
rect 40184 29192 41236 29220
rect 40184 29180 40190 29192
rect 41230 29180 41236 29192
rect 41288 29180 41294 29232
rect 38933 29155 38991 29161
rect 38933 29121 38945 29155
rect 38979 29121 38991 29155
rect 38933 29115 38991 29121
rect 39114 29112 39120 29164
rect 39172 29112 39178 29164
rect 40865 29155 40923 29161
rect 40865 29121 40877 29155
rect 40911 29152 40923 29155
rect 40954 29152 40960 29164
rect 40911 29124 40960 29152
rect 40911 29121 40923 29124
rect 40865 29115 40923 29121
rect 40954 29112 40960 29124
rect 41012 29112 41018 29164
rect 41049 29155 41107 29161
rect 41049 29121 41061 29155
rect 41095 29152 41107 29155
rect 41138 29152 41144 29164
rect 41095 29124 41144 29152
rect 41095 29121 41107 29124
rect 41049 29115 41107 29121
rect 41138 29112 41144 29124
rect 41196 29112 41202 29164
rect 41506 29112 41512 29164
rect 41564 29112 41570 29164
rect 41616 29158 41644 29260
rect 41966 29248 41972 29300
rect 42024 29288 42030 29300
rect 42024 29260 46520 29288
rect 42024 29248 42030 29260
rect 43070 29220 43076 29232
rect 41800 29192 42104 29220
rect 41705 29158 41763 29161
rect 41616 29155 41763 29158
rect 41616 29130 41717 29155
rect 41705 29121 41717 29130
rect 41751 29121 41763 29155
rect 41705 29115 41763 29121
rect 38672 29056 39988 29084
rect 37734 29016 37740 29028
rect 36740 28988 37740 29016
rect 34977 28979 35035 28985
rect 37734 28976 37740 28988
rect 37792 28976 37798 29028
rect 38841 29019 38899 29025
rect 38841 28985 38853 29019
rect 38887 29016 38899 29019
rect 39022 29016 39028 29028
rect 38887 28988 39028 29016
rect 38887 28985 38899 28988
rect 38841 28979 38899 28985
rect 39022 28976 39028 28988
rect 39080 28976 39086 29028
rect 39960 29016 39988 29056
rect 40034 29044 40040 29096
rect 40092 29084 40098 29096
rect 41322 29084 41328 29096
rect 40092 29056 41328 29084
rect 40092 29044 40098 29056
rect 41322 29044 41328 29056
rect 41380 29044 41386 29096
rect 41601 29087 41659 29093
rect 41601 29053 41613 29087
rect 41647 29084 41659 29087
rect 41800 29084 41828 29192
rect 42076 29164 42104 29192
rect 42812 29192 43076 29220
rect 41874 29112 41880 29164
rect 41932 29112 41938 29164
rect 42058 29112 42064 29164
rect 42116 29112 42122 29164
rect 42150 29112 42156 29164
rect 42208 29152 42214 29164
rect 42610 29152 42616 29164
rect 42208 29124 42616 29152
rect 42208 29112 42214 29124
rect 42610 29112 42616 29124
rect 42668 29112 42674 29164
rect 42812 29161 42840 29192
rect 43070 29180 43076 29192
rect 43128 29180 43134 29232
rect 42797 29155 42855 29161
rect 42797 29121 42809 29155
rect 42843 29121 42855 29155
rect 42797 29115 42855 29121
rect 42889 29155 42947 29161
rect 42889 29121 42901 29155
rect 42935 29152 42947 29155
rect 43162 29152 43168 29164
rect 42935 29124 43168 29152
rect 42935 29121 42947 29124
rect 42889 29115 42947 29121
rect 43162 29112 43168 29124
rect 43220 29112 43226 29164
rect 46492 29161 46520 29260
rect 46658 29248 46664 29300
rect 46716 29248 46722 29300
rect 46477 29155 46535 29161
rect 46477 29121 46489 29155
rect 46523 29121 46535 29155
rect 46477 29115 46535 29121
rect 43714 29084 43720 29096
rect 41647 29056 41828 29084
rect 41984 29056 43720 29084
rect 41647 29053 41659 29056
rect 41601 29047 41659 29053
rect 41984 29016 42012 29056
rect 43714 29044 43720 29056
rect 43772 29084 43778 29096
rect 44726 29084 44732 29096
rect 43772 29056 44732 29084
rect 43772 29044 43778 29056
rect 44726 29044 44732 29056
rect 44784 29084 44790 29096
rect 45002 29084 45008 29096
rect 44784 29056 45008 29084
rect 44784 29044 44790 29056
rect 45002 29044 45008 29056
rect 45060 29044 45066 29096
rect 39960 28988 42012 29016
rect 42061 29019 42119 29025
rect 42061 28985 42073 29019
rect 42107 29016 42119 29019
rect 42150 29016 42156 29028
rect 42107 28988 42156 29016
rect 42107 28985 42119 28988
rect 42061 28979 42119 28985
rect 42150 28976 42156 28988
rect 42208 28976 42214 29028
rect 33468 28920 34560 28948
rect 33468 28908 33474 28920
rect 37826 28908 37832 28960
rect 37884 28908 37890 28960
rect 41414 28908 41420 28960
rect 41472 28948 41478 28960
rect 41598 28948 41604 28960
rect 41472 28920 41604 28948
rect 41472 28908 41478 28920
rect 41598 28908 41604 28920
rect 41656 28908 41662 28960
rect 41966 28908 41972 28960
rect 42024 28948 42030 28960
rect 42429 28951 42487 28957
rect 42429 28948 42441 28951
rect 42024 28920 42441 28948
rect 42024 28908 42030 28920
rect 42429 28917 42441 28920
rect 42475 28917 42487 28951
rect 42429 28911 42487 28917
rect 1104 28858 47104 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 47104 28858
rect 1104 28784 47104 28806
rect 7834 28704 7840 28756
rect 7892 28744 7898 28756
rect 8021 28747 8079 28753
rect 8021 28744 8033 28747
rect 7892 28716 8033 28744
rect 7892 28704 7898 28716
rect 8021 28713 8033 28716
rect 8067 28713 8079 28747
rect 8021 28707 8079 28713
rect 9769 28747 9827 28753
rect 9769 28713 9781 28747
rect 9815 28744 9827 28747
rect 11054 28744 11060 28756
rect 9815 28716 11060 28744
rect 9815 28713 9827 28716
rect 9769 28707 9827 28713
rect 11054 28704 11060 28716
rect 11112 28704 11118 28756
rect 14090 28704 14096 28756
rect 14148 28704 14154 28756
rect 15197 28747 15255 28753
rect 15197 28713 15209 28747
rect 15243 28713 15255 28747
rect 15197 28707 15255 28713
rect 18233 28747 18291 28753
rect 18233 28713 18245 28747
rect 18279 28744 18291 28747
rect 19242 28744 19248 28756
rect 18279 28716 19248 28744
rect 18279 28713 18291 28716
rect 18233 28707 18291 28713
rect 5902 28636 5908 28688
rect 5960 28676 5966 28688
rect 6730 28676 6736 28688
rect 5960 28648 6736 28676
rect 5960 28636 5966 28648
rect 6730 28636 6736 28648
rect 6788 28636 6794 28688
rect 10962 28636 10968 28688
rect 11020 28636 11026 28688
rect 13998 28636 14004 28688
rect 14056 28676 14062 28688
rect 15212 28676 15240 28707
rect 19242 28704 19248 28716
rect 19300 28704 19306 28756
rect 19705 28747 19763 28753
rect 19705 28713 19717 28747
rect 19751 28744 19763 28747
rect 20254 28744 20260 28756
rect 19751 28716 20260 28744
rect 19751 28713 19763 28716
rect 19705 28707 19763 28713
rect 20254 28704 20260 28716
rect 20312 28744 20318 28756
rect 20806 28744 20812 28756
rect 20312 28716 20812 28744
rect 20312 28704 20318 28716
rect 20806 28704 20812 28716
rect 20864 28704 20870 28756
rect 29273 28747 29331 28753
rect 22066 28716 27200 28744
rect 14056 28648 15240 28676
rect 14056 28636 14062 28648
rect 19794 28636 19800 28688
rect 19852 28676 19858 28688
rect 22066 28676 22094 28716
rect 19852 28648 22094 28676
rect 19852 28636 19858 28648
rect 22186 28636 22192 28688
rect 22244 28676 22250 28688
rect 24394 28676 24400 28688
rect 22244 28648 24400 28676
rect 22244 28636 22250 28648
rect 24394 28636 24400 28648
rect 24452 28676 24458 28688
rect 24670 28676 24676 28688
rect 24452 28648 24676 28676
rect 24452 28636 24458 28648
rect 24670 28636 24676 28648
rect 24728 28636 24734 28688
rect 3234 28568 3240 28620
rect 3292 28608 3298 28620
rect 7098 28608 7104 28620
rect 3292 28580 4660 28608
rect 3292 28568 3298 28580
rect 4430 28500 4436 28552
rect 4488 28500 4494 28552
rect 4522 28500 4528 28552
rect 4580 28500 4586 28552
rect 4632 28540 4660 28580
rect 6472 28580 7104 28608
rect 6472 28552 6500 28580
rect 7098 28568 7104 28580
rect 7156 28568 7162 28620
rect 7282 28568 7288 28620
rect 7340 28568 7346 28620
rect 7466 28568 7472 28620
rect 7524 28568 7530 28620
rect 7576 28580 9076 28608
rect 6454 28540 6460 28552
rect 4632 28512 6460 28540
rect 6454 28500 6460 28512
rect 6512 28500 6518 28552
rect 6730 28500 6736 28552
rect 6788 28540 6794 28552
rect 7193 28543 7251 28549
rect 7193 28540 7205 28543
rect 6788 28512 7205 28540
rect 6788 28500 6794 28512
rect 7193 28509 7205 28512
rect 7239 28540 7251 28543
rect 7576 28540 7604 28580
rect 7239 28512 7604 28540
rect 8205 28543 8263 28549
rect 7239 28509 7251 28512
rect 7193 28503 7251 28509
rect 8205 28509 8217 28543
rect 8251 28540 8263 28543
rect 9048 28540 9076 28580
rect 9398 28568 9404 28620
rect 9456 28608 9462 28620
rect 9493 28611 9551 28617
rect 9493 28608 9505 28611
rect 9456 28580 9505 28608
rect 9456 28568 9462 28580
rect 9493 28577 9505 28580
rect 9539 28577 9551 28611
rect 9493 28571 9551 28577
rect 9858 28568 9864 28620
rect 9916 28608 9922 28620
rect 10229 28611 10287 28617
rect 10229 28608 10241 28611
rect 9916 28580 10241 28608
rect 9916 28568 9922 28580
rect 10229 28577 10241 28580
rect 10275 28577 10287 28611
rect 10229 28571 10287 28577
rect 10413 28611 10471 28617
rect 10413 28577 10425 28611
rect 10459 28608 10471 28611
rect 10870 28608 10876 28620
rect 10459 28580 10876 28608
rect 10459 28577 10471 28580
rect 10413 28571 10471 28577
rect 10870 28568 10876 28580
rect 10928 28568 10934 28620
rect 10980 28608 11008 28636
rect 11149 28611 11207 28617
rect 11149 28608 11161 28611
rect 10980 28580 11161 28608
rect 11149 28577 11161 28580
rect 11195 28577 11207 28611
rect 11149 28571 11207 28577
rect 11330 28568 11336 28620
rect 11388 28608 11394 28620
rect 11701 28611 11759 28617
rect 11701 28608 11713 28611
rect 11388 28580 11713 28608
rect 11388 28568 11394 28580
rect 11701 28577 11713 28580
rect 11747 28577 11759 28611
rect 11701 28571 11759 28577
rect 12618 28568 12624 28620
rect 12676 28568 12682 28620
rect 19334 28608 19340 28620
rect 14568 28580 19340 28608
rect 10965 28543 11023 28549
rect 10965 28540 10977 28543
rect 8251 28512 8984 28540
rect 9048 28512 10977 28540
rect 8251 28509 8263 28512
rect 8205 28503 8263 28509
rect 4770 28475 4828 28481
rect 4770 28472 4782 28475
rect 4264 28444 4782 28472
rect 2314 28364 2320 28416
rect 2372 28404 2378 28416
rect 2593 28407 2651 28413
rect 2593 28404 2605 28407
rect 2372 28376 2605 28404
rect 2372 28364 2378 28376
rect 2593 28373 2605 28376
rect 2639 28373 2651 28407
rect 2593 28367 2651 28373
rect 2958 28364 2964 28416
rect 3016 28364 3022 28416
rect 3053 28407 3111 28413
rect 3053 28373 3065 28407
rect 3099 28404 3111 28407
rect 4062 28404 4068 28416
rect 3099 28376 4068 28404
rect 3099 28373 3111 28376
rect 3053 28367 3111 28373
rect 4062 28364 4068 28376
rect 4120 28364 4126 28416
rect 4264 28413 4292 28444
rect 4770 28441 4782 28444
rect 4816 28441 4828 28475
rect 4770 28435 4828 28441
rect 4249 28407 4307 28413
rect 4249 28373 4261 28407
rect 4295 28373 4307 28407
rect 4249 28367 4307 28373
rect 6822 28364 6828 28416
rect 6880 28364 6886 28416
rect 8956 28413 8984 28512
rect 10965 28509 10977 28512
rect 11011 28509 11023 28543
rect 10965 28503 11023 28509
rect 11977 28543 12035 28549
rect 11977 28509 11989 28543
rect 12023 28509 12035 28543
rect 11977 28503 12035 28509
rect 9398 28432 9404 28484
rect 9456 28432 9462 28484
rect 10137 28475 10195 28481
rect 10137 28441 10149 28475
rect 10183 28472 10195 28475
rect 11992 28472 12020 28503
rect 12894 28500 12900 28552
rect 12952 28540 12958 28552
rect 13630 28540 13636 28552
rect 12952 28512 13636 28540
rect 12952 28500 12958 28512
rect 13630 28500 13636 28512
rect 13688 28540 13694 28552
rect 13688 28512 13860 28540
rect 13688 28500 13694 28512
rect 13832 28484 13860 28512
rect 14274 28500 14280 28552
rect 14332 28500 14338 28552
rect 14568 28549 14596 28580
rect 19334 28568 19340 28580
rect 19392 28568 19398 28620
rect 19426 28568 19432 28620
rect 19484 28608 19490 28620
rect 22370 28608 22376 28620
rect 19484 28580 22376 28608
rect 19484 28568 19490 28580
rect 22370 28568 22376 28580
rect 22428 28568 22434 28620
rect 25958 28608 25964 28620
rect 22480 28580 25964 28608
rect 14553 28543 14611 28549
rect 14553 28509 14565 28543
rect 14599 28509 14611 28543
rect 14553 28503 14611 28509
rect 18414 28500 18420 28552
rect 18472 28500 18478 28552
rect 19521 28543 19579 28549
rect 19521 28509 19533 28543
rect 19567 28509 19579 28543
rect 19521 28503 19579 28509
rect 10183 28444 10824 28472
rect 10183 28441 10195 28444
rect 10137 28435 10195 28441
rect 8941 28407 8999 28413
rect 8941 28373 8953 28407
rect 8987 28373 8999 28407
rect 8941 28367 8999 28373
rect 9306 28364 9312 28416
rect 9364 28364 9370 28416
rect 10594 28364 10600 28416
rect 10652 28364 10658 28416
rect 10796 28404 10824 28444
rect 10960 28444 12020 28472
rect 10960 28404 10988 28444
rect 10796 28376 10988 28404
rect 11054 28364 11060 28416
rect 11112 28364 11118 28416
rect 11992 28404 12020 28444
rect 13814 28432 13820 28484
rect 13872 28472 13878 28484
rect 15013 28475 15071 28481
rect 15013 28472 15025 28475
rect 13872 28444 15025 28472
rect 13872 28432 13878 28444
rect 15013 28441 15025 28444
rect 15059 28441 15071 28475
rect 15013 28435 15071 28441
rect 15102 28432 15108 28484
rect 15160 28472 15166 28484
rect 15213 28475 15271 28481
rect 15213 28472 15225 28475
rect 15160 28444 15225 28472
rect 15160 28432 15166 28444
rect 15213 28441 15225 28444
rect 15259 28441 15271 28475
rect 19536 28472 19564 28503
rect 21266 28500 21272 28552
rect 21324 28500 21330 28552
rect 21729 28543 21787 28549
rect 21729 28509 21741 28543
rect 21775 28540 21787 28543
rect 21818 28540 21824 28552
rect 21775 28512 21824 28540
rect 21775 28509 21787 28512
rect 21729 28503 21787 28509
rect 21818 28500 21824 28512
rect 21876 28500 21882 28552
rect 20162 28472 20168 28484
rect 19536 28444 20168 28472
rect 15213 28435 15271 28441
rect 20162 28432 20168 28444
rect 20220 28432 20226 28484
rect 20533 28475 20591 28481
rect 20533 28441 20545 28475
rect 20579 28472 20591 28475
rect 20714 28472 20720 28484
rect 20579 28444 20720 28472
rect 20579 28441 20591 28444
rect 20533 28435 20591 28441
rect 20714 28432 20720 28444
rect 20772 28472 20778 28484
rect 22480 28472 22508 28580
rect 25958 28568 25964 28580
rect 26016 28568 26022 28620
rect 27172 28608 27200 28716
rect 29273 28713 29285 28747
rect 29319 28744 29331 28747
rect 29454 28744 29460 28756
rect 29319 28716 29460 28744
rect 29319 28713 29331 28716
rect 29273 28707 29331 28713
rect 29454 28704 29460 28716
rect 29512 28744 29518 28756
rect 30190 28744 30196 28756
rect 29512 28716 30196 28744
rect 29512 28704 29518 28716
rect 30190 28704 30196 28716
rect 30248 28704 30254 28756
rect 30558 28704 30564 28756
rect 30616 28744 30622 28756
rect 32490 28744 32496 28756
rect 30616 28716 32496 28744
rect 30616 28704 30622 28716
rect 32490 28704 32496 28716
rect 32548 28704 32554 28756
rect 32674 28704 32680 28756
rect 32732 28744 32738 28756
rect 32732 28716 33640 28744
rect 32732 28704 32738 28716
rect 27246 28636 27252 28688
rect 27304 28676 27310 28688
rect 27304 28648 28304 28676
rect 27304 28636 27310 28648
rect 27522 28608 27528 28620
rect 27172 28580 27528 28608
rect 27522 28568 27528 28580
rect 27580 28608 27586 28620
rect 28169 28611 28227 28617
rect 28169 28608 28181 28611
rect 27580 28580 28181 28608
rect 27580 28568 27586 28580
rect 28169 28577 28181 28580
rect 28215 28577 28227 28611
rect 28276 28608 28304 28648
rect 28534 28636 28540 28688
rect 28592 28676 28598 28688
rect 28592 28648 29592 28676
rect 28592 28636 28598 28648
rect 29564 28617 29592 28648
rect 32508 28648 33548 28676
rect 29549 28611 29607 28617
rect 28276 28580 29500 28608
rect 28169 28571 28227 28577
rect 22554 28500 22560 28552
rect 22612 28540 22618 28552
rect 23290 28540 23296 28552
rect 22612 28512 23296 28540
rect 22612 28500 22618 28512
rect 23290 28500 23296 28512
rect 23348 28500 23354 28552
rect 24854 28500 24860 28552
rect 24912 28540 24918 28552
rect 26142 28540 26148 28552
rect 24912 28512 26148 28540
rect 24912 28500 24918 28512
rect 26142 28500 26148 28512
rect 26200 28500 26206 28552
rect 27985 28543 28043 28549
rect 27985 28540 27997 28543
rect 26252 28512 27997 28540
rect 20772 28444 22508 28472
rect 20772 28432 20778 28444
rect 22922 28432 22928 28484
rect 22980 28472 22986 28484
rect 26252 28472 26280 28512
rect 22980 28444 26280 28472
rect 26412 28475 26470 28481
rect 22980 28432 22986 28444
rect 26412 28441 26424 28475
rect 26458 28472 26470 28475
rect 26602 28472 26608 28484
rect 26458 28444 26608 28472
rect 26458 28441 26470 28444
rect 26412 28435 26470 28441
rect 26602 28432 26608 28444
rect 26660 28432 26666 28484
rect 13446 28404 13452 28416
rect 11992 28376 13452 28404
rect 13446 28364 13452 28376
rect 13504 28404 13510 28416
rect 13998 28404 14004 28416
rect 13504 28376 14004 28404
rect 13504 28364 13510 28376
rect 13998 28364 14004 28376
rect 14056 28364 14062 28416
rect 14458 28364 14464 28416
rect 14516 28364 14522 28416
rect 15378 28364 15384 28416
rect 15436 28364 15442 28416
rect 20346 28364 20352 28416
rect 20404 28404 20410 28416
rect 21085 28407 21143 28413
rect 21085 28404 21097 28407
rect 20404 28376 21097 28404
rect 20404 28364 20410 28376
rect 21085 28373 21097 28376
rect 21131 28373 21143 28407
rect 21085 28367 21143 28373
rect 21542 28364 21548 28416
rect 21600 28364 21606 28416
rect 21726 28364 21732 28416
rect 21784 28404 21790 28416
rect 27246 28404 27252 28416
rect 21784 28376 27252 28404
rect 21784 28364 21790 28376
rect 27246 28364 27252 28376
rect 27304 28364 27310 28416
rect 27540 28413 27568 28512
rect 27985 28509 27997 28512
rect 28031 28509 28043 28543
rect 27985 28503 28043 28509
rect 28721 28543 28779 28549
rect 28721 28509 28733 28543
rect 28767 28540 28779 28543
rect 29086 28540 29092 28552
rect 28767 28512 29092 28540
rect 28767 28509 28779 28512
rect 28721 28503 28779 28509
rect 29086 28500 29092 28512
rect 29144 28500 29150 28552
rect 29472 28540 29500 28580
rect 29549 28577 29561 28611
rect 29595 28577 29607 28611
rect 29549 28571 29607 28577
rect 31570 28568 31576 28620
rect 31628 28608 31634 28620
rect 32508 28617 32536 28648
rect 33520 28620 33548 28648
rect 32493 28611 32551 28617
rect 32493 28608 32505 28611
rect 31628 28580 32505 28608
rect 31628 28568 31634 28580
rect 32493 28577 32505 28580
rect 32539 28577 32551 28611
rect 32493 28571 32551 28577
rect 32582 28568 32588 28620
rect 32640 28568 32646 28620
rect 33318 28608 33324 28620
rect 33152 28580 33324 28608
rect 33152 28540 33180 28580
rect 33318 28568 33324 28580
rect 33376 28568 33382 28620
rect 33502 28568 33508 28620
rect 33560 28568 33566 28620
rect 33612 28617 33640 28716
rect 33870 28704 33876 28756
rect 33928 28704 33934 28756
rect 35802 28704 35808 28756
rect 35860 28744 35866 28756
rect 37001 28747 37059 28753
rect 37001 28744 37013 28747
rect 35860 28716 37013 28744
rect 35860 28704 35866 28716
rect 37001 28713 37013 28716
rect 37047 28713 37059 28747
rect 37001 28707 37059 28713
rect 37642 28704 37648 28756
rect 37700 28744 37706 28756
rect 38654 28744 38660 28756
rect 37700 28716 38660 28744
rect 37700 28704 37706 28716
rect 38654 28704 38660 28716
rect 38712 28744 38718 28756
rect 38749 28747 38807 28753
rect 38749 28744 38761 28747
rect 38712 28716 38761 28744
rect 38712 28704 38718 28716
rect 38749 28713 38761 28716
rect 38795 28713 38807 28747
rect 38749 28707 38807 28713
rect 40770 28704 40776 28756
rect 40828 28744 40834 28756
rect 44542 28744 44548 28756
rect 40828 28716 44548 28744
rect 40828 28704 40834 28716
rect 44542 28704 44548 28716
rect 44600 28704 44606 28756
rect 44177 28679 44235 28685
rect 44177 28676 44189 28679
rect 41386 28648 44189 28676
rect 33597 28611 33655 28617
rect 33597 28577 33609 28611
rect 33643 28577 33655 28611
rect 33597 28571 33655 28577
rect 29472 28512 33180 28540
rect 33336 28540 33364 28568
rect 33870 28540 33876 28552
rect 33336 28512 33876 28540
rect 33870 28500 33876 28512
rect 33928 28500 33934 28552
rect 34057 28543 34115 28549
rect 34057 28509 34069 28543
rect 34103 28509 34115 28543
rect 34057 28503 34115 28509
rect 37185 28543 37243 28549
rect 37185 28509 37197 28543
rect 37231 28540 37243 28543
rect 37826 28540 37832 28552
rect 37231 28512 37832 28540
rect 37231 28509 37243 28512
rect 37185 28503 37243 28509
rect 28994 28432 29000 28484
rect 29052 28432 29058 28484
rect 29178 28432 29184 28484
rect 29236 28472 29242 28484
rect 29794 28475 29852 28481
rect 29794 28472 29806 28475
rect 29236 28444 29806 28472
rect 29236 28432 29242 28444
rect 29794 28441 29806 28444
rect 29840 28441 29852 28475
rect 29794 28435 29852 28441
rect 32674 28432 32680 28484
rect 32732 28472 32738 28484
rect 33410 28472 33416 28484
rect 32732 28444 33416 28472
rect 32732 28432 32738 28444
rect 33410 28432 33416 28444
rect 33468 28432 33474 28484
rect 27525 28407 27583 28413
rect 27525 28373 27537 28407
rect 27571 28373 27583 28407
rect 27525 28367 27583 28373
rect 27614 28364 27620 28416
rect 27672 28364 27678 28416
rect 28077 28407 28135 28413
rect 28077 28373 28089 28407
rect 28123 28404 28135 28407
rect 29638 28404 29644 28416
rect 28123 28376 29644 28404
rect 28123 28373 28135 28376
rect 28077 28367 28135 28373
rect 29638 28364 29644 28376
rect 29696 28364 29702 28416
rect 29914 28364 29920 28416
rect 29972 28404 29978 28416
rect 30929 28407 30987 28413
rect 30929 28404 30941 28407
rect 29972 28376 30941 28404
rect 29972 28364 29978 28376
rect 30929 28373 30941 28376
rect 30975 28373 30987 28407
rect 30929 28367 30987 28373
rect 31938 28364 31944 28416
rect 31996 28404 32002 28416
rect 32033 28407 32091 28413
rect 32033 28404 32045 28407
rect 31996 28376 32045 28404
rect 31996 28364 32002 28376
rect 32033 28373 32045 28376
rect 32079 28373 32091 28407
rect 32033 28367 32091 28373
rect 32401 28407 32459 28413
rect 32401 28373 32413 28407
rect 32447 28404 32459 28407
rect 32858 28404 32864 28416
rect 32447 28376 32864 28404
rect 32447 28373 32459 28376
rect 32401 28367 32459 28373
rect 32858 28364 32864 28376
rect 32916 28364 32922 28416
rect 33045 28407 33103 28413
rect 33045 28373 33057 28407
rect 33091 28404 33103 28407
rect 34072 28404 34100 28503
rect 37826 28500 37832 28512
rect 37884 28500 37890 28552
rect 41386 28540 41414 28648
rect 44177 28645 44189 28648
rect 44223 28645 44235 28679
rect 44177 28639 44235 28645
rect 42058 28568 42064 28620
rect 42116 28568 42122 28620
rect 42426 28568 42432 28620
rect 42484 28608 42490 28620
rect 44453 28611 44511 28617
rect 44453 28608 44465 28611
rect 42484 28580 44465 28608
rect 42484 28568 42490 28580
rect 44453 28577 44465 28580
rect 44499 28577 44511 28611
rect 44453 28571 44511 28577
rect 44545 28611 44603 28617
rect 44545 28577 44557 28611
rect 44591 28608 44603 28611
rect 45462 28608 45468 28620
rect 44591 28580 45468 28608
rect 44591 28577 44603 28580
rect 44545 28571 44603 28577
rect 45462 28568 45468 28580
rect 45520 28568 45526 28620
rect 38580 28512 41414 28540
rect 36998 28432 37004 28484
rect 37056 28472 37062 28484
rect 37461 28475 37519 28481
rect 37461 28472 37473 28475
rect 37056 28444 37473 28472
rect 37056 28432 37062 28444
rect 37461 28441 37473 28444
rect 37507 28441 37519 28475
rect 37461 28435 37519 28441
rect 33091 28376 34100 28404
rect 37369 28407 37427 28413
rect 33091 28373 33103 28376
rect 33045 28367 33103 28373
rect 37369 28373 37381 28407
rect 37415 28404 37427 28407
rect 38580 28404 38608 28512
rect 41782 28500 41788 28552
rect 41840 28500 41846 28552
rect 41877 28543 41935 28549
rect 41877 28509 41889 28543
rect 41923 28540 41935 28543
rect 41966 28540 41972 28552
rect 41923 28512 41972 28540
rect 41923 28509 41935 28512
rect 41877 28503 41935 28509
rect 41966 28500 41972 28512
rect 42024 28500 42030 28552
rect 43714 28500 43720 28552
rect 43772 28500 43778 28552
rect 44174 28500 44180 28552
rect 44232 28540 44238 28552
rect 44361 28543 44419 28549
rect 44361 28540 44373 28543
rect 44232 28512 44373 28540
rect 44232 28500 44238 28512
rect 44361 28509 44373 28512
rect 44407 28509 44419 28543
rect 44361 28503 44419 28509
rect 44637 28543 44695 28549
rect 44637 28509 44649 28543
rect 44683 28540 44695 28543
rect 44910 28540 44916 28552
rect 44683 28512 44916 28540
rect 44683 28509 44695 28512
rect 44637 28503 44695 28509
rect 44910 28500 44916 28512
rect 44968 28500 44974 28552
rect 45002 28500 45008 28552
rect 45060 28500 45066 28552
rect 45094 28500 45100 28552
rect 45152 28540 45158 28552
rect 45189 28543 45247 28549
rect 45189 28540 45201 28543
rect 45152 28512 45201 28540
rect 45152 28500 45158 28512
rect 45189 28509 45201 28512
rect 45235 28509 45247 28543
rect 45189 28503 45247 28509
rect 38657 28475 38715 28481
rect 38657 28441 38669 28475
rect 38703 28472 38715 28475
rect 39022 28472 39028 28484
rect 38703 28444 39028 28472
rect 38703 28441 38715 28444
rect 38657 28435 38715 28441
rect 39022 28432 39028 28444
rect 39080 28432 39086 28484
rect 43901 28475 43959 28481
rect 43901 28441 43913 28475
rect 43947 28472 43959 28475
rect 45112 28472 45140 28500
rect 43947 28444 45140 28472
rect 43947 28441 43959 28444
rect 43901 28435 43959 28441
rect 37415 28376 38608 28404
rect 42061 28407 42119 28413
rect 37415 28373 37427 28376
rect 37369 28367 37427 28373
rect 42061 28373 42073 28407
rect 42107 28404 42119 28407
rect 42610 28404 42616 28416
rect 42107 28376 42616 28404
rect 42107 28373 42119 28376
rect 42061 28367 42119 28373
rect 42610 28364 42616 28376
rect 42668 28364 42674 28416
rect 43990 28364 43996 28416
rect 44048 28404 44054 28416
rect 44085 28407 44143 28413
rect 44085 28404 44097 28407
rect 44048 28376 44097 28404
rect 44048 28364 44054 28376
rect 44085 28373 44097 28376
rect 44131 28373 44143 28407
rect 44085 28367 44143 28373
rect 45186 28364 45192 28416
rect 45244 28364 45250 28416
rect 1104 28314 47104 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 47104 28314
rect 1104 28240 47104 28262
rect 11885 28203 11943 28209
rect 11885 28169 11897 28203
rect 11931 28200 11943 28203
rect 11974 28200 11980 28212
rect 11931 28172 11980 28200
rect 11931 28169 11943 28172
rect 11885 28163 11943 28169
rect 11974 28160 11980 28172
rect 12032 28160 12038 28212
rect 12345 28203 12403 28209
rect 12345 28169 12357 28203
rect 12391 28200 12403 28203
rect 12710 28200 12716 28212
rect 12391 28172 12716 28200
rect 12391 28169 12403 28172
rect 12345 28163 12403 28169
rect 12710 28160 12716 28172
rect 12768 28160 12774 28212
rect 14274 28200 14280 28212
rect 13740 28172 14280 28200
rect 1670 28092 1676 28144
rect 1728 28132 1734 28144
rect 4522 28132 4528 28144
rect 1728 28104 4528 28132
rect 1728 28092 1734 28104
rect 2314 28024 2320 28076
rect 2372 28024 2378 28076
rect 2608 28073 2636 28104
rect 4522 28092 4528 28104
rect 4580 28132 4586 28144
rect 4580 28104 4936 28132
rect 4580 28092 4586 28104
rect 2593 28067 2651 28073
rect 2593 28033 2605 28067
rect 2639 28033 2651 28067
rect 2593 28027 2651 28033
rect 2860 28067 2918 28073
rect 2860 28033 2872 28067
rect 2906 28064 2918 28067
rect 3142 28064 3148 28076
rect 2906 28036 3148 28064
rect 2906 28033 2918 28036
rect 2860 28027 2918 28033
rect 3142 28024 3148 28036
rect 3200 28024 3206 28076
rect 4614 28024 4620 28076
rect 4672 28024 4678 28076
rect 4908 28073 4936 28104
rect 6822 28092 6828 28144
rect 6880 28132 6886 28144
rect 12253 28135 12311 28141
rect 6880 28104 7696 28132
rect 6880 28092 6886 28104
rect 4893 28067 4951 28073
rect 4893 28033 4905 28067
rect 4939 28033 4951 28067
rect 4893 28027 4951 28033
rect 6914 28024 6920 28076
rect 6972 28064 6978 28076
rect 7668 28073 7696 28104
rect 12253 28101 12265 28135
rect 12299 28132 12311 28135
rect 12894 28132 12900 28144
rect 12299 28104 12900 28132
rect 12299 28101 12311 28104
rect 12253 28095 12311 28101
rect 12894 28092 12900 28104
rect 12952 28092 12958 28144
rect 7377 28067 7435 28073
rect 7377 28064 7389 28067
rect 6972 28036 7389 28064
rect 6972 28024 6978 28036
rect 7377 28033 7389 28036
rect 7423 28033 7435 28067
rect 7377 28027 7435 28033
rect 7653 28067 7711 28073
rect 7653 28033 7665 28067
rect 7699 28033 7711 28067
rect 7653 28027 7711 28033
rect 12618 28024 12624 28076
rect 12676 28064 12682 28076
rect 12713 28067 12771 28073
rect 12713 28064 12725 28067
rect 12676 28036 12725 28064
rect 12676 28024 12682 28036
rect 12713 28033 12725 28036
rect 12759 28033 12771 28067
rect 12713 28027 12771 28033
rect 10962 27956 10968 28008
rect 11020 27996 11026 28008
rect 12529 27999 12587 28005
rect 12529 27996 12541 27999
rect 11020 27968 12541 27996
rect 11020 27956 11026 27968
rect 12529 27965 12541 27968
rect 12575 27996 12587 27999
rect 13740 27996 13768 28172
rect 14274 28160 14280 28172
rect 14332 28160 14338 28212
rect 15010 28160 15016 28212
rect 15068 28200 15074 28212
rect 18233 28203 18291 28209
rect 18233 28200 18245 28203
rect 15068 28172 18245 28200
rect 15068 28160 15074 28172
rect 18233 28169 18245 28172
rect 18279 28169 18291 28203
rect 18233 28163 18291 28169
rect 21545 28203 21603 28209
rect 21545 28169 21557 28203
rect 21591 28200 21603 28203
rect 21726 28200 21732 28212
rect 21591 28172 21732 28200
rect 21591 28169 21603 28172
rect 21545 28163 21603 28169
rect 21726 28160 21732 28172
rect 21784 28160 21790 28212
rect 21818 28160 21824 28212
rect 21876 28160 21882 28212
rect 26602 28160 26608 28212
rect 26660 28160 26666 28212
rect 27801 28203 27859 28209
rect 27801 28169 27813 28203
rect 27847 28200 27859 28203
rect 27982 28200 27988 28212
rect 27847 28172 27988 28200
rect 27847 28169 27859 28172
rect 27801 28163 27859 28169
rect 27982 28160 27988 28172
rect 28040 28160 28046 28212
rect 28813 28203 28871 28209
rect 28813 28169 28825 28203
rect 28859 28200 28871 28203
rect 29178 28200 29184 28212
rect 28859 28172 29184 28200
rect 28859 28169 28871 28172
rect 28813 28163 28871 28169
rect 29178 28160 29184 28172
rect 29236 28160 29242 28212
rect 29365 28203 29423 28209
rect 29365 28169 29377 28203
rect 29411 28169 29423 28203
rect 29365 28163 29423 28169
rect 13814 28092 13820 28144
rect 13872 28092 13878 28144
rect 13906 28092 13912 28144
rect 13964 28132 13970 28144
rect 14093 28135 14151 28141
rect 14093 28132 14105 28135
rect 13964 28104 14105 28132
rect 13964 28092 13970 28104
rect 14093 28101 14105 28104
rect 14139 28101 14151 28135
rect 14093 28095 14151 28101
rect 14185 28135 14243 28141
rect 14185 28101 14197 28135
rect 14231 28132 14243 28135
rect 14366 28132 14372 28144
rect 14231 28104 14372 28132
rect 14231 28101 14243 28104
rect 14185 28095 14243 28101
rect 14366 28092 14372 28104
rect 14424 28132 14430 28144
rect 15933 28135 15991 28141
rect 14424 28104 14964 28132
rect 14424 28092 14430 28104
rect 13998 28024 14004 28076
rect 14056 28024 14062 28076
rect 14458 28024 14464 28076
rect 14516 28064 14522 28076
rect 14936 28073 14964 28104
rect 15933 28101 15945 28135
rect 15979 28132 15991 28135
rect 16298 28132 16304 28144
rect 15979 28104 16304 28132
rect 15979 28101 15991 28104
rect 15933 28095 15991 28101
rect 16298 28092 16304 28104
rect 16356 28092 16362 28144
rect 17129 28135 17187 28141
rect 17129 28101 17141 28135
rect 17175 28132 17187 28135
rect 19426 28132 19432 28144
rect 17175 28104 19432 28132
rect 17175 28101 17187 28104
rect 17129 28095 17187 28101
rect 14645 28067 14703 28073
rect 14645 28064 14657 28067
rect 14516 28036 14657 28064
rect 14516 28024 14522 28036
rect 14645 28033 14657 28036
rect 14691 28033 14703 28067
rect 14645 28027 14703 28033
rect 14829 28067 14887 28073
rect 14829 28033 14841 28067
rect 14875 28033 14887 28067
rect 14829 28027 14887 28033
rect 14921 28067 14979 28073
rect 14921 28033 14933 28067
rect 14967 28033 14979 28067
rect 14921 28027 14979 28033
rect 15565 28067 15623 28073
rect 15565 28033 15577 28067
rect 15611 28064 15623 28067
rect 16390 28064 16396 28076
rect 15611 28036 16396 28064
rect 15611 28033 15623 28036
rect 15565 28027 15623 28033
rect 12575 27968 13768 27996
rect 12575 27965 12587 27968
rect 12529 27959 12587 27965
rect 14550 27956 14556 28008
rect 14608 27956 14614 28008
rect 14844 27996 14872 28027
rect 16390 28024 16396 28036
rect 16448 28024 16454 28076
rect 16482 28024 16488 28076
rect 16540 28064 16546 28076
rect 16761 28067 16819 28073
rect 16761 28064 16773 28067
rect 16540 28036 16773 28064
rect 16540 28024 16546 28036
rect 16761 28033 16773 28036
rect 16807 28033 16819 28067
rect 16761 28027 16819 28033
rect 15194 27996 15200 28008
rect 14844 27968 15200 27996
rect 11330 27888 11336 27940
rect 11388 27928 11394 27940
rect 12989 27931 13047 27937
rect 12989 27928 13001 27931
rect 11388 27900 13001 27928
rect 11388 27888 11394 27900
rect 12989 27897 13001 27900
rect 13035 27897 13047 27931
rect 12989 27891 13047 27897
rect 13173 27931 13231 27937
rect 13173 27897 13185 27931
rect 13219 27928 13231 27931
rect 14844 27928 14872 27968
rect 15194 27956 15200 27968
rect 15252 27956 15258 28008
rect 15381 27999 15439 28005
rect 15381 27965 15393 27999
rect 15427 27996 15439 27999
rect 15470 27996 15476 28008
rect 15427 27968 15476 27996
rect 15427 27965 15439 27968
rect 15381 27959 15439 27965
rect 15470 27956 15476 27968
rect 15528 27956 15534 28008
rect 15838 27956 15844 28008
rect 15896 27956 15902 28008
rect 16022 27956 16028 28008
rect 16080 27956 16086 28008
rect 16206 27956 16212 28008
rect 16264 27996 16270 28008
rect 17144 27996 17172 28095
rect 19426 28092 19432 28104
rect 19484 28092 19490 28144
rect 20990 28092 20996 28144
rect 21048 28132 21054 28144
rect 21269 28135 21327 28141
rect 21269 28132 21281 28135
rect 21048 28104 21281 28132
rect 21048 28092 21054 28104
rect 21269 28101 21281 28104
rect 21315 28101 21327 28135
rect 21269 28095 21327 28101
rect 22186 28092 22192 28144
rect 22244 28092 22250 28144
rect 18141 28067 18199 28073
rect 18141 28033 18153 28067
rect 18187 28064 18199 28067
rect 18601 28067 18659 28073
rect 18601 28064 18613 28067
rect 18187 28036 18613 28064
rect 18187 28033 18199 28036
rect 18141 28027 18199 28033
rect 18601 28033 18613 28036
rect 18647 28064 18659 28067
rect 19061 28067 19119 28073
rect 19061 28064 19073 28067
rect 18647 28036 19073 28064
rect 18647 28033 18659 28036
rect 18601 28027 18659 28033
rect 19061 28033 19073 28036
rect 19107 28064 19119 28067
rect 19613 28067 19671 28073
rect 19613 28064 19625 28067
rect 19107 28036 19625 28064
rect 19107 28033 19119 28036
rect 19061 28027 19119 28033
rect 19613 28033 19625 28036
rect 19659 28064 19671 28067
rect 20162 28064 20168 28076
rect 19659 28036 20168 28064
rect 19659 28033 19671 28036
rect 19613 28027 19671 28033
rect 20162 28024 20168 28036
rect 20220 28064 20226 28076
rect 20349 28067 20407 28073
rect 20349 28064 20361 28067
rect 20220 28036 20361 28064
rect 20220 28024 20226 28036
rect 20349 28033 20361 28036
rect 20395 28033 20407 28067
rect 20349 28027 20407 28033
rect 16264 27968 17172 27996
rect 16264 27956 16270 27968
rect 17586 27956 17592 28008
rect 17644 27996 17650 28008
rect 19978 27996 19984 28008
rect 17644 27968 19984 27996
rect 17644 27956 17650 27968
rect 19978 27956 19984 27968
rect 20036 27956 20042 28008
rect 20073 27999 20131 28005
rect 20073 27965 20085 27999
rect 20119 27996 20131 27999
rect 20622 27996 20628 28008
rect 20119 27968 20628 27996
rect 20119 27965 20131 27968
rect 20073 27959 20131 27965
rect 20622 27956 20628 27968
rect 20680 27996 20686 28008
rect 21008 27996 21036 28092
rect 22281 28067 22339 28073
rect 22281 28033 22293 28067
rect 22327 28064 22339 28067
rect 22738 28064 22744 28076
rect 22327 28036 22744 28064
rect 22327 28033 22339 28036
rect 22281 28027 22339 28033
rect 22738 28024 22744 28036
rect 22796 28024 22802 28076
rect 23106 28064 23112 28076
rect 22848 28036 23112 28064
rect 20680 27968 21036 27996
rect 20680 27956 20686 27968
rect 22462 27956 22468 28008
rect 22520 27996 22526 28008
rect 22848 27996 22876 28036
rect 23106 28024 23112 28036
rect 23164 28024 23170 28076
rect 26789 28067 26847 28073
rect 26789 28033 26801 28067
rect 26835 28064 26847 28067
rect 27614 28064 27620 28076
rect 26835 28036 27620 28064
rect 26835 28033 26847 28036
rect 26789 28027 26847 28033
rect 27614 28024 27620 28036
rect 27672 28024 27678 28076
rect 27709 28067 27767 28073
rect 27709 28033 27721 28067
rect 27755 28064 27767 28067
rect 28442 28064 28448 28076
rect 27755 28036 28448 28064
rect 27755 28033 27767 28036
rect 27709 28027 27767 28033
rect 28442 28024 28448 28036
rect 28500 28024 28506 28076
rect 28997 28067 29055 28073
rect 28997 28033 29009 28067
rect 29043 28064 29055 28067
rect 29380 28064 29408 28163
rect 29638 28160 29644 28212
rect 29696 28200 29702 28212
rect 29733 28203 29791 28209
rect 29733 28200 29745 28203
rect 29696 28172 29745 28200
rect 29696 28160 29702 28172
rect 29733 28169 29745 28172
rect 29779 28169 29791 28203
rect 29733 28163 29791 28169
rect 29825 28203 29883 28209
rect 29825 28169 29837 28203
rect 29871 28200 29883 28203
rect 29914 28200 29920 28212
rect 29871 28172 29920 28200
rect 29871 28169 29883 28172
rect 29825 28163 29883 28169
rect 29748 28132 29776 28163
rect 29914 28160 29920 28172
rect 29972 28160 29978 28212
rect 31570 28200 31576 28212
rect 30300 28172 31576 28200
rect 30300 28132 30328 28172
rect 31570 28160 31576 28172
rect 31628 28160 31634 28212
rect 31757 28203 31815 28209
rect 31757 28169 31769 28203
rect 31803 28169 31815 28203
rect 31757 28163 31815 28169
rect 31772 28132 31800 28163
rect 32490 28160 32496 28212
rect 32548 28200 32554 28212
rect 33505 28203 33563 28209
rect 32548 28172 32812 28200
rect 32548 28160 32554 28172
rect 32370 28135 32428 28141
rect 32370 28132 32382 28135
rect 29748 28104 30328 28132
rect 30392 28104 30696 28132
rect 31772 28104 32382 28132
rect 30392 28064 30420 28104
rect 29043 28036 29408 28064
rect 29472 28036 30420 28064
rect 29043 28033 29055 28036
rect 28997 28027 29055 28033
rect 22520 27968 22876 27996
rect 22520 27956 22526 27968
rect 22922 27956 22928 28008
rect 22980 27996 22986 28008
rect 23201 27999 23259 28005
rect 23201 27996 23213 27999
rect 22980 27968 23213 27996
rect 22980 27956 22986 27968
rect 23201 27965 23213 27968
rect 23247 27965 23259 27999
rect 23201 27959 23259 27965
rect 23382 27956 23388 28008
rect 23440 27956 23446 28008
rect 23934 27996 23940 28008
rect 23492 27968 23940 27996
rect 13219 27900 14872 27928
rect 13219 27897 13231 27900
rect 13173 27891 13231 27897
rect 1946 27820 1952 27872
rect 2004 27860 2010 27872
rect 2133 27863 2191 27869
rect 2133 27860 2145 27863
rect 2004 27832 2145 27860
rect 2004 27820 2010 27832
rect 2133 27829 2145 27832
rect 2179 27829 2191 27863
rect 2133 27823 2191 27829
rect 3970 27820 3976 27872
rect 4028 27820 4034 27872
rect 7193 27863 7251 27869
rect 7193 27829 7205 27863
rect 7239 27860 7251 27863
rect 7374 27860 7380 27872
rect 7239 27832 7380 27860
rect 7239 27829 7251 27832
rect 7193 27823 7251 27829
rect 7374 27820 7380 27832
rect 7432 27820 7438 27872
rect 7469 27863 7527 27869
rect 7469 27829 7481 27863
rect 7515 27860 7527 27863
rect 8386 27860 8392 27872
rect 7515 27832 8392 27860
rect 7515 27829 7527 27832
rect 7469 27823 7527 27829
rect 8386 27820 8392 27832
rect 8444 27820 8450 27872
rect 12710 27820 12716 27872
rect 12768 27860 12774 27872
rect 13188 27860 13216 27891
rect 19518 27888 19524 27940
rect 19576 27928 19582 27940
rect 19576 27900 22784 27928
rect 19576 27888 19582 27900
rect 12768 27832 13216 27860
rect 16209 27863 16267 27869
rect 12768 27820 12774 27832
rect 16209 27829 16221 27863
rect 16255 27860 16267 27863
rect 16482 27860 16488 27872
rect 16255 27832 16488 27860
rect 16255 27829 16267 27832
rect 16209 27823 16267 27829
rect 16482 27820 16488 27832
rect 16540 27820 16546 27872
rect 18046 27820 18052 27872
rect 18104 27860 18110 27872
rect 18785 27863 18843 27869
rect 18785 27860 18797 27863
rect 18104 27832 18797 27860
rect 18104 27820 18110 27832
rect 18785 27829 18797 27832
rect 18831 27860 18843 27863
rect 18874 27860 18880 27872
rect 18831 27832 18880 27860
rect 18831 27829 18843 27832
rect 18785 27823 18843 27829
rect 18874 27820 18880 27832
rect 18932 27820 18938 27872
rect 19334 27820 19340 27872
rect 19392 27860 19398 27872
rect 19610 27860 19616 27872
rect 19392 27832 19616 27860
rect 19392 27820 19398 27832
rect 19610 27820 19616 27832
rect 19668 27820 19674 27872
rect 19886 27820 19892 27872
rect 19944 27820 19950 27872
rect 20806 27820 20812 27872
rect 20864 27860 20870 27872
rect 22094 27860 22100 27872
rect 20864 27832 22100 27860
rect 20864 27820 20870 27832
rect 22094 27820 22100 27832
rect 22152 27820 22158 27872
rect 22756 27860 22784 27900
rect 22830 27888 22836 27940
rect 22888 27928 22894 27940
rect 23492 27928 23520 27968
rect 23934 27956 23940 27968
rect 23992 27996 23998 28008
rect 24302 28005 24308 28008
rect 24121 27999 24179 28005
rect 24121 27996 24133 27999
rect 23992 27968 24133 27996
rect 23992 27956 23998 27968
rect 24121 27965 24133 27968
rect 24167 27965 24179 27999
rect 24121 27959 24179 27965
rect 24259 27999 24308 28005
rect 24259 27965 24271 27999
rect 24305 27965 24308 27999
rect 24259 27959 24308 27965
rect 24302 27956 24308 27959
rect 24360 27956 24366 28008
rect 24394 27956 24400 28008
rect 24452 27956 24458 28008
rect 25133 27999 25191 28005
rect 25133 27965 25145 27999
rect 25179 27996 25191 27999
rect 25222 27996 25228 28008
rect 25179 27968 25228 27996
rect 25179 27965 25191 27968
rect 25133 27959 25191 27965
rect 25222 27956 25228 27968
rect 25280 27956 25286 28008
rect 27893 27999 27951 28005
rect 27893 27965 27905 27999
rect 27939 27965 27951 27999
rect 27893 27959 27951 27965
rect 22888 27900 23520 27928
rect 22888 27888 22894 27900
rect 23842 27888 23848 27940
rect 23900 27888 23906 27940
rect 25041 27931 25099 27937
rect 25041 27897 25053 27931
rect 25087 27928 25099 27931
rect 25409 27931 25467 27937
rect 25409 27928 25421 27931
rect 25087 27900 25421 27928
rect 25087 27897 25099 27900
rect 25041 27891 25099 27897
rect 25409 27897 25421 27900
rect 25455 27897 25467 27931
rect 25409 27891 25467 27897
rect 26878 27888 26884 27940
rect 26936 27928 26942 27940
rect 27908 27928 27936 27959
rect 28258 27956 28264 28008
rect 28316 27996 28322 28008
rect 29472 27996 29500 28036
rect 30558 28024 30564 28076
rect 30616 28024 30622 28076
rect 30668 28064 30696 28104
rect 32370 28101 32382 28104
rect 32416 28101 32428 28135
rect 32370 28095 32428 28101
rect 32582 28092 32588 28144
rect 32640 28092 32646 28144
rect 30668 28036 31754 28064
rect 28316 27968 29500 27996
rect 28316 27956 28322 27968
rect 30006 27956 30012 28008
rect 30064 27956 30070 28008
rect 30653 27999 30711 28005
rect 30653 27965 30665 27999
rect 30699 27965 30711 27999
rect 30653 27959 30711 27965
rect 26936 27900 27936 27928
rect 26936 27888 26942 27900
rect 27982 27888 27988 27940
rect 28040 27928 28046 27940
rect 30466 27928 30472 27940
rect 28040 27900 30472 27928
rect 28040 27888 28046 27900
rect 30466 27888 30472 27900
rect 30524 27888 30530 27940
rect 23860 27860 23888 27888
rect 22756 27832 23888 27860
rect 25590 27820 25596 27872
rect 25648 27820 25654 27872
rect 27341 27863 27399 27869
rect 27341 27829 27353 27863
rect 27387 27860 27399 27863
rect 28718 27860 28724 27872
rect 27387 27832 28724 27860
rect 27387 27829 27399 27832
rect 27341 27823 27399 27829
rect 28718 27820 28724 27832
rect 28776 27820 28782 27872
rect 28994 27820 29000 27872
rect 29052 27860 29058 27872
rect 30193 27863 30251 27869
rect 30193 27860 30205 27863
rect 29052 27832 30205 27860
rect 29052 27820 29058 27832
rect 30193 27829 30205 27832
rect 30239 27829 30251 27863
rect 30668 27860 30696 27959
rect 30742 27956 30748 28008
rect 30800 27956 30806 28008
rect 31726 27928 31754 28036
rect 31938 28024 31944 28076
rect 31996 28024 32002 28076
rect 32600 28064 32628 28092
rect 32048 28036 32628 28064
rect 32784 28064 32812 28172
rect 33505 28169 33517 28203
rect 33551 28169 33563 28203
rect 33505 28163 33563 28169
rect 32858 28092 32864 28144
rect 32916 28132 32922 28144
rect 33520 28132 33548 28163
rect 39114 28160 39120 28212
rect 39172 28200 39178 28212
rect 39761 28203 39819 28209
rect 39761 28200 39773 28203
rect 39172 28172 39773 28200
rect 39172 28160 39178 28172
rect 39761 28169 39773 28172
rect 39807 28169 39819 28203
rect 39761 28163 39819 28169
rect 41693 28203 41751 28209
rect 41693 28169 41705 28203
rect 41739 28200 41751 28203
rect 41782 28200 41788 28212
rect 41739 28172 41788 28200
rect 41739 28169 41751 28172
rect 41693 28163 41751 28169
rect 41782 28160 41788 28172
rect 41840 28160 41846 28212
rect 42153 28203 42211 28209
rect 42153 28169 42165 28203
rect 42199 28200 42211 28203
rect 42199 28172 42472 28200
rect 42199 28169 42211 28172
rect 42153 28163 42211 28169
rect 33594 28132 33600 28144
rect 32916 28104 33600 28132
rect 32916 28092 32922 28104
rect 33594 28092 33600 28104
rect 33652 28092 33658 28144
rect 39206 28092 39212 28144
rect 39264 28132 39270 28144
rect 39393 28135 39451 28141
rect 39393 28132 39405 28135
rect 39264 28104 39405 28132
rect 39264 28092 39270 28104
rect 39393 28101 39405 28104
rect 39439 28101 39451 28135
rect 40494 28132 40500 28144
rect 39393 28095 39451 28101
rect 40144 28104 40500 28132
rect 40144 28076 40172 28104
rect 40494 28092 40500 28104
rect 40552 28092 40558 28144
rect 42444 28141 42472 28172
rect 42610 28160 42616 28212
rect 42668 28209 42674 28212
rect 42668 28203 42687 28209
rect 42675 28169 42687 28203
rect 44269 28203 44327 28209
rect 44269 28200 44281 28203
rect 42668 28163 42687 28169
rect 42812 28172 44281 28200
rect 42668 28160 42674 28163
rect 42429 28135 42487 28141
rect 41386 28104 41920 28132
rect 38197 28067 38255 28073
rect 32784 28036 33640 28064
rect 32048 27928 32076 28036
rect 32122 27956 32128 28008
rect 32180 27956 32186 28008
rect 33612 28005 33640 28036
rect 38197 28033 38209 28067
rect 38243 28064 38255 28067
rect 38746 28064 38752 28076
rect 38243 28036 38752 28064
rect 38243 28033 38255 28036
rect 38197 28027 38255 28033
rect 38746 28024 38752 28036
rect 38804 28024 38810 28076
rect 39942 28024 39948 28076
rect 40000 28024 40006 28076
rect 40037 28067 40095 28073
rect 40037 28033 40049 28067
rect 40083 28064 40095 28067
rect 40126 28064 40132 28076
rect 40083 28036 40132 28064
rect 40083 28033 40095 28036
rect 40037 28027 40095 28033
rect 40126 28024 40132 28036
rect 40184 28024 40190 28076
rect 40218 28024 40224 28076
rect 40276 28024 40282 28076
rect 40313 28067 40371 28073
rect 40313 28033 40325 28067
rect 40359 28064 40371 28067
rect 41386 28064 41414 28104
rect 40359 28036 41414 28064
rect 40359 28033 40371 28036
rect 40313 28027 40371 28033
rect 41506 28024 41512 28076
rect 41564 28024 41570 28076
rect 41785 28067 41843 28073
rect 41785 28033 41797 28067
rect 41831 28033 41843 28067
rect 41892 28064 41920 28104
rect 42429 28101 42441 28135
rect 42475 28101 42487 28135
rect 42429 28095 42487 28101
rect 42812 28064 42840 28172
rect 44269 28169 44281 28172
rect 44315 28169 44327 28203
rect 44269 28163 44327 28169
rect 44910 28160 44916 28212
rect 44968 28160 44974 28212
rect 46658 28160 46664 28212
rect 46716 28160 46722 28212
rect 43901 28135 43959 28141
rect 43901 28101 43913 28135
rect 43947 28132 43959 28135
rect 43990 28132 43996 28144
rect 43947 28104 43996 28132
rect 43947 28101 43959 28104
rect 43901 28095 43959 28101
rect 41892 28036 42840 28064
rect 41785 28027 41843 28033
rect 33597 27999 33655 28005
rect 33597 27965 33609 27999
rect 33643 27996 33655 27999
rect 35434 27996 35440 28008
rect 33643 27968 35440 27996
rect 33643 27965 33655 27968
rect 33597 27959 33655 27965
rect 35434 27956 35440 27968
rect 35492 27956 35498 28008
rect 38378 27956 38384 28008
rect 38436 27956 38442 28008
rect 41322 27956 41328 28008
rect 41380 27956 41386 28008
rect 34514 27928 34520 27940
rect 31726 27900 32076 27928
rect 33428 27900 34520 27928
rect 33428 27860 33456 27900
rect 34514 27888 34520 27900
rect 34572 27888 34578 27940
rect 39577 27931 39635 27937
rect 39577 27897 39589 27931
rect 39623 27928 39635 27931
rect 39758 27928 39764 27940
rect 39623 27900 39764 27928
rect 39623 27897 39635 27900
rect 39577 27891 39635 27897
rect 39758 27888 39764 27900
rect 39816 27888 39822 27940
rect 30668 27832 33456 27860
rect 30193 27823 30251 27829
rect 33502 27820 33508 27872
rect 33560 27860 33566 27872
rect 33827 27863 33885 27869
rect 33827 27860 33839 27863
rect 33560 27832 33839 27860
rect 33560 27820 33566 27832
rect 33827 27829 33839 27832
rect 33873 27829 33885 27863
rect 33827 27823 33885 27829
rect 38194 27820 38200 27872
rect 38252 27860 38258 27872
rect 38562 27860 38568 27872
rect 38252 27832 38568 27860
rect 38252 27820 38258 27832
rect 38562 27820 38568 27832
rect 38620 27820 38626 27872
rect 38654 27820 38660 27872
rect 38712 27820 38718 27872
rect 40954 27820 40960 27872
rect 41012 27860 41018 27872
rect 41340 27860 41368 27956
rect 41800 27928 41828 28027
rect 43530 28024 43536 28076
rect 43588 28024 43594 28076
rect 41874 27956 41880 28008
rect 41932 27956 41938 28008
rect 42426 27956 42432 28008
rect 42484 27996 42490 28008
rect 43916 27996 43944 28095
rect 43990 28092 43996 28104
rect 44048 28092 44054 28144
rect 44082 28092 44088 28144
rect 44140 28141 44146 28144
rect 44140 28135 44159 28141
rect 44147 28101 44159 28135
rect 44140 28095 44159 28101
rect 44140 28092 44146 28095
rect 44542 28092 44548 28144
rect 44600 28092 44606 28144
rect 46014 28132 46020 28144
rect 44744 28104 46020 28132
rect 44361 28067 44419 28073
rect 44361 28033 44373 28067
rect 44407 28064 44419 28067
rect 44450 28064 44456 28076
rect 44407 28036 44456 28064
rect 44407 28033 44419 28036
rect 44361 28027 44419 28033
rect 44450 28024 44456 28036
rect 44508 28024 44514 28076
rect 44634 28024 44640 28076
rect 44692 28024 44698 28076
rect 44744 28073 44772 28104
rect 46014 28092 46020 28104
rect 46072 28092 46078 28144
rect 44729 28067 44787 28073
rect 44729 28033 44741 28067
rect 44775 28033 44787 28067
rect 44729 28027 44787 28033
rect 45186 28024 45192 28076
rect 45244 28024 45250 28076
rect 45373 28067 45431 28073
rect 45373 28033 45385 28067
rect 45419 28064 45431 28067
rect 45649 28067 45707 28073
rect 45649 28064 45661 28067
rect 45419 28036 45661 28064
rect 45419 28033 45431 28036
rect 45373 28027 45431 28033
rect 45649 28033 45661 28036
rect 45695 28033 45707 28067
rect 45649 28027 45707 28033
rect 46566 28024 46572 28076
rect 46624 28024 46630 28076
rect 45005 27999 45063 28005
rect 45005 27996 45017 27999
rect 42484 27968 43760 27996
rect 43916 27968 45017 27996
rect 42484 27956 42490 27968
rect 41966 27928 41972 27940
rect 41800 27900 41972 27928
rect 41966 27888 41972 27900
rect 42024 27928 42030 27940
rect 42518 27928 42524 27940
rect 42024 27900 42524 27928
rect 42024 27888 42030 27900
rect 42518 27888 42524 27900
rect 42576 27888 42582 27940
rect 42886 27928 42892 27940
rect 42628 27900 42892 27928
rect 42628 27872 42656 27900
rect 42886 27888 42892 27900
rect 42944 27928 42950 27940
rect 43530 27928 43536 27940
rect 42944 27900 43536 27928
rect 42944 27888 42950 27900
rect 43530 27888 43536 27900
rect 43588 27888 43594 27940
rect 43732 27937 43760 27968
rect 45005 27965 45017 27968
rect 45051 27965 45063 27999
rect 45005 27959 45063 27965
rect 43717 27931 43775 27937
rect 43717 27897 43729 27931
rect 43763 27897 43775 27931
rect 45204 27928 45232 28024
rect 43717 27891 43775 27897
rect 44100 27900 45232 27928
rect 41782 27860 41788 27872
rect 41012 27832 41788 27860
rect 41012 27820 41018 27832
rect 41782 27820 41788 27832
rect 41840 27820 41846 27872
rect 41877 27863 41935 27869
rect 41877 27829 41889 27863
rect 41923 27860 41935 27863
rect 42058 27860 42064 27872
rect 41923 27832 42064 27860
rect 41923 27829 41935 27832
rect 41877 27823 41935 27829
rect 42058 27820 42064 27832
rect 42116 27820 42122 27872
rect 42610 27820 42616 27872
rect 42668 27820 42674 27872
rect 42794 27820 42800 27872
rect 42852 27820 42858 27872
rect 43548 27860 43576 27888
rect 43990 27860 43996 27872
rect 43548 27832 43996 27860
rect 43990 27820 43996 27832
rect 44048 27820 44054 27872
rect 44100 27869 44128 27900
rect 44085 27863 44143 27869
rect 44085 27829 44097 27863
rect 44131 27829 44143 27863
rect 44085 27823 44143 27829
rect 45462 27820 45468 27872
rect 45520 27820 45526 27872
rect 1104 27770 47104 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 47104 27770
rect 1104 27696 47104 27718
rect 2958 27616 2964 27668
rect 3016 27656 3022 27668
rect 3053 27659 3111 27665
rect 3053 27656 3065 27659
rect 3016 27628 3065 27656
rect 3016 27616 3022 27628
rect 3053 27625 3065 27628
rect 3099 27625 3111 27659
rect 3053 27619 3111 27625
rect 3142 27616 3148 27668
rect 3200 27616 3206 27668
rect 4614 27616 4620 27668
rect 4672 27656 4678 27668
rect 5445 27659 5503 27665
rect 5445 27656 5457 27659
rect 4672 27628 5457 27656
rect 4672 27616 4678 27628
rect 5445 27625 5457 27628
rect 5491 27625 5503 27659
rect 5445 27619 5503 27625
rect 6454 27616 6460 27668
rect 6512 27616 6518 27668
rect 10962 27616 10968 27668
rect 11020 27616 11026 27668
rect 13814 27616 13820 27668
rect 13872 27656 13878 27668
rect 14967 27659 15025 27665
rect 14967 27656 14979 27659
rect 13872 27628 14979 27656
rect 13872 27616 13878 27628
rect 14967 27625 14979 27628
rect 15013 27656 15025 27659
rect 16298 27656 16304 27668
rect 15013 27628 16304 27656
rect 15013 27625 15025 27628
rect 14967 27619 15025 27625
rect 16298 27616 16304 27628
rect 16356 27616 16362 27668
rect 16574 27616 16580 27668
rect 16632 27656 16638 27668
rect 17586 27656 17592 27668
rect 16632 27628 17592 27656
rect 16632 27616 16638 27628
rect 17586 27616 17592 27628
rect 17644 27616 17650 27668
rect 17678 27616 17684 27668
rect 17736 27656 17742 27668
rect 22462 27656 22468 27668
rect 17736 27628 22468 27656
rect 17736 27616 17742 27628
rect 22462 27616 22468 27628
rect 22520 27616 22526 27668
rect 22649 27659 22707 27665
rect 22649 27656 22661 27659
rect 22572 27628 22661 27656
rect 8389 27591 8447 27597
rect 8389 27588 8401 27591
rect 4448 27560 8401 27588
rect 1670 27480 1676 27532
rect 1728 27480 1734 27532
rect 3050 27480 3056 27532
rect 3108 27520 3114 27532
rect 3602 27520 3608 27532
rect 3108 27492 3608 27520
rect 3108 27480 3114 27492
rect 3602 27480 3608 27492
rect 3660 27520 3666 27532
rect 4448 27529 4476 27560
rect 8389 27557 8401 27560
rect 8435 27588 8447 27591
rect 8662 27588 8668 27600
rect 8435 27560 8668 27588
rect 8435 27557 8447 27560
rect 8389 27551 8447 27557
rect 8662 27548 8668 27560
rect 8720 27548 8726 27600
rect 10980 27588 11008 27616
rect 12345 27591 12403 27597
rect 10336 27560 11100 27588
rect 4433 27523 4491 27529
rect 3660 27492 4384 27520
rect 3660 27480 3666 27492
rect 1946 27461 1952 27464
rect 1940 27452 1952 27461
rect 1907 27424 1952 27452
rect 1940 27415 1952 27424
rect 1946 27412 1952 27415
rect 2004 27412 2010 27464
rect 3329 27455 3387 27461
rect 3329 27421 3341 27455
rect 3375 27452 3387 27455
rect 3375 27424 3832 27452
rect 3375 27421 3387 27424
rect 3329 27415 3387 27421
rect 3804 27325 3832 27424
rect 3970 27412 3976 27464
rect 4028 27452 4034 27464
rect 4157 27455 4215 27461
rect 4157 27452 4169 27455
rect 4028 27424 4169 27452
rect 4028 27412 4034 27424
rect 4157 27421 4169 27424
rect 4203 27421 4215 27455
rect 4356 27452 4384 27492
rect 4433 27489 4445 27523
rect 4479 27489 4491 27523
rect 5997 27523 6055 27529
rect 5997 27520 6009 27523
rect 4433 27483 4491 27489
rect 4540 27492 6009 27520
rect 4540 27452 4568 27492
rect 5997 27489 6009 27492
rect 6043 27489 6055 27523
rect 5997 27483 6055 27489
rect 7466 27480 7472 27532
rect 7524 27520 7530 27532
rect 7929 27523 7987 27529
rect 7929 27520 7941 27523
rect 7524 27492 7941 27520
rect 7524 27480 7530 27492
rect 7929 27489 7941 27492
rect 7975 27520 7987 27523
rect 8018 27520 8024 27532
rect 7975 27492 8024 27520
rect 7975 27489 7987 27492
rect 7929 27483 7987 27489
rect 8018 27480 8024 27492
rect 8076 27480 8082 27532
rect 9122 27520 9128 27532
rect 8128 27492 9128 27520
rect 4356 27424 4568 27452
rect 5813 27455 5871 27461
rect 4157 27415 4215 27421
rect 5813 27421 5825 27455
rect 5859 27452 5871 27455
rect 5902 27452 5908 27464
rect 5859 27424 5908 27452
rect 5859 27421 5871 27424
rect 5813 27415 5871 27421
rect 5902 27412 5908 27424
rect 5960 27412 5966 27464
rect 6273 27455 6331 27461
rect 6273 27421 6285 27455
rect 6319 27452 6331 27455
rect 7006 27452 7012 27464
rect 6319 27424 7012 27452
rect 6319 27421 6331 27424
rect 6273 27415 6331 27421
rect 7006 27412 7012 27424
rect 7064 27452 7070 27464
rect 8128 27452 8156 27492
rect 9122 27480 9128 27492
rect 9180 27480 9186 27532
rect 10134 27480 10140 27532
rect 10192 27480 10198 27532
rect 10336 27529 10364 27560
rect 10321 27523 10379 27529
rect 10321 27489 10333 27523
rect 10367 27489 10379 27523
rect 10321 27483 10379 27489
rect 10594 27480 10600 27532
rect 10652 27520 10658 27532
rect 11072 27529 11100 27560
rect 12345 27557 12357 27591
rect 12391 27588 12403 27591
rect 12618 27588 12624 27600
rect 12391 27560 12624 27588
rect 12391 27557 12403 27560
rect 12345 27551 12403 27557
rect 12618 27548 12624 27560
rect 12676 27548 12682 27600
rect 13906 27548 13912 27600
rect 13964 27588 13970 27600
rect 17034 27588 17040 27600
rect 13964 27560 17040 27588
rect 13964 27548 13970 27560
rect 17034 27548 17040 27560
rect 17092 27548 17098 27600
rect 18601 27591 18659 27597
rect 18601 27557 18613 27591
rect 18647 27588 18659 27591
rect 18690 27588 18696 27600
rect 18647 27560 18696 27588
rect 18647 27557 18659 27560
rect 18601 27551 18659 27557
rect 18690 27548 18696 27560
rect 18748 27548 18754 27600
rect 18966 27548 18972 27600
rect 19024 27548 19030 27600
rect 19613 27591 19671 27597
rect 19613 27557 19625 27591
rect 19659 27588 19671 27591
rect 19794 27588 19800 27600
rect 19659 27560 19800 27588
rect 19659 27557 19671 27560
rect 19613 27551 19671 27557
rect 19794 27548 19800 27560
rect 19852 27548 19858 27600
rect 10965 27523 11023 27529
rect 10965 27520 10977 27523
rect 10652 27492 10977 27520
rect 10652 27480 10658 27492
rect 10965 27489 10977 27492
rect 11011 27489 11023 27523
rect 10965 27483 11023 27489
rect 11057 27523 11115 27529
rect 11057 27489 11069 27523
rect 11103 27489 11115 27523
rect 11057 27483 11115 27489
rect 11974 27480 11980 27532
rect 12032 27520 12038 27532
rect 12437 27523 12495 27529
rect 12437 27520 12449 27523
rect 12032 27492 12449 27520
rect 12032 27480 12038 27492
rect 12437 27489 12449 27492
rect 12483 27520 12495 27523
rect 14274 27520 14280 27532
rect 12483 27492 14280 27520
rect 12483 27489 12495 27492
rect 12437 27483 12495 27489
rect 14274 27480 14280 27492
rect 14332 27480 14338 27532
rect 14553 27523 14611 27529
rect 14553 27489 14565 27523
rect 14599 27520 14611 27523
rect 14642 27520 14648 27532
rect 14599 27492 14648 27520
rect 14599 27489 14611 27492
rect 14553 27483 14611 27489
rect 14642 27480 14648 27492
rect 14700 27480 14706 27532
rect 14737 27523 14795 27529
rect 14737 27489 14749 27523
rect 14783 27520 14795 27523
rect 15102 27520 15108 27532
rect 14783 27492 15108 27520
rect 14783 27489 14795 27492
rect 14737 27483 14795 27489
rect 15102 27480 15108 27492
rect 15160 27480 15166 27532
rect 16577 27523 16635 27529
rect 16577 27489 16589 27523
rect 16623 27520 16635 27523
rect 16623 27492 19380 27520
rect 16623 27489 16635 27492
rect 16577 27483 16635 27489
rect 7064 27424 8156 27452
rect 7064 27412 7070 27424
rect 8202 27412 8208 27464
rect 8260 27452 8266 27464
rect 8260 27424 12434 27452
rect 8260 27412 8266 27424
rect 7745 27387 7803 27393
rect 7745 27353 7757 27387
rect 7791 27384 7803 27387
rect 8294 27384 8300 27396
rect 7791 27356 8300 27384
rect 7791 27353 7803 27356
rect 7745 27347 7803 27353
rect 8294 27344 8300 27356
rect 8352 27384 8358 27396
rect 9306 27384 9312 27396
rect 8352 27356 9312 27384
rect 8352 27344 8358 27356
rect 9306 27344 9312 27356
rect 9364 27344 9370 27396
rect 11330 27344 11336 27396
rect 11388 27384 11394 27396
rect 11977 27387 12035 27393
rect 11977 27384 11989 27387
rect 11388 27356 11989 27384
rect 11388 27344 11394 27356
rect 11977 27353 11989 27356
rect 12023 27353 12035 27387
rect 12406 27384 12434 27424
rect 13262 27412 13268 27464
rect 13320 27452 13326 27464
rect 13320 27424 14780 27452
rect 13320 27412 13326 27424
rect 12894 27384 12900 27396
rect 12406 27356 12900 27384
rect 11977 27347 12035 27353
rect 12894 27344 12900 27356
rect 12952 27344 12958 27396
rect 14277 27387 14335 27393
rect 14277 27353 14289 27387
rect 14323 27384 14335 27387
rect 14642 27384 14648 27396
rect 14323 27356 14648 27384
rect 14323 27353 14335 27356
rect 14277 27347 14335 27353
rect 14642 27344 14648 27356
rect 14700 27344 14706 27396
rect 3789 27319 3847 27325
rect 3789 27285 3801 27319
rect 3835 27285 3847 27319
rect 3789 27279 3847 27285
rect 4062 27276 4068 27328
rect 4120 27316 4126 27328
rect 4249 27319 4307 27325
rect 4249 27316 4261 27319
rect 4120 27288 4261 27316
rect 4120 27276 4126 27288
rect 4249 27285 4261 27288
rect 4295 27285 4307 27319
rect 4249 27279 4307 27285
rect 5902 27276 5908 27328
rect 5960 27276 5966 27328
rect 7190 27276 7196 27328
rect 7248 27316 7254 27328
rect 7377 27319 7435 27325
rect 7377 27316 7389 27319
rect 7248 27288 7389 27316
rect 7248 27276 7254 27288
rect 7377 27285 7389 27288
rect 7423 27285 7435 27319
rect 7377 27279 7435 27285
rect 7837 27319 7895 27325
rect 7837 27285 7849 27319
rect 7883 27316 7895 27319
rect 7926 27316 7932 27328
rect 7883 27288 7932 27316
rect 7883 27285 7895 27288
rect 7837 27279 7895 27285
rect 7926 27276 7932 27288
rect 7984 27276 7990 27328
rect 9677 27319 9735 27325
rect 9677 27285 9689 27319
rect 9723 27316 9735 27319
rect 9950 27316 9956 27328
rect 9723 27288 9956 27316
rect 9723 27285 9735 27288
rect 9677 27279 9735 27285
rect 9950 27276 9956 27288
rect 10008 27276 10014 27328
rect 10042 27276 10048 27328
rect 10100 27276 10106 27328
rect 10505 27319 10563 27325
rect 10505 27285 10517 27319
rect 10551 27316 10563 27319
rect 10778 27316 10784 27328
rect 10551 27288 10784 27316
rect 10551 27285 10563 27288
rect 10505 27279 10563 27285
rect 10778 27276 10784 27288
rect 10836 27276 10842 27328
rect 10873 27319 10931 27325
rect 10873 27285 10885 27319
rect 10919 27316 10931 27319
rect 11790 27316 11796 27328
rect 10919 27288 11796 27316
rect 10919 27285 10931 27288
rect 10873 27279 10931 27285
rect 11790 27276 11796 27288
rect 11848 27316 11854 27328
rect 12526 27316 12532 27328
rect 11848 27288 12532 27316
rect 11848 27276 11854 27288
rect 12526 27276 12532 27288
rect 12584 27316 12590 27328
rect 13262 27316 13268 27328
rect 12584 27288 13268 27316
rect 12584 27276 12590 27288
rect 13262 27276 13268 27288
rect 13320 27276 13326 27328
rect 14752 27316 14780 27424
rect 15194 27412 15200 27464
rect 15252 27452 15258 27464
rect 16942 27452 16948 27464
rect 15252 27424 16948 27452
rect 15252 27412 15258 27424
rect 16942 27412 16948 27424
rect 17000 27412 17006 27464
rect 17034 27412 17040 27464
rect 17092 27412 17098 27464
rect 18325 27455 18383 27461
rect 18325 27421 18337 27455
rect 18371 27452 18383 27455
rect 18414 27452 18420 27464
rect 18371 27424 18420 27452
rect 18371 27421 18383 27424
rect 18325 27415 18383 27421
rect 18414 27412 18420 27424
rect 18472 27412 18478 27464
rect 18690 27412 18696 27464
rect 18748 27452 18754 27464
rect 19352 27461 19380 27492
rect 21542 27461 21548 27464
rect 18785 27455 18843 27461
rect 18785 27452 18797 27455
rect 18748 27424 18797 27452
rect 18748 27412 18754 27424
rect 18785 27421 18797 27424
rect 18831 27421 18843 27455
rect 18785 27415 18843 27421
rect 19337 27455 19395 27461
rect 19337 27421 19349 27455
rect 19383 27421 19395 27455
rect 19337 27415 19395 27421
rect 19797 27455 19855 27461
rect 19797 27421 19809 27455
rect 19843 27452 19855 27455
rect 21269 27455 21327 27461
rect 21269 27452 21281 27455
rect 19843 27424 21281 27452
rect 19843 27421 19855 27424
rect 19797 27415 19855 27421
rect 21269 27421 21281 27424
rect 21315 27421 21327 27455
rect 21536 27452 21548 27461
rect 21503 27424 21548 27452
rect 21269 27415 21327 27421
rect 21536 27415 21548 27424
rect 16390 27344 16396 27396
rect 16448 27384 16454 27396
rect 16485 27387 16543 27393
rect 16485 27384 16497 27387
rect 16448 27356 16497 27384
rect 16448 27344 16454 27356
rect 16485 27353 16497 27356
rect 16531 27353 16543 27387
rect 17129 27387 17187 27393
rect 17129 27384 17141 27387
rect 16485 27347 16543 27353
rect 16592 27356 17141 27384
rect 15838 27316 15844 27328
rect 14752 27288 15844 27316
rect 15838 27276 15844 27288
rect 15896 27316 15902 27328
rect 16592 27316 16620 27356
rect 17129 27353 17141 27356
rect 17175 27353 17187 27387
rect 17129 27347 17187 27353
rect 17497 27387 17555 27393
rect 17497 27353 17509 27387
rect 17543 27353 17555 27387
rect 17497 27347 17555 27353
rect 15896 27288 16620 27316
rect 15896 27276 15902 27288
rect 16666 27276 16672 27328
rect 16724 27316 16730 27328
rect 17512 27316 17540 27347
rect 16724 27288 17540 27316
rect 19352 27316 19380 27415
rect 20064 27387 20122 27393
rect 20064 27353 20076 27387
rect 20110 27384 20122 27387
rect 20346 27384 20352 27396
rect 20110 27356 20352 27384
rect 20110 27353 20122 27356
rect 20064 27347 20122 27353
rect 20346 27344 20352 27356
rect 20404 27344 20410 27396
rect 21284 27384 21312 27415
rect 21542 27412 21548 27415
rect 21600 27412 21606 27464
rect 22094 27412 22100 27464
rect 22152 27452 22158 27464
rect 22572 27452 22600 27628
rect 22649 27625 22661 27628
rect 22695 27625 22707 27659
rect 22649 27619 22707 27625
rect 23198 27616 23204 27668
rect 23256 27656 23262 27668
rect 24026 27656 24032 27668
rect 23256 27628 24032 27656
rect 23256 27616 23262 27628
rect 24026 27616 24032 27628
rect 24084 27656 24090 27668
rect 24084 27628 25360 27656
rect 24084 27616 24090 27628
rect 22833 27591 22891 27597
rect 22833 27557 22845 27591
rect 22879 27588 22891 27591
rect 25332 27588 25360 27628
rect 28442 27616 28448 27668
rect 28500 27616 28506 27668
rect 29273 27659 29331 27665
rect 29273 27625 29285 27659
rect 29319 27656 29331 27659
rect 30006 27656 30012 27668
rect 29319 27628 30012 27656
rect 29319 27625 29331 27628
rect 29273 27619 29331 27625
rect 30006 27616 30012 27628
rect 30064 27616 30070 27668
rect 30558 27616 30564 27668
rect 30616 27656 30622 27668
rect 31389 27659 31447 27665
rect 31389 27656 31401 27659
rect 30616 27628 31401 27656
rect 30616 27616 30622 27628
rect 31389 27625 31401 27628
rect 31435 27625 31447 27659
rect 36630 27656 36636 27668
rect 31389 27619 31447 27625
rect 35268 27628 36636 27656
rect 26237 27591 26295 27597
rect 22879 27560 24440 27588
rect 25332 27560 26096 27588
rect 22879 27557 22891 27560
rect 22833 27551 22891 27557
rect 23382 27480 23388 27532
rect 23440 27520 23446 27532
rect 24121 27523 24179 27529
rect 23440 27492 23888 27520
rect 23440 27480 23446 27492
rect 22830 27452 22836 27464
rect 22152 27424 22836 27452
rect 22152 27412 22158 27424
rect 22830 27412 22836 27424
rect 22888 27412 22894 27464
rect 23017 27455 23075 27461
rect 23017 27421 23029 27455
rect 23063 27452 23075 27455
rect 23063 27424 23428 27452
rect 23063 27421 23075 27424
rect 23017 27415 23075 27421
rect 23106 27384 23112 27396
rect 21284 27356 23112 27384
rect 23106 27344 23112 27356
rect 23164 27344 23170 27396
rect 23198 27344 23204 27396
rect 23256 27344 23262 27396
rect 20162 27316 20168 27328
rect 19352 27288 20168 27316
rect 16724 27276 16730 27288
rect 20162 27276 20168 27288
rect 20220 27276 20226 27328
rect 21177 27319 21235 27325
rect 21177 27285 21189 27319
rect 21223 27316 21235 27319
rect 22186 27316 22192 27328
rect 21223 27288 22192 27316
rect 21223 27285 21235 27288
rect 21177 27279 21235 27285
rect 22186 27276 22192 27288
rect 22244 27276 22250 27328
rect 22462 27276 22468 27328
rect 22520 27316 22526 27328
rect 22738 27316 22744 27328
rect 22520 27288 22744 27316
rect 22520 27276 22526 27288
rect 22738 27276 22744 27288
rect 22796 27316 22802 27328
rect 23293 27319 23351 27325
rect 23293 27316 23305 27319
rect 22796 27288 23305 27316
rect 22796 27276 22802 27288
rect 23293 27285 23305 27288
rect 23339 27285 23351 27319
rect 23400 27316 23428 27424
rect 23860 27393 23888 27492
rect 24121 27489 24133 27523
rect 24167 27489 24179 27523
rect 24412 27520 24440 27560
rect 24412 27492 24532 27520
rect 24121 27483 24179 27489
rect 23937 27455 23995 27461
rect 23937 27421 23949 27455
rect 23983 27452 23995 27455
rect 24026 27452 24032 27464
rect 23983 27424 24032 27452
rect 23983 27421 23995 27424
rect 23937 27415 23995 27421
rect 24026 27412 24032 27424
rect 24084 27412 24090 27464
rect 23845 27387 23903 27393
rect 23845 27353 23857 27387
rect 23891 27384 23903 27387
rect 24136 27384 24164 27483
rect 24210 27412 24216 27464
rect 24268 27452 24274 27464
rect 24397 27455 24455 27461
rect 24397 27452 24409 27455
rect 24268 27424 24409 27452
rect 24268 27412 24274 27424
rect 24397 27421 24409 27424
rect 24443 27421 24455 27455
rect 24504 27452 24532 27492
rect 24653 27455 24711 27461
rect 24653 27452 24665 27455
rect 24504 27424 24665 27452
rect 24397 27415 24455 27421
rect 24653 27421 24665 27424
rect 24699 27421 24711 27455
rect 24653 27415 24711 27421
rect 24762 27384 24768 27396
rect 23891 27356 24072 27384
rect 24136 27356 24768 27384
rect 23891 27353 23903 27356
rect 23845 27347 23903 27353
rect 23477 27319 23535 27325
rect 23477 27316 23489 27319
rect 23400 27288 23489 27316
rect 23293 27279 23351 27285
rect 23477 27285 23489 27288
rect 23523 27285 23535 27319
rect 24044 27316 24072 27356
rect 24762 27344 24768 27356
rect 24820 27344 24826 27396
rect 26068 27384 26096 27560
rect 26237 27557 26249 27591
rect 26283 27557 26295 27591
rect 26237 27551 26295 27557
rect 26145 27455 26203 27461
rect 26145 27421 26157 27455
rect 26191 27452 26203 27455
rect 26252 27452 26280 27551
rect 26326 27480 26332 27532
rect 26384 27520 26390 27532
rect 26789 27523 26847 27529
rect 26789 27520 26801 27523
rect 26384 27492 26801 27520
rect 26384 27480 26390 27492
rect 26789 27489 26801 27492
rect 26835 27489 26847 27523
rect 28460 27520 28488 27616
rect 29638 27548 29644 27600
rect 29696 27588 29702 27600
rect 29696 27560 30328 27588
rect 29696 27548 29702 27560
rect 28460 27492 28948 27520
rect 26789 27483 26847 27489
rect 26191 27424 26280 27452
rect 27065 27455 27123 27461
rect 26191 27421 26203 27424
rect 26145 27415 26203 27421
rect 27065 27421 27077 27455
rect 27111 27452 27123 27455
rect 27614 27452 27620 27464
rect 27111 27424 27620 27452
rect 27111 27421 27123 27424
rect 27065 27415 27123 27421
rect 27614 27412 27620 27424
rect 27672 27452 27678 27464
rect 28534 27452 28540 27464
rect 27672 27424 28540 27452
rect 27672 27412 27678 27424
rect 28534 27412 28540 27424
rect 28592 27412 28598 27464
rect 28718 27412 28724 27464
rect 28776 27412 28782 27464
rect 27332 27387 27390 27393
rect 26068 27356 26740 27384
rect 25777 27319 25835 27325
rect 25777 27316 25789 27319
rect 24044 27288 25789 27316
rect 23477 27279 23535 27285
rect 25777 27285 25789 27288
rect 25823 27285 25835 27319
rect 25777 27279 25835 27285
rect 25961 27319 26019 27325
rect 25961 27285 25973 27319
rect 26007 27316 26019 27319
rect 26510 27316 26516 27328
rect 26007 27288 26516 27316
rect 26007 27285 26019 27288
rect 25961 27279 26019 27285
rect 26510 27276 26516 27288
rect 26568 27276 26574 27328
rect 26602 27276 26608 27328
rect 26660 27276 26666 27328
rect 26712 27325 26740 27356
rect 27332 27353 27344 27387
rect 27378 27384 27390 27387
rect 27378 27356 28580 27384
rect 27378 27353 27390 27356
rect 27332 27347 27390 27353
rect 26697 27319 26755 27325
rect 26697 27285 26709 27319
rect 26743 27316 26755 27319
rect 27982 27316 27988 27328
rect 26743 27288 27988 27316
rect 26743 27285 26755 27288
rect 26697 27279 26755 27285
rect 27982 27276 27988 27288
rect 28040 27276 28046 27328
rect 28552 27325 28580 27356
rect 28537 27319 28595 27325
rect 28537 27285 28549 27319
rect 28583 27285 28595 27319
rect 28920 27316 28948 27492
rect 29086 27480 29092 27532
rect 29144 27520 29150 27532
rect 29733 27523 29791 27529
rect 29733 27520 29745 27523
rect 29144 27492 29745 27520
rect 29144 27480 29150 27492
rect 29733 27489 29745 27492
rect 29779 27520 29791 27523
rect 29914 27520 29920 27532
rect 29779 27492 29920 27520
rect 29779 27489 29791 27492
rect 29733 27483 29791 27489
rect 29914 27480 29920 27492
rect 29972 27480 29978 27532
rect 30190 27480 30196 27532
rect 30248 27480 30254 27532
rect 30300 27520 30328 27560
rect 32600 27560 33456 27588
rect 30586 27523 30644 27529
rect 30586 27520 30598 27523
rect 30300 27492 30598 27520
rect 30586 27489 30598 27492
rect 30632 27489 30644 27523
rect 30586 27483 30644 27489
rect 30745 27523 30803 27529
rect 30745 27489 30757 27523
rect 30791 27520 30803 27523
rect 30926 27520 30932 27532
rect 30791 27492 30932 27520
rect 30791 27489 30803 27492
rect 30745 27483 30803 27489
rect 30926 27480 30932 27492
rect 30984 27480 30990 27532
rect 31294 27480 31300 27532
rect 31352 27520 31358 27532
rect 32401 27523 32459 27529
rect 32401 27520 32413 27523
rect 31352 27492 32413 27520
rect 31352 27480 31358 27492
rect 32401 27489 32413 27492
rect 32447 27489 32459 27523
rect 32401 27483 32459 27489
rect 29546 27412 29552 27464
rect 29604 27412 29610 27464
rect 30466 27412 30472 27464
rect 30524 27412 30530 27464
rect 32217 27455 32275 27461
rect 32217 27421 32229 27455
rect 32263 27452 32275 27455
rect 32600 27452 32628 27560
rect 32674 27480 32680 27532
rect 32732 27480 32738 27532
rect 33226 27480 33232 27532
rect 33284 27520 33290 27532
rect 33321 27523 33379 27529
rect 33321 27520 33333 27523
rect 33284 27492 33333 27520
rect 33284 27480 33290 27492
rect 33321 27489 33333 27492
rect 33367 27489 33379 27523
rect 33428 27520 33456 27560
rect 34514 27548 34520 27600
rect 34572 27548 34578 27600
rect 33714 27523 33772 27529
rect 33714 27520 33726 27523
rect 33428 27492 33726 27520
rect 33321 27483 33379 27489
rect 33714 27489 33726 27492
rect 33760 27520 33772 27523
rect 34054 27520 34060 27532
rect 33760 27492 34060 27520
rect 33760 27489 33772 27492
rect 33714 27483 33772 27489
rect 34054 27480 34060 27492
rect 34112 27480 34118 27532
rect 35268 27529 35296 27628
rect 36630 27616 36636 27628
rect 36688 27616 36694 27668
rect 37642 27616 37648 27668
rect 37700 27616 37706 27668
rect 38194 27656 38200 27668
rect 38028 27628 38200 27656
rect 37090 27588 37096 27600
rect 36924 27560 37096 27588
rect 35253 27523 35311 27529
rect 35253 27489 35265 27523
rect 35299 27489 35311 27523
rect 35253 27483 35311 27489
rect 32263 27424 32628 27452
rect 32263 27421 32275 27424
rect 32217 27415 32275 27421
rect 32858 27412 32864 27464
rect 32916 27412 32922 27464
rect 33594 27412 33600 27464
rect 33652 27412 33658 27464
rect 33870 27412 33876 27464
rect 33928 27412 33934 27464
rect 35158 27412 35164 27464
rect 35216 27412 35222 27464
rect 36078 27412 36084 27464
rect 36136 27452 36142 27464
rect 36924 27452 36952 27560
rect 37090 27548 37096 27560
rect 37148 27548 37154 27600
rect 37458 27520 37464 27532
rect 36136 27424 36952 27452
rect 37016 27492 37464 27520
rect 36136 27412 36142 27424
rect 28997 27387 29055 27393
rect 28997 27353 29009 27387
rect 29043 27384 29055 27387
rect 29178 27384 29184 27396
rect 29043 27356 29184 27384
rect 29043 27353 29055 27356
rect 28997 27347 29055 27353
rect 29178 27344 29184 27356
rect 29236 27344 29242 27396
rect 31570 27344 31576 27396
rect 31628 27384 31634 27396
rect 32309 27387 32367 27393
rect 32309 27384 32321 27387
rect 31628 27356 32321 27384
rect 31628 27344 31634 27356
rect 32309 27353 32321 27356
rect 32355 27353 32367 27387
rect 35498 27387 35556 27393
rect 35498 27384 35510 27387
rect 32309 27347 32367 27353
rect 34992 27356 35510 27384
rect 29914 27316 29920 27328
rect 28920 27288 29920 27316
rect 28537 27279 28595 27285
rect 29914 27276 29920 27288
rect 29972 27316 29978 27328
rect 30466 27316 30472 27328
rect 29972 27288 30472 27316
rect 29972 27276 29978 27288
rect 30466 27276 30472 27288
rect 30524 27276 30530 27328
rect 31846 27276 31852 27328
rect 31904 27276 31910 27328
rect 34992 27325 35020 27356
rect 35498 27353 35510 27356
rect 35544 27353 35556 27387
rect 35498 27347 35556 27353
rect 35618 27344 35624 27396
rect 35676 27384 35682 27396
rect 36725 27387 36783 27393
rect 36725 27384 36737 27387
rect 35676 27356 36737 27384
rect 35676 27344 35682 27356
rect 36725 27353 36737 27356
rect 36771 27353 36783 27387
rect 36725 27347 36783 27353
rect 36906 27344 36912 27396
rect 36964 27344 36970 27396
rect 34977 27319 35035 27325
rect 34977 27285 34989 27319
rect 35023 27285 35035 27319
rect 34977 27279 35035 27285
rect 36630 27276 36636 27328
rect 36688 27276 36694 27328
rect 37016 27325 37044 27492
rect 37458 27480 37464 27492
rect 37516 27480 37522 27532
rect 37090 27412 37096 27464
rect 37148 27452 37154 27464
rect 37277 27455 37335 27461
rect 37277 27452 37289 27455
rect 37148 27424 37289 27452
rect 37148 27412 37154 27424
rect 37277 27421 37289 27424
rect 37323 27421 37335 27455
rect 37277 27415 37335 27421
rect 37369 27455 37427 27461
rect 37369 27421 37381 27455
rect 37415 27452 37427 27455
rect 38028 27452 38056 27628
rect 38194 27616 38200 27628
rect 38252 27616 38258 27668
rect 38654 27656 38660 27668
rect 38580 27628 38660 27656
rect 38580 27588 38608 27628
rect 38654 27616 38660 27628
rect 38712 27616 38718 27668
rect 41782 27616 41788 27668
rect 41840 27616 41846 27668
rect 45646 27616 45652 27668
rect 45704 27656 45710 27668
rect 45833 27659 45891 27665
rect 45833 27656 45845 27659
rect 45704 27628 45845 27656
rect 45704 27616 45710 27628
rect 45833 27625 45845 27628
rect 45879 27625 45891 27659
rect 45833 27619 45891 27625
rect 39114 27588 39120 27600
rect 38120 27560 38608 27588
rect 38672 27560 39120 27588
rect 38120 27461 38148 27560
rect 38565 27523 38623 27529
rect 38565 27520 38577 27523
rect 38212 27492 38577 27520
rect 38212 27461 38240 27492
rect 38565 27489 38577 27492
rect 38611 27520 38623 27523
rect 38672 27520 38700 27560
rect 39114 27548 39120 27560
rect 39172 27548 39178 27600
rect 39206 27548 39212 27600
rect 39264 27588 39270 27600
rect 40129 27591 40187 27597
rect 40129 27588 40141 27591
rect 39264 27560 40141 27588
rect 39264 27548 39270 27560
rect 40129 27557 40141 27560
rect 40175 27557 40187 27591
rect 40129 27551 40187 27557
rect 40313 27591 40371 27597
rect 40313 27557 40325 27591
rect 40359 27588 40371 27591
rect 41414 27588 41420 27600
rect 40359 27560 41420 27588
rect 40359 27557 40371 27560
rect 40313 27551 40371 27557
rect 41414 27548 41420 27560
rect 41472 27548 41478 27600
rect 41693 27591 41751 27597
rect 41693 27557 41705 27591
rect 41739 27588 41751 27591
rect 41800 27588 41828 27616
rect 46106 27588 46112 27600
rect 41739 27560 46112 27588
rect 41739 27557 41751 27560
rect 41693 27551 41751 27557
rect 46106 27548 46112 27560
rect 46164 27548 46170 27600
rect 46198 27548 46204 27600
rect 46256 27548 46262 27600
rect 41782 27520 41788 27532
rect 38611 27492 38700 27520
rect 38764 27492 41788 27520
rect 38611 27489 38623 27492
rect 38565 27483 38623 27489
rect 37415 27424 38056 27452
rect 38105 27455 38163 27461
rect 37415 27421 37427 27424
rect 37369 27415 37427 27421
rect 38105 27421 38117 27455
rect 38151 27421 38163 27455
rect 38105 27415 38163 27421
rect 38197 27455 38255 27461
rect 38197 27421 38209 27455
rect 38243 27421 38255 27455
rect 38197 27415 38255 27421
rect 38381 27455 38439 27461
rect 38381 27421 38393 27455
rect 38427 27421 38439 27455
rect 38381 27415 38439 27421
rect 38483 27455 38541 27461
rect 38483 27421 38495 27455
rect 38529 27452 38541 27455
rect 38580 27452 38700 27454
rect 38764 27452 38792 27492
rect 41782 27480 41788 27492
rect 41840 27480 41846 27532
rect 41877 27523 41935 27529
rect 41877 27489 41889 27523
rect 41923 27489 41935 27523
rect 41877 27483 41935 27489
rect 38529 27426 38792 27452
rect 38529 27424 38608 27426
rect 38672 27424 38792 27426
rect 38841 27455 38899 27461
rect 38529 27421 38541 27424
rect 38483 27415 38541 27421
rect 38841 27421 38853 27455
rect 38887 27421 38899 27455
rect 38841 27415 38899 27421
rect 37921 27387 37979 27393
rect 37921 27384 37933 27387
rect 37476 27356 37933 27384
rect 37001 27319 37059 27325
rect 37001 27285 37013 27319
rect 37047 27285 37059 27319
rect 37001 27279 37059 27285
rect 37093 27319 37151 27325
rect 37093 27285 37105 27319
rect 37139 27316 37151 27319
rect 37476 27316 37504 27356
rect 37921 27353 37933 27356
rect 37967 27353 37979 27387
rect 37921 27347 37979 27353
rect 37139 27288 37504 27316
rect 37829 27319 37887 27325
rect 37139 27285 37151 27288
rect 37093 27279 37151 27285
rect 37829 27285 37841 27319
rect 37875 27316 37887 27319
rect 38286 27316 38292 27328
rect 37875 27288 38292 27316
rect 37875 27285 37887 27288
rect 37829 27279 37887 27285
rect 38286 27276 38292 27288
rect 38344 27276 38350 27328
rect 38396 27316 38424 27415
rect 38562 27344 38568 27396
rect 38620 27384 38626 27396
rect 38856 27384 38884 27415
rect 39114 27412 39120 27464
rect 39172 27452 39178 27464
rect 39172 27424 40080 27452
rect 39172 27412 39178 27424
rect 38620 27356 38884 27384
rect 38620 27344 38626 27356
rect 39390 27344 39396 27396
rect 39448 27384 39454 27396
rect 39853 27387 39911 27393
rect 39853 27384 39865 27387
rect 39448 27356 39865 27384
rect 39448 27344 39454 27356
rect 39853 27353 39865 27356
rect 39899 27384 39911 27387
rect 39942 27384 39948 27396
rect 39899 27356 39948 27384
rect 39899 27353 39911 27356
rect 39853 27347 39911 27353
rect 39942 27344 39948 27356
rect 40000 27344 40006 27396
rect 40052 27384 40080 27424
rect 40310 27412 40316 27464
rect 40368 27452 40374 27464
rect 40405 27455 40463 27461
rect 40405 27452 40417 27455
rect 40368 27424 40417 27452
rect 40368 27412 40374 27424
rect 40405 27421 40417 27424
rect 40451 27421 40463 27455
rect 40957 27455 41015 27461
rect 40405 27415 40463 27421
rect 40512 27424 40908 27452
rect 40512 27384 40540 27424
rect 40770 27384 40776 27396
rect 40052 27356 40540 27384
rect 40604 27356 40776 27384
rect 40034 27316 40040 27328
rect 38396 27288 40040 27316
rect 40034 27276 40040 27288
rect 40092 27276 40098 27328
rect 40604 27325 40632 27356
rect 40770 27344 40776 27356
rect 40828 27344 40834 27396
rect 40880 27384 40908 27424
rect 40957 27421 40969 27455
rect 41003 27452 41015 27455
rect 41417 27455 41475 27461
rect 41003 27424 41368 27452
rect 41003 27421 41015 27424
rect 40957 27415 41015 27421
rect 41046 27384 41052 27396
rect 40880 27356 41052 27384
rect 41046 27344 41052 27356
rect 41104 27344 41110 27396
rect 41138 27344 41144 27396
rect 41196 27344 41202 27396
rect 41340 27384 41368 27424
rect 41417 27421 41429 27455
rect 41463 27452 41475 27455
rect 41506 27452 41512 27464
rect 41463 27424 41512 27452
rect 41463 27421 41475 27424
rect 41417 27415 41475 27421
rect 41506 27412 41512 27424
rect 41564 27452 41570 27464
rect 41892 27452 41920 27483
rect 41966 27480 41972 27532
rect 42024 27520 42030 27532
rect 42794 27520 42800 27532
rect 42024 27492 42800 27520
rect 42024 27480 42030 27492
rect 42794 27480 42800 27492
rect 42852 27480 42858 27532
rect 45462 27480 45468 27532
rect 45520 27480 45526 27532
rect 42242 27452 42248 27464
rect 41564 27424 41644 27452
rect 41892 27424 42248 27452
rect 41564 27412 41570 27424
rect 41616 27384 41644 27424
rect 42242 27412 42248 27424
rect 42300 27412 42306 27464
rect 45646 27412 45652 27464
rect 45704 27412 45710 27464
rect 46198 27412 46204 27464
rect 46256 27452 46262 27464
rect 46385 27455 46443 27461
rect 46385 27452 46397 27455
rect 46256 27424 46397 27452
rect 46256 27412 46262 27424
rect 46385 27421 46397 27424
rect 46431 27421 46443 27455
rect 46385 27415 46443 27421
rect 41966 27384 41972 27396
rect 41340 27356 41460 27384
rect 41616 27356 41972 27384
rect 40589 27319 40647 27325
rect 40589 27285 40601 27319
rect 40635 27285 40647 27319
rect 40589 27279 40647 27285
rect 40678 27276 40684 27328
rect 40736 27316 40742 27328
rect 41325 27319 41383 27325
rect 41325 27316 41337 27319
rect 40736 27288 41337 27316
rect 40736 27276 40742 27288
rect 41325 27285 41337 27288
rect 41371 27285 41383 27319
rect 41432 27316 41460 27356
rect 41966 27344 41972 27356
rect 42024 27344 42030 27396
rect 41874 27316 41880 27328
rect 41432 27288 41880 27316
rect 41325 27279 41383 27285
rect 41874 27276 41880 27288
rect 41932 27276 41938 27328
rect 1104 27226 47104 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 47104 27226
rect 1104 27152 47104 27174
rect 2866 27072 2872 27124
rect 2924 27112 2930 27124
rect 4062 27112 4068 27124
rect 2924 27084 4068 27112
rect 2924 27072 2930 27084
rect 4062 27072 4068 27084
rect 4120 27112 4126 27124
rect 4801 27115 4859 27121
rect 4801 27112 4813 27115
rect 4120 27084 4813 27112
rect 4120 27072 4126 27084
rect 4801 27081 4813 27084
rect 4847 27112 4859 27115
rect 4847 27084 11744 27112
rect 4847 27081 4859 27084
rect 4801 27075 4859 27081
rect 8386 27053 8392 27056
rect 8380 27044 8392 27053
rect 6564 27016 8156 27044
rect 8347 27016 8392 27044
rect 1397 26979 1455 26985
rect 1397 26945 1409 26979
rect 1443 26976 1455 26979
rect 2498 26976 2504 26988
rect 1443 26948 2504 26976
rect 1443 26945 1455 26948
rect 1397 26939 1455 26945
rect 2498 26936 2504 26948
rect 2556 26936 2562 26988
rect 4614 26936 4620 26988
rect 4672 26976 4678 26988
rect 6564 26985 6592 27016
rect 6822 26985 6828 26988
rect 4709 26979 4767 26985
rect 4709 26976 4721 26979
rect 4672 26948 4721 26976
rect 4672 26936 4678 26948
rect 4709 26945 4721 26948
rect 4755 26945 4767 26979
rect 4709 26939 4767 26945
rect 6549 26979 6607 26985
rect 6549 26945 6561 26979
rect 6595 26945 6607 26979
rect 6549 26939 6607 26945
rect 6816 26939 6828 26985
rect 6822 26936 6828 26939
rect 6880 26936 6886 26988
rect 8128 26985 8156 27016
rect 8380 27007 8392 27016
rect 8386 27004 8392 27007
rect 8444 27004 8450 27056
rect 9858 27044 9864 27056
rect 8956 27016 9864 27044
rect 8113 26979 8171 26985
rect 8113 26945 8125 26979
rect 8159 26976 8171 26979
rect 8956 26976 8984 27016
rect 9858 27004 9864 27016
rect 9916 27004 9922 27056
rect 10042 27004 10048 27056
rect 10100 27044 10106 27056
rect 11609 27047 11667 27053
rect 11609 27044 11621 27047
rect 10100 27016 11621 27044
rect 10100 27004 10106 27016
rect 11609 27013 11621 27016
rect 11655 27013 11667 27047
rect 11609 27007 11667 27013
rect 8159 26948 8984 26976
rect 8159 26945 8171 26948
rect 8113 26939 8171 26945
rect 9674 26936 9680 26988
rect 9732 26936 9738 26988
rect 9950 26936 9956 26988
rect 10008 26976 10014 26988
rect 10229 26979 10287 26985
rect 10229 26976 10241 26979
rect 10008 26948 10241 26976
rect 10008 26936 10014 26948
rect 10229 26945 10241 26948
rect 10275 26945 10287 26979
rect 10229 26939 10287 26945
rect 10778 26936 10784 26988
rect 10836 26936 10842 26988
rect 4985 26911 5043 26917
rect 4985 26877 4997 26911
rect 5031 26908 5043 26911
rect 5031 26880 6592 26908
rect 5031 26877 5043 26880
rect 4985 26871 5043 26877
rect 2958 26800 2964 26852
rect 3016 26840 3022 26852
rect 5074 26840 5080 26852
rect 3016 26812 5080 26840
rect 3016 26800 3022 26812
rect 5074 26800 5080 26812
rect 5132 26800 5138 26852
rect 934 26732 940 26784
rect 992 26772 998 26784
rect 1581 26775 1639 26781
rect 1581 26772 1593 26775
rect 992 26744 1593 26772
rect 992 26732 998 26744
rect 1581 26741 1593 26744
rect 1627 26741 1639 26775
rect 1581 26735 1639 26741
rect 3970 26732 3976 26784
rect 4028 26772 4034 26784
rect 4341 26775 4399 26781
rect 4341 26772 4353 26775
rect 4028 26744 4353 26772
rect 4028 26732 4034 26744
rect 4341 26741 4353 26744
rect 4387 26741 4399 26775
rect 6564 26772 6592 26880
rect 9122 26868 9128 26920
rect 9180 26908 9186 26920
rect 11624 26908 11652 27007
rect 11716 26976 11744 27084
rect 11790 27072 11796 27124
rect 11848 27072 11854 27124
rect 11974 27072 11980 27124
rect 12032 27072 12038 27124
rect 12894 27072 12900 27124
rect 12952 27072 12958 27124
rect 13446 27072 13452 27124
rect 13504 27112 13510 27124
rect 14550 27112 14556 27124
rect 13504 27084 14556 27112
rect 13504 27072 13510 27084
rect 14550 27072 14556 27084
rect 14608 27072 14614 27124
rect 14734 27072 14740 27124
rect 14792 27112 14798 27124
rect 16758 27112 16764 27124
rect 14792 27084 16764 27112
rect 14792 27072 14798 27084
rect 16758 27072 16764 27084
rect 16816 27072 16822 27124
rect 18414 27112 18420 27124
rect 16868 27084 18420 27112
rect 11885 27047 11943 27053
rect 11885 27013 11897 27047
rect 11931 27044 11943 27047
rect 11931 27016 12480 27044
rect 11931 27013 11943 27016
rect 11885 27007 11943 27013
rect 12250 26976 12256 26988
rect 11716 26948 12256 26976
rect 12250 26936 12256 26948
rect 12308 26936 12314 26988
rect 12452 26976 12480 27016
rect 12526 27004 12532 27056
rect 12584 27004 12590 27056
rect 12710 27004 12716 27056
rect 12768 27004 12774 27056
rect 15197 27047 15255 27053
rect 13372 27016 14044 27044
rect 12621 26979 12679 26985
rect 12621 26976 12633 26979
rect 12452 26948 12633 26976
rect 12621 26945 12633 26948
rect 12667 26976 12679 26979
rect 13372 26976 13400 27016
rect 12667 26948 13400 26976
rect 12667 26945 12679 26948
rect 12621 26939 12679 26945
rect 13446 26936 13452 26988
rect 13504 26936 13510 26988
rect 13630 26936 13636 26988
rect 13688 26936 13694 26988
rect 14016 26985 14044 27016
rect 15197 27013 15209 27047
rect 15243 27044 15255 27047
rect 15378 27044 15384 27056
rect 15243 27016 15384 27044
rect 15243 27013 15255 27016
rect 15197 27007 15255 27013
rect 15378 27004 15384 27016
rect 15436 27004 15442 27056
rect 15657 27047 15715 27053
rect 15657 27013 15669 27047
rect 15703 27044 15715 27047
rect 16574 27044 16580 27056
rect 15703 27016 16580 27044
rect 15703 27013 15715 27016
rect 15657 27007 15715 27013
rect 16574 27004 16580 27016
rect 16632 27004 16638 27056
rect 16868 27053 16896 27084
rect 18414 27072 18420 27084
rect 18472 27072 18478 27124
rect 19058 27072 19064 27124
rect 19116 27072 19122 27124
rect 21266 27072 21272 27124
rect 21324 27112 21330 27124
rect 21821 27115 21879 27121
rect 21821 27112 21833 27115
rect 21324 27084 21833 27112
rect 21324 27072 21330 27084
rect 21821 27081 21833 27084
rect 21867 27081 21879 27115
rect 21821 27075 21879 27081
rect 22066 27084 25820 27112
rect 16853 27047 16911 27053
rect 16853 27013 16865 27047
rect 16899 27013 16911 27047
rect 16853 27007 16911 27013
rect 16942 27004 16948 27056
rect 17000 27044 17006 27056
rect 17313 27047 17371 27053
rect 17313 27044 17325 27047
rect 17000 27016 17325 27044
rect 17000 27004 17006 27016
rect 17313 27013 17325 27016
rect 17359 27013 17371 27047
rect 17313 27007 17371 27013
rect 18230 27004 18236 27056
rect 18288 27004 18294 27056
rect 18782 27004 18788 27056
rect 18840 27004 18846 27056
rect 21085 27047 21143 27053
rect 21085 27013 21097 27047
rect 21131 27044 21143 27047
rect 22066 27044 22094 27084
rect 21131 27016 22094 27044
rect 22281 27047 22339 27053
rect 21131 27013 21143 27016
rect 21085 27007 21143 27013
rect 22281 27013 22293 27047
rect 22327 27044 22339 27047
rect 22462 27044 22468 27056
rect 22327 27016 22468 27044
rect 22327 27013 22339 27016
rect 22281 27007 22339 27013
rect 22462 27004 22468 27016
rect 22520 27004 22526 27056
rect 25314 27004 25320 27056
rect 25372 27004 25378 27056
rect 14001 26979 14059 26985
rect 14001 26945 14013 26979
rect 14047 26976 14059 26979
rect 14458 26976 14464 26988
rect 14047 26948 14464 26976
rect 14047 26945 14059 26948
rect 14001 26939 14059 26945
rect 14458 26936 14464 26948
rect 14516 26976 14522 26988
rect 14734 26976 14740 26988
rect 14516 26948 14740 26976
rect 14516 26936 14522 26948
rect 14734 26936 14740 26948
rect 14792 26936 14798 26988
rect 15289 26979 15347 26985
rect 15289 26945 15301 26979
rect 15335 26945 15347 26979
rect 15289 26939 15347 26945
rect 11790 26908 11796 26920
rect 9180 26880 11100 26908
rect 11624 26880 11796 26908
rect 9180 26868 9186 26880
rect 7926 26800 7932 26852
rect 7984 26800 7990 26852
rect 9493 26843 9551 26849
rect 9493 26809 9505 26843
rect 9539 26840 9551 26843
rect 10962 26840 10968 26852
rect 9539 26812 10968 26840
rect 9539 26809 9551 26812
rect 9493 26803 9551 26809
rect 10962 26800 10968 26812
rect 11020 26800 11026 26852
rect 11072 26840 11100 26880
rect 11790 26868 11796 26880
rect 11848 26908 11854 26920
rect 12342 26908 12348 26920
rect 11848 26880 12348 26908
rect 11848 26868 11854 26880
rect 12342 26868 12348 26880
rect 12400 26868 12406 26920
rect 12894 26868 12900 26920
rect 12952 26908 12958 26920
rect 13725 26911 13783 26917
rect 13725 26908 13737 26911
rect 12952 26880 13737 26908
rect 12952 26868 12958 26880
rect 13725 26877 13737 26880
rect 13771 26908 13783 26911
rect 13814 26908 13820 26920
rect 13771 26880 13820 26908
rect 13771 26877 13783 26880
rect 13725 26871 13783 26877
rect 13814 26868 13820 26880
rect 13872 26868 13878 26920
rect 15194 26868 15200 26920
rect 15252 26908 15258 26920
rect 15304 26908 15332 26939
rect 16390 26936 16396 26988
rect 16448 26976 16454 26988
rect 17218 26976 17224 26988
rect 16448 26948 17224 26976
rect 16448 26936 16454 26948
rect 17218 26936 17224 26948
rect 17276 26936 17282 26988
rect 17402 26936 17408 26988
rect 17460 26936 17466 26988
rect 17865 26979 17923 26985
rect 17865 26945 17877 26979
rect 17911 26945 17923 26979
rect 17865 26939 17923 26945
rect 18417 26979 18475 26985
rect 18417 26945 18429 26979
rect 18463 26976 18475 26979
rect 18598 26976 18604 26988
rect 18463 26948 18604 26976
rect 18463 26945 18475 26948
rect 18417 26939 18475 26945
rect 15252 26880 15332 26908
rect 15749 26911 15807 26917
rect 15252 26868 15258 26880
rect 15749 26877 15761 26911
rect 15795 26908 15807 26911
rect 16758 26908 16764 26920
rect 15795 26880 16764 26908
rect 15795 26877 15807 26880
rect 15749 26871 15807 26877
rect 16758 26868 16764 26880
rect 16816 26868 16822 26920
rect 16942 26868 16948 26920
rect 17000 26908 17006 26920
rect 17880 26908 17908 26939
rect 18598 26936 18604 26948
rect 18656 26976 18662 26988
rect 18969 26979 19027 26985
rect 18969 26976 18981 26979
rect 18656 26948 18981 26976
rect 18656 26936 18662 26948
rect 18969 26945 18981 26948
rect 19015 26976 19027 26979
rect 19521 26979 19579 26985
rect 19521 26976 19533 26979
rect 19015 26948 19533 26976
rect 19015 26945 19027 26948
rect 18969 26939 19027 26945
rect 19521 26945 19533 26948
rect 19567 26976 19579 26979
rect 20257 26979 20315 26985
rect 20257 26976 20269 26979
rect 19567 26948 20269 26976
rect 19567 26945 19579 26948
rect 19521 26939 19579 26945
rect 20257 26945 20269 26948
rect 20303 26945 20315 26979
rect 21269 26979 21327 26985
rect 21269 26976 21281 26979
rect 20257 26939 20315 26945
rect 21100 26948 21281 26976
rect 21100 26920 21128 26948
rect 21269 26945 21281 26948
rect 21315 26976 21327 26979
rect 21358 26976 21364 26988
rect 21315 26948 21364 26976
rect 21315 26945 21327 26948
rect 21269 26939 21327 26945
rect 21358 26936 21364 26948
rect 21416 26936 21422 26988
rect 21450 26936 21456 26988
rect 21508 26936 21514 26988
rect 21545 26979 21603 26985
rect 21545 26945 21557 26979
rect 21591 26976 21603 26979
rect 21726 26976 21732 26988
rect 21591 26948 21732 26976
rect 21591 26945 21603 26948
rect 21545 26939 21603 26945
rect 21726 26936 21732 26948
rect 21784 26936 21790 26988
rect 22186 26936 22192 26988
rect 22244 26976 22250 26988
rect 23109 26979 23167 26985
rect 22244 26948 22600 26976
rect 22244 26936 22250 26948
rect 17000 26880 17908 26908
rect 19981 26911 20039 26917
rect 17000 26868 17006 26880
rect 19981 26877 19993 26911
rect 20027 26908 20039 26911
rect 20990 26908 20996 26920
rect 20027 26880 20996 26908
rect 20027 26877 20039 26880
rect 19981 26871 20039 26877
rect 20990 26868 20996 26880
rect 21048 26868 21054 26920
rect 21082 26868 21088 26920
rect 21140 26868 21146 26920
rect 22370 26868 22376 26920
rect 22428 26868 22434 26920
rect 11072 26812 12204 26840
rect 9766 26772 9772 26784
rect 6564 26744 9772 26772
rect 4341 26735 4399 26741
rect 9766 26732 9772 26744
rect 9824 26772 9830 26784
rect 9861 26775 9919 26781
rect 9861 26772 9873 26775
rect 9824 26744 9873 26772
rect 9824 26732 9830 26744
rect 9861 26741 9873 26744
rect 9907 26741 9919 26775
rect 9861 26735 9919 26741
rect 10042 26732 10048 26784
rect 10100 26732 10106 26784
rect 10597 26775 10655 26781
rect 10597 26741 10609 26775
rect 10643 26772 10655 26775
rect 10778 26772 10784 26784
rect 10643 26744 10784 26772
rect 10643 26741 10655 26744
rect 10597 26735 10655 26741
rect 10778 26732 10784 26744
rect 10836 26732 10842 26784
rect 12176 26781 12204 26812
rect 12250 26800 12256 26852
rect 12308 26840 12314 26852
rect 22462 26840 22468 26852
rect 12308 26812 22468 26840
rect 12308 26800 12314 26812
rect 22462 26800 22468 26812
rect 22520 26800 22526 26852
rect 12161 26775 12219 26781
rect 12161 26741 12173 26775
rect 12207 26741 12219 26775
rect 12161 26735 12219 26741
rect 13449 26775 13507 26781
rect 13449 26741 13461 26775
rect 13495 26772 13507 26775
rect 13630 26772 13636 26784
rect 13495 26744 13636 26772
rect 13495 26741 13507 26744
rect 13449 26735 13507 26741
rect 13630 26732 13636 26744
rect 13688 26732 13694 26784
rect 14274 26732 14280 26784
rect 14332 26772 14338 26784
rect 16022 26772 16028 26784
rect 14332 26744 16028 26772
rect 14332 26732 14338 26744
rect 16022 26732 16028 26744
rect 16080 26732 16086 26784
rect 19613 26775 19671 26781
rect 19613 26741 19625 26775
rect 19659 26772 19671 26775
rect 19702 26772 19708 26784
rect 19659 26744 19708 26772
rect 19659 26741 19671 26744
rect 19613 26735 19671 26741
rect 19702 26732 19708 26744
rect 19760 26732 19766 26784
rect 20806 26732 20812 26784
rect 20864 26772 20870 26784
rect 20990 26772 20996 26784
rect 20864 26744 20996 26772
rect 20864 26732 20870 26744
rect 20990 26732 20996 26744
rect 21048 26732 21054 26784
rect 22572 26772 22600 26948
rect 23109 26945 23121 26979
rect 23155 26976 23167 26979
rect 23290 26976 23296 26988
rect 23155 26948 23296 26976
rect 23155 26945 23167 26948
rect 23109 26939 23167 26945
rect 23290 26936 23296 26948
rect 23348 26936 23354 26988
rect 24026 26985 24032 26988
rect 23983 26979 24032 26985
rect 23983 26945 23995 26979
rect 24029 26945 24032 26979
rect 23983 26939 24032 26945
rect 24026 26936 24032 26939
rect 24084 26936 24090 26988
rect 25038 26936 25044 26988
rect 25096 26976 25102 26988
rect 25332 26976 25360 27004
rect 25792 26985 25820 27084
rect 26602 27072 26608 27124
rect 26660 27112 26666 27124
rect 28353 27115 28411 27121
rect 28353 27112 28365 27115
rect 26660 27084 28365 27112
rect 26660 27072 26666 27084
rect 28353 27081 28365 27084
rect 28399 27112 28411 27115
rect 28399 27084 29040 27112
rect 28399 27081 28411 27084
rect 28353 27075 28411 27081
rect 26510 27004 26516 27056
rect 26568 27044 26574 27056
rect 27218 27047 27276 27053
rect 27218 27044 27230 27047
rect 26568 27016 27230 27044
rect 26568 27004 26574 27016
rect 27218 27013 27230 27016
rect 27264 27013 27276 27047
rect 27218 27007 27276 27013
rect 25409 26979 25467 26985
rect 25409 26976 25421 26979
rect 25096 26948 25421 26976
rect 25096 26936 25102 26948
rect 25409 26945 25421 26948
rect 25455 26945 25467 26979
rect 25409 26939 25467 26945
rect 25501 26979 25559 26985
rect 25501 26945 25513 26979
rect 25547 26945 25559 26979
rect 25501 26939 25559 26945
rect 25777 26979 25835 26985
rect 25777 26945 25789 26979
rect 25823 26945 25835 26979
rect 25777 26939 25835 26945
rect 22922 26868 22928 26920
rect 22980 26868 22986 26920
rect 23842 26868 23848 26920
rect 23900 26868 23906 26920
rect 24118 26868 24124 26920
rect 24176 26868 24182 26920
rect 23566 26800 23572 26852
rect 23624 26800 23630 26852
rect 25516 26840 25544 26939
rect 25958 26936 25964 26988
rect 26016 26936 26022 26988
rect 26329 26979 26387 26985
rect 26329 26945 26341 26979
rect 26375 26976 26387 26979
rect 26878 26976 26884 26988
rect 26375 26948 26884 26976
rect 26375 26945 26387 26948
rect 26329 26939 26387 26945
rect 26878 26936 26884 26948
rect 26936 26936 26942 26988
rect 26973 26979 27031 26985
rect 26973 26945 26985 26979
rect 27019 26976 27031 26979
rect 27614 26976 27620 26988
rect 27019 26948 27620 26976
rect 27019 26945 27031 26948
rect 26973 26939 27031 26945
rect 27614 26936 27620 26948
rect 27672 26936 27678 26988
rect 25590 26868 25596 26920
rect 25648 26908 25654 26920
rect 25685 26911 25743 26917
rect 25685 26908 25697 26911
rect 25648 26880 25697 26908
rect 25648 26868 25654 26880
rect 25685 26877 25697 26880
rect 25731 26877 25743 26911
rect 25685 26871 25743 26877
rect 28905 26911 28963 26917
rect 28905 26877 28917 26911
rect 28951 26877 28963 26911
rect 29012 26908 29040 27084
rect 29270 27072 29276 27124
rect 29328 27112 29334 27124
rect 29730 27112 29736 27124
rect 29328 27084 29736 27112
rect 29328 27072 29334 27084
rect 29730 27072 29736 27084
rect 29788 27112 29794 27124
rect 30190 27112 30196 27124
rect 29788 27084 30196 27112
rect 29788 27072 29794 27084
rect 30190 27072 30196 27084
rect 30248 27072 30254 27124
rect 32858 27072 32864 27124
rect 32916 27112 32922 27124
rect 32916 27084 34744 27112
rect 32916 27072 32922 27084
rect 29086 26936 29092 26988
rect 29144 26936 29150 26988
rect 29822 26936 29828 26988
rect 29880 26936 29886 26988
rect 31846 26936 31852 26988
rect 31904 26976 31910 26988
rect 32309 26979 32367 26985
rect 32309 26976 32321 26979
rect 31904 26948 32321 26976
rect 31904 26936 31910 26948
rect 32309 26945 32321 26948
rect 32355 26945 32367 26979
rect 32309 26939 32367 26945
rect 32674 26936 32680 26988
rect 32732 26976 32738 26988
rect 33244 26985 33272 27084
rect 34716 27044 34744 27084
rect 35158 27072 35164 27124
rect 35216 27112 35222 27124
rect 35253 27115 35311 27121
rect 35253 27112 35265 27115
rect 35216 27084 35265 27112
rect 35216 27072 35222 27084
rect 35253 27081 35265 27084
rect 35299 27081 35311 27115
rect 35253 27075 35311 27081
rect 35621 27115 35679 27121
rect 35621 27081 35633 27115
rect 35667 27112 35679 27115
rect 36630 27112 36636 27124
rect 35667 27084 36636 27112
rect 35667 27081 35679 27084
rect 35621 27075 35679 27081
rect 35636 27044 35664 27075
rect 36630 27072 36636 27084
rect 36688 27072 36694 27124
rect 38105 27115 38163 27121
rect 38105 27081 38117 27115
rect 38151 27112 38163 27115
rect 38378 27112 38384 27124
rect 38151 27084 38384 27112
rect 38151 27081 38163 27084
rect 38105 27075 38163 27081
rect 38378 27072 38384 27084
rect 38436 27072 38442 27124
rect 38746 27072 38752 27124
rect 38804 27072 38810 27124
rect 40129 27115 40187 27121
rect 40129 27112 40141 27115
rect 38856 27084 40141 27112
rect 34716 27016 35664 27044
rect 36096 27016 36492 27044
rect 33045 26979 33103 26985
rect 33045 26976 33057 26979
rect 32732 26948 33057 26976
rect 32732 26936 32738 26948
rect 33045 26945 33057 26948
rect 33091 26945 33103 26979
rect 33045 26939 33103 26945
rect 33229 26979 33287 26985
rect 33229 26945 33241 26979
rect 33275 26945 33287 26979
rect 33229 26939 33287 26945
rect 34054 26936 34060 26988
rect 34112 26985 34118 26988
rect 34112 26979 34140 26985
rect 34128 26945 34140 26979
rect 34112 26939 34140 26945
rect 34112 26936 34118 26939
rect 35434 26936 35440 26988
rect 35492 26976 35498 26988
rect 36096 26985 36124 27016
rect 35713 26979 35771 26985
rect 35713 26976 35725 26979
rect 35492 26948 35725 26976
rect 35492 26936 35498 26948
rect 35713 26945 35725 26948
rect 35759 26945 35771 26979
rect 35713 26939 35771 26945
rect 36081 26979 36139 26985
rect 36081 26945 36093 26979
rect 36127 26945 36139 26979
rect 36081 26939 36139 26945
rect 36354 26936 36360 26988
rect 36412 26936 36418 26988
rect 36464 26976 36492 27016
rect 36906 27004 36912 27056
rect 36964 27044 36970 27056
rect 38856 27044 38884 27084
rect 40129 27081 40141 27084
rect 40175 27081 40187 27115
rect 40129 27075 40187 27081
rect 41138 27072 41144 27124
rect 41196 27112 41202 27124
rect 41325 27115 41383 27121
rect 41325 27112 41337 27115
rect 41196 27084 41337 27112
rect 41196 27072 41202 27084
rect 41325 27081 41337 27084
rect 41371 27081 41383 27115
rect 42058 27112 42064 27124
rect 41325 27075 41383 27081
rect 41524 27084 42064 27112
rect 40678 27044 40684 27056
rect 36964 27016 38884 27044
rect 38948 27016 40684 27044
rect 36964 27004 36970 27016
rect 37366 26976 37372 26988
rect 36464 26948 37372 26976
rect 37366 26936 37372 26948
rect 37424 26976 37430 26988
rect 38102 26976 38108 26988
rect 37424 26948 38108 26976
rect 37424 26936 37430 26948
rect 38102 26936 38108 26948
rect 38160 26936 38166 26988
rect 38286 26936 38292 26988
rect 38344 26936 38350 26988
rect 38948 26985 38976 27016
rect 40678 27004 40684 27016
rect 40736 27004 40742 27056
rect 38933 26979 38991 26985
rect 38933 26945 38945 26979
rect 38979 26945 38991 26979
rect 38933 26939 38991 26945
rect 39390 26936 39396 26988
rect 39448 26936 39454 26988
rect 39577 26979 39635 26985
rect 39577 26945 39589 26979
rect 39623 26976 39635 26979
rect 39758 26976 39764 26988
rect 39623 26948 39764 26976
rect 39623 26945 39635 26948
rect 39577 26939 39635 26945
rect 39758 26936 39764 26948
rect 39816 26936 39822 26988
rect 39942 26936 39948 26988
rect 40000 26976 40006 26988
rect 41524 26985 41552 27084
rect 42058 27072 42064 27084
rect 42116 27072 42122 27124
rect 45646 27072 45652 27124
rect 45704 27112 45710 27124
rect 46385 27115 46443 27121
rect 46385 27112 46397 27115
rect 45704 27084 46397 27112
rect 45704 27072 45710 27084
rect 46385 27081 46397 27084
rect 46431 27081 46443 27115
rect 46385 27075 46443 27081
rect 41782 27004 41788 27056
rect 41840 27044 41846 27056
rect 42426 27044 42432 27056
rect 41840 27016 42432 27044
rect 41840 27004 41846 27016
rect 42426 27004 42432 27016
rect 42484 27004 42490 27056
rect 43346 27044 43352 27056
rect 42904 27016 43352 27044
rect 40221 26979 40279 26985
rect 40221 26976 40233 26979
rect 40000 26948 40233 26976
rect 40000 26936 40006 26948
rect 40221 26945 40233 26948
rect 40267 26945 40279 26979
rect 40221 26939 40279 26945
rect 41509 26979 41567 26985
rect 41509 26945 41521 26979
rect 41555 26945 41567 26979
rect 41509 26939 41567 26945
rect 41693 26979 41751 26985
rect 41693 26945 41705 26979
rect 41739 26976 41751 26979
rect 41877 26979 41935 26985
rect 41877 26976 41889 26979
rect 41739 26948 41889 26976
rect 41739 26945 41751 26948
rect 41693 26939 41751 26945
rect 41877 26945 41889 26948
rect 41923 26976 41935 26979
rect 42242 26976 42248 26988
rect 41923 26948 42248 26976
rect 41923 26945 41935 26948
rect 41877 26939 41935 26945
rect 42242 26936 42248 26948
rect 42300 26936 42306 26988
rect 42610 26936 42616 26988
rect 42668 26936 42674 26988
rect 42904 26985 42932 27016
rect 43346 27004 43352 27016
rect 43404 27004 43410 27056
rect 42889 26979 42947 26985
rect 42889 26945 42901 26979
rect 42935 26945 42947 26979
rect 42889 26939 42947 26945
rect 43073 26979 43131 26985
rect 43073 26945 43085 26979
rect 43119 26945 43131 26979
rect 43073 26939 43131 26945
rect 29638 26908 29644 26920
rect 29012 26880 29644 26908
rect 28905 26871 28963 26877
rect 28920 26840 28948 26871
rect 29638 26868 29644 26880
rect 29696 26908 29702 26920
rect 29942 26911 30000 26917
rect 29942 26908 29954 26911
rect 29696 26880 29954 26908
rect 29696 26868 29702 26880
rect 29942 26877 29954 26880
rect 29988 26877 30000 26911
rect 29942 26871 30000 26877
rect 30111 26911 30169 26917
rect 30111 26877 30123 26911
rect 30157 26908 30169 26911
rect 30834 26908 30840 26920
rect 30157 26880 30840 26908
rect 30157 26877 30169 26880
rect 30111 26871 30169 26877
rect 30834 26868 30840 26880
rect 30892 26868 30898 26920
rect 33594 26868 33600 26920
rect 33652 26908 33658 26920
rect 33965 26911 34023 26917
rect 33965 26908 33977 26911
rect 33652 26880 33977 26908
rect 33652 26868 33658 26880
rect 33965 26877 33977 26880
rect 34011 26877 34023 26911
rect 33965 26871 34023 26877
rect 34238 26868 34244 26920
rect 34296 26868 34302 26920
rect 35342 26868 35348 26920
rect 35400 26908 35406 26920
rect 35805 26911 35863 26917
rect 35805 26908 35817 26911
rect 35400 26880 35817 26908
rect 35400 26868 35406 26880
rect 35805 26877 35817 26880
rect 35851 26877 35863 26911
rect 35805 26871 35863 26877
rect 38562 26868 38568 26920
rect 38620 26908 38626 26920
rect 39853 26911 39911 26917
rect 39853 26908 39865 26911
rect 38620 26880 39865 26908
rect 38620 26868 38626 26880
rect 39853 26877 39865 26880
rect 39899 26877 39911 26911
rect 39853 26871 39911 26877
rect 41598 26868 41604 26920
rect 41656 26908 41662 26920
rect 41785 26911 41843 26917
rect 41785 26908 41797 26911
rect 41656 26880 41797 26908
rect 41656 26868 41662 26880
rect 41785 26877 41797 26880
rect 41831 26908 41843 26911
rect 42153 26911 42211 26917
rect 42153 26908 42165 26911
rect 41831 26880 42165 26908
rect 41831 26877 41843 26880
rect 41785 26871 41843 26877
rect 42153 26877 42165 26880
rect 42199 26908 42211 26911
rect 42426 26908 42432 26920
rect 42199 26880 42432 26908
rect 42199 26877 42211 26880
rect 42153 26871 42211 26877
rect 42426 26868 42432 26880
rect 42484 26868 42490 26920
rect 42978 26868 42984 26920
rect 43036 26908 43042 26920
rect 43088 26908 43116 26939
rect 43254 26936 43260 26988
rect 43312 26936 43318 26988
rect 45554 26936 45560 26988
rect 45612 26936 45618 26988
rect 45649 26979 45707 26985
rect 45649 26945 45661 26979
rect 45695 26976 45707 26979
rect 45738 26976 45744 26988
rect 45695 26948 45744 26976
rect 45695 26945 45707 26948
rect 45649 26939 45707 26945
rect 45738 26936 45744 26948
rect 45796 26936 45802 26988
rect 46569 26979 46627 26985
rect 46569 26945 46581 26979
rect 46615 26976 46627 26979
rect 46750 26976 46756 26988
rect 46615 26948 46756 26976
rect 46615 26945 46627 26948
rect 46569 26939 46627 26945
rect 46750 26936 46756 26948
rect 46808 26936 46814 26988
rect 43036 26880 43116 26908
rect 45833 26911 45891 26917
rect 43036 26868 43042 26880
rect 45833 26877 45845 26911
rect 45879 26877 45891 26911
rect 45833 26871 45891 26877
rect 29454 26840 29460 26852
rect 25516 26812 26188 26840
rect 28920 26812 29460 26840
rect 24026 26772 24032 26784
rect 22572 26744 24032 26772
rect 24026 26732 24032 26744
rect 24084 26772 24090 26784
rect 24302 26772 24308 26784
rect 24084 26744 24308 26772
rect 24084 26732 24090 26744
rect 24302 26732 24308 26744
rect 24360 26732 24366 26784
rect 24762 26732 24768 26784
rect 24820 26732 24826 26784
rect 25222 26732 25228 26784
rect 25280 26732 25286 26784
rect 26160 26772 26188 26812
rect 29454 26800 29460 26812
rect 29512 26800 29518 26852
rect 29549 26843 29607 26849
rect 29549 26809 29561 26843
rect 29595 26809 29607 26843
rect 29549 26803 29607 26809
rect 28994 26772 29000 26784
rect 26160 26744 29000 26772
rect 28994 26732 29000 26744
rect 29052 26732 29058 26784
rect 29564 26772 29592 26803
rect 33686 26800 33692 26852
rect 33744 26800 33750 26852
rect 39577 26843 39635 26849
rect 39577 26809 39589 26843
rect 39623 26840 39635 26843
rect 40310 26840 40316 26852
rect 39623 26812 40316 26840
rect 39623 26809 39635 26812
rect 39577 26803 39635 26809
rect 40310 26800 40316 26812
rect 40368 26800 40374 26852
rect 41874 26800 41880 26852
rect 41932 26800 41938 26852
rect 41969 26843 42027 26849
rect 41969 26809 41981 26843
rect 42015 26840 42027 26843
rect 42058 26840 42064 26852
rect 42015 26812 42064 26840
rect 42015 26809 42027 26812
rect 41969 26803 42027 26809
rect 42058 26800 42064 26812
rect 42116 26840 42122 26852
rect 43349 26843 43407 26849
rect 43349 26840 43361 26843
rect 42116 26812 43361 26840
rect 42116 26800 42122 26812
rect 43349 26809 43361 26812
rect 43395 26809 43407 26843
rect 43349 26803 43407 26809
rect 45373 26843 45431 26849
rect 45373 26809 45385 26843
rect 45419 26840 45431 26843
rect 45848 26840 45876 26871
rect 45419 26812 45876 26840
rect 45419 26809 45431 26812
rect 45373 26803 45431 26809
rect 46014 26800 46020 26852
rect 46072 26800 46078 26852
rect 30282 26772 30288 26784
rect 29564 26744 30288 26772
rect 30282 26732 30288 26744
rect 30340 26732 30346 26784
rect 30558 26732 30564 26784
rect 30616 26772 30622 26784
rect 30745 26775 30803 26781
rect 30745 26772 30757 26775
rect 30616 26744 30757 26772
rect 30616 26732 30622 26744
rect 30745 26741 30757 26744
rect 30791 26741 30803 26775
rect 30745 26735 30803 26741
rect 32030 26732 32036 26784
rect 32088 26772 32094 26784
rect 32125 26775 32183 26781
rect 32125 26772 32137 26775
rect 32088 26744 32137 26772
rect 32088 26732 32094 26744
rect 32125 26741 32137 26744
rect 32171 26741 32183 26775
rect 32125 26735 32183 26741
rect 33318 26732 33324 26784
rect 33376 26772 33382 26784
rect 34885 26775 34943 26781
rect 34885 26772 34897 26775
rect 33376 26744 34897 26772
rect 33376 26732 33382 26744
rect 34885 26741 34897 26744
rect 34931 26741 34943 26775
rect 34885 26735 34943 26741
rect 37090 26732 37096 26784
rect 37148 26732 37154 26784
rect 38746 26732 38752 26784
rect 38804 26772 38810 26784
rect 39114 26772 39120 26784
rect 38804 26744 39120 26772
rect 38804 26732 38810 26744
rect 39114 26732 39120 26744
rect 39172 26732 39178 26784
rect 39945 26775 40003 26781
rect 39945 26741 39957 26775
rect 39991 26772 40003 26775
rect 40405 26775 40463 26781
rect 40405 26772 40417 26775
rect 39991 26744 40417 26772
rect 39991 26741 40003 26744
rect 39945 26735 40003 26741
rect 40405 26741 40417 26744
rect 40451 26772 40463 26775
rect 41230 26772 41236 26784
rect 40451 26744 41236 26772
rect 40451 26741 40463 26744
rect 40405 26735 40463 26741
rect 41230 26732 41236 26744
rect 41288 26772 41294 26784
rect 44634 26772 44640 26784
rect 41288 26744 44640 26772
rect 41288 26732 41294 26744
rect 44634 26732 44640 26744
rect 44692 26732 44698 26784
rect 1104 26682 47104 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 47104 26682
rect 1104 26608 47104 26630
rect 2774 26528 2780 26580
rect 2832 26568 2838 26580
rect 2961 26571 3019 26577
rect 2961 26568 2973 26571
rect 2832 26540 2973 26568
rect 2832 26528 2838 26540
rect 2961 26537 2973 26540
rect 3007 26568 3019 26571
rect 4522 26568 4528 26580
rect 3007 26540 4528 26568
rect 3007 26537 3019 26540
rect 2961 26531 3019 26537
rect 4522 26528 4528 26540
rect 4580 26568 4586 26580
rect 4580 26540 4844 26568
rect 4580 26528 4586 26540
rect 4062 26392 4068 26444
rect 4120 26392 4126 26444
rect 4614 26432 4620 26444
rect 4264 26404 4620 26432
rect 4264 26376 4292 26404
rect 4614 26392 4620 26404
rect 4672 26392 4678 26444
rect 4706 26392 4712 26444
rect 4764 26392 4770 26444
rect 4816 26432 4844 26540
rect 5626 26528 5632 26580
rect 5684 26568 5690 26580
rect 6086 26568 6092 26580
rect 5684 26540 6092 26568
rect 5684 26528 5690 26540
rect 6086 26528 6092 26540
rect 6144 26528 6150 26580
rect 6270 26528 6276 26580
rect 6328 26568 6334 26580
rect 6365 26571 6423 26577
rect 6365 26568 6377 26571
rect 6328 26540 6377 26568
rect 6328 26528 6334 26540
rect 6365 26537 6377 26540
rect 6411 26537 6423 26571
rect 6365 26531 6423 26537
rect 6822 26528 6828 26580
rect 6880 26568 6886 26580
rect 7009 26571 7067 26577
rect 7009 26568 7021 26571
rect 6880 26540 7021 26568
rect 6880 26528 6886 26540
rect 7009 26537 7021 26540
rect 7055 26537 7067 26571
rect 9858 26568 9864 26580
rect 7009 26531 7067 26537
rect 9232 26540 9864 26568
rect 5718 26460 5724 26512
rect 5776 26460 5782 26512
rect 7745 26503 7803 26509
rect 7745 26469 7757 26503
rect 7791 26500 7803 26503
rect 8570 26500 8576 26512
rect 7791 26472 8576 26500
rect 7791 26469 7803 26472
rect 7745 26463 7803 26469
rect 8570 26460 8576 26472
rect 8628 26460 8634 26512
rect 4985 26435 5043 26441
rect 4985 26432 4997 26435
rect 4816 26404 4997 26432
rect 4985 26401 4997 26404
rect 5031 26401 5043 26435
rect 4985 26395 5043 26401
rect 5074 26392 5080 26444
rect 5132 26441 5138 26444
rect 5132 26435 5160 26441
rect 5148 26401 5160 26435
rect 5132 26395 5160 26401
rect 5261 26435 5319 26441
rect 5261 26401 5273 26435
rect 5307 26432 5319 26435
rect 5736 26432 5764 26460
rect 5307 26404 7328 26432
rect 5307 26401 5319 26404
rect 5261 26395 5319 26401
rect 5132 26392 5138 26395
rect 1581 26367 1639 26373
rect 1581 26333 1593 26367
rect 1627 26364 1639 26367
rect 1670 26364 1676 26376
rect 1627 26336 1676 26364
rect 1627 26333 1639 26336
rect 1581 26327 1639 26333
rect 1670 26324 1676 26336
rect 1728 26324 1734 26376
rect 3970 26324 3976 26376
rect 4028 26324 4034 26376
rect 4246 26324 4252 26376
rect 4304 26324 4310 26376
rect 6178 26324 6184 26376
rect 6236 26324 6242 26376
rect 7190 26324 7196 26376
rect 7248 26324 7254 26376
rect 1848 26299 1906 26305
rect 1848 26265 1860 26299
rect 1894 26296 1906 26299
rect 2038 26296 2044 26308
rect 1894 26268 2044 26296
rect 1894 26265 1906 26268
rect 1848 26259 1906 26265
rect 2038 26256 2044 26268
rect 2096 26256 2102 26308
rect 5905 26299 5963 26305
rect 5905 26265 5917 26299
rect 5951 26296 5963 26299
rect 6822 26296 6828 26308
rect 5951 26268 6828 26296
rect 5951 26265 5963 26268
rect 5905 26259 5963 26265
rect 6822 26256 6828 26268
rect 6880 26256 6886 26308
rect 7300 26296 7328 26404
rect 7926 26392 7932 26444
rect 7984 26432 7990 26444
rect 9232 26441 9260 26540
rect 9858 26528 9864 26540
rect 9916 26568 9922 26580
rect 12069 26571 12127 26577
rect 9916 26540 10272 26568
rect 9916 26528 9922 26540
rect 8205 26435 8263 26441
rect 8205 26432 8217 26435
rect 7984 26404 8217 26432
rect 7984 26392 7990 26404
rect 8205 26401 8217 26404
rect 8251 26401 8263 26435
rect 8205 26395 8263 26401
rect 8297 26435 8355 26441
rect 8297 26401 8309 26435
rect 8343 26401 8355 26435
rect 8297 26395 8355 26401
rect 9217 26435 9275 26441
rect 9217 26401 9229 26435
rect 9263 26401 9275 26435
rect 10244 26432 10272 26540
rect 12069 26537 12081 26571
rect 12115 26568 12127 26571
rect 12345 26571 12403 26577
rect 12345 26568 12357 26571
rect 12115 26540 12357 26568
rect 12115 26537 12127 26540
rect 12069 26531 12127 26537
rect 12345 26537 12357 26540
rect 12391 26568 12403 26571
rect 12986 26568 12992 26580
rect 12391 26540 12992 26568
rect 12391 26537 12403 26540
rect 12345 26531 12403 26537
rect 12986 26528 12992 26540
rect 13044 26528 13050 26580
rect 14277 26571 14335 26577
rect 13096 26540 14228 26568
rect 12529 26503 12587 26509
rect 12529 26469 12541 26503
rect 12575 26469 12587 26503
rect 12529 26463 12587 26469
rect 10689 26435 10747 26441
rect 10689 26432 10701 26435
rect 10244 26404 10701 26432
rect 9217 26395 9275 26401
rect 10689 26401 10701 26404
rect 10735 26401 10747 26435
rect 10689 26395 10747 26401
rect 8018 26324 8024 26376
rect 8076 26364 8082 26376
rect 8312 26364 8340 26395
rect 12342 26392 12348 26444
rect 12400 26432 12406 26444
rect 12400 26404 12480 26432
rect 12400 26392 12406 26404
rect 8076 26336 8340 26364
rect 9484 26367 9542 26373
rect 8076 26324 8082 26336
rect 9484 26333 9496 26367
rect 9530 26364 9542 26367
rect 10042 26364 10048 26376
rect 9530 26336 10048 26364
rect 9530 26333 9542 26336
rect 9484 26327 9542 26333
rect 10042 26324 10048 26336
rect 10100 26324 10106 26376
rect 10778 26324 10784 26376
rect 10836 26364 10842 26376
rect 10945 26367 11003 26373
rect 10945 26364 10957 26367
rect 10836 26336 10957 26364
rect 10836 26324 10842 26336
rect 10945 26333 10957 26336
rect 10991 26333 11003 26367
rect 10945 26327 11003 26333
rect 8113 26299 8171 26305
rect 7300 26268 8064 26296
rect 3789 26231 3847 26237
rect 3789 26197 3801 26231
rect 3835 26228 3847 26231
rect 3878 26228 3884 26240
rect 3835 26200 3884 26228
rect 3835 26197 3847 26200
rect 3789 26191 3847 26197
rect 3878 26188 3884 26200
rect 3936 26188 3942 26240
rect 4614 26188 4620 26240
rect 4672 26228 4678 26240
rect 4982 26228 4988 26240
rect 4672 26200 4988 26228
rect 4672 26188 4678 26200
rect 4982 26188 4988 26200
rect 5040 26188 5046 26240
rect 8036 26228 8064 26268
rect 8113 26265 8125 26299
rect 8159 26296 8171 26299
rect 8294 26296 8300 26308
rect 8159 26268 8300 26296
rect 8159 26265 8171 26268
rect 8113 26259 8171 26265
rect 8294 26256 8300 26268
rect 8352 26256 8358 26308
rect 10410 26296 10416 26308
rect 8404 26268 10416 26296
rect 8404 26228 8432 26268
rect 10410 26256 10416 26268
rect 10468 26256 10474 26308
rect 12161 26299 12219 26305
rect 12161 26265 12173 26299
rect 12207 26265 12219 26299
rect 12452 26296 12480 26404
rect 12544 26376 12572 26463
rect 12526 26324 12532 26376
rect 12584 26324 12590 26376
rect 12621 26367 12679 26373
rect 12621 26333 12633 26367
rect 12667 26364 12679 26367
rect 12710 26364 12716 26376
rect 12667 26336 12716 26364
rect 12667 26333 12679 26336
rect 12621 26327 12679 26333
rect 12710 26324 12716 26336
rect 12768 26324 12774 26376
rect 13096 26364 13124 26540
rect 13173 26503 13231 26509
rect 13173 26469 13185 26503
rect 13219 26469 13231 26503
rect 13173 26463 13231 26469
rect 13188 26432 13216 26463
rect 13814 26460 13820 26512
rect 13872 26460 13878 26512
rect 14200 26500 14228 26540
rect 14277 26537 14289 26571
rect 14323 26568 14335 26571
rect 14550 26568 14556 26580
rect 14323 26540 14556 26568
rect 14323 26537 14335 26540
rect 14277 26531 14335 26537
rect 14550 26528 14556 26540
rect 14608 26528 14614 26580
rect 15102 26528 15108 26580
rect 15160 26568 15166 26580
rect 18693 26571 18751 26577
rect 18693 26568 18705 26571
rect 15160 26540 18705 26568
rect 15160 26528 15166 26540
rect 18693 26537 18705 26540
rect 18739 26537 18751 26571
rect 18693 26531 18751 26537
rect 25222 26528 25228 26580
rect 25280 26568 25286 26580
rect 33137 26571 33195 26577
rect 25280 26540 33088 26568
rect 25280 26528 25286 26540
rect 15194 26500 15200 26512
rect 14200 26472 15200 26500
rect 15194 26460 15200 26472
rect 15252 26460 15258 26512
rect 15289 26503 15347 26509
rect 15289 26469 15301 26503
rect 15335 26500 15347 26503
rect 15470 26500 15476 26512
rect 15335 26472 15476 26500
rect 15335 26469 15347 26472
rect 15289 26463 15347 26469
rect 15470 26460 15476 26472
rect 15528 26500 15534 26512
rect 15528 26472 16620 26500
rect 15528 26460 15534 26472
rect 15228 26432 15256 26460
rect 15381 26435 15439 26441
rect 15381 26432 15393 26435
rect 13188 26404 14320 26432
rect 15228 26404 15393 26432
rect 13265 26367 13323 26373
rect 13265 26364 13277 26367
rect 12820 26336 13277 26364
rect 12820 26296 12848 26336
rect 13265 26333 13277 26336
rect 13311 26333 13323 26367
rect 13265 26327 13323 26333
rect 13538 26324 13544 26376
rect 13596 26364 13602 26376
rect 13596 26336 14136 26364
rect 13596 26324 13602 26336
rect 12452 26268 12848 26296
rect 12161 26259 12219 26265
rect 8036 26200 8432 26228
rect 10594 26188 10600 26240
rect 10652 26228 10658 26240
rect 12176 26228 12204 26259
rect 12894 26256 12900 26308
rect 12952 26296 12958 26308
rect 12989 26299 13047 26305
rect 12989 26296 13001 26299
rect 12952 26268 13001 26296
rect 12952 26256 12958 26268
rect 12989 26265 13001 26268
rect 13035 26265 13047 26299
rect 12989 26259 13047 26265
rect 13630 26256 13636 26308
rect 13688 26296 13694 26308
rect 14108 26305 14136 26336
rect 14292 26305 14320 26404
rect 15381 26401 15393 26404
rect 15427 26401 15439 26435
rect 15381 26395 15439 26401
rect 15746 26392 15752 26444
rect 15804 26432 15810 26444
rect 16114 26432 16120 26444
rect 15804 26404 16120 26432
rect 15804 26392 15810 26404
rect 16114 26392 16120 26404
rect 16172 26392 16178 26444
rect 16592 26441 16620 26472
rect 17034 26460 17040 26512
rect 17092 26460 17098 26512
rect 20346 26460 20352 26512
rect 20404 26460 20410 26512
rect 20806 26460 20812 26512
rect 20864 26460 20870 26512
rect 21177 26503 21235 26509
rect 21177 26469 21189 26503
rect 21223 26500 21235 26503
rect 23753 26503 23811 26509
rect 21223 26472 23428 26500
rect 21223 26469 21235 26472
rect 21177 26463 21235 26469
rect 16577 26435 16635 26441
rect 16577 26401 16589 26435
rect 16623 26432 16635 26435
rect 16758 26432 16764 26444
rect 16623 26404 16764 26432
rect 16623 26401 16635 26404
rect 16577 26395 16635 26401
rect 16758 26392 16764 26404
rect 16816 26392 16822 26444
rect 17052 26432 17080 26460
rect 17402 26432 17408 26444
rect 17052 26404 17408 26432
rect 14553 26367 14611 26373
rect 14553 26333 14565 26367
rect 14599 26364 14611 26367
rect 14642 26364 14648 26376
rect 14599 26336 14648 26364
rect 14599 26333 14611 26336
rect 14553 26327 14611 26333
rect 14642 26324 14648 26336
rect 14700 26324 14706 26376
rect 14734 26324 14740 26376
rect 14792 26364 14798 26376
rect 14829 26367 14887 26373
rect 14829 26364 14841 26367
rect 14792 26336 14841 26364
rect 14792 26324 14798 26336
rect 14829 26333 14841 26336
rect 14875 26333 14887 26367
rect 14829 26327 14887 26333
rect 14921 26367 14979 26373
rect 14921 26333 14933 26367
rect 14967 26364 14979 26367
rect 16206 26364 16212 26376
rect 14967 26336 16212 26364
rect 14967 26333 14979 26336
rect 14921 26327 14979 26333
rect 14093 26299 14151 26305
rect 13688 26268 14044 26296
rect 13688 26256 13694 26268
rect 12250 26228 12256 26240
rect 10652 26200 12256 26228
rect 10652 26188 10658 26200
rect 12250 26188 12256 26200
rect 12308 26188 12314 26240
rect 12371 26231 12429 26237
rect 12371 26197 12383 26231
rect 12417 26228 12429 26231
rect 12912 26228 12940 26256
rect 12417 26200 12940 26228
rect 12417 26197 12429 26200
rect 12371 26191 12429 26197
rect 13262 26188 13268 26240
rect 13320 26228 13326 26240
rect 13449 26231 13507 26237
rect 13449 26228 13461 26231
rect 13320 26200 13461 26228
rect 13320 26188 13326 26200
rect 13449 26197 13461 26200
rect 13495 26197 13507 26231
rect 13449 26191 13507 26197
rect 13541 26231 13599 26237
rect 13541 26197 13553 26231
rect 13587 26228 13599 26231
rect 13906 26228 13912 26240
rect 13587 26200 13912 26228
rect 13587 26197 13599 26200
rect 13541 26191 13599 26197
rect 13906 26188 13912 26200
rect 13964 26188 13970 26240
rect 14016 26228 14044 26268
rect 14093 26265 14105 26299
rect 14139 26265 14151 26299
rect 14093 26259 14151 26265
rect 14277 26299 14335 26305
rect 14277 26265 14289 26299
rect 14323 26265 14335 26299
rect 14277 26259 14335 26265
rect 14936 26228 14964 26327
rect 16206 26324 16212 26336
rect 16264 26324 16270 26376
rect 17034 26324 17040 26376
rect 17092 26324 17098 26376
rect 17236 26373 17264 26404
rect 17402 26392 17408 26404
rect 17460 26392 17466 26444
rect 20530 26392 20536 26444
rect 20588 26432 20594 26444
rect 20588 26404 22094 26432
rect 20588 26392 20594 26404
rect 17221 26367 17279 26373
rect 17221 26333 17233 26367
rect 17267 26364 17279 26367
rect 17773 26367 17831 26373
rect 17773 26364 17785 26367
rect 17267 26336 17785 26364
rect 17267 26333 17279 26336
rect 17221 26327 17279 26333
rect 17773 26333 17785 26336
rect 17819 26333 17831 26367
rect 17773 26327 17831 26333
rect 18598 26324 18604 26376
rect 18656 26364 18662 26376
rect 19521 26367 19579 26373
rect 19521 26364 19533 26367
rect 18656 26336 19533 26364
rect 18656 26324 18662 26336
rect 19521 26333 19533 26336
rect 19567 26364 19579 26367
rect 20165 26367 20223 26373
rect 20165 26364 20177 26367
rect 19567 26336 20177 26364
rect 19567 26333 19579 26336
rect 19521 26327 19579 26333
rect 20165 26333 20177 26336
rect 20211 26333 20223 26367
rect 20165 26327 20223 26333
rect 20622 26324 20628 26376
rect 20680 26324 20686 26376
rect 20993 26367 21051 26373
rect 20993 26333 21005 26367
rect 21039 26364 21051 26367
rect 21174 26364 21180 26376
rect 21039 26336 21180 26364
rect 21039 26333 21051 26336
rect 20993 26327 21051 26333
rect 21174 26324 21180 26336
rect 21232 26324 21238 26376
rect 16022 26256 16028 26308
rect 16080 26296 16086 26308
rect 16669 26299 16727 26305
rect 16080 26268 16620 26296
rect 16080 26256 16086 26268
rect 14016 26200 14964 26228
rect 16592 26228 16620 26268
rect 16669 26265 16681 26299
rect 16715 26296 16727 26299
rect 16850 26296 16856 26308
rect 16715 26268 16856 26296
rect 16715 26265 16727 26268
rect 16669 26259 16727 26265
rect 16850 26256 16856 26268
rect 16908 26256 16914 26308
rect 17129 26299 17187 26305
rect 17129 26296 17141 26299
rect 16960 26268 17141 26296
rect 16960 26228 16988 26268
rect 17129 26265 17141 26268
rect 17175 26265 17187 26299
rect 17129 26259 17187 26265
rect 17586 26256 17592 26308
rect 17644 26256 17650 26308
rect 19610 26256 19616 26308
rect 19668 26296 19674 26308
rect 19889 26299 19947 26305
rect 19889 26296 19901 26299
rect 19668 26268 19901 26296
rect 19668 26256 19674 26268
rect 19889 26265 19901 26268
rect 19935 26296 19947 26299
rect 19978 26296 19984 26308
rect 19935 26268 19984 26296
rect 19935 26265 19947 26268
rect 19889 26259 19947 26265
rect 19978 26256 19984 26268
rect 20036 26256 20042 26308
rect 22066 26296 22094 26404
rect 23400 26364 23428 26472
rect 23753 26469 23765 26503
rect 23799 26500 23811 26503
rect 24762 26500 24768 26512
rect 23799 26472 24768 26500
rect 23799 26469 23811 26472
rect 23753 26463 23811 26469
rect 24762 26460 24768 26472
rect 24820 26460 24826 26512
rect 26326 26460 26332 26512
rect 26384 26500 26390 26512
rect 26421 26503 26479 26509
rect 26421 26500 26433 26503
rect 26384 26472 26433 26500
rect 26384 26460 26390 26472
rect 26421 26469 26433 26472
rect 26467 26469 26479 26503
rect 26421 26463 26479 26469
rect 30193 26503 30251 26509
rect 30193 26469 30205 26503
rect 30239 26469 30251 26503
rect 33060 26500 33088 26540
rect 33137 26537 33149 26571
rect 33183 26568 33195 26571
rect 34054 26568 34060 26580
rect 33183 26540 34060 26568
rect 33183 26537 33195 26540
rect 33137 26531 33195 26537
rect 34054 26528 34060 26540
rect 34112 26528 34118 26580
rect 35342 26528 35348 26580
rect 35400 26568 35406 26580
rect 35621 26571 35679 26577
rect 35621 26568 35633 26571
rect 35400 26540 35633 26568
rect 35400 26528 35406 26540
rect 35621 26537 35633 26540
rect 35667 26537 35679 26571
rect 35621 26531 35679 26537
rect 37642 26528 37648 26580
rect 37700 26568 37706 26580
rect 38289 26571 38347 26577
rect 38289 26568 38301 26571
rect 37700 26540 38301 26568
rect 37700 26528 37706 26540
rect 38289 26537 38301 26540
rect 38335 26568 38347 26571
rect 38841 26571 38899 26577
rect 38841 26568 38853 26571
rect 38335 26540 38853 26568
rect 38335 26537 38347 26540
rect 38289 26531 38347 26537
rect 38841 26537 38853 26540
rect 38887 26537 38899 26571
rect 38841 26531 38899 26537
rect 42610 26528 42616 26580
rect 42668 26568 42674 26580
rect 43162 26568 43168 26580
rect 42668 26540 43168 26568
rect 42668 26528 42674 26540
rect 43162 26528 43168 26540
rect 43220 26528 43226 26580
rect 46014 26528 46020 26580
rect 46072 26528 46078 26580
rect 46198 26528 46204 26580
rect 46256 26528 46262 26580
rect 46385 26571 46443 26577
rect 46385 26537 46397 26571
rect 46431 26537 46443 26571
rect 46385 26531 46443 26537
rect 36354 26500 36360 26512
rect 33060 26472 36360 26500
rect 30193 26463 30251 26469
rect 23474 26392 23480 26444
rect 23532 26432 23538 26444
rect 30208 26432 30236 26463
rect 36354 26460 36360 26472
rect 36412 26460 36418 26512
rect 38378 26460 38384 26512
rect 38436 26500 38442 26512
rect 40954 26500 40960 26512
rect 38436 26472 40960 26500
rect 38436 26460 38442 26472
rect 40954 26460 40960 26472
rect 41012 26460 41018 26512
rect 42153 26503 42211 26509
rect 42153 26469 42165 26503
rect 42199 26500 42211 26503
rect 42794 26500 42800 26512
rect 42199 26472 42800 26500
rect 42199 26469 42211 26472
rect 42153 26463 42211 26469
rect 42794 26460 42800 26472
rect 42852 26460 42858 26512
rect 46032 26500 46060 26528
rect 46400 26500 46428 26531
rect 46750 26528 46756 26580
rect 46808 26528 46814 26580
rect 46032 26472 46428 26500
rect 23532 26404 30236 26432
rect 30837 26435 30895 26441
rect 23532 26392 23538 26404
rect 30837 26401 30849 26435
rect 30883 26432 30895 26435
rect 31570 26432 31576 26444
rect 30883 26404 31576 26432
rect 30883 26401 30895 26404
rect 30837 26395 30895 26401
rect 31570 26392 31576 26404
rect 31628 26392 31634 26444
rect 38562 26392 38568 26444
rect 38620 26432 38626 26444
rect 42610 26432 42616 26444
rect 38620 26404 42616 26432
rect 38620 26392 38626 26404
rect 23400 26336 23888 26364
rect 22922 26296 22928 26308
rect 22066 26268 22928 26296
rect 22922 26256 22928 26268
rect 22980 26296 22986 26308
rect 23385 26299 23443 26305
rect 23385 26296 23397 26299
rect 22980 26268 23397 26296
rect 22980 26256 22986 26268
rect 23385 26265 23397 26268
rect 23431 26265 23443 26299
rect 23860 26296 23888 26336
rect 23934 26324 23940 26376
rect 23992 26364 23998 26376
rect 26050 26364 26056 26376
rect 23992 26336 26056 26364
rect 23992 26324 23998 26336
rect 26050 26324 26056 26336
rect 26108 26324 26114 26376
rect 26142 26324 26148 26376
rect 26200 26364 26206 26376
rect 28534 26364 28540 26376
rect 26200 26336 28540 26364
rect 26200 26324 26206 26336
rect 28534 26324 28540 26336
rect 28592 26324 28598 26376
rect 30558 26324 30564 26376
rect 30616 26324 30622 26376
rect 31757 26367 31815 26373
rect 31757 26333 31769 26367
rect 31803 26364 31815 26367
rect 31846 26364 31852 26376
rect 31803 26336 31852 26364
rect 31803 26333 31815 26336
rect 31757 26327 31815 26333
rect 31846 26324 31852 26336
rect 31904 26324 31910 26376
rect 32030 26373 32036 26376
rect 32024 26364 32036 26373
rect 31991 26336 32036 26364
rect 32024 26327 32036 26336
rect 32030 26324 32036 26327
rect 32088 26324 32094 26376
rect 32766 26324 32772 26376
rect 32824 26364 32830 26376
rect 33962 26364 33968 26376
rect 32824 26336 33968 26364
rect 32824 26324 32830 26336
rect 33962 26324 33968 26336
rect 34020 26324 34026 26376
rect 34146 26324 34152 26376
rect 34204 26364 34210 26376
rect 35529 26367 35587 26373
rect 35529 26364 35541 26367
rect 34204 26336 35541 26364
rect 34204 26324 34210 26336
rect 35529 26333 35541 26336
rect 35575 26364 35587 26367
rect 37366 26364 37372 26376
rect 35575 26336 37372 26364
rect 35575 26333 35587 26336
rect 35529 26327 35587 26333
rect 37366 26324 37372 26336
rect 37424 26324 37430 26376
rect 38194 26364 38200 26376
rect 38155 26336 38200 26364
rect 38194 26324 38200 26336
rect 38252 26364 38258 26376
rect 41616 26373 41644 26404
rect 42610 26392 42616 26404
rect 42668 26392 42674 26444
rect 42705 26435 42763 26441
rect 42705 26401 42717 26435
rect 42751 26401 42763 26435
rect 43254 26432 43260 26444
rect 42705 26395 42763 26401
rect 42812 26404 43260 26432
rect 38749 26367 38807 26373
rect 38749 26364 38761 26367
rect 38252 26336 38761 26364
rect 38252 26324 38258 26336
rect 38749 26333 38761 26336
rect 38795 26333 38807 26367
rect 38749 26327 38807 26333
rect 41601 26367 41659 26373
rect 41601 26333 41613 26367
rect 41647 26333 41659 26367
rect 41601 26327 41659 26333
rect 41690 26324 41696 26376
rect 41748 26364 41754 26376
rect 41877 26367 41935 26373
rect 41877 26364 41889 26367
rect 41748 26336 41889 26364
rect 41748 26324 41754 26336
rect 41877 26333 41889 26336
rect 41923 26333 41935 26367
rect 41877 26327 41935 26333
rect 41966 26324 41972 26376
rect 42024 26324 42030 26376
rect 42242 26324 42248 26376
rect 42300 26324 42306 26376
rect 42426 26324 42432 26376
rect 42484 26364 42490 26376
rect 42521 26367 42579 26373
rect 42521 26364 42533 26367
rect 42484 26336 42533 26364
rect 42484 26324 42490 26336
rect 42521 26333 42533 26336
rect 42567 26333 42579 26367
rect 42521 26327 42579 26333
rect 23860 26268 23980 26296
rect 23385 26259 23443 26265
rect 16592 26200 16988 26228
rect 17034 26188 17040 26240
rect 17092 26228 17098 26240
rect 17218 26228 17224 26240
rect 17092 26200 17224 26228
rect 17092 26188 17098 26200
rect 17218 26188 17224 26200
rect 17276 26188 17282 26240
rect 23750 26188 23756 26240
rect 23808 26228 23814 26240
rect 23845 26231 23903 26237
rect 23845 26228 23857 26231
rect 23808 26200 23857 26228
rect 23808 26188 23814 26200
rect 23845 26197 23857 26200
rect 23891 26197 23903 26231
rect 23952 26228 23980 26268
rect 26234 26256 26240 26308
rect 26292 26256 26298 26308
rect 30653 26299 30711 26305
rect 30653 26265 30665 26299
rect 30699 26296 30711 26299
rect 33318 26296 33324 26308
rect 30699 26268 33324 26296
rect 30699 26265 30711 26268
rect 30653 26259 30711 26265
rect 33318 26256 33324 26268
rect 33376 26256 33382 26308
rect 37090 26256 37096 26308
rect 37148 26296 37154 26308
rect 41785 26299 41843 26305
rect 41785 26296 41797 26299
rect 37148 26268 41797 26296
rect 37148 26256 37154 26268
rect 41785 26265 41797 26268
rect 41831 26265 41843 26299
rect 42720 26296 42748 26395
rect 42812 26373 42840 26404
rect 43254 26392 43260 26404
rect 43312 26432 43318 26444
rect 43533 26435 43591 26441
rect 43533 26432 43545 26435
rect 43312 26404 43545 26432
rect 43312 26392 43318 26404
rect 43533 26401 43545 26404
rect 43579 26401 43591 26435
rect 43533 26395 43591 26401
rect 42797 26367 42855 26373
rect 42797 26333 42809 26367
rect 42843 26333 42855 26367
rect 42797 26327 42855 26333
rect 42978 26324 42984 26376
rect 43036 26324 43042 26376
rect 43162 26324 43168 26376
rect 43220 26324 43226 26376
rect 43346 26324 43352 26376
rect 43404 26324 43410 26376
rect 45738 26324 45744 26376
rect 45796 26364 45802 26376
rect 46293 26367 46351 26373
rect 46293 26364 46305 26367
rect 45796 26336 46305 26364
rect 45796 26324 45802 26336
rect 46293 26333 46305 26336
rect 46339 26333 46351 26367
rect 46293 26327 46351 26333
rect 43990 26296 43996 26308
rect 41785 26259 41843 26265
rect 41984 26268 42656 26296
rect 42720 26268 43996 26296
rect 26050 26228 26056 26240
rect 23952 26200 26056 26228
rect 23845 26191 23903 26197
rect 26050 26188 26056 26200
rect 26108 26188 26114 26240
rect 38657 26231 38715 26237
rect 38657 26197 38669 26231
rect 38703 26228 38715 26231
rect 39114 26228 39120 26240
rect 38703 26200 39120 26228
rect 38703 26197 38715 26200
rect 38657 26191 38715 26197
rect 39114 26188 39120 26200
rect 39172 26188 39178 26240
rect 39209 26231 39267 26237
rect 39209 26197 39221 26231
rect 39255 26228 39267 26231
rect 39666 26228 39672 26240
rect 39255 26200 39672 26228
rect 39255 26197 39267 26200
rect 39209 26191 39267 26197
rect 39666 26188 39672 26200
rect 39724 26188 39730 26240
rect 41800 26228 41828 26259
rect 41984 26228 42012 26268
rect 41800 26200 42012 26228
rect 42628 26228 42656 26268
rect 43990 26256 43996 26268
rect 44048 26256 44054 26308
rect 43254 26228 43260 26240
rect 42628 26200 43260 26228
rect 43254 26188 43260 26200
rect 43312 26188 43318 26240
rect 1104 26138 47104 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 47104 26138
rect 1104 26064 47104 26086
rect 2038 25984 2044 26036
rect 2096 25984 2102 26036
rect 2409 26027 2467 26033
rect 2409 25993 2421 26027
rect 2455 25993 2467 26027
rect 2409 25987 2467 25993
rect 2225 25891 2283 25897
rect 2225 25857 2237 25891
rect 2271 25888 2283 25891
rect 2424 25888 2452 25987
rect 2774 25984 2780 26036
rect 2832 25984 2838 26036
rect 2866 25984 2872 26036
rect 2924 25984 2930 26036
rect 6270 26024 6276 26036
rect 3896 25996 6276 26024
rect 2271 25860 2452 25888
rect 2271 25857 2283 25860
rect 2225 25851 2283 25857
rect 3053 25823 3111 25829
rect 3053 25789 3065 25823
rect 3099 25820 3111 25823
rect 3896 25820 3924 25996
rect 6270 25984 6276 25996
rect 6328 25984 6334 26036
rect 12526 25984 12532 26036
rect 12584 26024 12590 26036
rect 13541 26027 13599 26033
rect 13541 26024 13553 26027
rect 12584 25996 13553 26024
rect 12584 25984 12590 25996
rect 13541 25993 13553 25996
rect 13587 25993 13599 26027
rect 13541 25987 13599 25993
rect 14826 25984 14832 26036
rect 14884 26024 14890 26036
rect 15746 26024 15752 26036
rect 14884 25996 15752 26024
rect 14884 25984 14890 25996
rect 15746 25984 15752 25996
rect 15804 25984 15810 26036
rect 17405 26027 17463 26033
rect 17405 25993 17417 26027
rect 17451 26024 17463 26027
rect 22002 26024 22008 26036
rect 17451 25996 22008 26024
rect 17451 25993 17463 25996
rect 17405 25987 17463 25993
rect 22002 25984 22008 25996
rect 22060 25984 22066 26036
rect 23106 25984 23112 26036
rect 23164 26024 23170 26036
rect 23937 26027 23995 26033
rect 23937 26024 23949 26027
rect 23164 25996 23949 26024
rect 23164 25984 23170 25996
rect 23937 25993 23949 25996
rect 23983 25993 23995 26027
rect 23937 25987 23995 25993
rect 25866 25984 25872 26036
rect 25924 26024 25930 26036
rect 29454 26024 29460 26036
rect 25924 25996 29460 26024
rect 25924 25984 25930 25996
rect 29454 25984 29460 25996
rect 29512 25984 29518 26036
rect 42886 26024 42892 26036
rect 42444 25996 42892 26024
rect 5813 25959 5871 25965
rect 5813 25925 5825 25959
rect 5859 25956 5871 25959
rect 9858 25956 9864 25968
rect 5859 25928 9864 25956
rect 5859 25925 5871 25928
rect 5813 25919 5871 25925
rect 9858 25916 9864 25928
rect 9916 25916 9922 25968
rect 13262 25956 13268 25968
rect 9968 25928 13268 25956
rect 3973 25891 4031 25897
rect 3973 25857 3985 25891
rect 4019 25888 4031 25891
rect 4062 25888 4068 25900
rect 4019 25860 4068 25888
rect 4019 25857 4031 25860
rect 3973 25851 4031 25857
rect 4062 25848 4068 25860
rect 4120 25848 4126 25900
rect 4890 25848 4896 25900
rect 4948 25848 4954 25900
rect 5074 25897 5080 25900
rect 5031 25891 5080 25897
rect 5031 25857 5043 25891
rect 5077 25857 5080 25891
rect 5031 25851 5080 25857
rect 5074 25848 5080 25851
rect 5132 25848 5138 25900
rect 7377 25891 7435 25897
rect 7377 25857 7389 25891
rect 7423 25888 7435 25891
rect 7650 25888 7656 25900
rect 7423 25860 7656 25888
rect 7423 25857 7435 25860
rect 7377 25851 7435 25857
rect 7650 25848 7656 25860
rect 7708 25848 7714 25900
rect 8570 25848 8576 25900
rect 8628 25848 8634 25900
rect 9033 25891 9091 25897
rect 9033 25857 9045 25891
rect 9079 25888 9091 25891
rect 9398 25888 9404 25900
rect 9079 25860 9404 25888
rect 9079 25857 9091 25860
rect 9033 25851 9091 25857
rect 9398 25848 9404 25860
rect 9456 25848 9462 25900
rect 9968 25897 9996 25928
rect 13262 25916 13268 25928
rect 13320 25916 13326 25968
rect 13357 25959 13415 25965
rect 13357 25925 13369 25959
rect 13403 25956 13415 25959
rect 13446 25956 13452 25968
rect 13403 25928 13452 25956
rect 13403 25925 13415 25928
rect 13357 25919 13415 25925
rect 13446 25916 13452 25928
rect 13504 25916 13510 25968
rect 14734 25956 14740 25968
rect 14200 25928 14740 25956
rect 9953 25891 10011 25897
rect 9953 25857 9965 25891
rect 9999 25857 10011 25891
rect 9953 25851 10011 25857
rect 10594 25848 10600 25900
rect 10652 25888 10658 25900
rect 14200 25897 14228 25928
rect 14734 25916 14740 25928
rect 14792 25916 14798 25968
rect 16298 25916 16304 25968
rect 16356 25956 16362 25968
rect 17586 25956 17592 25968
rect 16356 25928 17592 25956
rect 16356 25916 16362 25928
rect 17586 25916 17592 25928
rect 17644 25916 17650 25968
rect 20714 25956 20720 25968
rect 18156 25928 20720 25956
rect 11517 25891 11575 25897
rect 11517 25888 11529 25891
rect 10652 25860 11529 25888
rect 10652 25848 10658 25860
rect 11517 25857 11529 25860
rect 11563 25857 11575 25891
rect 13817 25891 13875 25897
rect 13817 25888 13829 25891
rect 11517 25851 11575 25857
rect 11624 25860 13829 25888
rect 3099 25792 3924 25820
rect 4157 25823 4215 25829
rect 3099 25789 3111 25792
rect 3053 25783 3111 25789
rect 4157 25789 4169 25823
rect 4203 25820 4215 25823
rect 4246 25820 4252 25832
rect 4203 25792 4252 25820
rect 4203 25789 4215 25792
rect 4157 25783 4215 25789
rect 4246 25780 4252 25792
rect 4304 25820 4310 25832
rect 5169 25823 5227 25829
rect 4304 25792 4568 25820
rect 4304 25780 4310 25792
rect 4540 25684 4568 25792
rect 5169 25789 5181 25823
rect 5215 25820 5227 25823
rect 5350 25820 5356 25832
rect 5215 25792 5356 25820
rect 5215 25789 5227 25792
rect 5169 25783 5227 25789
rect 5350 25780 5356 25792
rect 5408 25780 5414 25832
rect 7466 25780 7472 25832
rect 7524 25780 7530 25832
rect 7561 25823 7619 25829
rect 7561 25789 7573 25823
rect 7607 25820 7619 25823
rect 8018 25820 8024 25832
rect 7607 25792 8024 25820
rect 7607 25789 7619 25792
rect 7561 25783 7619 25789
rect 8018 25780 8024 25792
rect 8076 25780 8082 25832
rect 9122 25780 9128 25832
rect 9180 25820 9186 25832
rect 9309 25823 9367 25829
rect 9309 25820 9321 25823
rect 9180 25792 9321 25820
rect 9180 25780 9186 25792
rect 9309 25789 9321 25792
rect 9355 25789 9367 25823
rect 9309 25783 9367 25789
rect 9766 25780 9772 25832
rect 9824 25820 9830 25832
rect 10229 25823 10287 25829
rect 10229 25820 10241 25823
rect 9824 25792 10241 25820
rect 9824 25780 9830 25792
rect 10229 25789 10241 25792
rect 10275 25789 10287 25823
rect 10229 25783 10287 25789
rect 4617 25755 4675 25761
rect 4617 25721 4629 25755
rect 4663 25752 4675 25755
rect 4706 25752 4712 25764
rect 4663 25724 4712 25752
rect 4663 25721 4675 25724
rect 4617 25715 4675 25721
rect 4706 25712 4712 25724
rect 4764 25712 4770 25764
rect 6178 25712 6184 25764
rect 6236 25752 6242 25764
rect 6454 25752 6460 25764
rect 6236 25724 6460 25752
rect 6236 25712 6242 25724
rect 6454 25712 6460 25724
rect 6512 25752 6518 25764
rect 11624 25752 11652 25860
rect 13817 25857 13829 25860
rect 13863 25857 13875 25891
rect 13817 25851 13875 25857
rect 14185 25891 14243 25897
rect 14185 25857 14197 25891
rect 14231 25857 14243 25891
rect 14185 25851 14243 25857
rect 14274 25848 14280 25900
rect 14332 25848 14338 25900
rect 14366 25848 14372 25900
rect 14424 25848 14430 25900
rect 15470 25848 15476 25900
rect 15528 25848 15534 25900
rect 18156 25897 18184 25928
rect 20714 25916 20720 25928
rect 20772 25916 20778 25968
rect 20806 25916 20812 25968
rect 20864 25956 20870 25968
rect 34146 25956 34152 25968
rect 20864 25928 34152 25956
rect 20864 25916 20870 25928
rect 34146 25916 34152 25928
rect 34204 25916 34210 25968
rect 36725 25959 36783 25965
rect 36725 25925 36737 25959
rect 36771 25956 36783 25959
rect 41138 25956 41144 25968
rect 36771 25928 41144 25956
rect 36771 25925 36783 25928
rect 36725 25919 36783 25925
rect 41138 25916 41144 25928
rect 41196 25916 41202 25968
rect 17221 25891 17279 25897
rect 17221 25857 17233 25891
rect 17267 25888 17279 25891
rect 17865 25891 17923 25897
rect 17267 25860 17816 25888
rect 17267 25857 17279 25860
rect 17221 25851 17279 25857
rect 11790 25780 11796 25832
rect 11848 25780 11854 25832
rect 12437 25823 12495 25829
rect 12437 25789 12449 25823
rect 12483 25789 12495 25823
rect 12437 25783 12495 25789
rect 6512 25724 11652 25752
rect 12452 25752 12480 25783
rect 12618 25780 12624 25832
rect 12676 25820 12682 25832
rect 12713 25823 12771 25829
rect 12713 25820 12725 25823
rect 12676 25792 12725 25820
rect 12676 25780 12682 25792
rect 12713 25789 12725 25792
rect 12759 25789 12771 25823
rect 12986 25820 12992 25832
rect 12713 25783 12771 25789
rect 12820 25792 12992 25820
rect 12820 25752 12848 25792
rect 12986 25780 12992 25792
rect 13044 25820 13050 25832
rect 14090 25820 14096 25832
rect 13044 25792 14096 25820
rect 13044 25780 13050 25792
rect 14090 25780 14096 25792
rect 14148 25820 14154 25832
rect 15197 25823 15255 25829
rect 15197 25820 15209 25823
rect 14148 25792 15209 25820
rect 14148 25780 14154 25792
rect 15197 25789 15209 25792
rect 15243 25789 15255 25823
rect 15197 25783 15255 25789
rect 17236 25752 17264 25851
rect 17788 25820 17816 25860
rect 17865 25857 17877 25891
rect 17911 25888 17923 25891
rect 18141 25891 18199 25897
rect 18141 25888 18153 25891
rect 17911 25860 18153 25888
rect 17911 25857 17923 25860
rect 17865 25851 17923 25857
rect 18141 25857 18153 25860
rect 18187 25857 18199 25891
rect 18141 25851 18199 25857
rect 19061 25891 19119 25897
rect 19061 25857 19073 25891
rect 19107 25857 19119 25891
rect 19061 25851 19119 25857
rect 19076 25820 19104 25851
rect 23014 25848 23020 25900
rect 23072 25888 23078 25900
rect 23290 25888 23296 25900
rect 23072 25860 23296 25888
rect 23072 25848 23078 25860
rect 23290 25848 23296 25860
rect 23348 25848 23354 25900
rect 23382 25848 23388 25900
rect 23440 25848 23446 25900
rect 23661 25891 23719 25897
rect 23661 25888 23673 25891
rect 23492 25860 23673 25888
rect 17788 25792 19104 25820
rect 22002 25780 22008 25832
rect 22060 25820 22066 25832
rect 22830 25820 22836 25832
rect 22060 25792 22836 25820
rect 22060 25780 22066 25792
rect 22830 25780 22836 25792
rect 22888 25780 22894 25832
rect 12452 25724 12848 25752
rect 13464 25724 17264 25752
rect 6512 25712 6518 25724
rect 5166 25684 5172 25696
rect 4540 25656 5172 25684
rect 5166 25644 5172 25656
rect 5224 25644 5230 25696
rect 6822 25644 6828 25696
rect 6880 25684 6886 25696
rect 7009 25687 7067 25693
rect 7009 25684 7021 25687
rect 6880 25656 7021 25684
rect 6880 25644 6886 25656
rect 7009 25653 7021 25656
rect 7055 25653 7067 25687
rect 7009 25647 7067 25653
rect 8386 25644 8392 25696
rect 8444 25644 8450 25696
rect 10962 25644 10968 25696
rect 11020 25684 11026 25696
rect 13464 25684 13492 25724
rect 17310 25712 17316 25764
rect 17368 25752 17374 25764
rect 23492 25752 23520 25860
rect 23661 25857 23673 25860
rect 23707 25857 23719 25891
rect 23661 25851 23719 25857
rect 23845 25891 23903 25897
rect 23845 25857 23857 25891
rect 23891 25857 23903 25891
rect 23845 25851 23903 25857
rect 23569 25823 23627 25829
rect 23569 25789 23581 25823
rect 23615 25820 23627 25823
rect 23750 25820 23756 25832
rect 23615 25792 23756 25820
rect 23615 25789 23627 25792
rect 23569 25783 23627 25789
rect 23750 25780 23756 25792
rect 23808 25780 23814 25832
rect 17368 25724 23520 25752
rect 23860 25752 23888 25851
rect 25682 25848 25688 25900
rect 25740 25888 25746 25900
rect 25958 25888 25964 25900
rect 25740 25860 25964 25888
rect 25740 25848 25746 25860
rect 25958 25848 25964 25860
rect 26016 25848 26022 25900
rect 33042 25848 33048 25900
rect 33100 25888 33106 25900
rect 33781 25891 33839 25897
rect 33781 25888 33793 25891
rect 33100 25860 33793 25888
rect 33100 25848 33106 25860
rect 33781 25857 33793 25860
rect 33827 25857 33839 25891
rect 33781 25851 33839 25857
rect 36538 25848 36544 25900
rect 36596 25848 36602 25900
rect 36817 25891 36875 25897
rect 36817 25857 36829 25891
rect 36863 25888 36875 25891
rect 36998 25888 37004 25900
rect 36863 25860 37004 25888
rect 36863 25857 36875 25860
rect 36817 25851 36875 25857
rect 36998 25848 37004 25860
rect 37056 25888 37062 25900
rect 37918 25888 37924 25900
rect 37056 25860 37924 25888
rect 37056 25848 37062 25860
rect 37918 25848 37924 25860
rect 37976 25848 37982 25900
rect 39666 25848 39672 25900
rect 39724 25848 39730 25900
rect 42444 25897 42472 25996
rect 42886 25984 42892 25996
rect 42944 26024 42950 26036
rect 44082 26024 44088 26036
rect 42944 25996 44088 26024
rect 42944 25984 42950 25996
rect 44082 25984 44088 25996
rect 44140 25984 44146 26036
rect 45554 25984 45560 26036
rect 45612 26024 45618 26036
rect 46201 26027 46259 26033
rect 46201 26024 46213 26027
rect 45612 25996 46213 26024
rect 45612 25984 45618 25996
rect 46201 25993 46213 25996
rect 46247 25993 46259 26027
rect 46201 25987 46259 25993
rect 43990 25916 43996 25968
rect 44048 25956 44054 25968
rect 44048 25928 44404 25956
rect 44048 25916 44054 25928
rect 42429 25891 42487 25897
rect 42429 25857 42441 25891
rect 42475 25857 42487 25891
rect 42429 25851 42487 25857
rect 42518 25848 42524 25900
rect 42576 25888 42582 25900
rect 42889 25891 42947 25897
rect 42889 25888 42901 25891
rect 42576 25860 42901 25888
rect 42576 25848 42582 25860
rect 42889 25857 42901 25860
rect 42935 25857 42947 25891
rect 42889 25851 42947 25857
rect 43254 25848 43260 25900
rect 43312 25848 43318 25900
rect 44376 25897 44404 25928
rect 43533 25891 43591 25897
rect 43533 25857 43545 25891
rect 43579 25857 43591 25891
rect 44085 25891 44143 25897
rect 44085 25888 44097 25891
rect 43533 25851 43591 25857
rect 44008 25860 44097 25888
rect 30558 25780 30564 25832
rect 30616 25820 30622 25832
rect 33502 25820 33508 25832
rect 30616 25792 33508 25820
rect 30616 25780 30622 25792
rect 33502 25780 33508 25792
rect 33560 25780 33566 25832
rect 34422 25780 34428 25832
rect 34480 25820 34486 25832
rect 34698 25820 34704 25832
rect 34480 25792 34704 25820
rect 34480 25780 34486 25792
rect 34698 25780 34704 25792
rect 34756 25780 34762 25832
rect 42058 25780 42064 25832
rect 42116 25820 42122 25832
rect 42610 25820 42616 25832
rect 42116 25792 42616 25820
rect 42116 25780 42122 25792
rect 42610 25780 42616 25792
rect 42668 25780 42674 25832
rect 42794 25780 42800 25832
rect 42852 25780 42858 25832
rect 43162 25780 43168 25832
rect 43220 25820 43226 25832
rect 43548 25820 43576 25851
rect 43220 25792 43576 25820
rect 43220 25780 43226 25792
rect 36078 25752 36084 25764
rect 23860 25724 36084 25752
rect 17368 25712 17374 25724
rect 36078 25712 36084 25724
rect 36136 25712 36142 25764
rect 11020 25656 13492 25684
rect 11020 25644 11026 25656
rect 13538 25644 13544 25696
rect 13596 25644 13602 25696
rect 14182 25644 14188 25696
rect 14240 25684 14246 25696
rect 14553 25687 14611 25693
rect 14553 25684 14565 25687
rect 14240 25656 14565 25684
rect 14240 25644 14246 25656
rect 14553 25653 14565 25656
rect 14599 25684 14611 25687
rect 17494 25684 17500 25696
rect 14599 25656 17500 25684
rect 14599 25653 14611 25656
rect 14553 25647 14611 25653
rect 17494 25644 17500 25656
rect 17552 25644 17558 25696
rect 18046 25644 18052 25696
rect 18104 25684 18110 25696
rect 18371 25687 18429 25693
rect 18371 25684 18383 25687
rect 18104 25656 18383 25684
rect 18104 25644 18110 25656
rect 18371 25653 18383 25656
rect 18417 25653 18429 25687
rect 18371 25647 18429 25653
rect 19245 25687 19303 25693
rect 19245 25653 19257 25687
rect 19291 25684 19303 25687
rect 19794 25684 19800 25696
rect 19291 25656 19800 25684
rect 19291 25653 19303 25656
rect 19245 25647 19303 25653
rect 19794 25644 19800 25656
rect 19852 25644 19858 25696
rect 23109 25687 23167 25693
rect 23109 25653 23121 25687
rect 23155 25684 23167 25687
rect 23382 25684 23388 25696
rect 23155 25656 23388 25684
rect 23155 25653 23167 25656
rect 23109 25647 23167 25653
rect 23382 25644 23388 25656
rect 23440 25644 23446 25696
rect 26237 25687 26295 25693
rect 26237 25653 26249 25687
rect 26283 25684 26295 25687
rect 31110 25684 31116 25696
rect 26283 25656 31116 25684
rect 26283 25653 26295 25656
rect 26237 25647 26295 25653
rect 31110 25644 31116 25656
rect 31168 25684 31174 25696
rect 33594 25684 33600 25696
rect 31168 25656 33600 25684
rect 31168 25644 31174 25656
rect 33594 25644 33600 25656
rect 33652 25644 33658 25696
rect 36170 25644 36176 25696
rect 36228 25684 36234 25696
rect 36357 25687 36415 25693
rect 36357 25684 36369 25687
rect 36228 25656 36369 25684
rect 36228 25644 36234 25656
rect 36357 25653 36369 25656
rect 36403 25653 36415 25687
rect 36357 25647 36415 25653
rect 39485 25687 39543 25693
rect 39485 25653 39497 25687
rect 39531 25684 39543 25687
rect 40310 25684 40316 25696
rect 39531 25656 40316 25684
rect 39531 25653 39543 25656
rect 39485 25647 39543 25653
rect 40310 25644 40316 25656
rect 40368 25644 40374 25696
rect 42518 25644 42524 25696
rect 42576 25644 42582 25696
rect 43254 25644 43260 25696
rect 43312 25684 43318 25696
rect 43625 25687 43683 25693
rect 43625 25684 43637 25687
rect 43312 25656 43637 25684
rect 43312 25644 43318 25656
rect 43625 25653 43637 25656
rect 43671 25653 43683 25687
rect 43625 25647 43683 25653
rect 43898 25644 43904 25696
rect 43956 25684 43962 25696
rect 44008 25693 44036 25860
rect 44085 25857 44097 25860
rect 44131 25857 44143 25891
rect 44085 25851 44143 25857
rect 44269 25891 44327 25897
rect 44269 25857 44281 25891
rect 44315 25857 44327 25891
rect 44269 25851 44327 25857
rect 44361 25891 44419 25897
rect 44361 25857 44373 25891
rect 44407 25857 44419 25891
rect 44361 25851 44419 25857
rect 44082 25712 44088 25764
rect 44140 25752 44146 25764
rect 44284 25752 44312 25851
rect 45738 25848 45744 25900
rect 45796 25888 45802 25900
rect 46198 25888 46204 25900
rect 45796 25860 46204 25888
rect 45796 25848 45802 25860
rect 46198 25848 46204 25860
rect 46256 25848 46262 25900
rect 44140 25724 44312 25752
rect 44140 25712 44146 25724
rect 43993 25687 44051 25693
rect 43993 25684 44005 25687
rect 43956 25656 44005 25684
rect 43956 25644 43962 25656
rect 43993 25653 44005 25656
rect 44039 25653 44051 25687
rect 43993 25647 44051 25653
rect 44361 25687 44419 25693
rect 44361 25653 44373 25687
rect 44407 25684 44419 25687
rect 45278 25684 45284 25696
rect 44407 25656 45284 25684
rect 44407 25653 44419 25656
rect 44361 25647 44419 25653
rect 45278 25644 45284 25656
rect 45336 25644 45342 25696
rect 46014 25644 46020 25696
rect 46072 25684 46078 25696
rect 46290 25684 46296 25696
rect 46072 25656 46296 25684
rect 46072 25644 46078 25656
rect 46290 25644 46296 25656
rect 46348 25644 46354 25696
rect 1104 25594 47104 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 47104 25594
rect 1104 25520 47104 25542
rect 5166 25440 5172 25492
rect 5224 25440 5230 25492
rect 13078 25480 13084 25492
rect 9048 25452 13084 25480
rect 7466 25304 7472 25356
rect 7524 25344 7530 25356
rect 7745 25347 7803 25353
rect 7745 25344 7757 25347
rect 7524 25316 7757 25344
rect 7524 25304 7530 25316
rect 7745 25313 7757 25316
rect 7791 25313 7803 25347
rect 7745 25307 7803 25313
rect 7929 25347 7987 25353
rect 7929 25313 7941 25347
rect 7975 25344 7987 25347
rect 8018 25344 8024 25356
rect 7975 25316 8024 25344
rect 7975 25313 7987 25316
rect 7929 25307 7987 25313
rect 8018 25304 8024 25316
rect 8076 25304 8082 25356
rect 1670 25236 1676 25288
rect 1728 25276 1734 25288
rect 1857 25279 1915 25285
rect 1857 25276 1869 25279
rect 1728 25248 1869 25276
rect 1728 25236 1734 25248
rect 1857 25245 1869 25248
rect 1903 25276 1915 25279
rect 3789 25279 3847 25285
rect 3789 25276 3801 25279
rect 1903 25248 3801 25276
rect 1903 25245 1915 25248
rect 1857 25239 1915 25245
rect 3789 25245 3801 25248
rect 3835 25245 3847 25279
rect 3789 25239 3847 25245
rect 3878 25236 3884 25288
rect 3936 25276 3942 25288
rect 4045 25279 4103 25285
rect 4045 25276 4057 25279
rect 3936 25248 4057 25276
rect 3936 25236 3942 25248
rect 4045 25245 4057 25248
rect 4091 25245 4103 25279
rect 4045 25239 4103 25245
rect 6822 25236 6828 25288
rect 6880 25236 6886 25288
rect 7650 25236 7656 25288
rect 7708 25276 7714 25288
rect 9048 25276 9076 25452
rect 13078 25440 13084 25452
rect 13136 25440 13142 25492
rect 14093 25483 14151 25489
rect 14093 25449 14105 25483
rect 14139 25480 14151 25483
rect 14366 25480 14372 25492
rect 14139 25452 14372 25480
rect 14139 25449 14151 25452
rect 14093 25443 14151 25449
rect 14366 25440 14372 25452
rect 14424 25440 14430 25492
rect 18690 25480 18696 25492
rect 15856 25452 18696 25480
rect 12710 25372 12716 25424
rect 12768 25372 12774 25424
rect 9125 25347 9183 25353
rect 9125 25313 9137 25347
rect 9171 25344 9183 25347
rect 9766 25344 9772 25356
rect 9171 25316 9772 25344
rect 9171 25313 9183 25316
rect 9125 25307 9183 25313
rect 9766 25304 9772 25316
rect 9824 25304 9830 25356
rect 9858 25304 9864 25356
rect 9916 25344 9922 25356
rect 12437 25347 12495 25353
rect 12437 25344 12449 25347
rect 9916 25316 12449 25344
rect 9916 25304 9922 25316
rect 12437 25313 12449 25316
rect 12483 25313 12495 25347
rect 12437 25307 12495 25313
rect 12802 25304 12808 25356
rect 12860 25344 12866 25356
rect 15856 25353 15884 25452
rect 18690 25440 18696 25452
rect 18748 25440 18754 25492
rect 21729 25483 21787 25489
rect 21729 25449 21741 25483
rect 21775 25480 21787 25483
rect 28902 25480 28908 25492
rect 21775 25452 28908 25480
rect 21775 25449 21787 25452
rect 21729 25443 21787 25449
rect 28902 25440 28908 25452
rect 28960 25440 28966 25492
rect 33870 25480 33876 25492
rect 31726 25452 33876 25480
rect 16206 25372 16212 25424
rect 16264 25412 16270 25424
rect 17310 25412 17316 25424
rect 16264 25384 17316 25412
rect 16264 25372 16270 25384
rect 17310 25372 17316 25384
rect 17368 25372 17374 25424
rect 17494 25372 17500 25424
rect 17552 25412 17558 25424
rect 17552 25384 21496 25412
rect 17552 25372 17558 25384
rect 14737 25347 14795 25353
rect 14737 25344 14749 25347
rect 12860 25316 14749 25344
rect 12860 25304 12866 25316
rect 7708 25248 9076 25276
rect 7708 25236 7714 25248
rect 9398 25236 9404 25288
rect 9456 25236 9462 25288
rect 12158 25236 12164 25288
rect 12216 25276 12222 25288
rect 12529 25279 12587 25285
rect 12529 25276 12541 25279
rect 12216 25248 12541 25276
rect 12216 25236 12222 25248
rect 12529 25245 12541 25248
rect 12575 25276 12587 25279
rect 12618 25276 12624 25288
rect 12575 25248 12624 25276
rect 12575 25245 12587 25248
rect 12529 25239 12587 25245
rect 12618 25236 12624 25248
rect 12676 25236 12682 25288
rect 14090 25236 14096 25288
rect 14148 25236 14154 25288
rect 14292 25285 14320 25316
rect 14737 25313 14749 25316
rect 14783 25313 14795 25347
rect 14737 25307 14795 25313
rect 15013 25347 15071 25353
rect 15013 25313 15025 25347
rect 15059 25344 15071 25347
rect 15749 25347 15807 25353
rect 15749 25344 15761 25347
rect 15059 25316 15761 25344
rect 15059 25313 15071 25316
rect 15013 25307 15071 25313
rect 15749 25313 15761 25316
rect 15795 25313 15807 25347
rect 15749 25307 15807 25313
rect 15841 25347 15899 25353
rect 15841 25313 15853 25347
rect 15887 25313 15899 25347
rect 15841 25307 15899 25313
rect 14277 25279 14335 25285
rect 14277 25245 14289 25279
rect 14323 25245 14335 25279
rect 14277 25239 14335 25245
rect 2124 25211 2182 25217
rect 2124 25177 2136 25211
rect 2170 25208 2182 25211
rect 2774 25208 2780 25220
rect 2170 25180 2780 25208
rect 2170 25177 2182 25180
rect 2124 25171 2182 25177
rect 2774 25168 2780 25180
rect 2832 25168 2838 25220
rect 8938 25168 8944 25220
rect 8996 25208 9002 25220
rect 9416 25208 9444 25236
rect 8996 25180 9444 25208
rect 8996 25168 9002 25180
rect 3234 25100 3240 25152
rect 3292 25100 3298 25152
rect 6546 25100 6552 25152
rect 6604 25140 6610 25152
rect 6641 25143 6699 25149
rect 6641 25140 6653 25143
rect 6604 25112 6653 25140
rect 6604 25100 6610 25112
rect 6641 25109 6653 25112
rect 6687 25109 6699 25143
rect 6641 25103 6699 25109
rect 7282 25100 7288 25152
rect 7340 25100 7346 25152
rect 12066 25100 12072 25152
rect 12124 25100 12130 25152
rect 15764 25140 15792 25307
rect 16224 25285 16252 25372
rect 16758 25344 16764 25356
rect 16408 25316 16764 25344
rect 16209 25279 16267 25285
rect 16209 25245 16221 25279
rect 16255 25245 16267 25279
rect 16209 25239 16267 25245
rect 16298 25236 16304 25288
rect 16356 25236 16362 25288
rect 16408 25285 16436 25316
rect 16758 25304 16764 25316
rect 16816 25304 16822 25356
rect 16853 25347 16911 25353
rect 16853 25313 16865 25347
rect 16899 25344 16911 25347
rect 20806 25344 20812 25356
rect 16899 25316 20812 25344
rect 16899 25313 16911 25316
rect 16853 25307 16911 25313
rect 20806 25304 20812 25316
rect 20864 25304 20870 25356
rect 21266 25304 21272 25356
rect 21324 25304 21330 25356
rect 16393 25279 16451 25285
rect 16393 25245 16405 25279
rect 16439 25245 16451 25279
rect 17034 25276 17040 25288
rect 16393 25239 16451 25245
rect 16500 25248 17040 25276
rect 16500 25140 16528 25248
rect 17034 25236 17040 25248
rect 17092 25276 17098 25288
rect 17221 25279 17279 25285
rect 17221 25276 17233 25279
rect 17092 25248 17233 25276
rect 17092 25236 17098 25248
rect 17221 25245 17233 25248
rect 17267 25245 17279 25279
rect 17221 25239 17279 25245
rect 17310 25236 17316 25288
rect 17368 25236 17374 25288
rect 17402 25236 17408 25288
rect 17460 25236 17466 25288
rect 17957 25279 18015 25285
rect 17957 25245 17969 25279
rect 18003 25245 18015 25279
rect 17957 25239 18015 25245
rect 17972 25208 18000 25239
rect 18046 25236 18052 25288
rect 18104 25236 18110 25288
rect 18230 25236 18236 25288
rect 18288 25276 18294 25288
rect 18325 25279 18383 25285
rect 18325 25276 18337 25279
rect 18288 25248 18337 25276
rect 18288 25236 18294 25248
rect 18325 25245 18337 25248
rect 18371 25245 18383 25279
rect 18325 25239 18383 25245
rect 18248 25208 18276 25236
rect 17972 25180 18276 25208
rect 21468 25208 21496 25384
rect 21542 25372 21548 25424
rect 21600 25372 21606 25424
rect 24118 25372 24124 25424
rect 24176 25372 24182 25424
rect 26329 25415 26387 25421
rect 26329 25381 26341 25415
rect 26375 25412 26387 25415
rect 30650 25412 30656 25424
rect 26375 25384 30656 25412
rect 26375 25381 26387 25384
rect 26329 25375 26387 25381
rect 30650 25372 30656 25384
rect 30708 25412 30714 25424
rect 31726 25412 31754 25452
rect 33870 25440 33876 25452
rect 33928 25440 33934 25492
rect 37369 25483 37427 25489
rect 37369 25449 37381 25483
rect 37415 25480 37427 25483
rect 38378 25480 38384 25492
rect 37415 25452 38384 25480
rect 37415 25449 37427 25452
rect 37369 25443 37427 25449
rect 38378 25440 38384 25452
rect 38436 25440 38442 25492
rect 30708 25384 31754 25412
rect 37553 25415 37611 25421
rect 30708 25372 30714 25384
rect 37553 25381 37565 25415
rect 37599 25381 37611 25415
rect 37553 25375 37611 25381
rect 36262 25344 36268 25356
rect 27172 25316 33272 25344
rect 22094 25236 22100 25288
rect 22152 25276 22158 25288
rect 23106 25276 23112 25288
rect 22152 25248 23112 25276
rect 22152 25236 22158 25248
rect 23106 25236 23112 25248
rect 23164 25236 23170 25288
rect 23382 25236 23388 25288
rect 23440 25236 23446 25288
rect 26234 25276 26240 25288
rect 23492 25248 26240 25276
rect 23492 25208 23520 25248
rect 26234 25236 26240 25248
rect 26292 25236 26298 25288
rect 27172 25285 27200 25316
rect 27157 25279 27215 25285
rect 27157 25245 27169 25279
rect 27203 25245 27215 25279
rect 27157 25239 27215 25245
rect 29914 25236 29920 25288
rect 29972 25276 29978 25288
rect 30834 25276 30840 25288
rect 29972 25248 30840 25276
rect 29972 25236 29978 25248
rect 30834 25236 30840 25248
rect 30892 25236 30898 25288
rect 31018 25236 31024 25288
rect 31076 25236 31082 25288
rect 31754 25236 31760 25288
rect 31812 25276 31818 25288
rect 33042 25276 33048 25288
rect 31812 25248 33048 25276
rect 31812 25236 31818 25248
rect 33042 25236 33048 25248
rect 33100 25276 33106 25288
rect 33137 25279 33195 25285
rect 33137 25276 33149 25279
rect 33100 25248 33149 25276
rect 33100 25236 33106 25248
rect 33137 25245 33149 25248
rect 33183 25245 33195 25279
rect 33244 25276 33272 25316
rect 34900 25316 36268 25344
rect 34900 25276 34928 25316
rect 36262 25304 36268 25316
rect 36320 25304 36326 25356
rect 37274 25304 37280 25356
rect 37332 25304 37338 25356
rect 37568 25344 37596 25375
rect 38838 25372 38844 25424
rect 38896 25412 38902 25424
rect 39025 25415 39083 25421
rect 39025 25412 39037 25415
rect 38896 25384 39037 25412
rect 38896 25372 38902 25384
rect 39025 25381 39037 25384
rect 39071 25381 39083 25415
rect 39025 25375 39083 25381
rect 45278 25372 45284 25424
rect 45336 25372 45342 25424
rect 40129 25347 40187 25353
rect 37568 25316 38884 25344
rect 33244 25248 34928 25276
rect 34977 25279 35035 25285
rect 33137 25239 33195 25245
rect 34977 25245 34989 25279
rect 35023 25276 35035 25279
rect 35342 25276 35348 25288
rect 35023 25248 35348 25276
rect 35023 25245 35035 25248
rect 34977 25239 35035 25245
rect 35342 25236 35348 25248
rect 35400 25236 35406 25288
rect 36538 25236 36544 25288
rect 36596 25236 36602 25288
rect 37090 25236 37096 25288
rect 37148 25276 37154 25288
rect 37185 25279 37243 25285
rect 37185 25276 37197 25279
rect 37148 25248 37197 25276
rect 37148 25236 37154 25248
rect 37185 25245 37197 25248
rect 37231 25245 37243 25279
rect 37185 25239 37243 25245
rect 37921 25279 37979 25285
rect 37921 25245 37933 25279
rect 37967 25245 37979 25279
rect 37921 25239 37979 25245
rect 38381 25279 38439 25285
rect 38381 25245 38393 25279
rect 38427 25245 38439 25279
rect 38381 25239 38439 25245
rect 21468 25180 23520 25208
rect 26050 25168 26056 25220
rect 26108 25168 26114 25220
rect 28166 25208 28172 25220
rect 26896 25180 28172 25208
rect 15764 25112 16528 25140
rect 17770 25100 17776 25152
rect 17828 25100 17834 25152
rect 25222 25100 25228 25152
rect 25280 25140 25286 25152
rect 26896 25140 26924 25180
rect 28166 25168 28172 25180
rect 28224 25168 28230 25220
rect 33226 25168 33232 25220
rect 33284 25208 33290 25220
rect 33382 25211 33440 25217
rect 33382 25208 33394 25211
rect 33284 25180 33394 25208
rect 33284 25168 33290 25180
rect 33382 25177 33394 25180
rect 33428 25177 33440 25211
rect 33382 25171 33440 25177
rect 25280 25112 26924 25140
rect 25280 25100 25286 25112
rect 26970 25100 26976 25152
rect 27028 25100 27034 25152
rect 30834 25100 30840 25152
rect 30892 25100 30898 25152
rect 34330 25100 34336 25152
rect 34388 25140 34394 25152
rect 34514 25140 34520 25152
rect 34388 25112 34520 25140
rect 34388 25100 34394 25112
rect 34514 25100 34520 25112
rect 34572 25100 34578 25152
rect 34793 25143 34851 25149
rect 34793 25109 34805 25143
rect 34839 25140 34851 25143
rect 35434 25140 35440 25152
rect 34839 25112 35440 25140
rect 34839 25109 34851 25112
rect 34793 25103 34851 25109
rect 35434 25100 35440 25112
rect 35492 25100 35498 25152
rect 37936 25140 37964 25239
rect 38396 25208 38424 25239
rect 38470 25236 38476 25288
rect 38528 25236 38534 25288
rect 38856 25285 38884 25316
rect 40129 25313 40141 25347
rect 40175 25344 40187 25347
rect 43714 25344 43720 25356
rect 40175 25316 43720 25344
rect 40175 25313 40187 25316
rect 40129 25307 40187 25313
rect 43714 25304 43720 25316
rect 43772 25304 43778 25356
rect 43898 25304 43904 25356
rect 43956 25304 43962 25356
rect 45830 25304 45836 25356
rect 45888 25344 45894 25356
rect 46201 25347 46259 25353
rect 46201 25344 46213 25347
rect 45888 25316 46213 25344
rect 45888 25304 45894 25316
rect 46201 25313 46213 25316
rect 46247 25313 46259 25347
rect 46201 25307 46259 25313
rect 38841 25279 38899 25285
rect 38841 25245 38853 25279
rect 38887 25245 38899 25279
rect 38841 25239 38899 25245
rect 39114 25236 39120 25288
rect 39172 25276 39178 25288
rect 40037 25279 40095 25285
rect 40037 25276 40049 25279
rect 39172 25248 40049 25276
rect 39172 25236 39178 25248
rect 40037 25245 40049 25248
rect 40083 25245 40095 25279
rect 40037 25239 40095 25245
rect 40310 25236 40316 25288
rect 40368 25236 40374 25288
rect 43990 25236 43996 25288
rect 44048 25236 44054 25288
rect 44450 25236 44456 25288
rect 44508 25236 44514 25288
rect 44542 25236 44548 25288
rect 44600 25276 44606 25288
rect 44729 25279 44787 25285
rect 44729 25276 44741 25279
rect 44600 25248 44741 25276
rect 44600 25236 44606 25248
rect 44729 25245 44741 25248
rect 44775 25245 44787 25279
rect 44729 25239 44787 25245
rect 45922 25236 45928 25288
rect 45980 25236 45986 25288
rect 38746 25208 38752 25220
rect 38396 25180 38752 25208
rect 38746 25168 38752 25180
rect 38804 25168 38810 25220
rect 39298 25168 39304 25220
rect 39356 25168 39362 25220
rect 44269 25211 44327 25217
rect 44269 25177 44281 25211
rect 44315 25208 44327 25211
rect 45005 25211 45063 25217
rect 45005 25208 45017 25211
rect 44315 25180 45017 25208
rect 44315 25177 44327 25180
rect 44269 25171 44327 25177
rect 45005 25177 45017 25180
rect 45051 25208 45063 25211
rect 45738 25208 45744 25220
rect 45051 25180 45744 25208
rect 45051 25177 45063 25180
rect 45005 25171 45063 25177
rect 45738 25168 45744 25180
rect 45796 25168 45802 25220
rect 38838 25140 38844 25152
rect 37936 25112 38844 25140
rect 38838 25100 38844 25112
rect 38896 25100 38902 25152
rect 38930 25100 38936 25152
rect 38988 25140 38994 25152
rect 39393 25143 39451 25149
rect 39393 25140 39405 25143
rect 38988 25112 39405 25140
rect 38988 25100 38994 25112
rect 39393 25109 39405 25112
rect 39439 25109 39451 25143
rect 39393 25103 39451 25109
rect 39853 25143 39911 25149
rect 39853 25109 39865 25143
rect 39899 25140 39911 25143
rect 40034 25140 40040 25152
rect 39899 25112 40040 25140
rect 39899 25109 39911 25112
rect 39853 25103 39911 25109
rect 40034 25100 40040 25112
rect 40092 25100 40098 25152
rect 40773 25143 40831 25149
rect 40773 25109 40785 25143
rect 40819 25140 40831 25143
rect 40862 25140 40868 25152
rect 40819 25112 40868 25140
rect 40819 25109 40831 25112
rect 40773 25103 40831 25109
rect 40862 25100 40868 25112
rect 40920 25100 40926 25152
rect 44726 25100 44732 25152
rect 44784 25140 44790 25152
rect 45465 25143 45523 25149
rect 45465 25140 45477 25143
rect 44784 25112 45477 25140
rect 44784 25100 44790 25112
rect 45465 25109 45477 25112
rect 45511 25109 45523 25143
rect 45465 25103 45523 25109
rect 1104 25050 47104 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 47104 25050
rect 1104 24976 47104 24998
rect 2774 24896 2780 24948
rect 2832 24896 2838 24948
rect 5258 24896 5264 24948
rect 5316 24936 5322 24948
rect 5626 24936 5632 24948
rect 5316 24908 5632 24936
rect 5316 24896 5322 24908
rect 5626 24896 5632 24908
rect 5684 24896 5690 24948
rect 13262 24896 13268 24948
rect 13320 24936 13326 24948
rect 18046 24936 18052 24948
rect 13320 24908 18052 24936
rect 13320 24896 13326 24908
rect 18046 24896 18052 24908
rect 18104 24936 18110 24948
rect 18598 24936 18604 24948
rect 18104 24908 18604 24936
rect 18104 24896 18110 24908
rect 18598 24896 18604 24908
rect 18656 24896 18662 24948
rect 19245 24939 19303 24945
rect 19245 24936 19257 24939
rect 19168 24908 19257 24936
rect 2317 24871 2375 24877
rect 2317 24837 2329 24871
rect 2363 24868 2375 24871
rect 5534 24868 5540 24880
rect 2363 24840 5540 24868
rect 2363 24837 2375 24840
rect 2317 24831 2375 24837
rect 5534 24828 5540 24840
rect 5592 24868 5598 24880
rect 5994 24868 6000 24880
rect 5592 24840 6000 24868
rect 5592 24828 5598 24840
rect 5994 24828 6000 24840
rect 6052 24828 6058 24880
rect 8386 24828 8392 24880
rect 8444 24868 8450 24880
rect 9278 24871 9336 24877
rect 9278 24868 9290 24871
rect 8444 24840 9290 24868
rect 8444 24828 8450 24840
rect 9278 24837 9290 24840
rect 9324 24837 9336 24871
rect 18230 24868 18236 24880
rect 9278 24831 9336 24837
rect 16684 24840 18236 24868
rect 934 24760 940 24812
rect 992 24800 998 24812
rect 1397 24803 1455 24809
rect 1397 24800 1409 24803
rect 992 24772 1409 24800
rect 992 24760 998 24772
rect 1397 24769 1409 24772
rect 1443 24769 1455 24803
rect 2961 24803 3019 24809
rect 2961 24800 2973 24803
rect 1397 24763 1455 24769
rect 2746 24772 2973 24800
rect 2406 24692 2412 24744
rect 2464 24692 2470 24744
rect 2498 24692 2504 24744
rect 2556 24692 2562 24744
rect 1949 24667 2007 24673
rect 1949 24633 1961 24667
rect 1995 24664 2007 24667
rect 2746 24664 2774 24772
rect 2961 24769 2973 24772
rect 3007 24769 3019 24803
rect 2961 24763 3019 24769
rect 7374 24760 7380 24812
rect 7432 24800 7438 24812
rect 7817 24803 7875 24809
rect 7817 24800 7829 24803
rect 7432 24772 7829 24800
rect 7432 24760 7438 24772
rect 7817 24769 7829 24772
rect 7863 24769 7875 24803
rect 9122 24800 9128 24812
rect 7817 24763 7875 24769
rect 9048 24772 9128 24800
rect 7190 24692 7196 24744
rect 7248 24732 7254 24744
rect 9048 24741 9076 24772
rect 9122 24760 9128 24772
rect 9180 24760 9186 24812
rect 9674 24760 9680 24812
rect 9732 24800 9738 24812
rect 12161 24803 12219 24809
rect 12161 24800 12173 24803
rect 9732 24772 12173 24800
rect 9732 24760 9738 24772
rect 12161 24769 12173 24772
rect 12207 24769 12219 24803
rect 12161 24763 12219 24769
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24800 12311 24803
rect 12434 24800 12440 24812
rect 12299 24772 12440 24800
rect 12299 24769 12311 24772
rect 12253 24763 12311 24769
rect 12434 24760 12440 24772
rect 12492 24760 12498 24812
rect 16684 24809 16712 24840
rect 18230 24828 18236 24840
rect 18288 24828 18294 24880
rect 16669 24803 16727 24809
rect 16669 24769 16681 24803
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 18040 24803 18098 24809
rect 18040 24769 18052 24803
rect 18086 24800 18098 24803
rect 19168 24800 19196 24908
rect 19245 24905 19257 24908
rect 19291 24905 19303 24939
rect 19245 24899 19303 24905
rect 19886 24896 19892 24948
rect 19944 24936 19950 24948
rect 25222 24936 25228 24948
rect 19944 24908 25228 24936
rect 19944 24896 19950 24908
rect 25222 24896 25228 24908
rect 25280 24896 25286 24948
rect 26970 24936 26976 24948
rect 25424 24908 26976 24936
rect 19352 24840 19564 24868
rect 19352 24800 19380 24840
rect 18086 24772 19196 24800
rect 19306 24772 19380 24800
rect 18086 24769 18098 24772
rect 18040 24763 18098 24769
rect 7561 24735 7619 24741
rect 7561 24732 7573 24735
rect 7248 24704 7573 24732
rect 7248 24692 7254 24704
rect 7561 24701 7573 24704
rect 7607 24701 7619 24735
rect 9033 24735 9091 24741
rect 9033 24732 9045 24735
rect 7561 24695 7619 24701
rect 8588 24704 9045 24732
rect 1995 24636 2774 24664
rect 1995 24633 2007 24636
rect 1949 24627 2007 24633
rect 1578 24556 1584 24608
rect 1636 24556 1642 24608
rect 7576 24596 7604 24695
rect 8588 24596 8616 24704
rect 9033 24701 9045 24704
rect 9079 24701 9091 24735
rect 9033 24695 9091 24701
rect 11514 24692 11520 24744
rect 11572 24732 11578 24744
rect 11793 24735 11851 24741
rect 11793 24732 11805 24735
rect 11572 24704 11805 24732
rect 11572 24692 11578 24704
rect 11793 24701 11805 24704
rect 11839 24701 11851 24735
rect 11793 24695 11851 24701
rect 16022 24692 16028 24744
rect 16080 24732 16086 24744
rect 16945 24735 17003 24741
rect 16945 24732 16957 24735
rect 16080 24704 16957 24732
rect 16080 24692 16086 24704
rect 16945 24701 16957 24704
rect 16991 24701 17003 24735
rect 16945 24695 17003 24701
rect 17770 24692 17776 24744
rect 17828 24692 17834 24744
rect 18966 24692 18972 24744
rect 19024 24732 19030 24744
rect 19306 24732 19334 24772
rect 19426 24760 19432 24812
rect 19484 24760 19490 24812
rect 19536 24800 19564 24840
rect 21266 24828 21272 24880
rect 21324 24868 21330 24880
rect 23201 24871 23259 24877
rect 23201 24868 23213 24871
rect 21324 24840 23213 24868
rect 21324 24828 21330 24840
rect 23201 24837 23213 24840
rect 23247 24868 23259 24871
rect 24486 24868 24492 24880
rect 23247 24840 24492 24868
rect 23247 24837 23259 24840
rect 23201 24831 23259 24837
rect 24486 24828 24492 24840
rect 24544 24828 24550 24880
rect 19536 24772 19932 24800
rect 19024 24704 19334 24732
rect 19024 24692 19030 24704
rect 19518 24692 19524 24744
rect 19576 24692 19582 24744
rect 19705 24735 19763 24741
rect 19705 24701 19717 24735
rect 19751 24701 19763 24735
rect 19705 24695 19763 24701
rect 14090 24664 14096 24676
rect 10336 24636 14096 24664
rect 7576 24568 8616 24596
rect 8941 24599 8999 24605
rect 8941 24565 8953 24599
rect 8987 24596 8999 24599
rect 10336 24596 10364 24636
rect 14090 24624 14096 24636
rect 14148 24624 14154 24676
rect 19610 24664 19616 24676
rect 19076 24636 19616 24664
rect 8987 24568 10364 24596
rect 10413 24599 10471 24605
rect 8987 24565 8999 24568
rect 8941 24559 8999 24565
rect 10413 24565 10425 24599
rect 10459 24596 10471 24599
rect 10594 24596 10600 24608
rect 10459 24568 10600 24596
rect 10459 24565 10471 24568
rect 10413 24559 10471 24565
rect 10594 24556 10600 24568
rect 10652 24556 10658 24608
rect 12437 24599 12495 24605
rect 12437 24565 12449 24599
rect 12483 24596 12495 24599
rect 19076 24596 19104 24636
rect 19610 24624 19616 24636
rect 19668 24624 19674 24676
rect 12483 24568 19104 24596
rect 12483 24565 12495 24568
rect 12437 24559 12495 24565
rect 19150 24556 19156 24608
rect 19208 24596 19214 24608
rect 19720 24596 19748 24695
rect 19208 24568 19748 24596
rect 19904 24596 19932 24772
rect 22370 24760 22376 24812
rect 22428 24760 22434 24812
rect 24949 24803 25007 24809
rect 24949 24769 24961 24803
rect 24995 24800 25007 24803
rect 25222 24800 25228 24812
rect 24995 24772 25228 24800
rect 24995 24769 25007 24772
rect 24949 24763 25007 24769
rect 25222 24760 25228 24772
rect 25280 24760 25286 24812
rect 25424 24809 25452 24908
rect 26970 24896 26976 24908
rect 27028 24896 27034 24948
rect 33137 24939 33195 24945
rect 33137 24905 33149 24939
rect 33183 24936 33195 24939
rect 33226 24936 33232 24948
rect 33183 24908 33232 24936
rect 33183 24905 33195 24908
rect 33137 24899 33195 24905
rect 33226 24896 33232 24908
rect 33284 24896 33290 24948
rect 36170 24896 36176 24948
rect 36228 24896 36234 24948
rect 36262 24896 36268 24948
rect 36320 24936 36326 24948
rect 36906 24936 36912 24948
rect 36320 24908 36912 24936
rect 36320 24896 36326 24908
rect 36906 24896 36912 24908
rect 36964 24936 36970 24948
rect 37001 24939 37059 24945
rect 37001 24936 37013 24939
rect 36964 24908 37013 24936
rect 36964 24896 36970 24908
rect 37001 24905 37013 24908
rect 37047 24905 37059 24939
rect 37001 24899 37059 24905
rect 41138 24896 41144 24948
rect 41196 24896 41202 24948
rect 41690 24936 41696 24948
rect 41248 24908 41696 24936
rect 30377 24871 30435 24877
rect 25608 24840 26188 24868
rect 25409 24803 25467 24809
rect 25409 24769 25421 24803
rect 25455 24769 25467 24803
rect 25409 24763 25467 24769
rect 25498 24760 25504 24812
rect 25556 24800 25562 24812
rect 25608 24800 25636 24840
rect 25556 24772 25636 24800
rect 25676 24803 25734 24809
rect 25556 24760 25562 24772
rect 25676 24769 25688 24803
rect 25722 24800 25734 24803
rect 26050 24800 26056 24812
rect 25722 24772 26056 24800
rect 25722 24769 25734 24772
rect 25676 24763 25734 24769
rect 26050 24760 26056 24772
rect 26108 24760 26114 24812
rect 26160 24800 26188 24840
rect 27172 24840 27384 24868
rect 27172 24800 27200 24840
rect 27246 24809 27252 24812
rect 26160 24772 27200 24800
rect 27240 24763 27252 24809
rect 27246 24760 27252 24763
rect 27304 24760 27310 24812
rect 27356 24800 27384 24840
rect 30377 24837 30389 24871
rect 30423 24868 30435 24871
rect 30650 24868 30656 24880
rect 30423 24840 30656 24868
rect 30423 24837 30435 24840
rect 30377 24831 30435 24837
rect 30650 24828 30656 24840
rect 30708 24828 30714 24880
rect 30834 24877 30840 24880
rect 30828 24868 30840 24877
rect 30795 24840 30840 24868
rect 30828 24831 30840 24840
rect 30834 24828 30840 24831
rect 30892 24828 30898 24880
rect 28718 24800 28724 24812
rect 27356 24772 28724 24800
rect 28718 24760 28724 24772
rect 28776 24760 28782 24812
rect 30190 24760 30196 24812
rect 30248 24760 30254 24812
rect 30466 24760 30472 24812
rect 30524 24760 30530 24812
rect 32398 24760 32404 24812
rect 32456 24760 32462 24812
rect 33318 24760 33324 24812
rect 33376 24760 33382 24812
rect 34330 24760 34336 24812
rect 34388 24760 34394 24812
rect 34606 24760 34612 24812
rect 34664 24760 34670 24812
rect 36188 24744 36216 24896
rect 37274 24828 37280 24880
rect 37332 24868 37338 24880
rect 38381 24871 38439 24877
rect 38381 24868 38393 24871
rect 37332 24840 38393 24868
rect 37332 24828 37338 24840
rect 38381 24837 38393 24840
rect 38427 24837 38439 24871
rect 38381 24831 38439 24837
rect 38838 24828 38844 24880
rect 38896 24868 38902 24880
rect 41248 24868 41276 24908
rect 41690 24896 41696 24908
rect 41748 24896 41754 24948
rect 43993 24939 44051 24945
rect 43993 24905 44005 24939
rect 44039 24936 44051 24939
rect 44174 24936 44180 24948
rect 44039 24908 44180 24936
rect 44039 24905 44051 24908
rect 43993 24899 44051 24905
rect 44174 24896 44180 24908
rect 44232 24896 44238 24948
rect 41782 24868 41788 24880
rect 38896 24840 41276 24868
rect 41340 24840 41788 24868
rect 38896 24828 38902 24840
rect 36354 24760 36360 24812
rect 36412 24800 36418 24812
rect 36449 24803 36507 24809
rect 36449 24800 36461 24803
rect 36412 24772 36461 24800
rect 36412 24760 36418 24772
rect 36449 24769 36461 24772
rect 36495 24800 36507 24803
rect 36909 24803 36967 24809
rect 36909 24800 36921 24803
rect 36495 24772 36921 24800
rect 36495 24769 36507 24772
rect 36449 24763 36507 24769
rect 36909 24769 36921 24772
rect 36955 24769 36967 24803
rect 36909 24763 36967 24769
rect 38562 24760 38568 24812
rect 38620 24760 38626 24812
rect 38933 24803 38991 24809
rect 38933 24769 38945 24803
rect 38979 24769 38991 24803
rect 38933 24763 38991 24769
rect 20438 24692 20444 24744
rect 20496 24692 20502 24744
rect 20530 24692 20536 24744
rect 20588 24741 20594 24744
rect 20588 24735 20616 24741
rect 20604 24701 20616 24735
rect 20588 24695 20616 24701
rect 20717 24735 20775 24741
rect 20717 24701 20729 24735
rect 20763 24732 20775 24735
rect 21450 24732 21456 24744
rect 20763 24704 21456 24732
rect 20763 24701 20775 24704
rect 20717 24695 20775 24701
rect 20588 24692 20594 24695
rect 21450 24692 21456 24704
rect 21508 24692 21514 24744
rect 22094 24692 22100 24744
rect 22152 24692 22158 24744
rect 26970 24692 26976 24744
rect 27028 24692 27034 24744
rect 29086 24692 29092 24744
rect 29144 24732 29150 24744
rect 29144 24704 29776 24732
rect 29144 24692 29150 24704
rect 20165 24667 20223 24673
rect 20165 24633 20177 24667
rect 20211 24664 20223 24667
rect 20254 24664 20260 24676
rect 20211 24636 20260 24664
rect 20211 24633 20223 24636
rect 20165 24627 20223 24633
rect 20254 24624 20260 24636
rect 20312 24624 20318 24676
rect 23569 24667 23627 24673
rect 22756 24636 23244 24664
rect 20714 24596 20720 24608
rect 19904 24568 20720 24596
rect 19208 24556 19214 24568
rect 20714 24556 20720 24568
rect 20772 24556 20778 24608
rect 21361 24599 21419 24605
rect 21361 24565 21373 24599
rect 21407 24596 21419 24599
rect 21910 24596 21916 24608
rect 21407 24568 21916 24596
rect 21407 24565 21419 24568
rect 21361 24559 21419 24565
rect 21910 24556 21916 24568
rect 21968 24556 21974 24608
rect 22462 24556 22468 24608
rect 22520 24596 22526 24608
rect 22756 24596 22784 24636
rect 22520 24568 22784 24596
rect 22520 24556 22526 24568
rect 23106 24556 23112 24608
rect 23164 24556 23170 24608
rect 23216 24596 23244 24636
rect 23569 24633 23581 24667
rect 23615 24664 23627 24667
rect 29362 24664 29368 24676
rect 23615 24636 25452 24664
rect 23615 24633 23627 24636
rect 23569 24627 23627 24633
rect 23661 24599 23719 24605
rect 23661 24596 23673 24599
rect 23216 24568 23673 24596
rect 23661 24565 23673 24568
rect 23707 24565 23719 24599
rect 23661 24559 23719 24565
rect 24670 24556 24676 24608
rect 24728 24596 24734 24608
rect 24765 24599 24823 24605
rect 24765 24596 24777 24599
rect 24728 24568 24777 24596
rect 24728 24556 24734 24568
rect 24765 24565 24777 24568
rect 24811 24565 24823 24599
rect 25424 24596 25452 24636
rect 28276 24636 29368 24664
rect 26602 24596 26608 24608
rect 25424 24568 26608 24596
rect 24765 24559 24823 24565
rect 26602 24556 26608 24568
rect 26660 24556 26666 24608
rect 26694 24556 26700 24608
rect 26752 24596 26758 24608
rect 26789 24599 26847 24605
rect 26789 24596 26801 24599
rect 26752 24568 26801 24596
rect 26752 24556 26758 24568
rect 26789 24565 26801 24568
rect 26835 24565 26847 24599
rect 26789 24559 26847 24565
rect 26970 24556 26976 24608
rect 27028 24596 27034 24608
rect 28276 24596 28304 24636
rect 29362 24624 29368 24636
rect 29420 24624 29426 24676
rect 29457 24667 29515 24673
rect 29457 24633 29469 24667
rect 29503 24664 29515 24667
rect 29638 24664 29644 24676
rect 29503 24636 29644 24664
rect 29503 24633 29515 24636
rect 29457 24627 29515 24633
rect 29638 24624 29644 24636
rect 29696 24624 29702 24676
rect 29748 24664 29776 24704
rect 30006 24692 30012 24744
rect 30064 24732 30070 24744
rect 30558 24732 30564 24744
rect 30064 24704 30564 24732
rect 30064 24692 30070 24704
rect 30558 24692 30564 24704
rect 30616 24692 30622 24744
rect 33410 24692 33416 24744
rect 33468 24692 33474 24744
rect 33597 24735 33655 24741
rect 33597 24701 33609 24735
rect 33643 24732 33655 24735
rect 33778 24732 33784 24744
rect 33643 24704 33784 24732
rect 33643 24701 33655 24704
rect 33597 24695 33655 24701
rect 33778 24692 33784 24704
rect 33836 24692 33842 24744
rect 33962 24692 33968 24744
rect 34020 24732 34026 24744
rect 34057 24735 34115 24741
rect 34057 24732 34069 24735
rect 34020 24704 34069 24732
rect 34020 24692 34026 24704
rect 34057 24701 34069 24704
rect 34103 24701 34115 24735
rect 34057 24695 34115 24701
rect 34146 24692 34152 24744
rect 34204 24732 34210 24744
rect 34450 24735 34508 24741
rect 34450 24732 34462 24735
rect 34204 24704 34462 24732
rect 34204 24692 34210 24704
rect 34450 24701 34462 24704
rect 34496 24701 34508 24735
rect 34450 24695 34508 24701
rect 36170 24692 36176 24744
rect 36228 24692 36234 24744
rect 38948 24732 38976 24763
rect 39206 24760 39212 24812
rect 39264 24800 39270 24812
rect 39301 24803 39359 24809
rect 39301 24800 39313 24803
rect 39264 24772 39313 24800
rect 39264 24760 39270 24772
rect 39301 24769 39313 24772
rect 39347 24769 39359 24803
rect 39301 24763 39359 24769
rect 39574 24760 39580 24812
rect 39632 24760 39638 24812
rect 40512 24809 40540 24840
rect 40497 24803 40555 24809
rect 40497 24769 40509 24803
rect 40543 24769 40555 24803
rect 40497 24763 40555 24769
rect 40678 24760 40684 24812
rect 40736 24760 40742 24812
rect 40773 24803 40831 24809
rect 40773 24769 40785 24803
rect 40819 24769 40831 24803
rect 40773 24763 40831 24769
rect 39390 24732 39396 24744
rect 38948 24704 39396 24732
rect 39390 24692 39396 24704
rect 39448 24732 39454 24744
rect 39853 24735 39911 24741
rect 39853 24732 39865 24735
rect 39448 24704 39865 24732
rect 39448 24692 39454 24704
rect 39853 24701 39865 24704
rect 39899 24701 39911 24735
rect 40788 24732 40816 24763
rect 40862 24760 40868 24812
rect 40920 24760 40926 24812
rect 41340 24809 41368 24840
rect 41782 24828 41788 24840
rect 41840 24828 41846 24880
rect 44542 24868 44548 24880
rect 43916 24840 44548 24868
rect 41325 24803 41383 24809
rect 41325 24769 41337 24803
rect 41371 24769 41383 24803
rect 41325 24763 41383 24769
rect 41414 24760 41420 24812
rect 41472 24800 41478 24812
rect 42518 24800 42524 24812
rect 41472 24772 42524 24800
rect 41472 24760 41478 24772
rect 42518 24760 42524 24772
rect 42576 24760 42582 24812
rect 43916 24809 43944 24840
rect 44542 24828 44548 24840
rect 44600 24828 44606 24880
rect 43901 24803 43959 24809
rect 43901 24769 43913 24803
rect 43947 24800 43959 24803
rect 43990 24800 43996 24812
rect 43947 24772 43996 24800
rect 43947 24769 43959 24772
rect 43901 24763 43959 24769
rect 43990 24760 43996 24772
rect 44048 24760 44054 24812
rect 44085 24803 44143 24809
rect 44085 24769 44097 24803
rect 44131 24800 44143 24803
rect 44450 24800 44456 24812
rect 44131 24772 44456 24800
rect 44131 24769 44143 24772
rect 44085 24763 44143 24769
rect 44450 24760 44456 24772
rect 44508 24760 44514 24812
rect 44726 24760 44732 24812
rect 44784 24760 44790 24812
rect 46382 24760 46388 24812
rect 46440 24800 46446 24812
rect 46477 24803 46535 24809
rect 46477 24800 46489 24803
rect 46440 24772 46489 24800
rect 46440 24760 46446 24772
rect 46477 24769 46489 24772
rect 46523 24769 46535 24803
rect 46477 24763 46535 24769
rect 41230 24732 41236 24744
rect 40788 24704 41236 24732
rect 39853 24695 39911 24701
rect 41230 24692 41236 24704
rect 41288 24692 41294 24744
rect 41506 24692 41512 24744
rect 41564 24692 41570 24744
rect 41601 24735 41659 24741
rect 41601 24701 41613 24735
rect 41647 24701 41659 24735
rect 41601 24695 41659 24701
rect 30374 24664 30380 24676
rect 29748 24636 30380 24664
rect 30374 24624 30380 24636
rect 30432 24624 30438 24676
rect 32950 24624 32956 24676
rect 33008 24664 33014 24676
rect 33980 24664 34008 24692
rect 40126 24664 40132 24676
rect 33008 24636 34008 24664
rect 39224 24636 40132 24664
rect 33008 24624 33014 24636
rect 39224 24608 39252 24636
rect 40126 24624 40132 24636
rect 40184 24624 40190 24676
rect 41049 24667 41107 24673
rect 41049 24633 41061 24667
rect 41095 24664 41107 24667
rect 41616 24664 41644 24695
rect 41095 24636 41644 24664
rect 41095 24633 41107 24636
rect 41049 24627 41107 24633
rect 43714 24624 43720 24676
rect 43772 24664 43778 24676
rect 44545 24667 44603 24673
rect 44545 24664 44557 24667
rect 43772 24636 44557 24664
rect 43772 24624 43778 24636
rect 44545 24633 44557 24636
rect 44591 24633 44603 24667
rect 44545 24627 44603 24633
rect 27028 24568 28304 24596
rect 27028 24556 27034 24568
rect 28350 24556 28356 24608
rect 28408 24556 28414 24608
rect 29549 24599 29607 24605
rect 29549 24565 29561 24599
rect 29595 24596 29607 24599
rect 29730 24596 29736 24608
rect 29595 24568 29736 24596
rect 29595 24565 29607 24568
rect 29549 24559 29607 24565
rect 29730 24556 29736 24568
rect 29788 24556 29794 24608
rect 29822 24556 29828 24608
rect 29880 24596 29886 24608
rect 30009 24599 30067 24605
rect 30009 24596 30021 24599
rect 29880 24568 30021 24596
rect 29880 24556 29886 24568
rect 30009 24565 30021 24568
rect 30055 24565 30067 24599
rect 30009 24559 30067 24565
rect 31662 24556 31668 24608
rect 31720 24596 31726 24608
rect 31941 24599 31999 24605
rect 31941 24596 31953 24599
rect 31720 24568 31953 24596
rect 31720 24556 31726 24568
rect 31941 24565 31953 24568
rect 31987 24565 31999 24599
rect 31941 24559 31999 24565
rect 32214 24556 32220 24608
rect 32272 24556 32278 24608
rect 33226 24556 33232 24608
rect 33284 24596 33290 24608
rect 35253 24599 35311 24605
rect 35253 24596 35265 24599
rect 33284 24568 35265 24596
rect 33284 24556 33290 24568
rect 35253 24565 35265 24568
rect 35299 24565 35311 24599
rect 35253 24559 35311 24565
rect 39025 24599 39083 24605
rect 39025 24565 39037 24599
rect 39071 24596 39083 24599
rect 39206 24596 39212 24608
rect 39071 24568 39212 24596
rect 39071 24565 39083 24568
rect 39025 24559 39083 24565
rect 39206 24556 39212 24568
rect 39264 24556 39270 24608
rect 39393 24599 39451 24605
rect 39393 24565 39405 24599
rect 39439 24596 39451 24599
rect 39482 24596 39488 24608
rect 39439 24568 39488 24596
rect 39439 24565 39451 24568
rect 39393 24559 39451 24565
rect 39482 24556 39488 24568
rect 39540 24556 39546 24608
rect 46566 24556 46572 24608
rect 46624 24556 46630 24608
rect 1104 24506 47104 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 47104 24506
rect 1104 24432 47104 24454
rect 6288 24364 7236 24392
rect 6288 24268 6316 24364
rect 7208 24324 7236 24364
rect 7466 24352 7472 24404
rect 7524 24392 7530 24404
rect 7653 24395 7711 24401
rect 7653 24392 7665 24395
rect 7524 24364 7665 24392
rect 7524 24352 7530 24364
rect 7653 24361 7665 24364
rect 7699 24361 7711 24395
rect 12713 24395 12771 24401
rect 12713 24392 12725 24395
rect 7653 24355 7711 24361
rect 11164 24364 12725 24392
rect 8938 24324 8944 24336
rect 7208 24296 8944 24324
rect 8938 24284 8944 24296
rect 8996 24284 9002 24336
rect 5169 24259 5227 24265
rect 5169 24225 5181 24259
rect 5215 24225 5227 24259
rect 5169 24219 5227 24225
rect 4522 24148 4528 24200
rect 4580 24188 4586 24200
rect 4798 24188 4804 24200
rect 4580 24160 4804 24188
rect 4580 24148 4586 24160
rect 4798 24148 4804 24160
rect 4856 24188 4862 24200
rect 4856 24160 5145 24188
rect 4856 24148 4862 24160
rect 3694 24080 3700 24132
rect 3752 24120 3758 24132
rect 4985 24123 5043 24129
rect 4985 24120 4997 24123
rect 3752 24092 4997 24120
rect 3752 24080 3758 24092
rect 4985 24089 4997 24092
rect 5031 24089 5043 24123
rect 4985 24083 5043 24089
rect 4525 24055 4583 24061
rect 4525 24021 4537 24055
rect 4571 24052 4583 24055
rect 4614 24052 4620 24064
rect 4571 24024 4620 24052
rect 4571 24021 4583 24024
rect 4525 24015 4583 24021
rect 4614 24012 4620 24024
rect 4672 24012 4678 24064
rect 4798 24012 4804 24064
rect 4856 24052 4862 24064
rect 4893 24055 4951 24061
rect 4893 24052 4905 24055
rect 4856 24024 4905 24052
rect 4856 24012 4862 24024
rect 4893 24021 4905 24024
rect 4939 24021 4951 24055
rect 5117 24052 5145 24160
rect 5184 24120 5212 24219
rect 6270 24216 6276 24268
rect 6328 24216 6334 24268
rect 6546 24197 6552 24200
rect 6540 24188 6552 24197
rect 6507 24160 6552 24188
rect 6540 24151 6552 24160
rect 6546 24148 6552 24151
rect 6604 24148 6610 24200
rect 7282 24148 7288 24200
rect 7340 24188 7346 24200
rect 11164 24197 11192 24364
rect 12713 24361 12725 24364
rect 12759 24361 12771 24395
rect 12713 24355 12771 24361
rect 14366 24352 14372 24404
rect 14424 24392 14430 24404
rect 14645 24395 14703 24401
rect 14645 24392 14657 24395
rect 14424 24364 14657 24392
rect 14424 24352 14430 24364
rect 14645 24361 14657 24364
rect 14691 24392 14703 24395
rect 14691 24364 17080 24392
rect 14691 24361 14703 24364
rect 14645 24355 14703 24361
rect 12621 24327 12679 24333
rect 12621 24293 12633 24327
rect 12667 24324 12679 24327
rect 13078 24324 13084 24336
rect 12667 24296 13084 24324
rect 12667 24293 12679 24296
rect 12621 24287 12679 24293
rect 13078 24284 13084 24296
rect 13136 24284 13142 24336
rect 13630 24284 13636 24336
rect 13688 24324 13694 24336
rect 13688 24296 16068 24324
rect 13688 24284 13694 24296
rect 13096 24197 13124 24284
rect 16040 24268 16068 24296
rect 13170 24216 13176 24268
rect 13228 24256 13234 24268
rect 13265 24259 13323 24265
rect 13265 24256 13277 24259
rect 13228 24228 13277 24256
rect 13228 24216 13234 24228
rect 13265 24225 13277 24228
rect 13311 24225 13323 24259
rect 13265 24219 13323 24225
rect 14108 24228 14964 24256
rect 14108 24200 14136 24228
rect 7929 24191 7987 24197
rect 7929 24188 7941 24191
rect 7340 24160 7941 24188
rect 7340 24148 7346 24160
rect 7929 24157 7941 24160
rect 7975 24157 7987 24191
rect 7929 24151 7987 24157
rect 11149 24191 11207 24197
rect 11149 24157 11161 24191
rect 11195 24157 11207 24191
rect 11149 24151 11207 24157
rect 11241 24191 11299 24197
rect 11241 24157 11253 24191
rect 11287 24188 11299 24191
rect 13081 24191 13139 24197
rect 11287 24160 12434 24188
rect 11287 24157 11299 24160
rect 11241 24151 11299 24157
rect 9306 24120 9312 24132
rect 5184 24092 9312 24120
rect 9306 24080 9312 24092
rect 9364 24080 9370 24132
rect 11486 24123 11544 24129
rect 11486 24120 11498 24123
rect 10980 24092 11498 24120
rect 7374 24052 7380 24064
rect 5117 24024 7380 24052
rect 4893 24015 4951 24021
rect 7374 24012 7380 24024
rect 7432 24012 7438 24064
rect 7745 24055 7803 24061
rect 7745 24021 7757 24055
rect 7791 24052 7803 24055
rect 8294 24052 8300 24064
rect 7791 24024 8300 24052
rect 7791 24021 7803 24024
rect 7745 24015 7803 24021
rect 8294 24012 8300 24024
rect 8352 24012 8358 24064
rect 10980 24061 11008 24092
rect 11486 24089 11498 24092
rect 11532 24089 11544 24123
rect 12406 24120 12434 24160
rect 13081 24157 13093 24191
rect 13127 24157 13139 24191
rect 13081 24151 13139 24157
rect 14090 24148 14096 24200
rect 14148 24148 14154 24200
rect 14936 24197 14964 24228
rect 16022 24216 16028 24268
rect 16080 24216 16086 24268
rect 14461 24191 14519 24197
rect 14461 24188 14473 24191
rect 14292 24160 14473 24188
rect 12802 24120 12808 24132
rect 12406 24092 12808 24120
rect 11486 24083 11544 24089
rect 12802 24080 12808 24092
rect 12860 24120 12866 24132
rect 13630 24120 13636 24132
rect 12860 24092 13636 24120
rect 12860 24080 12866 24092
rect 13630 24080 13636 24092
rect 13688 24080 13694 24132
rect 10965 24055 11023 24061
rect 10965 24021 10977 24055
rect 11011 24021 11023 24055
rect 10965 24015 11023 24021
rect 13173 24055 13231 24061
rect 13173 24021 13185 24055
rect 13219 24052 13231 24055
rect 13262 24052 13268 24064
rect 13219 24024 13268 24052
rect 13219 24021 13231 24024
rect 13173 24015 13231 24021
rect 13262 24012 13268 24024
rect 13320 24012 13326 24064
rect 13354 24012 13360 24064
rect 13412 24052 13418 24064
rect 14292 24061 14320 24160
rect 14461 24157 14473 24160
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 14921 24191 14979 24197
rect 14921 24157 14933 24191
rect 14967 24157 14979 24191
rect 14921 24151 14979 24157
rect 15930 24148 15936 24200
rect 15988 24148 15994 24200
rect 16270 24123 16328 24129
rect 16270 24120 16282 24123
rect 15764 24092 16282 24120
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 13412 24024 14289 24052
rect 13412 24012 13418 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 14277 24015 14335 24021
rect 14550 24012 14556 24064
rect 14608 24052 14614 24064
rect 15010 24052 15016 24064
rect 14608 24024 15016 24052
rect 14608 24012 14614 24024
rect 15010 24012 15016 24024
rect 15068 24012 15074 24064
rect 15105 24055 15163 24061
rect 15105 24021 15117 24055
rect 15151 24052 15163 24055
rect 15470 24052 15476 24064
rect 15151 24024 15476 24052
rect 15151 24021 15163 24024
rect 15105 24015 15163 24021
rect 15470 24012 15476 24024
rect 15528 24012 15534 24064
rect 15764 24061 15792 24092
rect 16270 24089 16282 24092
rect 16316 24089 16328 24123
rect 17052 24120 17080 24364
rect 17586 24352 17592 24404
rect 17644 24352 17650 24404
rect 18141 24395 18199 24401
rect 18141 24361 18153 24395
rect 18187 24392 18199 24395
rect 19426 24392 19432 24404
rect 18187 24364 19432 24392
rect 18187 24361 18199 24364
rect 18141 24355 18199 24361
rect 19426 24352 19432 24364
rect 19484 24352 19490 24404
rect 19610 24352 19616 24404
rect 19668 24392 19674 24404
rect 21361 24395 21419 24401
rect 19668 24364 21312 24392
rect 19668 24352 19674 24364
rect 17604 24324 17632 24352
rect 17604 24296 20300 24324
rect 18785 24259 18843 24265
rect 18785 24225 18797 24259
rect 18831 24256 18843 24259
rect 18874 24256 18880 24268
rect 18831 24228 18880 24256
rect 18831 24225 18843 24228
rect 18785 24219 18843 24225
rect 18874 24216 18880 24228
rect 18932 24216 18938 24268
rect 19705 24259 19763 24265
rect 19705 24256 19717 24259
rect 19444 24228 19717 24256
rect 18509 24191 18567 24197
rect 18509 24157 18521 24191
rect 18555 24188 18567 24191
rect 19150 24188 19156 24200
rect 18555 24160 19156 24188
rect 18555 24157 18567 24160
rect 18509 24151 18567 24157
rect 19150 24148 19156 24160
rect 19208 24188 19214 24200
rect 19444 24188 19472 24228
rect 19705 24225 19717 24228
rect 19751 24225 19763 24259
rect 19705 24219 19763 24225
rect 20162 24216 20168 24268
rect 20220 24216 20226 24268
rect 20272 24256 20300 24296
rect 20530 24256 20536 24268
rect 20588 24265 20594 24268
rect 20588 24259 20616 24265
rect 20272 24228 20536 24256
rect 20530 24216 20536 24228
rect 20604 24225 20616 24259
rect 20588 24219 20616 24225
rect 20588 24216 20594 24219
rect 20714 24216 20720 24268
rect 20772 24216 20778 24268
rect 19208 24160 19472 24188
rect 19208 24148 19214 24160
rect 19518 24148 19524 24200
rect 19576 24148 19582 24200
rect 20438 24148 20444 24200
rect 20496 24148 20502 24200
rect 19702 24120 19708 24132
rect 17052 24092 19708 24120
rect 16270 24083 16328 24089
rect 19702 24080 19708 24092
rect 19760 24080 19766 24132
rect 15749 24055 15807 24061
rect 15749 24021 15761 24055
rect 15795 24021 15807 24055
rect 15749 24015 15807 24021
rect 17402 24012 17408 24064
rect 17460 24012 17466 24064
rect 17586 24012 17592 24064
rect 17644 24052 17650 24064
rect 18601 24055 18659 24061
rect 18601 24052 18613 24055
rect 17644 24024 18613 24052
rect 17644 24012 17650 24024
rect 18601 24021 18613 24024
rect 18647 24052 18659 24055
rect 20162 24052 20168 24064
rect 18647 24024 20168 24052
rect 18647 24021 18659 24024
rect 18601 24015 18659 24021
rect 20162 24012 20168 24024
rect 20220 24012 20226 24064
rect 21284 24052 21312 24364
rect 21361 24361 21373 24395
rect 21407 24392 21419 24395
rect 21542 24392 21548 24404
rect 21407 24364 21548 24392
rect 21407 24361 21419 24364
rect 21361 24355 21419 24361
rect 21542 24352 21548 24364
rect 21600 24352 21606 24404
rect 22189 24395 22247 24401
rect 22189 24361 22201 24395
rect 22235 24392 22247 24395
rect 22370 24392 22376 24404
rect 22235 24364 22376 24392
rect 22235 24361 22247 24364
rect 22189 24355 22247 24361
rect 22370 24352 22376 24364
rect 22428 24352 22434 24404
rect 23106 24352 23112 24404
rect 23164 24392 23170 24404
rect 23164 24364 26004 24392
rect 23164 24352 23170 24364
rect 21910 24284 21916 24336
rect 21968 24284 21974 24336
rect 22830 24284 22836 24336
rect 22888 24324 22894 24336
rect 25976 24324 26004 24364
rect 26050 24352 26056 24404
rect 26108 24352 26114 24404
rect 26970 24392 26976 24404
rect 26620 24364 26976 24392
rect 26620 24324 26648 24364
rect 26970 24352 26976 24364
rect 27028 24352 27034 24404
rect 27157 24395 27215 24401
rect 27157 24361 27169 24395
rect 27203 24392 27215 24395
rect 27246 24392 27252 24404
rect 27203 24364 27252 24392
rect 27203 24361 27215 24364
rect 27157 24355 27215 24361
rect 27246 24352 27252 24364
rect 27304 24352 27310 24404
rect 27890 24352 27896 24404
rect 27948 24392 27954 24404
rect 28626 24392 28632 24404
rect 27948 24364 28632 24392
rect 27948 24352 27954 24364
rect 28626 24352 28632 24364
rect 28684 24352 28690 24404
rect 28718 24352 28724 24404
rect 28776 24392 28782 24404
rect 30009 24395 30067 24401
rect 30009 24392 30021 24395
rect 28776 24364 30021 24392
rect 28776 24352 28782 24364
rect 30009 24361 30021 24364
rect 30055 24361 30067 24395
rect 30009 24355 30067 24361
rect 30837 24395 30895 24401
rect 30837 24361 30849 24395
rect 30883 24392 30895 24395
rect 31018 24392 31024 24404
rect 30883 24364 31024 24392
rect 30883 24361 30895 24364
rect 30837 24355 30895 24361
rect 31018 24352 31024 24364
rect 31076 24352 31082 24404
rect 33226 24392 33232 24404
rect 31726 24364 33232 24392
rect 22888 24296 23060 24324
rect 25976 24296 26648 24324
rect 22888 24284 22894 24296
rect 22097 24259 22155 24265
rect 22097 24225 22109 24259
rect 22143 24256 22155 24259
rect 22649 24259 22707 24265
rect 22143 24228 22600 24256
rect 22143 24225 22155 24228
rect 22097 24219 22155 24225
rect 22370 24148 22376 24200
rect 22428 24148 22434 24200
rect 22465 24191 22523 24197
rect 22465 24157 22477 24191
rect 22511 24157 22523 24191
rect 22572 24188 22600 24228
rect 22649 24225 22661 24259
rect 22695 24256 22707 24259
rect 23032 24256 23060 24296
rect 26694 24284 26700 24336
rect 26752 24324 26758 24336
rect 26752 24296 28212 24324
rect 26752 24284 26758 24296
rect 23382 24256 23388 24268
rect 22695 24228 22968 24256
rect 22695 24225 22707 24228
rect 22649 24219 22707 24225
rect 22741 24191 22799 24197
rect 22741 24188 22753 24191
rect 22572 24160 22753 24188
rect 22465 24151 22523 24157
rect 22741 24157 22753 24160
rect 22787 24157 22799 24191
rect 22741 24151 22799 24157
rect 21634 24080 21640 24132
rect 21692 24080 21698 24132
rect 22480 24120 22508 24151
rect 22833 24123 22891 24129
rect 22833 24120 22845 24123
rect 22480 24092 22845 24120
rect 22833 24089 22845 24092
rect 22879 24089 22891 24123
rect 22833 24083 22891 24089
rect 22940 24052 22968 24228
rect 23032 24228 23388 24256
rect 23032 24197 23060 24228
rect 23382 24216 23388 24228
rect 23440 24216 23446 24268
rect 26970 24216 26976 24268
rect 27028 24216 27034 24268
rect 27433 24259 27491 24265
rect 27433 24225 27445 24259
rect 27479 24256 27491 24259
rect 27522 24256 27528 24268
rect 27479 24228 27528 24256
rect 27479 24225 27491 24228
rect 27433 24219 27491 24225
rect 27522 24216 27528 24228
rect 27580 24216 27586 24268
rect 28074 24216 28080 24268
rect 28132 24216 28138 24268
rect 28184 24256 28212 24296
rect 29086 24284 29092 24336
rect 29144 24324 29150 24336
rect 31726 24324 31754 24364
rect 33226 24352 33232 24364
rect 33284 24352 33290 24404
rect 33318 24352 33324 24404
rect 33376 24392 33382 24404
rect 33597 24395 33655 24401
rect 33597 24392 33609 24395
rect 33376 24364 33609 24392
rect 33376 24352 33382 24364
rect 33597 24361 33609 24364
rect 33643 24361 33655 24395
rect 33597 24355 33655 24361
rect 33778 24352 33784 24404
rect 33836 24392 33842 24404
rect 36814 24392 36820 24404
rect 33836 24364 36820 24392
rect 33836 24352 33842 24364
rect 36814 24352 36820 24364
rect 36872 24352 36878 24404
rect 36998 24352 37004 24404
rect 37056 24392 37062 24404
rect 39485 24395 39543 24401
rect 37056 24364 38884 24392
rect 37056 24352 37062 24364
rect 29144 24296 31754 24324
rect 29144 24284 29150 24296
rect 33502 24284 33508 24336
rect 33560 24324 33566 24336
rect 33560 24296 35388 24324
rect 33560 24284 33566 24296
rect 28470 24259 28528 24265
rect 28470 24256 28482 24259
rect 28184 24228 28482 24256
rect 28470 24225 28482 24228
rect 28516 24256 28528 24259
rect 28994 24256 29000 24268
rect 28516 24228 29000 24256
rect 28516 24225 28528 24228
rect 28470 24219 28528 24225
rect 28994 24216 29000 24228
rect 29052 24216 29058 24268
rect 29178 24216 29184 24268
rect 29236 24256 29242 24268
rect 29236 24228 29960 24256
rect 29236 24216 29242 24228
rect 23017 24191 23075 24197
rect 23017 24157 23029 24191
rect 23063 24157 23075 24191
rect 23017 24151 23075 24157
rect 23198 24148 23204 24200
rect 23256 24188 23262 24200
rect 23293 24191 23351 24197
rect 23293 24188 23305 24191
rect 23256 24160 23305 24188
rect 23256 24148 23262 24160
rect 23293 24157 23305 24160
rect 23339 24188 23351 24191
rect 23750 24188 23756 24200
rect 23339 24160 23756 24188
rect 23339 24157 23351 24160
rect 23293 24151 23351 24157
rect 23750 24148 23756 24160
rect 23808 24188 23814 24200
rect 23934 24188 23940 24200
rect 23808 24160 23940 24188
rect 23808 24148 23814 24160
rect 23934 24148 23940 24160
rect 23992 24148 23998 24200
rect 24302 24148 24308 24200
rect 24360 24188 24366 24200
rect 24670 24197 24676 24200
rect 24397 24191 24455 24197
rect 24397 24188 24409 24191
rect 24360 24160 24409 24188
rect 24360 24148 24366 24160
rect 24397 24157 24409 24160
rect 24443 24157 24455 24191
rect 24664 24188 24676 24197
rect 24631 24160 24676 24188
rect 24397 24151 24455 24157
rect 24664 24151 24676 24160
rect 24670 24148 24676 24151
rect 24728 24148 24734 24200
rect 25774 24188 25780 24200
rect 25700 24160 25780 24188
rect 24026 24080 24032 24132
rect 24084 24080 24090 24132
rect 21284 24024 22968 24052
rect 23198 24012 23204 24064
rect 23256 24012 23262 24064
rect 23934 24012 23940 24064
rect 23992 24052 23998 24064
rect 24121 24055 24179 24061
rect 24121 24052 24133 24055
rect 23992 24024 24133 24052
rect 23992 24012 23998 24024
rect 24121 24021 24133 24024
rect 24167 24052 24179 24055
rect 25700 24052 25728 24160
rect 25774 24148 25780 24160
rect 25832 24148 25838 24200
rect 26237 24191 26295 24197
rect 26237 24157 26249 24191
rect 26283 24188 26295 24191
rect 26283 24160 26372 24188
rect 26283 24157 26295 24160
rect 26237 24151 26295 24157
rect 24167 24024 25728 24052
rect 25777 24055 25835 24061
rect 24167 24021 24179 24024
rect 24121 24015 24179 24021
rect 25777 24021 25789 24055
rect 25823 24052 25835 24055
rect 26050 24052 26056 24064
rect 25823 24024 26056 24052
rect 25823 24021 25835 24024
rect 25777 24015 25835 24021
rect 26050 24012 26056 24024
rect 26108 24012 26114 24064
rect 26344 24061 26372 24160
rect 26694 24148 26700 24200
rect 26752 24148 26758 24200
rect 26789 24191 26847 24197
rect 26789 24157 26801 24191
rect 26835 24188 26847 24191
rect 26835 24160 27016 24188
rect 26835 24157 26847 24160
rect 26789 24151 26847 24157
rect 26602 24080 26608 24132
rect 26660 24120 26666 24132
rect 26988 24120 27016 24160
rect 27062 24148 27068 24200
rect 27120 24188 27126 24200
rect 27341 24191 27399 24197
rect 27341 24188 27353 24191
rect 27120 24160 27353 24188
rect 27120 24148 27126 24160
rect 27341 24157 27353 24160
rect 27387 24157 27399 24191
rect 27341 24151 27399 24157
rect 27617 24191 27675 24197
rect 27617 24157 27629 24191
rect 27663 24188 27675 24191
rect 27798 24188 27804 24200
rect 27663 24160 27804 24188
rect 27663 24157 27675 24160
rect 27617 24151 27675 24157
rect 27798 24148 27804 24160
rect 27856 24148 27862 24200
rect 28350 24148 28356 24200
rect 28408 24148 28414 24200
rect 28626 24148 28632 24200
rect 28684 24148 28690 24200
rect 29730 24148 29736 24200
rect 29788 24148 29794 24200
rect 29822 24148 29828 24200
rect 29880 24148 29886 24200
rect 29932 24188 29960 24228
rect 30466 24216 30472 24268
rect 30524 24256 30530 24268
rect 30834 24256 30840 24268
rect 30524 24228 30840 24256
rect 30524 24216 30530 24228
rect 30834 24216 30840 24228
rect 30892 24216 30898 24268
rect 31386 24216 31392 24268
rect 31444 24216 31450 24268
rect 34238 24216 34244 24268
rect 34296 24216 34302 24268
rect 35360 24265 35388 24296
rect 37826 24284 37832 24336
rect 37884 24324 37890 24336
rect 38562 24324 38568 24336
rect 37884 24296 38568 24324
rect 37884 24284 37890 24296
rect 38562 24284 38568 24296
rect 38620 24324 38626 24336
rect 38620 24296 38792 24324
rect 38620 24284 38626 24296
rect 35345 24259 35403 24265
rect 35345 24225 35357 24259
rect 35391 24225 35403 24259
rect 35345 24219 35403 24225
rect 30101 24191 30159 24197
rect 30101 24188 30113 24191
rect 29932 24160 30113 24188
rect 30101 24157 30113 24160
rect 30147 24157 30159 24191
rect 30101 24151 30159 24157
rect 31202 24148 31208 24200
rect 31260 24148 31266 24200
rect 31754 24148 31760 24200
rect 31812 24188 31818 24200
rect 32214 24197 32220 24200
rect 31941 24191 31999 24197
rect 31941 24188 31953 24191
rect 31812 24160 31953 24188
rect 31812 24148 31818 24160
rect 31941 24157 31953 24160
rect 31987 24157 31999 24191
rect 32208 24188 32220 24197
rect 32175 24160 32220 24188
rect 31941 24151 31999 24157
rect 32208 24151 32220 24160
rect 32214 24148 32220 24151
rect 32272 24148 32278 24200
rect 33502 24148 33508 24200
rect 33560 24188 33566 24200
rect 33870 24188 33876 24200
rect 33560 24160 33876 24188
rect 33560 24148 33566 24160
rect 33870 24148 33876 24160
rect 33928 24148 33934 24200
rect 33965 24191 34023 24197
rect 33965 24157 33977 24191
rect 34011 24188 34023 24191
rect 34514 24188 34520 24200
rect 34011 24160 34520 24188
rect 34011 24157 34023 24160
rect 33965 24151 34023 24157
rect 27522 24120 27528 24132
rect 26660 24092 26924 24120
rect 26988 24092 27528 24120
rect 26660 24080 26666 24092
rect 26329 24055 26387 24061
rect 26329 24021 26341 24055
rect 26375 24021 26387 24055
rect 26896 24052 26924 24092
rect 27522 24080 27528 24092
rect 27580 24080 27586 24132
rect 29546 24080 29552 24132
rect 29604 24080 29610 24132
rect 31220 24120 31248 24148
rect 34348 24132 34376 24160
rect 34514 24148 34520 24160
rect 34572 24148 34578 24200
rect 31297 24123 31355 24129
rect 31297 24120 31309 24123
rect 31220 24092 31309 24120
rect 31297 24089 31309 24092
rect 31343 24089 31355 24123
rect 34146 24120 34152 24132
rect 31297 24083 31355 24089
rect 33336 24092 34152 24120
rect 29273 24055 29331 24061
rect 29273 24052 29285 24055
rect 26896 24024 29285 24052
rect 26329 24015 26387 24021
rect 29273 24021 29285 24024
rect 29319 24021 29331 24055
rect 29273 24015 29331 24021
rect 29362 24012 29368 24064
rect 29420 24052 29426 24064
rect 31205 24055 31263 24061
rect 31205 24052 31217 24055
rect 29420 24024 31217 24052
rect 29420 24012 29426 24024
rect 31205 24021 31217 24024
rect 31251 24052 31263 24055
rect 31662 24052 31668 24064
rect 31251 24024 31668 24052
rect 31251 24021 31263 24024
rect 31205 24015 31263 24021
rect 31662 24012 31668 24024
rect 31720 24012 31726 24064
rect 32766 24012 32772 24064
rect 32824 24052 32830 24064
rect 33336 24061 33364 24092
rect 34146 24080 34152 24092
rect 34204 24080 34210 24132
rect 34330 24080 34336 24132
rect 34388 24080 34394 24132
rect 35360 24120 35388 24219
rect 36446 24216 36452 24268
rect 36504 24256 36510 24268
rect 36722 24256 36728 24268
rect 36504 24228 36728 24256
rect 36504 24216 36510 24228
rect 36722 24216 36728 24228
rect 36780 24256 36786 24268
rect 36780 24228 36952 24256
rect 36780 24216 36786 24228
rect 35434 24148 35440 24200
rect 35492 24188 35498 24200
rect 35601 24191 35659 24197
rect 35601 24188 35613 24191
rect 35492 24160 35613 24188
rect 35492 24148 35498 24160
rect 35601 24157 35613 24160
rect 35647 24157 35659 24191
rect 36817 24191 36875 24197
rect 36817 24188 36829 24191
rect 35601 24151 35659 24157
rect 36372 24160 36829 24188
rect 36372 24132 36400 24160
rect 36817 24157 36829 24160
rect 36863 24157 36875 24191
rect 36924 24188 36952 24228
rect 36924 24160 37228 24188
rect 36817 24151 36875 24157
rect 36354 24120 36360 24132
rect 35360 24092 36360 24120
rect 36354 24080 36360 24092
rect 36412 24080 36418 24132
rect 36630 24080 36636 24132
rect 36688 24120 36694 24132
rect 37062 24123 37120 24129
rect 37062 24120 37074 24123
rect 36688 24092 37074 24120
rect 36688 24080 36694 24092
rect 37062 24089 37074 24092
rect 37108 24089 37120 24123
rect 37200 24120 37228 24160
rect 38286 24148 38292 24200
rect 38344 24148 38350 24200
rect 38470 24197 38476 24200
rect 38437 24191 38476 24197
rect 38437 24157 38449 24191
rect 38437 24151 38476 24157
rect 38470 24148 38476 24151
rect 38528 24148 38534 24200
rect 38764 24197 38792 24296
rect 38657 24191 38715 24197
rect 38657 24157 38669 24191
rect 38703 24157 38715 24191
rect 38657 24151 38715 24157
rect 38754 24191 38812 24197
rect 38754 24157 38766 24191
rect 38800 24157 38812 24191
rect 38754 24151 38812 24157
rect 38565 24123 38623 24129
rect 38565 24120 38577 24123
rect 37200 24092 38577 24120
rect 37062 24083 37120 24089
rect 38565 24089 38577 24092
rect 38611 24089 38623 24123
rect 38672 24120 38700 24151
rect 38856 24120 38884 24364
rect 39485 24361 39497 24395
rect 39531 24392 39543 24395
rect 40221 24395 40279 24401
rect 40221 24392 40233 24395
rect 39531 24364 40233 24392
rect 39531 24361 39543 24364
rect 39485 24355 39543 24361
rect 40221 24361 40233 24364
rect 40267 24361 40279 24395
rect 40221 24355 40279 24361
rect 41506 24352 41512 24404
rect 41564 24392 41570 24404
rect 42429 24395 42487 24401
rect 42429 24392 42441 24395
rect 41564 24364 42441 24392
rect 41564 24352 41570 24364
rect 42429 24361 42441 24364
rect 42475 24361 42487 24395
rect 46385 24395 46443 24401
rect 46385 24392 46397 24395
rect 42429 24355 42487 24361
rect 42536 24364 46397 24392
rect 41877 24327 41935 24333
rect 41877 24293 41889 24327
rect 41923 24324 41935 24327
rect 42150 24324 42156 24336
rect 41923 24296 42156 24324
rect 41923 24293 41935 24296
rect 41877 24287 41935 24293
rect 42150 24284 42156 24296
rect 42208 24324 42214 24336
rect 42245 24327 42303 24333
rect 42245 24324 42257 24327
rect 42208 24296 42257 24324
rect 42208 24284 42214 24296
rect 42245 24293 42257 24296
rect 42291 24293 42303 24327
rect 42536 24324 42564 24364
rect 46385 24361 46397 24364
rect 46431 24361 46443 24395
rect 46385 24355 46443 24361
rect 44450 24324 44456 24336
rect 42245 24287 42303 24293
rect 42352 24296 42564 24324
rect 42628 24296 44456 24324
rect 39853 24259 39911 24265
rect 39853 24225 39865 24259
rect 39899 24256 39911 24259
rect 42352 24256 42380 24296
rect 39899 24228 42380 24256
rect 39899 24225 39911 24228
rect 39853 24219 39911 24225
rect 42426 24216 42432 24268
rect 42484 24216 42490 24268
rect 42518 24216 42524 24268
rect 42576 24216 42582 24268
rect 39209 24191 39267 24197
rect 39209 24157 39221 24191
rect 39255 24188 39267 24191
rect 39298 24188 39304 24200
rect 39255 24160 39304 24188
rect 39255 24157 39267 24160
rect 39209 24151 39267 24157
rect 39298 24148 39304 24160
rect 39356 24148 39362 24200
rect 40034 24148 40040 24200
rect 40092 24148 40098 24200
rect 41598 24148 41604 24200
rect 41656 24188 41662 24200
rect 41693 24191 41751 24197
rect 41693 24188 41705 24191
rect 41656 24160 41705 24188
rect 41656 24148 41662 24160
rect 41693 24157 41705 24160
rect 41739 24157 41751 24191
rect 41693 24151 41751 24157
rect 41785 24191 41843 24197
rect 41785 24157 41797 24191
rect 41831 24188 41843 24191
rect 41874 24188 41880 24200
rect 41831 24160 41880 24188
rect 41831 24157 41843 24160
rect 41785 24151 41843 24157
rect 41874 24148 41880 24160
rect 41932 24148 41938 24200
rect 41966 24148 41972 24200
rect 42024 24148 42030 24200
rect 42153 24191 42211 24197
rect 42153 24157 42165 24191
rect 42199 24157 42211 24191
rect 42153 24151 42211 24157
rect 38672 24092 38884 24120
rect 38565 24083 38623 24089
rect 42168 24064 42196 24151
rect 42536 24120 42564 24216
rect 42628 24197 42656 24296
rect 42613 24191 42671 24197
rect 42613 24157 42625 24191
rect 42659 24157 42671 24191
rect 43070 24188 43076 24200
rect 42613 24151 42671 24157
rect 42716 24160 43076 24188
rect 42716 24120 42744 24160
rect 43070 24148 43076 24160
rect 43128 24148 43134 24200
rect 43180 24197 43208 24296
rect 44450 24284 44456 24296
rect 44508 24284 44514 24336
rect 45649 24327 45707 24333
rect 45649 24293 45661 24327
rect 45695 24293 45707 24327
rect 45649 24287 45707 24293
rect 43346 24216 43352 24268
rect 43404 24216 43410 24268
rect 45664 24256 45692 24287
rect 45922 24256 45928 24268
rect 45664 24228 45928 24256
rect 45922 24216 45928 24228
rect 45980 24216 45986 24268
rect 46658 24256 46664 24268
rect 46124 24228 46664 24256
rect 43165 24191 43223 24197
rect 43165 24157 43177 24191
rect 43211 24157 43223 24191
rect 43165 24151 43223 24157
rect 43254 24148 43260 24200
rect 43312 24148 43318 24200
rect 44910 24148 44916 24200
rect 44968 24188 44974 24200
rect 45005 24191 45063 24197
rect 45005 24188 45017 24191
rect 44968 24160 45017 24188
rect 44968 24148 44974 24160
rect 45005 24157 45017 24160
rect 45051 24157 45063 24191
rect 45005 24151 45063 24157
rect 45186 24148 45192 24200
rect 45244 24148 45250 24200
rect 45373 24191 45431 24197
rect 45373 24157 45385 24191
rect 45419 24188 45431 24191
rect 45554 24188 45560 24200
rect 45419 24160 45560 24188
rect 45419 24157 45431 24160
rect 45373 24151 45431 24157
rect 45554 24148 45560 24160
rect 45612 24188 45618 24200
rect 45741 24191 45799 24197
rect 45741 24188 45753 24191
rect 45612 24160 45753 24188
rect 45612 24148 45618 24160
rect 45741 24157 45753 24160
rect 45787 24157 45799 24191
rect 45741 24151 45799 24157
rect 45833 24191 45891 24197
rect 45833 24157 45845 24191
rect 45879 24157 45891 24191
rect 45833 24151 45891 24157
rect 42536 24092 42744 24120
rect 42889 24123 42947 24129
rect 42889 24089 42901 24123
rect 42935 24120 42947 24123
rect 43530 24120 43536 24132
rect 42935 24092 43536 24120
rect 42935 24089 42947 24092
rect 42889 24083 42947 24089
rect 43530 24080 43536 24092
rect 43588 24080 43594 24132
rect 45462 24080 45468 24132
rect 45520 24080 45526 24132
rect 45646 24080 45652 24132
rect 45704 24120 45710 24132
rect 45848 24120 45876 24151
rect 46014 24148 46020 24200
rect 46072 24148 46078 24200
rect 46124 24197 46152 24228
rect 46658 24216 46664 24228
rect 46716 24216 46722 24268
rect 46109 24191 46167 24197
rect 46109 24157 46121 24191
rect 46155 24157 46167 24191
rect 46109 24151 46167 24157
rect 46385 24191 46443 24197
rect 46385 24157 46397 24191
rect 46431 24157 46443 24191
rect 46385 24151 46443 24157
rect 45704 24092 45876 24120
rect 45704 24080 45710 24092
rect 45922 24080 45928 24132
rect 45980 24120 45986 24132
rect 46293 24123 46351 24129
rect 46293 24120 46305 24123
rect 45980 24092 46305 24120
rect 45980 24080 45986 24092
rect 46293 24089 46305 24092
rect 46339 24089 46351 24123
rect 46293 24083 46351 24089
rect 33321 24055 33379 24061
rect 33321 24052 33333 24055
rect 32824 24024 33333 24052
rect 32824 24012 32830 24024
rect 33321 24021 33333 24024
rect 33367 24021 33379 24055
rect 33321 24015 33379 24021
rect 34057 24055 34115 24061
rect 34057 24021 34069 24055
rect 34103 24052 34115 24055
rect 34698 24052 34704 24064
rect 34103 24024 34704 24052
rect 34103 24021 34115 24024
rect 34057 24015 34115 24021
rect 34698 24012 34704 24024
rect 34756 24052 34762 24064
rect 35434 24052 35440 24064
rect 34756 24024 35440 24052
rect 34756 24012 34762 24024
rect 35434 24012 35440 24024
rect 35492 24012 35498 24064
rect 36078 24012 36084 24064
rect 36136 24052 36142 24064
rect 36725 24055 36783 24061
rect 36725 24052 36737 24055
rect 36136 24024 36737 24052
rect 36136 24012 36142 24024
rect 36725 24021 36737 24024
rect 36771 24021 36783 24055
rect 36725 24015 36783 24021
rect 36814 24012 36820 24064
rect 36872 24052 36878 24064
rect 38197 24055 38255 24061
rect 38197 24052 38209 24055
rect 36872 24024 38209 24052
rect 36872 24012 36878 24024
rect 38197 24021 38209 24024
rect 38243 24021 38255 24055
rect 38197 24015 38255 24021
rect 38378 24012 38384 24064
rect 38436 24052 38442 24064
rect 38933 24055 38991 24061
rect 38933 24052 38945 24055
rect 38436 24024 38945 24052
rect 38436 24012 38442 24024
rect 38933 24021 38945 24024
rect 38979 24021 38991 24055
rect 38933 24015 38991 24021
rect 39669 24055 39727 24061
rect 39669 24021 39681 24055
rect 39715 24052 39727 24055
rect 39758 24052 39764 24064
rect 39715 24024 39764 24052
rect 39715 24021 39727 24024
rect 39669 24015 39727 24021
rect 39758 24012 39764 24024
rect 39816 24012 39822 24064
rect 40586 24012 40592 24064
rect 40644 24052 40650 24064
rect 41509 24055 41567 24061
rect 41509 24052 41521 24055
rect 40644 24024 41521 24052
rect 40644 24012 40650 24024
rect 41509 24021 41521 24024
rect 41555 24021 41567 24055
rect 41509 24015 41567 24021
rect 42150 24012 42156 24064
rect 42208 24012 42214 24064
rect 45557 24055 45615 24061
rect 45557 24021 45569 24055
rect 45603 24052 45615 24055
rect 46400 24052 46428 24151
rect 46566 24148 46572 24200
rect 46624 24148 46630 24200
rect 45603 24024 46428 24052
rect 45603 24021 45615 24024
rect 45557 24015 45615 24021
rect 1104 23962 47104 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 47104 23962
rect 1104 23888 47104 23910
rect 11514 23808 11520 23860
rect 11572 23848 11578 23860
rect 12345 23851 12403 23857
rect 12345 23848 12357 23851
rect 11572 23820 12357 23848
rect 11572 23808 11578 23820
rect 12345 23817 12357 23820
rect 12391 23848 12403 23851
rect 12529 23851 12587 23857
rect 12529 23848 12541 23851
rect 12391 23820 12541 23848
rect 12391 23817 12403 23820
rect 12345 23811 12403 23817
rect 12529 23817 12541 23820
rect 12575 23817 12587 23851
rect 12529 23811 12587 23817
rect 12894 23808 12900 23860
rect 12952 23848 12958 23860
rect 13541 23851 13599 23857
rect 13541 23848 13553 23851
rect 12952 23820 13553 23848
rect 12952 23808 12958 23820
rect 13541 23817 13553 23820
rect 13587 23848 13599 23851
rect 13587 23820 15332 23848
rect 13587 23817 13599 23820
rect 13541 23811 13599 23817
rect 13992 23783 14050 23789
rect 13992 23749 14004 23783
rect 14038 23780 14050 23783
rect 15304 23780 15332 23820
rect 15930 23808 15936 23860
rect 15988 23848 15994 23860
rect 16669 23851 16727 23857
rect 16669 23848 16681 23851
rect 15988 23820 16681 23848
rect 15988 23808 15994 23820
rect 16669 23817 16681 23820
rect 16715 23817 16727 23851
rect 16669 23811 16727 23817
rect 17037 23851 17095 23857
rect 17037 23817 17049 23851
rect 17083 23848 17095 23851
rect 17402 23848 17408 23860
rect 17083 23820 17408 23848
rect 17083 23817 17095 23820
rect 17037 23811 17095 23817
rect 17402 23808 17408 23820
rect 17460 23808 17466 23860
rect 18782 23848 18788 23860
rect 17512 23820 18788 23848
rect 17512 23780 17540 23820
rect 18782 23808 18788 23820
rect 18840 23808 18846 23860
rect 19518 23808 19524 23860
rect 19576 23848 19582 23860
rect 23106 23848 23112 23860
rect 19576 23820 23112 23848
rect 19576 23808 19582 23820
rect 23106 23808 23112 23820
rect 23164 23808 23170 23860
rect 23198 23808 23204 23860
rect 23256 23848 23262 23860
rect 23256 23820 24900 23848
rect 23256 23808 23262 23820
rect 14038 23752 14780 23780
rect 15304 23752 17540 23780
rect 14038 23749 14050 23752
rect 13992 23743 14050 23749
rect 2409 23715 2467 23721
rect 2409 23681 2421 23715
rect 2455 23712 2467 23715
rect 3234 23712 3240 23724
rect 2455 23684 3240 23712
rect 2455 23681 2467 23684
rect 2409 23675 2467 23681
rect 3234 23672 3240 23684
rect 3292 23672 3298 23724
rect 5534 23672 5540 23724
rect 5592 23672 5598 23724
rect 9122 23672 9128 23724
rect 9180 23672 9186 23724
rect 10962 23672 10968 23724
rect 11020 23712 11026 23724
rect 12158 23712 12164 23724
rect 11020 23684 12164 23712
rect 11020 23672 11026 23684
rect 12158 23672 12164 23684
rect 12216 23712 12222 23724
rect 12253 23715 12311 23721
rect 12253 23712 12265 23715
rect 12216 23684 12265 23712
rect 12216 23672 12222 23684
rect 12253 23681 12265 23684
rect 12299 23681 12311 23715
rect 12253 23675 12311 23681
rect 12434 23672 12440 23724
rect 12492 23712 12498 23724
rect 12986 23712 12992 23724
rect 12492 23684 12992 23712
rect 12492 23672 12498 23684
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 13354 23672 13360 23724
rect 13412 23672 13418 23724
rect 13630 23672 13636 23724
rect 13688 23712 13694 23724
rect 13725 23715 13783 23721
rect 13725 23712 13737 23715
rect 13688 23684 13737 23712
rect 13688 23672 13694 23684
rect 13725 23681 13737 23684
rect 13771 23681 13783 23715
rect 13725 23675 13783 23681
rect 4341 23647 4399 23653
rect 4341 23613 4353 23647
rect 4387 23613 4399 23647
rect 4341 23607 4399 23613
rect 4525 23647 4583 23653
rect 4525 23613 4537 23647
rect 4571 23644 4583 23647
rect 5074 23644 5080 23656
rect 4571 23616 5080 23644
rect 4571 23613 4583 23616
rect 4525 23607 4583 23613
rect 4356 23576 4384 23607
rect 5074 23604 5080 23616
rect 5132 23604 5138 23656
rect 5258 23604 5264 23656
rect 5316 23604 5322 23656
rect 5399 23647 5457 23653
rect 5399 23613 5411 23647
rect 5445 23644 5457 23647
rect 5718 23644 5724 23656
rect 5445 23616 5724 23644
rect 5445 23613 5457 23616
rect 5399 23607 5457 23613
rect 5718 23604 5724 23616
rect 5776 23604 5782 23656
rect 6178 23604 6184 23656
rect 6236 23604 6242 23656
rect 9214 23604 9220 23656
rect 9272 23604 9278 23656
rect 9306 23604 9312 23656
rect 9364 23604 9370 23656
rect 12894 23604 12900 23656
rect 12952 23604 12958 23656
rect 14752 23644 14780 23752
rect 17586 23740 17592 23792
rect 17644 23740 17650 23792
rect 19426 23740 19432 23792
rect 19484 23780 19490 23792
rect 19794 23780 19800 23792
rect 19484 23752 19800 23780
rect 19484 23740 19490 23752
rect 19794 23740 19800 23752
rect 19852 23740 19858 23792
rect 20806 23780 20812 23792
rect 19904 23752 20812 23780
rect 15010 23672 15016 23724
rect 15068 23712 15074 23724
rect 15068 23684 15332 23712
rect 15068 23672 15074 23684
rect 15304 23644 15332 23684
rect 15378 23672 15384 23724
rect 15436 23672 15442 23724
rect 15470 23672 15476 23724
rect 15528 23712 15534 23724
rect 18509 23715 18567 23721
rect 18509 23712 18521 23715
rect 15528 23684 18521 23712
rect 15528 23672 15534 23684
rect 18509 23681 18521 23684
rect 18555 23712 18567 23715
rect 19904 23712 19932 23752
rect 20806 23740 20812 23752
rect 20864 23740 20870 23792
rect 20898 23740 20904 23792
rect 20956 23780 20962 23792
rect 20956 23752 21404 23780
rect 20956 23740 20962 23752
rect 18555 23684 19932 23712
rect 18555 23681 18567 23684
rect 18509 23675 18567 23681
rect 19978 23672 19984 23724
rect 20036 23672 20042 23724
rect 21082 23672 21088 23724
rect 21140 23672 21146 23724
rect 21266 23672 21272 23724
rect 21324 23672 21330 23724
rect 21376 23721 21404 23752
rect 21450 23740 21456 23792
rect 21508 23780 21514 23792
rect 24026 23780 24032 23792
rect 21508 23752 24032 23780
rect 21508 23740 21514 23752
rect 24026 23740 24032 23752
rect 24084 23780 24090 23792
rect 24765 23783 24823 23789
rect 24765 23780 24777 23783
rect 24084 23752 24777 23780
rect 24084 23740 24090 23752
rect 24765 23749 24777 23752
rect 24811 23749 24823 23783
rect 24872 23780 24900 23820
rect 25222 23808 25228 23860
rect 25280 23808 25286 23860
rect 27062 23808 27068 23860
rect 27120 23808 27126 23860
rect 29086 23848 29092 23860
rect 27172 23820 29092 23848
rect 27172 23780 27200 23820
rect 29086 23808 29092 23820
rect 29144 23808 29150 23860
rect 29638 23808 29644 23860
rect 29696 23848 29702 23860
rect 29733 23851 29791 23857
rect 29733 23848 29745 23851
rect 29696 23820 29745 23848
rect 29696 23808 29702 23820
rect 29733 23817 29745 23820
rect 29779 23817 29791 23851
rect 29733 23811 29791 23817
rect 32398 23808 32404 23860
rect 32456 23808 32462 23860
rect 32766 23808 32772 23860
rect 32824 23808 32830 23860
rect 33594 23808 33600 23860
rect 33652 23848 33658 23860
rect 34606 23848 34612 23860
rect 33652 23820 34612 23848
rect 33652 23808 33658 23820
rect 34606 23808 34612 23820
rect 34664 23808 34670 23860
rect 35250 23808 35256 23860
rect 35308 23808 35314 23860
rect 35342 23808 35348 23860
rect 35400 23808 35406 23860
rect 35434 23808 35440 23860
rect 35492 23848 35498 23860
rect 35805 23851 35863 23857
rect 35805 23848 35817 23851
rect 35492 23820 35817 23848
rect 35492 23808 35498 23820
rect 35805 23817 35817 23820
rect 35851 23817 35863 23851
rect 35805 23811 35863 23817
rect 38286 23808 38292 23860
rect 38344 23848 38350 23860
rect 40221 23851 40279 23857
rect 40221 23848 40233 23851
rect 38344 23820 40233 23848
rect 38344 23808 38350 23820
rect 40221 23817 40233 23820
rect 40267 23817 40279 23851
rect 40221 23811 40279 23817
rect 41417 23851 41475 23857
rect 41417 23817 41429 23851
rect 41463 23848 41475 23851
rect 41785 23851 41843 23857
rect 41785 23848 41797 23851
rect 41463 23820 41797 23848
rect 41463 23817 41475 23820
rect 41417 23811 41475 23817
rect 41785 23817 41797 23820
rect 41831 23848 41843 23851
rect 42150 23848 42156 23860
rect 41831 23820 42156 23848
rect 41831 23817 41843 23820
rect 41785 23811 41843 23817
rect 42150 23808 42156 23820
rect 42208 23808 42214 23860
rect 42334 23808 42340 23860
rect 42392 23848 42398 23860
rect 42613 23851 42671 23857
rect 42613 23848 42625 23851
rect 42392 23820 42625 23848
rect 42392 23808 42398 23820
rect 42613 23817 42625 23820
rect 42659 23817 42671 23851
rect 42613 23811 42671 23817
rect 43070 23808 43076 23860
rect 43128 23848 43134 23860
rect 43990 23848 43996 23860
rect 43128 23820 43996 23848
rect 43128 23808 43134 23820
rect 43990 23808 43996 23820
rect 44048 23808 44054 23860
rect 44450 23808 44456 23860
rect 44508 23848 44514 23860
rect 44545 23851 44603 23857
rect 44545 23848 44557 23851
rect 44508 23820 44557 23848
rect 44508 23808 44514 23820
rect 44545 23817 44557 23820
rect 44591 23817 44603 23851
rect 44545 23811 44603 23817
rect 45186 23808 45192 23860
rect 45244 23848 45250 23860
rect 46658 23848 46664 23860
rect 45244 23820 46664 23848
rect 45244 23808 45250 23820
rect 46658 23808 46664 23820
rect 46716 23808 46722 23860
rect 24872 23752 27200 23780
rect 27525 23783 27583 23789
rect 24765 23743 24823 23749
rect 27525 23749 27537 23783
rect 27571 23780 27583 23783
rect 27614 23780 27620 23792
rect 27571 23752 27620 23780
rect 27571 23749 27583 23752
rect 27525 23743 27583 23749
rect 27614 23740 27620 23752
rect 27672 23740 27678 23792
rect 31294 23740 31300 23792
rect 31352 23780 31358 23792
rect 32861 23783 32919 23789
rect 32861 23780 32873 23783
rect 31352 23752 32873 23780
rect 31352 23740 31358 23752
rect 32861 23749 32873 23752
rect 32907 23780 32919 23783
rect 33318 23780 33324 23792
rect 32907 23752 33324 23780
rect 32907 23749 32919 23752
rect 32861 23743 32919 23749
rect 33318 23740 33324 23752
rect 33376 23740 33382 23792
rect 39301 23783 39359 23789
rect 39301 23749 39313 23783
rect 39347 23780 39359 23783
rect 41233 23783 41291 23789
rect 39347 23752 40724 23780
rect 39347 23749 39359 23752
rect 39301 23743 39359 23749
rect 21361 23715 21419 23721
rect 21361 23681 21373 23715
rect 21407 23712 21419 23715
rect 21407 23684 21588 23712
rect 21407 23681 21419 23684
rect 21361 23675 21419 23681
rect 17129 23647 17187 23653
rect 17129 23644 17141 23647
rect 14752 23616 15240 23644
rect 15304 23616 17141 23644
rect 4890 23576 4896 23588
rect 4356 23548 4896 23576
rect 4890 23536 4896 23548
rect 4948 23536 4954 23588
rect 15212 23585 15240 23616
rect 17129 23613 17141 23616
rect 17175 23613 17187 23647
rect 17129 23607 17187 23613
rect 4985 23579 5043 23585
rect 4985 23545 4997 23579
rect 5031 23545 5043 23579
rect 4985 23539 5043 23545
rect 15197 23579 15255 23585
rect 15197 23545 15209 23579
rect 15243 23545 15255 23579
rect 17144 23576 17172 23607
rect 17218 23604 17224 23656
rect 17276 23604 17282 23656
rect 20438 23644 20444 23656
rect 18616 23616 20444 23644
rect 17773 23579 17831 23585
rect 17773 23576 17785 23579
rect 17144 23548 17785 23576
rect 15197 23539 15255 23545
rect 17773 23545 17785 23548
rect 17819 23545 17831 23579
rect 17773 23539 17831 23545
rect 2038 23468 2044 23520
rect 2096 23508 2102 23520
rect 2225 23511 2283 23517
rect 2225 23508 2237 23511
rect 2096 23480 2237 23508
rect 2096 23468 2102 23480
rect 2225 23477 2237 23480
rect 2271 23477 2283 23511
rect 2225 23471 2283 23477
rect 4522 23468 4528 23520
rect 4580 23508 4586 23520
rect 5000 23508 5028 23539
rect 4580 23480 5028 23508
rect 4580 23468 4586 23480
rect 5534 23468 5540 23520
rect 5592 23508 5598 23520
rect 8018 23508 8024 23520
rect 5592 23480 8024 23508
rect 5592 23468 5598 23480
rect 8018 23468 8024 23480
rect 8076 23468 8082 23520
rect 8754 23468 8760 23520
rect 8812 23468 8818 23520
rect 13170 23468 13176 23520
rect 13228 23468 13234 23520
rect 15102 23468 15108 23520
rect 15160 23508 15166 23520
rect 18616 23508 18644 23616
rect 20438 23604 20444 23616
rect 20496 23604 20502 23656
rect 21100 23644 21128 23672
rect 21450 23644 21456 23656
rect 21100 23616 21456 23644
rect 21450 23604 21456 23616
rect 21508 23604 21514 23656
rect 21560 23644 21588 23684
rect 21634 23672 21640 23724
rect 21692 23712 21698 23724
rect 23934 23712 23940 23724
rect 21692 23684 23940 23712
rect 21692 23672 21698 23684
rect 23934 23672 23940 23684
rect 23992 23672 23998 23724
rect 25593 23715 25651 23721
rect 25593 23681 25605 23715
rect 25639 23712 25651 23715
rect 26050 23712 26056 23724
rect 25639 23684 26056 23712
rect 25639 23681 25651 23684
rect 25593 23675 25651 23681
rect 26050 23672 26056 23684
rect 26108 23672 26114 23724
rect 27433 23715 27491 23721
rect 27433 23681 27445 23715
rect 27479 23712 27491 23715
rect 28258 23712 28264 23724
rect 27479 23684 28264 23712
rect 27479 23681 27491 23684
rect 27433 23675 27491 23681
rect 28258 23672 28264 23684
rect 28316 23672 28322 23724
rect 28902 23672 28908 23724
rect 28960 23721 28966 23724
rect 28960 23715 28988 23721
rect 28976 23681 28988 23715
rect 28960 23675 28988 23681
rect 28960 23672 28966 23675
rect 30466 23672 30472 23724
rect 30524 23672 30530 23724
rect 34330 23672 34336 23724
rect 34388 23672 34394 23724
rect 35713 23715 35771 23721
rect 35713 23681 35725 23715
rect 35759 23712 35771 23715
rect 36078 23712 36084 23724
rect 35759 23684 36084 23712
rect 35759 23681 35771 23684
rect 35713 23675 35771 23681
rect 21910 23644 21916 23656
rect 21560 23616 21916 23644
rect 21910 23604 21916 23616
rect 21968 23604 21974 23656
rect 25498 23644 25504 23656
rect 22066 23616 25504 23644
rect 18693 23579 18751 23585
rect 18693 23545 18705 23579
rect 18739 23576 18751 23579
rect 19242 23576 19248 23588
rect 18739 23548 19248 23576
rect 18739 23545 18751 23548
rect 18693 23539 18751 23545
rect 19242 23536 19248 23548
rect 19300 23576 19306 23588
rect 19702 23576 19708 23588
rect 19300 23548 19708 23576
rect 19300 23536 19306 23548
rect 19702 23536 19708 23548
rect 19760 23536 19766 23588
rect 19794 23536 19800 23588
rect 19852 23576 19858 23588
rect 20257 23579 20315 23585
rect 20257 23576 20269 23579
rect 19852 23548 20269 23576
rect 19852 23536 19858 23548
rect 20257 23545 20269 23548
rect 20303 23576 20315 23579
rect 20622 23576 20628 23588
rect 20303 23548 20628 23576
rect 20303 23545 20315 23548
rect 20257 23539 20315 23545
rect 20622 23536 20628 23548
rect 20680 23536 20686 23588
rect 20901 23579 20959 23585
rect 20901 23545 20913 23579
rect 20947 23576 20959 23579
rect 22066 23576 22094 23616
rect 25498 23604 25504 23616
rect 25556 23604 25562 23656
rect 25685 23647 25743 23653
rect 25685 23613 25697 23647
rect 25731 23613 25743 23647
rect 25685 23607 25743 23613
rect 25869 23647 25927 23653
rect 25869 23613 25881 23647
rect 25915 23613 25927 23647
rect 25869 23607 25927 23613
rect 27617 23647 27675 23653
rect 27617 23613 27629 23647
rect 27663 23613 27675 23647
rect 27617 23607 27675 23613
rect 25041 23579 25099 23585
rect 20947 23548 22094 23576
rect 24780 23548 24992 23576
rect 20947 23545 20959 23548
rect 20901 23539 20959 23545
rect 15160 23480 18644 23508
rect 15160 23468 15166 23480
rect 19518 23468 19524 23520
rect 19576 23508 19582 23520
rect 19978 23508 19984 23520
rect 19576 23480 19984 23508
rect 19576 23468 19582 23480
rect 19978 23468 19984 23480
rect 20036 23468 20042 23520
rect 20162 23468 20168 23520
rect 20220 23508 20226 23520
rect 24780 23508 24808 23548
rect 20220 23480 24808 23508
rect 24964 23508 24992 23548
rect 25041 23545 25053 23579
rect 25087 23576 25099 23579
rect 25222 23576 25228 23588
rect 25087 23548 25228 23576
rect 25087 23545 25099 23548
rect 25041 23539 25099 23545
rect 25222 23536 25228 23548
rect 25280 23536 25286 23588
rect 25590 23536 25596 23588
rect 25648 23576 25654 23588
rect 25700 23576 25728 23607
rect 25648 23548 25728 23576
rect 25884 23576 25912 23607
rect 27632 23576 27660 23607
rect 27706 23604 27712 23656
rect 27764 23644 27770 23656
rect 27893 23647 27951 23653
rect 27893 23644 27905 23647
rect 27764 23616 27905 23644
rect 27764 23604 27770 23616
rect 27893 23613 27905 23616
rect 27939 23644 27951 23647
rect 27982 23644 27988 23656
rect 27939 23616 27988 23644
rect 27939 23613 27951 23616
rect 27893 23607 27951 23613
rect 27982 23604 27988 23616
rect 28040 23604 28046 23656
rect 28077 23647 28135 23653
rect 28077 23613 28089 23647
rect 28123 23613 28135 23647
rect 28276 23644 28304 23672
rect 28813 23647 28871 23653
rect 28813 23644 28825 23647
rect 28276 23616 28825 23644
rect 28077 23607 28135 23613
rect 28813 23613 28825 23616
rect 28859 23613 28871 23647
rect 28813 23607 28871 23613
rect 25884 23548 27660 23576
rect 25648 23536 25654 23548
rect 27540 23520 27568 23548
rect 27798 23536 27804 23588
rect 27856 23576 27862 23588
rect 28092 23576 28120 23607
rect 29086 23604 29092 23656
rect 29144 23644 29150 23656
rect 29454 23644 29460 23656
rect 29144 23616 29460 23644
rect 29144 23604 29150 23616
rect 29454 23604 29460 23616
rect 29512 23604 29518 23656
rect 29822 23604 29828 23656
rect 29880 23644 29886 23656
rect 31386 23644 31392 23656
rect 29880 23616 31392 23644
rect 29880 23604 29886 23616
rect 31386 23604 31392 23616
rect 31444 23604 31450 23656
rect 33042 23604 33048 23656
rect 33100 23604 33106 23656
rect 33410 23604 33416 23656
rect 33468 23604 33474 23656
rect 33597 23647 33655 23653
rect 33597 23613 33609 23647
rect 33643 23613 33655 23647
rect 33597 23607 33655 23613
rect 27856 23548 28120 23576
rect 27856 23536 27862 23548
rect 27430 23508 27436 23520
rect 24964 23480 27436 23508
rect 20220 23468 20226 23480
rect 27430 23468 27436 23480
rect 27488 23468 27494 23520
rect 27522 23468 27528 23520
rect 27580 23468 27586 23520
rect 28092 23508 28120 23548
rect 28534 23536 28540 23588
rect 28592 23536 28598 23588
rect 31202 23576 31208 23588
rect 30116 23548 31208 23576
rect 30116 23508 30144 23548
rect 31202 23536 31208 23548
rect 31260 23536 31266 23588
rect 28092 23480 30144 23508
rect 30190 23468 30196 23520
rect 30248 23508 30254 23520
rect 30285 23511 30343 23517
rect 30285 23508 30297 23511
rect 30248 23480 30297 23508
rect 30248 23468 30254 23480
rect 30285 23477 30297 23480
rect 30331 23477 30343 23511
rect 33428 23508 33456 23604
rect 33612 23576 33640 23607
rect 34146 23604 34152 23656
rect 34204 23644 34210 23656
rect 34450 23647 34508 23653
rect 34450 23644 34462 23647
rect 34204 23616 34462 23644
rect 34204 23604 34210 23616
rect 34450 23613 34462 23616
rect 34496 23613 34508 23647
rect 34450 23607 34508 23613
rect 34606 23604 34612 23656
rect 34664 23604 34670 23656
rect 35728 23644 35756 23675
rect 36078 23672 36084 23684
rect 36136 23672 36142 23724
rect 36173 23715 36231 23721
rect 36173 23681 36185 23715
rect 36219 23712 36231 23715
rect 36538 23712 36544 23724
rect 36219 23684 36544 23712
rect 36219 23681 36231 23684
rect 36173 23675 36231 23681
rect 36538 23672 36544 23684
rect 36596 23672 36602 23724
rect 38102 23672 38108 23724
rect 38160 23672 38166 23724
rect 38286 23672 38292 23724
rect 38344 23712 38350 23724
rect 38381 23715 38439 23721
rect 38381 23712 38393 23715
rect 38344 23684 38393 23712
rect 38344 23672 38350 23684
rect 38381 23681 38393 23684
rect 38427 23681 38439 23715
rect 38381 23675 38439 23681
rect 39482 23672 39488 23724
rect 39540 23672 39546 23724
rect 39758 23672 39764 23724
rect 39816 23672 39822 23724
rect 39942 23672 39948 23724
rect 40000 23672 40006 23724
rect 40405 23715 40463 23721
rect 40405 23681 40417 23715
rect 40451 23712 40463 23715
rect 40494 23712 40500 23724
rect 40451 23684 40500 23712
rect 40451 23681 40463 23684
rect 40405 23675 40463 23681
rect 40494 23672 40500 23684
rect 40552 23672 40558 23724
rect 40586 23672 40592 23724
rect 40644 23672 40650 23724
rect 40696 23721 40724 23752
rect 41233 23749 41245 23783
rect 41279 23780 41291 23783
rect 41874 23780 41880 23792
rect 41279 23752 41880 23780
rect 41279 23749 41291 23752
rect 41233 23743 41291 23749
rect 41874 23740 41880 23752
rect 41932 23740 41938 23792
rect 42429 23783 42487 23789
rect 42429 23749 42441 23783
rect 42475 23780 42487 23783
rect 42794 23780 42800 23792
rect 42475 23752 42800 23780
rect 42475 23749 42487 23752
rect 42429 23743 42487 23749
rect 42794 23740 42800 23752
rect 42852 23780 42858 23792
rect 43346 23780 43352 23792
rect 42852 23752 43352 23780
rect 42852 23740 42858 23752
rect 43346 23740 43352 23752
rect 43404 23740 43410 23792
rect 45462 23740 45468 23792
rect 45520 23780 45526 23792
rect 45520 23752 45600 23780
rect 45520 23740 45526 23752
rect 40681 23715 40739 23721
rect 40681 23681 40693 23715
rect 40727 23681 40739 23715
rect 40681 23675 40739 23681
rect 41414 23672 41420 23724
rect 41472 23712 41478 23724
rect 41509 23715 41567 23721
rect 41509 23712 41521 23715
rect 41472 23684 41521 23712
rect 41472 23672 41478 23684
rect 41509 23681 41521 23684
rect 41555 23681 41567 23715
rect 41509 23675 41567 23681
rect 41598 23672 41604 23724
rect 41656 23672 41662 23724
rect 41690 23672 41696 23724
rect 41748 23712 41754 23724
rect 41785 23715 41843 23721
rect 41785 23712 41797 23715
rect 41748 23684 41797 23712
rect 41748 23672 41754 23684
rect 41785 23681 41797 23684
rect 41831 23681 41843 23715
rect 41785 23675 41843 23681
rect 42705 23715 42763 23721
rect 42705 23681 42717 23715
rect 42751 23712 42763 23715
rect 42751 23684 42840 23712
rect 42751 23681 42763 23684
rect 42705 23675 42763 23681
rect 34992 23616 35756 23644
rect 35897 23647 35955 23653
rect 33778 23576 33784 23588
rect 33612 23548 33784 23576
rect 33778 23536 33784 23548
rect 33836 23536 33842 23588
rect 33870 23536 33876 23588
rect 33928 23576 33934 23588
rect 34057 23579 34115 23585
rect 34057 23576 34069 23579
rect 33928 23548 34069 23576
rect 33928 23536 33934 23548
rect 34057 23545 34069 23548
rect 34103 23545 34115 23579
rect 34057 23539 34115 23545
rect 34992 23508 35020 23616
rect 35897 23613 35909 23647
rect 35943 23613 35955 23647
rect 35897 23607 35955 23613
rect 35342 23536 35348 23588
rect 35400 23576 35406 23588
rect 35912 23576 35940 23607
rect 36354 23604 36360 23656
rect 36412 23644 36418 23656
rect 36449 23647 36507 23653
rect 36449 23644 36461 23647
rect 36412 23616 36461 23644
rect 36412 23604 36418 23616
rect 36449 23613 36461 23616
rect 36495 23613 36507 23647
rect 41616 23644 41644 23672
rect 42812 23644 42840 23684
rect 43714 23672 43720 23724
rect 43772 23672 43778 23724
rect 43901 23715 43959 23721
rect 43901 23712 43913 23715
rect 43824 23684 43913 23712
rect 43070 23644 43076 23656
rect 36449 23607 36507 23613
rect 39132 23616 41558 23644
rect 41616 23616 42564 23644
rect 42812 23616 43076 23644
rect 35400 23548 35940 23576
rect 35400 23536 35406 23548
rect 36538 23536 36544 23588
rect 36596 23576 36602 23588
rect 37366 23576 37372 23588
rect 36596 23548 37372 23576
rect 36596 23536 36602 23548
rect 37366 23536 37372 23548
rect 37424 23536 37430 23588
rect 39132 23585 39160 23616
rect 39117 23579 39175 23585
rect 39117 23545 39129 23579
rect 39163 23545 39175 23579
rect 39117 23539 39175 23545
rect 39390 23536 39396 23588
rect 39448 23576 39454 23588
rect 39577 23579 39635 23585
rect 39577 23576 39589 23579
rect 39448 23548 39589 23576
rect 39448 23536 39454 23548
rect 39577 23545 39589 23548
rect 39623 23545 39635 23579
rect 39577 23539 39635 23545
rect 39669 23579 39727 23585
rect 39669 23545 39681 23579
rect 39715 23576 39727 23579
rect 39758 23576 39764 23588
rect 39715 23548 39764 23576
rect 39715 23545 39727 23548
rect 39669 23539 39727 23545
rect 39758 23536 39764 23548
rect 39816 23536 39822 23588
rect 40497 23579 40555 23585
rect 40497 23545 40509 23579
rect 40543 23545 40555 23579
rect 40497 23539 40555 23545
rect 33428 23480 35020 23508
rect 30285 23471 30343 23477
rect 39298 23468 39304 23520
rect 39356 23508 39362 23520
rect 39942 23508 39948 23520
rect 39356 23480 39948 23508
rect 39356 23468 39362 23480
rect 39942 23468 39948 23480
rect 40000 23468 40006 23520
rect 40512 23508 40540 23539
rect 41233 23511 41291 23517
rect 41233 23508 41245 23511
rect 40512 23480 41245 23508
rect 41233 23477 41245 23480
rect 41279 23477 41291 23511
rect 41530 23508 41558 23616
rect 42242 23536 42248 23588
rect 42300 23576 42306 23588
rect 42429 23579 42487 23585
rect 42429 23576 42441 23579
rect 42300 23548 42441 23576
rect 42300 23536 42306 23548
rect 42429 23545 42441 23548
rect 42475 23545 42487 23579
rect 42536 23576 42564 23616
rect 43070 23604 43076 23616
rect 43128 23604 43134 23656
rect 43824 23576 43852 23684
rect 43901 23681 43913 23684
rect 43947 23712 43959 23715
rect 44266 23712 44272 23724
rect 43947 23684 44272 23712
rect 43947 23681 43959 23684
rect 43901 23675 43959 23681
rect 44266 23672 44272 23684
rect 44324 23712 44330 23724
rect 44361 23715 44419 23721
rect 44361 23712 44373 23715
rect 44324 23684 44373 23712
rect 44324 23672 44330 23684
rect 44361 23681 44373 23684
rect 44407 23712 44419 23715
rect 44637 23715 44695 23721
rect 44637 23712 44649 23715
rect 44407 23684 44649 23712
rect 44407 23681 44419 23684
rect 44361 23675 44419 23681
rect 44637 23681 44649 23684
rect 44683 23681 44695 23715
rect 44637 23675 44695 23681
rect 44177 23647 44235 23653
rect 44177 23613 44189 23647
rect 44223 23644 44235 23647
rect 44450 23644 44456 23656
rect 44223 23616 44456 23644
rect 44223 23613 44235 23616
rect 44177 23607 44235 23613
rect 44450 23604 44456 23616
rect 44508 23644 44514 23656
rect 45370 23644 45376 23656
rect 44508 23616 45376 23644
rect 44508 23604 44514 23616
rect 45370 23604 45376 23616
rect 45428 23604 45434 23656
rect 44913 23579 44971 23585
rect 44913 23576 44925 23579
rect 42536 23548 43852 23576
rect 44192 23548 44925 23576
rect 42429 23539 42487 23545
rect 44192 23520 44220 23548
rect 44913 23545 44925 23548
rect 44959 23545 44971 23579
rect 44913 23539 44971 23545
rect 45097 23579 45155 23585
rect 45097 23545 45109 23579
rect 45143 23576 45155 23579
rect 45572 23576 45600 23752
rect 45646 23740 45652 23792
rect 45704 23780 45710 23792
rect 45704 23752 46336 23780
rect 45704 23740 45710 23752
rect 45833 23715 45891 23721
rect 45833 23681 45845 23715
rect 45879 23712 45891 23715
rect 45922 23712 45928 23724
rect 45879 23684 45928 23712
rect 45879 23681 45891 23684
rect 45833 23675 45891 23681
rect 45922 23672 45928 23684
rect 45980 23672 45986 23724
rect 46308 23721 46336 23752
rect 46293 23715 46351 23721
rect 46293 23681 46305 23715
rect 46339 23681 46351 23715
rect 46293 23675 46351 23681
rect 45738 23604 45744 23656
rect 45796 23604 45802 23656
rect 46201 23647 46259 23653
rect 46201 23613 46213 23647
rect 46247 23613 46259 23647
rect 46201 23607 46259 23613
rect 46216 23576 46244 23607
rect 45143 23548 46244 23576
rect 45143 23545 45155 23548
rect 45097 23539 45155 23545
rect 46382 23536 46388 23588
rect 46440 23536 46446 23588
rect 43714 23508 43720 23520
rect 41530 23480 43720 23508
rect 41233 23471 41291 23477
rect 43714 23468 43720 23480
rect 43772 23468 43778 23520
rect 44174 23468 44180 23520
rect 44232 23468 44238 23520
rect 1104 23418 47104 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 47104 23418
rect 1104 23344 47104 23366
rect 2130 23264 2136 23316
rect 2188 23304 2194 23316
rect 2188 23276 12434 23304
rect 2188 23264 2194 23276
rect 3145 23239 3203 23245
rect 3145 23205 3157 23239
rect 3191 23236 3203 23239
rect 3786 23236 3792 23248
rect 3191 23208 3792 23236
rect 3191 23205 3203 23208
rect 3145 23199 3203 23205
rect 3786 23196 3792 23208
rect 3844 23196 3850 23248
rect 12406 23236 12434 23276
rect 12986 23264 12992 23316
rect 13044 23304 13050 23316
rect 13633 23307 13691 23313
rect 13633 23304 13645 23307
rect 13044 23276 13645 23304
rect 13044 23264 13050 23276
rect 13633 23273 13645 23276
rect 13679 23273 13691 23307
rect 13633 23267 13691 23273
rect 14093 23307 14151 23313
rect 14093 23273 14105 23307
rect 14139 23304 14151 23307
rect 15378 23304 15384 23316
rect 14139 23276 15384 23304
rect 14139 23273 14151 23276
rect 14093 23267 14151 23273
rect 15378 23264 15384 23276
rect 15436 23264 15442 23316
rect 15672 23276 18736 23304
rect 15672 23236 15700 23276
rect 12406 23208 15700 23236
rect 17402 23196 17408 23248
rect 17460 23196 17466 23248
rect 4614 23168 4620 23180
rect 4448 23140 4620 23168
rect 1670 23060 1676 23112
rect 1728 23100 1734 23112
rect 2038 23109 2044 23112
rect 1765 23103 1823 23109
rect 1765 23100 1777 23103
rect 1728 23072 1777 23100
rect 1728 23060 1734 23072
rect 1765 23069 1777 23072
rect 1811 23069 1823 23103
rect 2032 23100 2044 23109
rect 1999 23072 2044 23100
rect 1765 23063 1823 23069
rect 2032 23063 2044 23072
rect 2038 23060 2044 23063
rect 2096 23060 2102 23112
rect 4448 23109 4476 23140
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 4709 23171 4767 23177
rect 4709 23137 4721 23171
rect 4755 23168 4767 23171
rect 5074 23168 5080 23180
rect 4755 23140 5080 23168
rect 4755 23137 4767 23140
rect 4709 23131 4767 23137
rect 5074 23128 5080 23140
rect 5132 23128 5138 23180
rect 5166 23128 5172 23180
rect 5224 23128 5230 23180
rect 5626 23177 5632 23180
rect 5583 23171 5632 23177
rect 5583 23137 5595 23171
rect 5629 23137 5632 23171
rect 5583 23131 5632 23137
rect 5626 23128 5632 23131
rect 5684 23128 5690 23180
rect 6365 23171 6423 23177
rect 6365 23137 6377 23171
rect 6411 23168 6423 23171
rect 6411 23140 9076 23168
rect 6411 23137 6423 23140
rect 6365 23131 6423 23137
rect 4433 23103 4491 23109
rect 4433 23069 4445 23103
rect 4479 23069 4491 23103
rect 4433 23063 4491 23069
rect 4522 23060 4528 23112
rect 4580 23100 4586 23112
rect 4890 23100 4896 23112
rect 4580 23072 4896 23100
rect 4580 23060 4586 23072
rect 4890 23060 4896 23072
rect 4948 23060 4954 23112
rect 5442 23060 5448 23112
rect 5500 23060 5506 23112
rect 5718 23060 5724 23112
rect 5776 23060 5782 23112
rect 8754 23060 8760 23112
rect 8812 23060 8818 23112
rect 8938 23060 8944 23112
rect 8996 23060 9002 23112
rect 9048 23100 9076 23140
rect 14734 23128 14740 23180
rect 14792 23128 14798 23180
rect 9674 23100 9680 23112
rect 9048 23072 9680 23100
rect 9674 23060 9680 23072
rect 9732 23060 9738 23112
rect 15562 23060 15568 23112
rect 15620 23060 15626 23112
rect 15654 23060 15660 23112
rect 15712 23060 15718 23112
rect 15924 23103 15982 23109
rect 15924 23100 15936 23103
rect 15764 23072 15936 23100
rect 9186 23035 9244 23041
rect 9186 23032 9198 23035
rect 8588 23004 9198 23032
rect 4249 22967 4307 22973
rect 4249 22933 4261 22967
rect 4295 22964 4307 22967
rect 4614 22964 4620 22976
rect 4295 22936 4620 22964
rect 4295 22933 4307 22936
rect 4249 22927 4307 22933
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 5626 22924 5632 22976
rect 5684 22964 5690 22976
rect 6270 22964 6276 22976
rect 5684 22936 6276 22964
rect 5684 22924 5690 22936
rect 6270 22924 6276 22936
rect 6328 22924 6334 22976
rect 8588 22973 8616 23004
rect 9186 23001 9198 23004
rect 9232 23001 9244 23035
rect 9186 22995 9244 23001
rect 9398 22992 9404 23044
rect 9456 23032 9462 23044
rect 11149 23035 11207 23041
rect 9456 23004 10456 23032
rect 9456 22992 9462 23004
rect 8573 22967 8631 22973
rect 8573 22933 8585 22967
rect 8619 22933 8631 22967
rect 8573 22927 8631 22933
rect 9490 22924 9496 22976
rect 9548 22964 9554 22976
rect 10321 22967 10379 22973
rect 10321 22964 10333 22967
rect 9548 22936 10333 22964
rect 9548 22924 9554 22936
rect 10321 22933 10333 22936
rect 10367 22933 10379 22967
rect 10428 22964 10456 23004
rect 11149 23001 11161 23035
rect 11195 23032 11207 23035
rect 11882 23032 11888 23044
rect 11195 23004 11888 23032
rect 11195 23001 11207 23004
rect 11149 22995 11207 23001
rect 11882 22992 11888 23004
rect 11940 22992 11946 23044
rect 13354 22992 13360 23044
rect 13412 23032 13418 23044
rect 13541 23035 13599 23041
rect 13541 23032 13553 23035
rect 13412 23004 13553 23032
rect 13412 22992 13418 23004
rect 13541 23001 13553 23004
rect 13587 23001 13599 23035
rect 13541 22995 13599 23001
rect 14461 23035 14519 23041
rect 14461 23001 14473 23035
rect 14507 23032 14519 23035
rect 15102 23032 15108 23044
rect 14507 23004 15108 23032
rect 14507 23001 14519 23004
rect 14461 22995 14519 23001
rect 15102 22992 15108 23004
rect 15160 22992 15166 23044
rect 11241 22967 11299 22973
rect 11241 22964 11253 22967
rect 10428 22936 11253 22964
rect 10321 22927 10379 22933
rect 11241 22933 11253 22936
rect 11287 22933 11299 22967
rect 11241 22927 11299 22933
rect 14550 22924 14556 22976
rect 14608 22924 14614 22976
rect 15381 22967 15439 22973
rect 15381 22933 15393 22967
rect 15427 22964 15439 22967
rect 15764 22964 15792 23072
rect 15924 23069 15936 23072
rect 15970 23069 15982 23103
rect 15924 23063 15982 23069
rect 17586 23060 17592 23112
rect 17644 23060 17650 23112
rect 17678 23060 17684 23112
rect 17736 23060 17742 23112
rect 18708 23100 18736 23276
rect 18782 23264 18788 23316
rect 18840 23304 18846 23316
rect 18840 23276 30972 23304
rect 18840 23264 18846 23276
rect 21542 23196 21548 23248
rect 21600 23236 21606 23248
rect 22097 23239 22155 23245
rect 22097 23236 22109 23239
rect 21600 23208 22109 23236
rect 21600 23196 21606 23208
rect 22097 23205 22109 23208
rect 22143 23205 22155 23239
rect 22097 23199 22155 23205
rect 22281 23239 22339 23245
rect 22281 23205 22293 23239
rect 22327 23236 22339 23239
rect 22327 23208 23152 23236
rect 22327 23205 22339 23208
rect 22281 23199 22339 23205
rect 21634 23128 21640 23180
rect 21692 23168 21698 23180
rect 21821 23171 21879 23177
rect 21821 23168 21833 23171
rect 21692 23140 21833 23168
rect 21692 23128 21698 23140
rect 21821 23137 21833 23140
rect 21867 23137 21879 23171
rect 21821 23131 21879 23137
rect 22002 23128 22008 23180
rect 22060 23168 22066 23180
rect 23017 23171 23075 23177
rect 23017 23168 23029 23171
rect 22060 23140 23029 23168
rect 22060 23128 22066 23140
rect 23017 23137 23029 23140
rect 23063 23137 23075 23171
rect 23017 23131 23075 23137
rect 18708 23072 21864 23100
rect 17402 22992 17408 23044
rect 17460 23032 17466 23044
rect 17926 23035 17984 23041
rect 17926 23032 17938 23035
rect 17460 23004 17938 23032
rect 17460 22992 17466 23004
rect 17926 23001 17938 23004
rect 17972 23001 17984 23035
rect 17926 22995 17984 23001
rect 18046 22992 18052 23044
rect 18104 23032 18110 23044
rect 21836 23032 21864 23072
rect 22738 23060 22744 23112
rect 22796 23060 22802 23112
rect 23124 23109 23152 23208
rect 24486 23196 24492 23248
rect 24544 23236 24550 23248
rect 25590 23236 25596 23248
rect 24544 23208 25596 23236
rect 24544 23196 24550 23208
rect 25590 23196 25596 23208
rect 25648 23196 25654 23248
rect 26234 23196 26240 23248
rect 26292 23236 26298 23248
rect 27706 23236 27712 23248
rect 26292 23208 27712 23236
rect 26292 23196 26298 23208
rect 27706 23196 27712 23208
rect 27764 23196 27770 23248
rect 23198 23128 23204 23180
rect 23256 23168 23262 23180
rect 24670 23168 24676 23180
rect 23256 23140 24676 23168
rect 23256 23128 23262 23140
rect 24670 23128 24676 23140
rect 24728 23168 24734 23180
rect 29822 23168 29828 23180
rect 24728 23140 29828 23168
rect 24728 23128 24734 23140
rect 29822 23128 29828 23140
rect 29880 23128 29886 23180
rect 22833 23103 22891 23109
rect 22833 23069 22845 23103
rect 22879 23069 22891 23103
rect 22833 23063 22891 23069
rect 23109 23103 23167 23109
rect 23109 23069 23121 23103
rect 23155 23069 23167 23103
rect 23109 23063 23167 23069
rect 22848 23032 22876 23063
rect 23382 23060 23388 23112
rect 23440 23060 23446 23112
rect 23661 23103 23719 23109
rect 23661 23069 23673 23103
rect 23707 23100 23719 23103
rect 23750 23100 23756 23112
rect 23707 23072 23756 23100
rect 23707 23069 23719 23072
rect 23661 23063 23719 23069
rect 23750 23060 23756 23072
rect 23808 23060 23814 23112
rect 25590 23060 25596 23112
rect 25648 23100 25654 23112
rect 29638 23100 29644 23112
rect 25648 23072 29644 23100
rect 25648 23060 25654 23072
rect 29638 23060 29644 23072
rect 29696 23060 29702 23112
rect 29917 23103 29975 23109
rect 29917 23069 29929 23103
rect 29963 23100 29975 23103
rect 30006 23100 30012 23112
rect 29963 23072 30012 23100
rect 29963 23069 29975 23072
rect 29917 23063 29975 23069
rect 30006 23060 30012 23072
rect 30064 23060 30070 23112
rect 30190 23109 30196 23112
rect 30184 23100 30196 23109
rect 30151 23072 30196 23100
rect 30184 23063 30196 23072
rect 30190 23060 30196 23063
rect 30248 23060 30254 23112
rect 30944 23100 30972 23276
rect 31202 23264 31208 23316
rect 31260 23304 31266 23316
rect 31297 23307 31355 23313
rect 31297 23304 31309 23307
rect 31260 23276 31309 23304
rect 31260 23264 31266 23276
rect 31297 23273 31309 23276
rect 31343 23273 31355 23307
rect 31297 23267 31355 23273
rect 31386 23264 31392 23316
rect 31444 23304 31450 23316
rect 32030 23304 32036 23316
rect 31444 23276 32036 23304
rect 31444 23264 31450 23276
rect 32030 23264 32036 23276
rect 32088 23264 32094 23316
rect 35897 23307 35955 23313
rect 35897 23273 35909 23307
rect 35943 23304 35955 23307
rect 36630 23304 36636 23316
rect 35943 23276 36636 23304
rect 35943 23273 35955 23276
rect 35897 23267 35955 23273
rect 36630 23264 36636 23276
rect 36688 23264 36694 23316
rect 38838 23264 38844 23316
rect 38896 23304 38902 23316
rect 39025 23307 39083 23313
rect 39025 23304 39037 23307
rect 38896 23276 39037 23304
rect 38896 23264 38902 23276
rect 39025 23273 39037 23276
rect 39071 23273 39083 23307
rect 39025 23267 39083 23273
rect 41874 23264 41880 23316
rect 41932 23304 41938 23316
rect 42426 23304 42432 23316
rect 41932 23276 42432 23304
rect 41932 23264 41938 23276
rect 42426 23264 42432 23276
rect 42484 23304 42490 23316
rect 46201 23307 46259 23313
rect 46201 23304 46213 23307
rect 42484 23276 46213 23304
rect 42484 23264 42490 23276
rect 46201 23273 46213 23276
rect 46247 23273 46259 23307
rect 46201 23267 46259 23273
rect 32950 23196 32956 23248
rect 33008 23236 33014 23248
rect 34054 23236 34060 23248
rect 33008 23208 34060 23236
rect 33008 23196 33014 23208
rect 34054 23196 34060 23208
rect 34112 23196 34118 23248
rect 36357 23239 36415 23245
rect 36357 23205 36369 23239
rect 36403 23205 36415 23239
rect 36357 23199 36415 23205
rect 41969 23239 42027 23245
rect 41969 23205 41981 23239
rect 42015 23236 42027 23239
rect 42058 23236 42064 23248
rect 42015 23208 42064 23236
rect 42015 23205 42027 23208
rect 41969 23199 42027 23205
rect 31018 23128 31024 23180
rect 31076 23168 31082 23180
rect 31076 23140 33088 23168
rect 31076 23128 31082 23140
rect 32950 23100 32956 23112
rect 30944 23072 32956 23100
rect 32950 23060 32956 23072
rect 33008 23060 33014 23112
rect 33060 23109 33088 23140
rect 33318 23128 33324 23180
rect 33376 23168 33382 23180
rect 34698 23168 34704 23180
rect 33376 23140 34704 23168
rect 33376 23128 33382 23140
rect 34698 23128 34704 23140
rect 34756 23128 34762 23180
rect 33045 23103 33103 23109
rect 33045 23069 33057 23103
rect 33091 23069 33103 23103
rect 33045 23063 33103 23069
rect 36081 23103 36139 23109
rect 36081 23069 36093 23103
rect 36127 23100 36139 23103
rect 36372 23100 36400 23199
rect 42058 23196 42064 23208
rect 42116 23236 42122 23248
rect 43070 23236 43076 23248
rect 42116 23208 43076 23236
rect 42116 23196 42122 23208
rect 36906 23128 36912 23180
rect 36964 23128 36970 23180
rect 38654 23128 38660 23180
rect 38712 23168 38718 23180
rect 39022 23168 39028 23180
rect 38712 23140 39028 23168
rect 38712 23128 38718 23140
rect 39022 23128 39028 23140
rect 39080 23128 39086 23180
rect 42518 23128 42524 23180
rect 42576 23128 42582 23180
rect 42996 23177 43024 23208
rect 43070 23196 43076 23208
rect 43128 23196 43134 23248
rect 44453 23239 44511 23245
rect 44453 23236 44465 23239
rect 43548 23208 44465 23236
rect 42981 23171 43039 23177
rect 42981 23137 42993 23171
rect 43027 23137 43039 23171
rect 43548 23168 43576 23208
rect 44453 23205 44465 23208
rect 44499 23205 44511 23239
rect 44453 23199 44511 23205
rect 44634 23196 44640 23248
rect 44692 23236 44698 23248
rect 45833 23239 45891 23245
rect 45833 23236 45845 23239
rect 44692 23208 45845 23236
rect 44692 23196 44698 23208
rect 45833 23205 45845 23208
rect 45879 23205 45891 23239
rect 45833 23199 45891 23205
rect 46382 23196 46388 23248
rect 46440 23196 46446 23248
rect 46753 23239 46811 23245
rect 46753 23205 46765 23239
rect 46799 23236 46811 23239
rect 46934 23236 46940 23248
rect 46799 23208 46940 23236
rect 46799 23205 46811 23208
rect 46753 23199 46811 23205
rect 46934 23196 46940 23208
rect 46992 23196 46998 23248
rect 42981 23131 43039 23137
rect 43456 23140 43576 23168
rect 36127 23072 36400 23100
rect 36725 23103 36783 23109
rect 36127 23069 36139 23072
rect 36081 23063 36139 23069
rect 36725 23069 36737 23103
rect 36771 23100 36783 23103
rect 36814 23100 36820 23112
rect 36771 23072 36820 23100
rect 36771 23069 36783 23072
rect 36725 23063 36783 23069
rect 23201 23035 23259 23041
rect 23201 23032 23213 23035
rect 18104 23004 21220 23032
rect 21836 23004 22692 23032
rect 22848 23004 23213 23032
rect 18104 22992 18110 23004
rect 15427 22936 15792 22964
rect 15427 22933 15439 22936
rect 15381 22927 15439 22933
rect 17034 22924 17040 22976
rect 17092 22924 17098 22976
rect 19061 22967 19119 22973
rect 19061 22933 19073 22967
rect 19107 22964 19119 22967
rect 19886 22964 19892 22976
rect 19107 22936 19892 22964
rect 19107 22933 19119 22936
rect 19061 22927 19119 22933
rect 19886 22924 19892 22936
rect 19944 22924 19950 22976
rect 21192 22964 21220 23004
rect 22002 22964 22008 22976
rect 21192 22936 22008 22964
rect 22002 22924 22008 22936
rect 22060 22924 22066 22976
rect 22554 22924 22560 22976
rect 22612 22924 22618 22976
rect 22664 22964 22692 23004
rect 23201 23001 23213 23004
rect 23247 23001 23259 23035
rect 32858 23032 32864 23044
rect 23201 22995 23259 23001
rect 23308 23004 32864 23032
rect 23308 22964 23336 23004
rect 32858 22992 32864 23004
rect 32916 22992 32922 23044
rect 22664 22936 23336 22964
rect 23569 22967 23627 22973
rect 23569 22933 23581 22967
rect 23615 22964 23627 22967
rect 24946 22964 24952 22976
rect 23615 22936 24952 22964
rect 23615 22933 23627 22936
rect 23569 22927 23627 22933
rect 24946 22924 24952 22936
rect 25004 22924 25010 22976
rect 27614 22924 27620 22976
rect 27672 22964 27678 22976
rect 31018 22964 31024 22976
rect 27672 22936 31024 22964
rect 27672 22924 27678 22936
rect 31018 22924 31024 22936
rect 31076 22924 31082 22976
rect 33060 22964 33088 23063
rect 36814 23060 36820 23072
rect 36872 23060 36878 23112
rect 38841 23103 38899 23109
rect 38841 23069 38853 23103
rect 38887 23100 38899 23103
rect 39666 23100 39672 23112
rect 38887 23072 39672 23100
rect 38887 23069 38899 23072
rect 38841 23063 38899 23069
rect 39666 23060 39672 23072
rect 39724 23060 39730 23112
rect 42337 23103 42395 23109
rect 42337 23069 42349 23103
rect 42383 23100 42395 23103
rect 42426 23100 42432 23112
rect 42383 23072 42432 23100
rect 42383 23069 42395 23072
rect 42337 23063 42395 23069
rect 42426 23060 42432 23072
rect 42484 23100 42490 23112
rect 42613 23103 42671 23109
rect 42613 23100 42625 23103
rect 42484 23072 42625 23100
rect 42484 23060 42490 23072
rect 42613 23069 42625 23072
rect 42659 23069 42671 23103
rect 42613 23063 42671 23069
rect 42705 23103 42763 23109
rect 42705 23069 42717 23103
rect 42751 23100 42763 23103
rect 42886 23100 42892 23112
rect 42751 23072 42892 23100
rect 42751 23069 42763 23072
rect 42705 23063 42763 23069
rect 42245 23035 42303 23041
rect 42245 23001 42257 23035
rect 42291 23032 42303 23035
rect 42720 23032 42748 23063
rect 42886 23060 42892 23072
rect 42944 23060 42950 23112
rect 43456 23109 43484 23140
rect 43714 23128 43720 23180
rect 43772 23128 43778 23180
rect 44910 23168 44916 23180
rect 43916 23140 44916 23168
rect 43441 23103 43499 23109
rect 43441 23069 43453 23103
rect 43487 23069 43499 23103
rect 43441 23063 43499 23069
rect 43530 23060 43536 23112
rect 43588 23060 43594 23112
rect 43622 23060 43628 23112
rect 43680 23100 43686 23112
rect 43916 23109 43944 23140
rect 43809 23103 43867 23109
rect 43809 23100 43821 23103
rect 43680 23072 43821 23100
rect 43680 23060 43686 23072
rect 43809 23069 43821 23072
rect 43855 23100 43867 23103
rect 43901 23103 43959 23109
rect 43901 23100 43913 23103
rect 43855 23072 43913 23100
rect 43855 23069 43867 23072
rect 43809 23063 43867 23069
rect 43901 23069 43913 23072
rect 43947 23069 43959 23103
rect 43901 23063 43959 23069
rect 44174 23060 44180 23112
rect 44232 23060 44238 23112
rect 44266 23060 44272 23112
rect 44324 23060 44330 23112
rect 44652 23109 44680 23140
rect 44910 23128 44916 23140
rect 44968 23128 44974 23180
rect 46400 23168 46428 23196
rect 45848 23140 46428 23168
rect 45848 23109 45876 23140
rect 44637 23103 44695 23109
rect 44637 23069 44649 23103
rect 44683 23069 44695 23103
rect 44637 23063 44695 23069
rect 44729 23103 44787 23109
rect 44729 23069 44741 23103
rect 44775 23100 44787 23103
rect 45005 23103 45063 23109
rect 45005 23100 45017 23103
rect 44775 23072 45017 23100
rect 44775 23069 44787 23072
rect 44729 23063 44787 23069
rect 45005 23069 45017 23072
rect 45051 23069 45063 23103
rect 45005 23063 45063 23069
rect 45373 23103 45431 23109
rect 45373 23069 45385 23103
rect 45419 23069 45431 23103
rect 45373 23063 45431 23069
rect 45833 23103 45891 23109
rect 45833 23069 45845 23103
rect 45879 23069 45891 23103
rect 45833 23063 45891 23069
rect 42291 23004 42748 23032
rect 42291 23001 42303 23004
rect 42245 22995 42303 23001
rect 43714 22992 43720 23044
rect 43772 23032 43778 23044
rect 44085 23035 44143 23041
rect 44085 23032 44097 23035
rect 43772 23004 44097 23032
rect 43772 22992 43778 23004
rect 44085 23001 44097 23004
rect 44131 23032 44143 23035
rect 45186 23032 45192 23044
rect 44131 23004 45192 23032
rect 44131 23001 44143 23004
rect 44085 22995 44143 23001
rect 45186 22992 45192 23004
rect 45244 23032 45250 23044
rect 45388 23032 45416 23063
rect 45922 23060 45928 23112
rect 45980 23100 45986 23112
rect 46201 23103 46259 23109
rect 46201 23100 46213 23103
rect 45980 23072 46213 23100
rect 45980 23060 45986 23072
rect 46201 23069 46213 23072
rect 46247 23069 46259 23103
rect 46201 23063 46259 23069
rect 46385 23103 46443 23109
rect 46385 23069 46397 23103
rect 46431 23069 46443 23103
rect 46385 23063 46443 23069
rect 45244 23004 45416 23032
rect 45244 22992 45250 23004
rect 45738 22992 45744 23044
rect 45796 23032 45802 23044
rect 46400 23032 46428 23063
rect 46566 23060 46572 23112
rect 46624 23060 46630 23112
rect 45796 23004 46428 23032
rect 45796 22992 45802 23004
rect 36817 22967 36875 22973
rect 36817 22964 36829 22967
rect 33060 22936 36829 22964
rect 36817 22933 36829 22936
rect 36863 22964 36875 22967
rect 38378 22964 38384 22976
rect 36863 22936 38384 22964
rect 36863 22933 36875 22936
rect 36817 22927 36875 22933
rect 38378 22924 38384 22936
rect 38436 22924 38442 22976
rect 42153 22967 42211 22973
rect 42153 22933 42165 22967
rect 42199 22964 42211 22967
rect 42610 22964 42616 22976
rect 42199 22936 42616 22964
rect 42199 22933 42211 22936
rect 42153 22927 42211 22933
rect 42610 22924 42616 22936
rect 42668 22964 42674 22976
rect 42797 22967 42855 22973
rect 42797 22964 42809 22967
rect 42668 22936 42809 22964
rect 42668 22924 42674 22936
rect 42797 22933 42809 22936
rect 42843 22933 42855 22967
rect 42797 22927 42855 22933
rect 42886 22924 42892 22976
rect 42944 22924 42950 22976
rect 43254 22924 43260 22976
rect 43312 22924 43318 22976
rect 1104 22874 47104 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 47104 22874
rect 1104 22800 47104 22822
rect 3234 22720 3240 22772
rect 3292 22720 3298 22772
rect 3605 22763 3663 22769
rect 3605 22729 3617 22763
rect 3651 22760 3663 22763
rect 3786 22760 3792 22772
rect 3651 22732 3792 22760
rect 3651 22729 3663 22732
rect 3605 22723 3663 22729
rect 3786 22720 3792 22732
rect 3844 22720 3850 22772
rect 4525 22763 4583 22769
rect 4525 22729 4537 22763
rect 4571 22729 4583 22763
rect 4525 22723 4583 22729
rect 3694 22652 3700 22704
rect 3752 22652 3758 22704
rect 4540 22692 4568 22723
rect 4798 22720 4804 22772
rect 4856 22760 4862 22772
rect 4856 22732 5212 22760
rect 4856 22720 4862 22732
rect 5046 22695 5104 22701
rect 5046 22692 5058 22695
rect 4540 22664 5058 22692
rect 5046 22661 5058 22664
rect 5092 22661 5104 22695
rect 5184 22692 5212 22732
rect 5350 22720 5356 22772
rect 5408 22760 5414 22772
rect 5718 22760 5724 22772
rect 5408 22732 5724 22760
rect 5408 22720 5414 22732
rect 5718 22720 5724 22732
rect 5776 22760 5782 22772
rect 6181 22763 6239 22769
rect 6181 22760 6193 22763
rect 5776 22732 6193 22760
rect 5776 22720 5782 22732
rect 6181 22729 6193 22732
rect 6227 22729 6239 22763
rect 6181 22723 6239 22729
rect 8113 22763 8171 22769
rect 8113 22729 8125 22763
rect 8159 22760 8171 22763
rect 8386 22760 8392 22772
rect 8159 22732 8392 22760
rect 8159 22729 8171 22732
rect 8113 22723 8171 22729
rect 8386 22720 8392 22732
rect 8444 22720 8450 22772
rect 8481 22763 8539 22769
rect 8481 22729 8493 22763
rect 8527 22729 8539 22763
rect 8481 22723 8539 22729
rect 5626 22692 5632 22704
rect 5184 22664 5632 22692
rect 5046 22655 5104 22661
rect 5626 22652 5632 22664
rect 5684 22652 5690 22704
rect 2038 22633 2044 22636
rect 2032 22587 2044 22633
rect 2038 22584 2044 22587
rect 2096 22584 2102 22636
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22624 4767 22627
rect 5350 22624 5356 22636
rect 4755 22596 5356 22624
rect 4755 22593 4767 22596
rect 4709 22587 4767 22593
rect 5350 22584 5356 22596
rect 5408 22584 5414 22636
rect 8021 22627 8079 22633
rect 8021 22593 8033 22627
rect 8067 22624 8079 22627
rect 8386 22624 8392 22636
rect 8067 22596 8392 22624
rect 8067 22593 8079 22596
rect 8021 22587 8079 22593
rect 8386 22584 8392 22596
rect 8444 22584 8450 22636
rect 8496 22568 8524 22723
rect 8570 22720 8576 22772
rect 8628 22760 8634 22772
rect 8941 22763 8999 22769
rect 8941 22760 8953 22763
rect 8628 22732 8953 22760
rect 8628 22720 8634 22732
rect 8941 22729 8953 22732
rect 8987 22760 8999 22763
rect 9214 22760 9220 22772
rect 8987 22732 9220 22760
rect 8987 22729 8999 22732
rect 8941 22723 8999 22729
rect 9214 22720 9220 22732
rect 9272 22760 9278 22772
rect 10778 22760 10784 22772
rect 9272 22732 10784 22760
rect 9272 22720 9278 22732
rect 10778 22720 10784 22732
rect 10836 22720 10842 22772
rect 11146 22720 11152 22772
rect 11204 22720 11210 22772
rect 11333 22763 11391 22769
rect 11333 22729 11345 22763
rect 11379 22760 11391 22763
rect 12894 22760 12900 22772
rect 11379 22732 12900 22760
rect 11379 22729 11391 22732
rect 11333 22723 11391 22729
rect 12894 22720 12900 22732
rect 12952 22720 12958 22772
rect 12986 22720 12992 22772
rect 13044 22760 13050 22772
rect 15286 22760 15292 22772
rect 13044 22732 15292 22760
rect 13044 22720 13050 22732
rect 15286 22720 15292 22732
rect 15344 22720 15350 22772
rect 15562 22720 15568 22772
rect 15620 22760 15626 22772
rect 16669 22763 16727 22769
rect 16669 22760 16681 22763
rect 15620 22732 16681 22760
rect 15620 22720 15626 22732
rect 16669 22729 16681 22732
rect 16715 22729 16727 22763
rect 16669 22723 16727 22729
rect 17586 22720 17592 22772
rect 17644 22760 17650 22772
rect 18325 22763 18383 22769
rect 18325 22760 18337 22763
rect 17644 22732 18337 22760
rect 17644 22720 17650 22732
rect 18325 22729 18337 22732
rect 18371 22729 18383 22763
rect 20714 22760 20720 22772
rect 18325 22723 18383 22729
rect 18892 22732 20720 22760
rect 9398 22652 9404 22704
rect 9456 22692 9462 22704
rect 11164 22692 11192 22720
rect 11793 22695 11851 22701
rect 11793 22692 11805 22695
rect 9456 22664 9720 22692
rect 11164 22664 11805 22692
rect 9456 22652 9462 22664
rect 8846 22584 8852 22636
rect 8904 22584 8910 22636
rect 9122 22584 9128 22636
rect 9180 22624 9186 22636
rect 9490 22624 9496 22636
rect 9180 22596 9496 22624
rect 9180 22584 9186 22596
rect 9490 22584 9496 22596
rect 9548 22584 9554 22636
rect 9692 22624 9720 22664
rect 11793 22661 11805 22664
rect 11839 22661 11851 22695
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 11793 22655 11851 22661
rect 14844 22664 17141 22692
rect 11517 22627 11575 22633
rect 9692 22596 9812 22624
rect 1670 22516 1676 22568
rect 1728 22556 1734 22568
rect 1765 22559 1823 22565
rect 1765 22556 1777 22559
rect 1728 22528 1777 22556
rect 1728 22516 1734 22528
rect 1765 22525 1777 22528
rect 1811 22525 1823 22559
rect 1765 22519 1823 22525
rect 3786 22516 3792 22568
rect 3844 22516 3850 22568
rect 4798 22516 4804 22568
rect 4856 22516 4862 22568
rect 8202 22516 8208 22568
rect 8260 22516 8266 22568
rect 8478 22516 8484 22568
rect 8536 22516 8542 22568
rect 9033 22559 9091 22565
rect 9033 22525 9045 22559
rect 9079 22525 9091 22559
rect 9033 22519 9091 22525
rect 6178 22448 6184 22500
rect 6236 22488 6242 22500
rect 6236 22460 7788 22488
rect 6236 22448 6242 22460
rect 2958 22380 2964 22432
rect 3016 22420 3022 22432
rect 3145 22423 3203 22429
rect 3145 22420 3157 22423
rect 3016 22392 3157 22420
rect 3016 22380 3022 22392
rect 3145 22389 3157 22392
rect 3191 22420 3203 22423
rect 5534 22420 5540 22432
rect 3191 22392 5540 22420
rect 3191 22389 3203 22392
rect 3145 22383 3203 22389
rect 5534 22380 5540 22392
rect 5592 22380 5598 22432
rect 7098 22380 7104 22432
rect 7156 22420 7162 22432
rect 7653 22423 7711 22429
rect 7653 22420 7665 22423
rect 7156 22392 7665 22420
rect 7156 22380 7162 22392
rect 7653 22389 7665 22392
rect 7699 22389 7711 22423
rect 7760 22420 7788 22460
rect 7834 22448 7840 22500
rect 7892 22488 7898 22500
rect 9048 22488 9076 22519
rect 9674 22516 9680 22568
rect 9732 22516 9738 22568
rect 9784 22556 9812 22596
rect 11517 22593 11529 22627
rect 11563 22624 11575 22627
rect 11882 22624 11888 22636
rect 11563 22596 11888 22624
rect 11563 22593 11575 22596
rect 11517 22587 11575 22593
rect 11882 22584 11888 22596
rect 11940 22584 11946 22636
rect 11974 22584 11980 22636
rect 12032 22624 12038 22636
rect 12069 22627 12127 22633
rect 12069 22624 12081 22627
rect 12032 22596 12081 22624
rect 12032 22584 12038 22596
rect 12069 22593 12081 22596
rect 12115 22593 12127 22627
rect 12069 22587 12127 22593
rect 12526 22584 12532 22636
rect 12584 22624 12590 22636
rect 12802 22624 12808 22636
rect 12584 22596 12808 22624
rect 12584 22584 12590 22596
rect 12802 22584 12808 22596
rect 12860 22624 12866 22636
rect 13170 22633 13176 22636
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12860 22596 12909 22624
rect 12860 22584 12866 22596
rect 12897 22593 12909 22596
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 13164 22587 13176 22633
rect 13170 22584 13176 22587
rect 13228 22584 13234 22636
rect 14737 22627 14795 22633
rect 14737 22593 14749 22627
rect 14783 22593 14795 22627
rect 14737 22587 14795 22593
rect 10137 22559 10195 22565
rect 10137 22556 10149 22559
rect 9784 22528 10149 22556
rect 10137 22525 10149 22528
rect 10183 22525 10195 22559
rect 10137 22519 10195 22525
rect 10410 22516 10416 22568
rect 10468 22516 10474 22568
rect 10502 22516 10508 22568
rect 10560 22565 10566 22568
rect 10560 22559 10588 22565
rect 10576 22525 10588 22559
rect 10560 22519 10588 22525
rect 10689 22559 10747 22565
rect 10689 22525 10701 22559
rect 10735 22556 10747 22559
rect 10735 22528 11100 22556
rect 10735 22525 10747 22528
rect 10689 22519 10747 22525
rect 10560 22516 10566 22519
rect 7892 22460 9076 22488
rect 11072 22488 11100 22528
rect 12253 22491 12311 22497
rect 12253 22488 12265 22491
rect 11072 22460 12265 22488
rect 7892 22448 7898 22460
rect 11072 22420 11100 22460
rect 12253 22457 12265 22460
rect 12299 22457 12311 22491
rect 12253 22451 12311 22457
rect 13906 22448 13912 22500
rect 13964 22488 13970 22500
rect 14369 22491 14427 22497
rect 14369 22488 14381 22491
rect 13964 22460 14381 22488
rect 13964 22448 13970 22460
rect 14369 22457 14381 22460
rect 14415 22457 14427 22491
rect 14369 22451 14427 22457
rect 14752 22488 14780 22587
rect 14844 22568 14872 22664
rect 17129 22661 17141 22664
rect 17175 22692 17187 22695
rect 17494 22692 17500 22704
rect 17175 22664 17500 22692
rect 17175 22661 17187 22664
rect 17129 22655 17187 22661
rect 17494 22652 17500 22664
rect 17552 22652 17558 22704
rect 18892 22692 18920 22732
rect 20714 22720 20720 22732
rect 20772 22720 20778 22772
rect 21542 22720 21548 22772
rect 21600 22720 21606 22772
rect 22281 22763 22339 22769
rect 22281 22729 22293 22763
rect 22327 22729 22339 22763
rect 22281 22723 22339 22729
rect 18616 22664 18920 22692
rect 16025 22627 16083 22633
rect 16025 22593 16037 22627
rect 16071 22624 16083 22627
rect 16482 22624 16488 22636
rect 16071 22596 16488 22624
rect 16071 22593 16083 22596
rect 16025 22587 16083 22593
rect 16482 22584 16488 22596
rect 16540 22584 16546 22636
rect 17034 22584 17040 22636
rect 17092 22624 17098 22636
rect 18616 22624 18644 22664
rect 17092 22596 18644 22624
rect 18693 22627 18751 22633
rect 17092 22584 17098 22596
rect 18693 22593 18705 22627
rect 18739 22624 18751 22627
rect 22296 22624 22324 22723
rect 22738 22720 22744 22772
rect 22796 22760 22802 22772
rect 23385 22763 23443 22769
rect 23385 22760 23397 22763
rect 22796 22732 23397 22760
rect 22796 22720 22802 22732
rect 23385 22729 23397 22732
rect 23431 22729 23443 22763
rect 23385 22723 23443 22729
rect 23934 22720 23940 22772
rect 23992 22760 23998 22772
rect 27709 22763 27767 22769
rect 27709 22760 27721 22763
rect 23992 22732 27721 22760
rect 23992 22720 23998 22732
rect 27709 22729 27721 22732
rect 27755 22760 27767 22763
rect 29365 22763 29423 22769
rect 29365 22760 29377 22763
rect 27755 22732 29377 22760
rect 27755 22729 27767 22732
rect 27709 22723 27767 22729
rect 29365 22729 29377 22732
rect 29411 22729 29423 22763
rect 29365 22723 29423 22729
rect 22554 22652 22560 22704
rect 22612 22692 22618 22704
rect 28534 22692 28540 22704
rect 22612 22664 28540 22692
rect 22612 22652 22618 22664
rect 28534 22652 28540 22664
rect 28592 22652 28598 22704
rect 29380 22692 29408 22723
rect 30466 22720 30472 22772
rect 30524 22720 30530 22772
rect 30929 22763 30987 22769
rect 30929 22729 30941 22763
rect 30975 22760 30987 22763
rect 31202 22760 31208 22772
rect 30975 22732 31208 22760
rect 30975 22729 30987 22732
rect 30929 22723 30987 22729
rect 31202 22720 31208 22732
rect 31260 22720 31266 22772
rect 32950 22760 32956 22772
rect 31726 22732 32956 22760
rect 31726 22692 31754 22732
rect 32950 22720 32956 22732
rect 33008 22720 33014 22772
rect 38746 22720 38752 22772
rect 38804 22720 38810 22772
rect 39666 22720 39672 22772
rect 39724 22760 39730 22772
rect 44450 22760 44456 22772
rect 39724 22732 44456 22760
rect 39724 22720 39730 22732
rect 44450 22720 44456 22732
rect 44508 22720 44514 22772
rect 29380 22664 31754 22692
rect 38194 22652 38200 22704
rect 38252 22692 38258 22704
rect 38657 22695 38715 22701
rect 38657 22692 38669 22695
rect 38252 22664 38669 22692
rect 38252 22652 38258 22664
rect 38657 22661 38669 22664
rect 38703 22661 38715 22695
rect 38657 22655 38715 22661
rect 22649 22627 22707 22633
rect 18739 22596 19932 22624
rect 22296 22596 22600 22624
rect 18739 22593 18751 22596
rect 18693 22587 18751 22593
rect 19904 22568 19932 22596
rect 14826 22516 14832 22568
rect 14884 22516 14890 22568
rect 14918 22516 14924 22568
rect 14976 22516 14982 22568
rect 16206 22516 16212 22568
rect 16264 22556 16270 22568
rect 17218 22556 17224 22568
rect 16264 22528 17224 22556
rect 16264 22516 16270 22528
rect 17218 22516 17224 22528
rect 17276 22516 17282 22568
rect 18782 22516 18788 22568
rect 18840 22516 18846 22568
rect 18874 22516 18880 22568
rect 18932 22516 18938 22568
rect 19702 22516 19708 22568
rect 19760 22516 19766 22568
rect 19886 22516 19892 22568
rect 19944 22516 19950 22568
rect 20254 22516 20260 22568
rect 20312 22556 20318 22568
rect 20349 22559 20407 22565
rect 20349 22556 20361 22559
rect 20312 22528 20361 22556
rect 20312 22516 20318 22528
rect 20349 22525 20361 22528
rect 20395 22525 20407 22559
rect 20622 22556 20628 22568
rect 20349 22519 20407 22525
rect 20456 22528 20628 22556
rect 20456 22488 20484 22528
rect 20622 22516 20628 22528
rect 20680 22516 20686 22568
rect 20714 22516 20720 22568
rect 20772 22565 20778 22568
rect 20772 22559 20800 22565
rect 20788 22525 20800 22559
rect 20772 22519 20800 22525
rect 20772 22516 20778 22519
rect 20898 22516 20904 22568
rect 20956 22556 20962 22568
rect 21266 22556 21272 22568
rect 20956 22528 21272 22556
rect 20956 22516 20962 22528
rect 21266 22516 21272 22528
rect 21324 22516 21330 22568
rect 21542 22516 21548 22568
rect 21600 22556 21606 22568
rect 21821 22559 21879 22565
rect 21821 22556 21833 22559
rect 21600 22528 21833 22556
rect 21600 22516 21606 22528
rect 21821 22525 21833 22528
rect 21867 22556 21879 22559
rect 22462 22556 22468 22568
rect 21867 22528 22468 22556
rect 21867 22525 21879 22528
rect 21821 22519 21879 22525
rect 22462 22516 22468 22528
rect 22520 22516 22526 22568
rect 22572 22556 22600 22596
rect 22649 22593 22661 22627
rect 22695 22624 22707 22627
rect 23474 22624 23480 22636
rect 22695 22596 23480 22624
rect 22695 22593 22707 22596
rect 22649 22587 22707 22593
rect 23474 22584 23480 22596
rect 23532 22584 23538 22636
rect 24394 22624 24400 22636
rect 24228 22596 24400 22624
rect 22738 22556 22744 22568
rect 22572 22528 22744 22556
rect 22738 22516 22744 22528
rect 22796 22516 22802 22568
rect 22922 22516 22928 22568
rect 22980 22516 22986 22568
rect 23658 22556 23664 22568
rect 23216 22528 23664 22556
rect 14752 22460 20484 22488
rect 7760 22392 11100 22420
rect 14277 22423 14335 22429
rect 7653 22383 7711 22389
rect 14277 22389 14289 22423
rect 14323 22420 14335 22423
rect 14752 22420 14780 22460
rect 22002 22448 22008 22500
rect 22060 22488 22066 22500
rect 22097 22491 22155 22497
rect 22097 22488 22109 22491
rect 22060 22460 22109 22488
rect 22060 22448 22066 22460
rect 22097 22457 22109 22460
rect 22143 22457 22155 22491
rect 23216 22488 23244 22528
rect 23658 22516 23664 22528
rect 23716 22556 23722 22568
rect 24228 22556 24256 22596
rect 24394 22584 24400 22596
rect 24452 22584 24458 22636
rect 24578 22633 24584 22636
rect 24572 22587 24584 22633
rect 24578 22584 24584 22587
rect 24636 22584 24642 22636
rect 25406 22584 25412 22636
rect 25464 22624 25470 22636
rect 27614 22624 27620 22636
rect 25464 22596 27620 22624
rect 25464 22584 25470 22596
rect 27614 22584 27620 22596
rect 27672 22584 27678 22636
rect 28077 22627 28135 22633
rect 28077 22624 28089 22627
rect 27816 22596 28089 22624
rect 23716 22528 24256 22556
rect 24305 22559 24363 22565
rect 23716 22516 23722 22528
rect 24305 22525 24317 22559
rect 24351 22525 24363 22559
rect 27062 22556 27068 22568
rect 24305 22519 24363 22525
rect 25332 22528 27068 22556
rect 22097 22451 22155 22457
rect 22204 22460 23244 22488
rect 23293 22491 23351 22497
rect 14323 22392 14780 22420
rect 14323 22389 14335 22392
rect 14277 22383 14335 22389
rect 16206 22380 16212 22432
rect 16264 22380 16270 22432
rect 20254 22380 20260 22432
rect 20312 22420 20318 22432
rect 22204 22420 22232 22460
rect 23293 22457 23305 22491
rect 23339 22488 23351 22491
rect 24026 22488 24032 22500
rect 23339 22460 24032 22488
rect 23339 22457 23351 22460
rect 23293 22451 23351 22457
rect 24026 22448 24032 22460
rect 24084 22448 24090 22500
rect 24320 22432 24348 22519
rect 20312 22392 22232 22420
rect 20312 22380 20318 22392
rect 22462 22380 22468 22432
rect 22520 22380 22526 22432
rect 24302 22380 24308 22432
rect 24360 22420 24366 22432
rect 25332 22420 25360 22528
rect 27062 22516 27068 22528
rect 27120 22516 27126 22568
rect 25590 22448 25596 22500
rect 25648 22488 25654 22500
rect 26970 22488 26976 22500
rect 25648 22460 26976 22488
rect 25648 22448 25654 22460
rect 26970 22448 26976 22460
rect 27028 22448 27034 22500
rect 27154 22448 27160 22500
rect 27212 22488 27218 22500
rect 27816 22488 27844 22596
rect 28077 22593 28089 22596
rect 28123 22624 28135 22627
rect 29086 22624 29092 22636
rect 28123 22596 29092 22624
rect 28123 22593 28135 22596
rect 28077 22587 28135 22593
rect 29086 22584 29092 22596
rect 29144 22584 29150 22636
rect 30285 22627 30343 22633
rect 30285 22593 30297 22627
rect 30331 22624 30343 22627
rect 30650 22624 30656 22636
rect 30331 22596 30656 22624
rect 30331 22593 30343 22596
rect 30285 22587 30343 22593
rect 30650 22584 30656 22596
rect 30708 22584 30714 22636
rect 30837 22627 30895 22633
rect 30837 22593 30849 22627
rect 30883 22624 30895 22627
rect 31294 22624 31300 22636
rect 30883 22596 31300 22624
rect 30883 22593 30895 22596
rect 30837 22587 30895 22593
rect 31294 22584 31300 22596
rect 31352 22584 31358 22636
rect 36262 22584 36268 22636
rect 36320 22624 36326 22636
rect 37277 22627 37335 22633
rect 37277 22624 37289 22627
rect 36320 22596 37289 22624
rect 36320 22584 36326 22596
rect 37277 22593 37289 22596
rect 37323 22593 37335 22627
rect 37277 22587 37335 22593
rect 38470 22584 38476 22636
rect 38528 22584 38534 22636
rect 38746 22584 38752 22636
rect 38804 22584 38810 22636
rect 39114 22584 39120 22636
rect 39172 22584 39178 22636
rect 42702 22584 42708 22636
rect 42760 22584 42766 22636
rect 42886 22584 42892 22636
rect 42944 22584 42950 22636
rect 27893 22559 27951 22565
rect 27893 22525 27905 22559
rect 27939 22525 27951 22559
rect 27893 22519 27951 22525
rect 27212 22460 27844 22488
rect 27908 22488 27936 22519
rect 28350 22516 28356 22568
rect 28408 22516 28414 22568
rect 29454 22516 29460 22568
rect 29512 22516 29518 22568
rect 29641 22559 29699 22565
rect 29641 22525 29653 22559
rect 29687 22525 29699 22559
rect 29641 22519 29699 22525
rect 31113 22559 31171 22565
rect 31113 22525 31125 22559
rect 31159 22525 31171 22559
rect 31113 22519 31171 22525
rect 28166 22488 28172 22500
rect 27908 22460 28172 22488
rect 27212 22448 27218 22460
rect 28166 22448 28172 22460
rect 28224 22448 28230 22500
rect 29362 22448 29368 22500
rect 29420 22488 29426 22500
rect 29656 22488 29684 22519
rect 31128 22488 31156 22519
rect 37366 22516 37372 22568
rect 37424 22556 37430 22568
rect 37553 22559 37611 22565
rect 37553 22556 37565 22559
rect 37424 22528 37565 22556
rect 37424 22516 37430 22528
rect 37553 22525 37565 22528
rect 37599 22525 37611 22559
rect 37553 22519 37611 22525
rect 42429 22559 42487 22565
rect 42429 22525 42441 22559
rect 42475 22556 42487 22559
rect 42610 22556 42616 22568
rect 42475 22528 42616 22556
rect 42475 22525 42487 22528
rect 42429 22519 42487 22525
rect 42610 22516 42616 22528
rect 42668 22556 42674 22568
rect 43254 22556 43260 22568
rect 42668 22528 43260 22556
rect 42668 22516 42674 22528
rect 43254 22516 43260 22528
rect 43312 22516 43318 22568
rect 29420 22460 31156 22488
rect 29420 22448 29426 22460
rect 39850 22448 39856 22500
rect 39908 22488 39914 22500
rect 43806 22488 43812 22500
rect 39908 22460 43812 22488
rect 39908 22448 39914 22460
rect 43806 22448 43812 22460
rect 43864 22448 43870 22500
rect 24360 22392 25360 22420
rect 25685 22423 25743 22429
rect 24360 22380 24366 22392
rect 25685 22389 25697 22423
rect 25731 22420 25743 22423
rect 25774 22420 25780 22432
rect 25731 22392 25780 22420
rect 25731 22389 25743 22392
rect 25685 22383 25743 22389
rect 25774 22380 25780 22392
rect 25832 22380 25838 22432
rect 27249 22423 27307 22429
rect 27249 22389 27261 22423
rect 27295 22420 27307 22423
rect 27982 22420 27988 22432
rect 27295 22392 27988 22420
rect 27295 22389 27307 22392
rect 27249 22383 27307 22389
rect 27982 22380 27988 22392
rect 28040 22380 28046 22432
rect 28902 22380 28908 22432
rect 28960 22420 28966 22432
rect 28997 22423 29055 22429
rect 28997 22420 29009 22423
rect 28960 22392 29009 22420
rect 28960 22380 28966 22392
rect 28997 22389 29009 22392
rect 29043 22389 29055 22423
rect 28997 22383 29055 22389
rect 30006 22380 30012 22432
rect 30064 22420 30070 22432
rect 30101 22423 30159 22429
rect 30101 22420 30113 22423
rect 30064 22392 30113 22420
rect 30064 22380 30070 22392
rect 30101 22389 30113 22392
rect 30147 22389 30159 22423
rect 30101 22383 30159 22389
rect 30650 22380 30656 22432
rect 30708 22420 30714 22432
rect 31202 22420 31208 22432
rect 30708 22392 31208 22420
rect 30708 22380 30714 22392
rect 31202 22380 31208 22392
rect 31260 22380 31266 22432
rect 32858 22380 32864 22432
rect 32916 22420 32922 22432
rect 38746 22420 38752 22432
rect 32916 22392 38752 22420
rect 32916 22380 32922 22392
rect 38746 22380 38752 22392
rect 38804 22420 38810 22432
rect 39209 22423 39267 22429
rect 39209 22420 39221 22423
rect 38804 22392 39221 22420
rect 38804 22380 38810 22392
rect 39209 22389 39221 22392
rect 39255 22389 39267 22423
rect 39209 22383 39267 22389
rect 42705 22423 42763 22429
rect 42705 22389 42717 22423
rect 42751 22420 42763 22423
rect 43254 22420 43260 22432
rect 42751 22392 43260 22420
rect 42751 22389 42763 22392
rect 42705 22383 42763 22389
rect 43254 22380 43260 22392
rect 43312 22380 43318 22432
rect 1104 22330 47104 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 47104 22330
rect 1104 22256 47104 22278
rect 2038 22176 2044 22228
rect 2096 22216 2102 22228
rect 2133 22219 2191 22225
rect 2133 22216 2145 22219
rect 2096 22188 2145 22216
rect 2096 22176 2102 22188
rect 2133 22185 2145 22188
rect 2179 22185 2191 22219
rect 4798 22216 4804 22228
rect 2133 22179 2191 22185
rect 3896 22188 4804 22216
rect 3252 22120 3832 22148
rect 3252 22092 3280 22120
rect 3234 22040 3240 22092
rect 3292 22040 3298 22092
rect 934 21972 940 22024
rect 992 22012 998 22024
rect 1581 22015 1639 22021
rect 1581 22012 1593 22015
rect 992 21984 1593 22012
rect 992 21972 998 21984
rect 1581 21981 1593 21984
rect 1627 21981 1639 22015
rect 1581 21975 1639 21981
rect 2317 22015 2375 22021
rect 2317 21981 2329 22015
rect 2363 22012 2375 22015
rect 2363 21984 2636 22012
rect 2363 21981 2375 21984
rect 2317 21975 2375 21981
rect 1397 21879 1455 21885
rect 1397 21845 1409 21879
rect 1443 21876 1455 21879
rect 2406 21876 2412 21888
rect 1443 21848 2412 21876
rect 1443 21845 1455 21848
rect 1397 21839 1455 21845
rect 2406 21836 2412 21848
rect 2464 21836 2470 21888
rect 2608 21885 2636 21984
rect 2958 21972 2964 22024
rect 3016 21972 3022 22024
rect 3804 22012 3832 22120
rect 3896 22089 3924 22188
rect 4798 22176 4804 22188
rect 4856 22176 4862 22228
rect 5258 22176 5264 22228
rect 5316 22176 5322 22228
rect 5350 22176 5356 22228
rect 5408 22176 5414 22228
rect 8202 22216 8208 22228
rect 5736 22188 8208 22216
rect 3881 22083 3939 22089
rect 3881 22049 3893 22083
rect 3927 22049 3939 22083
rect 5736 22080 5764 22188
rect 8202 22176 8208 22188
rect 8260 22176 8266 22228
rect 8386 22176 8392 22228
rect 8444 22216 8450 22228
rect 8573 22219 8631 22225
rect 8573 22216 8585 22219
rect 8444 22188 8585 22216
rect 8444 22176 8450 22188
rect 8573 22185 8585 22188
rect 8619 22216 8631 22219
rect 10502 22216 10508 22228
rect 8619 22188 10508 22216
rect 8619 22185 8631 22188
rect 8573 22179 8631 22185
rect 10502 22176 10508 22188
rect 10560 22176 10566 22228
rect 10778 22176 10784 22228
rect 10836 22216 10842 22228
rect 10836 22188 12434 22216
rect 10836 22176 10842 22188
rect 6270 22148 6276 22160
rect 6012 22120 6276 22148
rect 6012 22089 6040 22120
rect 6270 22108 6276 22120
rect 6328 22108 6334 22160
rect 8846 22108 8852 22160
rect 8904 22148 8910 22160
rect 12406 22148 12434 22188
rect 13170 22176 13176 22228
rect 13228 22216 13234 22228
rect 13265 22219 13323 22225
rect 13265 22216 13277 22219
rect 13228 22188 13277 22216
rect 13228 22176 13234 22188
rect 13265 22185 13277 22188
rect 13311 22185 13323 22219
rect 13265 22179 13323 22185
rect 15654 22176 15660 22228
rect 15712 22216 15718 22228
rect 15712 22188 16712 22216
rect 15712 22176 15718 22188
rect 14826 22148 14832 22160
rect 8904 22120 10272 22148
rect 12406 22120 14832 22148
rect 8904 22108 8910 22120
rect 3881 22043 3939 22049
rect 4908 22052 5764 22080
rect 5997 22083 6055 22089
rect 4148 22015 4206 22021
rect 3804 21984 3924 22012
rect 3896 21944 3924 21984
rect 4148 21981 4160 22015
rect 4194 22012 4206 22015
rect 4614 22012 4620 22024
rect 4194 21984 4620 22012
rect 4194 21981 4206 21984
rect 4148 21975 4206 21981
rect 4614 21972 4620 21984
rect 4672 21972 4678 22024
rect 4908 21944 4936 22052
rect 5997 22049 6009 22083
rect 6043 22049 6055 22083
rect 5997 22043 6055 22049
rect 7190 22040 7196 22092
rect 7248 22040 7254 22092
rect 9490 22040 9496 22092
rect 9548 22040 9554 22092
rect 10134 22040 10140 22092
rect 10192 22040 10198 22092
rect 10244 22080 10272 22120
rect 14826 22108 14832 22120
rect 14884 22108 14890 22160
rect 16684 22148 16712 22188
rect 17494 22176 17500 22228
rect 17552 22176 17558 22228
rect 18782 22176 18788 22228
rect 18840 22216 18846 22228
rect 18840 22188 23428 22216
rect 18840 22176 18846 22188
rect 17678 22148 17684 22160
rect 16684 22120 17684 22148
rect 17678 22108 17684 22120
rect 17736 22108 17742 22160
rect 20162 22108 20168 22160
rect 20220 22148 20226 22160
rect 20349 22151 20407 22157
rect 20349 22148 20361 22151
rect 20220 22120 20361 22148
rect 20220 22108 20226 22120
rect 20349 22117 20361 22120
rect 20395 22117 20407 22151
rect 21818 22148 21824 22160
rect 20349 22111 20407 22117
rect 21284 22120 21824 22148
rect 21284 22092 21312 22120
rect 21818 22108 21824 22120
rect 21876 22108 21882 22160
rect 22002 22108 22008 22160
rect 22060 22108 22066 22160
rect 23400 22148 23428 22188
rect 23474 22176 23480 22228
rect 23532 22176 23538 22228
rect 24854 22176 24860 22228
rect 24912 22216 24918 22228
rect 25774 22216 25780 22228
rect 24912 22188 25780 22216
rect 24912 22176 24918 22188
rect 25774 22176 25780 22188
rect 25832 22216 25838 22228
rect 26326 22216 26332 22228
rect 25832 22188 26332 22216
rect 25832 22176 25838 22188
rect 26326 22176 26332 22188
rect 26384 22176 26390 22228
rect 28166 22176 28172 22228
rect 28224 22216 28230 22228
rect 28224 22188 30696 22216
rect 28224 22176 28230 22188
rect 24486 22148 24492 22160
rect 23400 22120 24492 22148
rect 24486 22108 24492 22120
rect 24544 22148 24550 22160
rect 25590 22148 25596 22160
rect 24544 22120 24992 22148
rect 24544 22108 24550 22120
rect 10410 22080 10416 22092
rect 10244 22052 10416 22080
rect 10410 22040 10416 22052
rect 10468 22040 10474 22092
rect 10502 22040 10508 22092
rect 10560 22089 10566 22092
rect 10560 22083 10588 22089
rect 10576 22049 10588 22083
rect 11974 22080 11980 22092
rect 10560 22043 10588 22049
rect 11532 22052 11980 22080
rect 10560 22040 10566 22043
rect 5718 21972 5724 22024
rect 5776 21972 5782 22024
rect 5810 21972 5816 22024
rect 5868 22012 5874 22024
rect 6086 22012 6092 22024
rect 5868 21984 6092 22012
rect 5868 21972 5874 21984
rect 6086 21972 6092 21984
rect 6144 21972 6150 22024
rect 7098 21972 7104 22024
rect 7156 21972 7162 22024
rect 9674 21972 9680 22024
rect 9732 21972 9738 22024
rect 10686 21972 10692 22024
rect 10744 21972 10750 22024
rect 11532 22021 11560 22052
rect 11974 22040 11980 22052
rect 12032 22080 12038 22092
rect 12032 22052 16436 22080
rect 12032 22040 12038 22052
rect 11517 22015 11575 22021
rect 11517 21981 11529 22015
rect 11563 21981 11575 22015
rect 11517 21975 11575 21981
rect 13449 22015 13507 22021
rect 13449 21981 13461 22015
rect 13495 22012 13507 22015
rect 13906 22012 13912 22024
rect 13495 21984 13912 22012
rect 13495 21981 13507 21984
rect 13449 21975 13507 21981
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 14093 22015 14151 22021
rect 14093 21981 14105 22015
rect 14139 22012 14151 22015
rect 14642 22012 14648 22024
rect 14139 21984 14648 22012
rect 14139 21981 14151 21984
rect 14093 21975 14151 21981
rect 14642 21972 14648 21984
rect 14700 21972 14706 22024
rect 16408 22021 16436 22052
rect 18690 22040 18696 22092
rect 18748 22080 18754 22092
rect 19150 22080 19156 22092
rect 18748 22052 19156 22080
rect 18748 22040 18754 22052
rect 19150 22040 19156 22052
rect 19208 22040 19214 22092
rect 19886 22040 19892 22092
rect 19944 22040 19950 22092
rect 20622 22040 20628 22092
rect 20680 22040 20686 22092
rect 20714 22040 20720 22092
rect 20772 22089 20778 22092
rect 20772 22083 20800 22089
rect 20788 22049 20800 22083
rect 20772 22043 20800 22049
rect 20901 22083 20959 22089
rect 20901 22049 20913 22083
rect 20947 22080 20959 22083
rect 21082 22080 21088 22092
rect 20947 22052 21088 22080
rect 20947 22049 20959 22052
rect 20901 22043 20959 22049
rect 20772 22040 20778 22043
rect 21082 22040 21088 22052
rect 21140 22040 21146 22092
rect 21266 22040 21272 22092
rect 21324 22040 21330 22092
rect 21545 22083 21603 22089
rect 21545 22049 21557 22083
rect 21591 22080 21603 22083
rect 22020 22080 22048 22108
rect 21591 22052 22048 22080
rect 21591 22049 21603 22052
rect 21545 22043 21603 22049
rect 23934 22040 23940 22092
rect 23992 22040 23998 22092
rect 24121 22083 24179 22089
rect 24121 22049 24133 22083
rect 24167 22080 24179 22083
rect 24670 22080 24676 22092
rect 24167 22052 24676 22080
rect 24167 22049 24179 22052
rect 24121 22043 24179 22049
rect 24670 22040 24676 22052
rect 24728 22040 24734 22092
rect 24762 22040 24768 22092
rect 24820 22080 24826 22092
rect 24964 22089 24992 22120
rect 25148 22120 25596 22148
rect 25148 22089 25176 22120
rect 25590 22108 25596 22120
rect 25648 22108 25654 22160
rect 30668 22148 30696 22188
rect 31202 22176 31208 22228
rect 31260 22176 31266 22228
rect 34701 22219 34759 22225
rect 34701 22185 34713 22219
rect 34747 22216 34759 22219
rect 35710 22216 35716 22228
rect 34747 22188 35716 22216
rect 34747 22185 34759 22188
rect 34701 22179 34759 22185
rect 35710 22176 35716 22188
rect 35768 22176 35774 22228
rect 38470 22176 38476 22228
rect 38528 22216 38534 22228
rect 38657 22219 38715 22225
rect 38657 22216 38669 22219
rect 38528 22188 38669 22216
rect 38528 22176 38534 22188
rect 38657 22185 38669 22188
rect 38703 22185 38715 22219
rect 38657 22179 38715 22185
rect 38746 22176 38752 22228
rect 38804 22216 38810 22228
rect 38933 22219 38991 22225
rect 38933 22216 38945 22219
rect 38804 22188 38945 22216
rect 38804 22176 38810 22188
rect 38933 22185 38945 22188
rect 38979 22216 38991 22219
rect 43346 22216 43352 22228
rect 38979 22188 43352 22216
rect 38979 22185 38991 22188
rect 38933 22179 38991 22185
rect 43346 22176 43352 22188
rect 43404 22176 43410 22228
rect 30668 22120 31800 22148
rect 24949 22083 25007 22089
rect 24820 22052 24900 22080
rect 24820 22040 24826 22052
rect 16393 22015 16451 22021
rect 16393 21981 16405 22015
rect 16439 22012 16451 22015
rect 16758 22012 16764 22024
rect 16439 21984 16764 22012
rect 16439 21981 16451 21984
rect 16393 21975 16451 21981
rect 16758 21972 16764 21984
rect 16816 21972 16822 22024
rect 17405 22015 17463 22021
rect 17405 21981 17417 22015
rect 17451 22012 17463 22015
rect 18782 22012 18788 22024
rect 17451 21984 18788 22012
rect 17451 21981 17463 21984
rect 17405 21975 17463 21981
rect 18782 21972 18788 21984
rect 18840 21972 18846 22024
rect 19702 21972 19708 22024
rect 19760 21972 19766 22024
rect 22005 22015 22063 22021
rect 22005 21981 22017 22015
rect 22051 22012 22063 22015
rect 22830 22012 22836 22024
rect 22051 21984 22836 22012
rect 22051 21981 22063 21984
rect 22005 21975 22063 21981
rect 22830 21972 22836 21984
rect 22888 22012 22894 22024
rect 24302 22012 24308 22024
rect 22888 21984 24308 22012
rect 22888 21972 22894 21984
rect 24302 21972 24308 21984
rect 24360 21972 24366 22024
rect 24872 22021 24900 22052
rect 24949 22049 24961 22083
rect 24995 22049 25007 22083
rect 24949 22043 25007 22049
rect 25133 22083 25191 22089
rect 25133 22049 25145 22083
rect 25179 22049 25191 22083
rect 25133 22043 25191 22049
rect 25958 22040 25964 22092
rect 26016 22040 26022 22092
rect 26050 22040 26056 22092
rect 26108 22080 26114 22092
rect 26237 22083 26295 22089
rect 26237 22080 26249 22083
rect 26108 22052 26249 22080
rect 26108 22040 26114 22052
rect 26237 22049 26249 22052
rect 26283 22049 26295 22083
rect 26237 22043 26295 22049
rect 27062 22040 27068 22092
rect 27120 22040 27126 22092
rect 31294 22040 31300 22092
rect 31352 22080 31358 22092
rect 31772 22089 31800 22120
rect 34606 22108 34612 22160
rect 34664 22148 34670 22160
rect 35066 22148 35072 22160
rect 34664 22120 35072 22148
rect 34664 22108 34670 22120
rect 35066 22108 35072 22120
rect 35124 22108 35130 22160
rect 36262 22108 36268 22160
rect 36320 22148 36326 22160
rect 36906 22148 36912 22160
rect 36320 22120 36912 22148
rect 36320 22108 36326 22120
rect 36906 22108 36912 22120
rect 36964 22108 36970 22160
rect 39850 22148 39856 22160
rect 38856 22120 39856 22148
rect 31665 22083 31723 22089
rect 31665 22080 31677 22083
rect 31352 22052 31677 22080
rect 31352 22040 31358 22052
rect 31665 22049 31677 22052
rect 31711 22049 31723 22083
rect 31665 22043 31723 22049
rect 31757 22083 31815 22089
rect 31757 22049 31769 22083
rect 31803 22080 31815 22083
rect 31803 22052 31837 22080
rect 32324 22052 34100 22080
rect 31803 22049 31815 22052
rect 31757 22043 31815 22049
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 21981 24915 22015
rect 24857 21975 24915 21981
rect 25317 22015 25375 22021
rect 25317 21981 25329 22015
rect 25363 22012 25375 22015
rect 25406 22012 25412 22024
rect 25363 21984 25412 22012
rect 25363 21981 25375 21984
rect 25317 21975 25375 21981
rect 7438 21947 7496 21953
rect 7438 21944 7450 21947
rect 3896 21916 4936 21944
rect 6932 21916 7450 21944
rect 2593 21879 2651 21885
rect 2593 21845 2605 21879
rect 2639 21845 2651 21879
rect 2593 21839 2651 21845
rect 3053 21879 3111 21885
rect 3053 21845 3065 21879
rect 3099 21876 3111 21879
rect 3694 21876 3700 21888
rect 3099 21848 3700 21876
rect 3099 21845 3111 21848
rect 3053 21839 3111 21845
rect 3694 21836 3700 21848
rect 3752 21876 3758 21888
rect 5810 21876 5816 21888
rect 3752 21848 5816 21876
rect 3752 21836 3758 21848
rect 5810 21836 5816 21848
rect 5868 21836 5874 21888
rect 6932 21885 6960 21916
rect 7438 21913 7450 21916
rect 7484 21913 7496 21947
rect 7438 21907 7496 21913
rect 6917 21879 6975 21885
rect 6917 21845 6929 21879
rect 6963 21845 6975 21879
rect 9692 21876 9720 21972
rect 11882 21904 11888 21956
rect 11940 21944 11946 21956
rect 17310 21944 17316 21956
rect 11940 21916 17316 21944
rect 11940 21904 11946 21916
rect 17310 21904 17316 21916
rect 17368 21944 17374 21956
rect 17773 21947 17831 21953
rect 17773 21944 17785 21947
rect 17368 21916 17785 21944
rect 17368 21904 17374 21916
rect 17773 21913 17785 21916
rect 17819 21913 17831 21947
rect 18322 21944 18328 21956
rect 17773 21907 17831 21913
rect 17880 21916 18328 21944
rect 10686 21876 10692 21888
rect 9692 21848 10692 21876
rect 6917 21839 6975 21845
rect 10686 21836 10692 21848
rect 10744 21836 10750 21888
rect 11330 21836 11336 21888
rect 11388 21836 11394 21888
rect 11790 21836 11796 21888
rect 11848 21836 11854 21888
rect 13630 21836 13636 21888
rect 13688 21876 13694 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 13688 21848 14289 21876
rect 13688 21836 13694 21848
rect 14277 21845 14289 21848
rect 14323 21876 14335 21879
rect 14918 21876 14924 21888
rect 14323 21848 14924 21876
rect 14323 21845 14335 21848
rect 14277 21839 14335 21845
rect 14918 21836 14924 21848
rect 14976 21836 14982 21888
rect 16577 21879 16635 21885
rect 16577 21845 16589 21879
rect 16623 21876 16635 21879
rect 17880 21876 17908 21916
rect 18322 21904 18328 21916
rect 18380 21904 18386 21956
rect 16623 21848 17908 21876
rect 16623 21845 16635 21848
rect 16577 21839 16635 21845
rect 17954 21836 17960 21888
rect 18012 21876 18018 21888
rect 18049 21879 18107 21885
rect 18049 21876 18061 21879
rect 18012 21848 18061 21876
rect 18012 21836 18018 21848
rect 18049 21845 18061 21848
rect 18095 21876 18107 21879
rect 18138 21876 18144 21888
rect 18095 21848 18144 21876
rect 18095 21845 18107 21848
rect 18049 21839 18107 21845
rect 18138 21836 18144 21848
rect 18196 21876 18202 21888
rect 18690 21876 18696 21888
rect 18196 21848 18696 21876
rect 18196 21836 18202 21848
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 19720 21876 19748 21972
rect 22272 21947 22330 21953
rect 22272 21913 22284 21947
rect 22318 21944 22330 21947
rect 22462 21944 22468 21956
rect 22318 21916 22468 21944
rect 22318 21913 22330 21916
rect 22272 21907 22330 21913
rect 22462 21904 22468 21916
rect 22520 21904 22526 21956
rect 23566 21904 23572 21956
rect 23624 21944 23630 21956
rect 23934 21944 23940 21956
rect 23624 21916 23940 21944
rect 23624 21904 23630 21916
rect 23934 21904 23940 21916
rect 23992 21904 23998 21956
rect 24026 21904 24032 21956
rect 24084 21944 24090 21956
rect 24762 21944 24768 21956
rect 24084 21916 24768 21944
rect 24084 21904 24090 21916
rect 24762 21904 24768 21916
rect 24820 21904 24826 21956
rect 25332 21944 25360 21975
rect 25406 21972 25412 21984
rect 25464 21972 25470 22024
rect 25501 22015 25559 22021
rect 25501 21981 25513 22015
rect 25547 21981 25559 22015
rect 25501 21975 25559 21981
rect 24872 21916 25360 21944
rect 23385 21879 23443 21885
rect 23385 21876 23397 21879
rect 19720 21848 23397 21876
rect 23385 21845 23397 21848
rect 23431 21876 23443 21879
rect 23845 21879 23903 21885
rect 23845 21876 23857 21879
rect 23431 21848 23857 21876
rect 23431 21845 23443 21848
rect 23385 21839 23443 21845
rect 23845 21845 23857 21848
rect 23891 21845 23903 21879
rect 23845 21839 23903 21845
rect 24486 21836 24492 21888
rect 24544 21836 24550 21888
rect 24670 21836 24676 21888
rect 24728 21876 24734 21888
rect 24872 21876 24900 21916
rect 24728 21848 24900 21876
rect 24728 21836 24734 21848
rect 24946 21836 24952 21888
rect 25004 21876 25010 21888
rect 25516 21876 25544 21975
rect 26326 21972 26332 22024
rect 26384 22021 26390 22024
rect 26384 22015 26412 22021
rect 26400 21981 26412 22015
rect 26384 21975 26412 21981
rect 26384 21972 26390 21975
rect 26510 21972 26516 22024
rect 26568 21972 26574 22024
rect 27080 22012 27108 22040
rect 27249 22015 27307 22021
rect 27249 22012 27261 22015
rect 27080 21984 27261 22012
rect 27249 21981 27261 21984
rect 27295 22012 27307 22015
rect 28074 22012 28080 22024
rect 27295 21984 28080 22012
rect 27295 21981 27307 21984
rect 27249 21975 27307 21981
rect 28074 21972 28080 21984
rect 28132 22012 28138 22024
rect 28350 22012 28356 22024
rect 28132 21984 28356 22012
rect 28132 21972 28138 21984
rect 28350 21972 28356 21984
rect 28408 21972 28414 22024
rect 28902 21972 28908 22024
rect 28960 21972 28966 22024
rect 29730 21972 29736 22024
rect 29788 21972 29794 22024
rect 30006 22021 30012 22024
rect 30000 21975 30012 22021
rect 30006 21972 30012 21975
rect 30064 21972 30070 22024
rect 27516 21947 27574 21953
rect 27516 21913 27528 21947
rect 27562 21944 27574 21947
rect 27798 21944 27804 21956
rect 27562 21916 27804 21944
rect 27562 21913 27574 21916
rect 27516 21907 27574 21913
rect 27798 21904 27804 21916
rect 27856 21904 27862 21956
rect 28534 21904 28540 21956
rect 28592 21944 28598 21956
rect 32324 21944 32352 22052
rect 33778 21972 33784 22024
rect 33836 22012 33842 22024
rect 33962 22012 33968 22024
rect 33836 21984 33968 22012
rect 33836 21972 33842 21984
rect 33962 21972 33968 21984
rect 34020 21972 34026 22024
rect 34072 22012 34100 22052
rect 35250 22040 35256 22092
rect 35308 22040 35314 22092
rect 35342 22040 35348 22092
rect 35400 22080 35406 22092
rect 36354 22080 36360 22092
rect 35400 22052 36360 22080
rect 35400 22040 35406 22052
rect 36354 22040 36360 22052
rect 36412 22040 36418 22092
rect 36924 22080 36952 22108
rect 38856 22089 38884 22120
rect 39850 22108 39856 22120
rect 39908 22108 39914 22160
rect 42518 22108 42524 22160
rect 42576 22148 42582 22160
rect 42797 22151 42855 22157
rect 42576 22120 42748 22148
rect 42576 22108 42582 22120
rect 37001 22083 37059 22089
rect 37001 22080 37013 22083
rect 36924 22052 37013 22080
rect 37001 22049 37013 22052
rect 37047 22049 37059 22083
rect 37001 22043 37059 22049
rect 38841 22083 38899 22089
rect 38841 22049 38853 22083
rect 38887 22049 38899 22083
rect 39482 22080 39488 22092
rect 38841 22043 38899 22049
rect 39132 22052 39488 22080
rect 39132 22046 39160 22052
rect 35069 22015 35127 22021
rect 34072 21984 34744 22012
rect 28592 21916 32352 21944
rect 28592 21904 28598 21916
rect 32398 21904 32404 21956
rect 32456 21944 32462 21956
rect 34606 21944 34612 21956
rect 32456 21916 34612 21944
rect 32456 21904 32462 21916
rect 34606 21904 34612 21916
rect 34664 21904 34670 21956
rect 34716 21944 34744 21984
rect 35069 21981 35081 22015
rect 35115 22012 35127 22015
rect 35158 22012 35164 22024
rect 35115 21984 35164 22012
rect 35115 21981 35127 21984
rect 35069 21975 35127 21981
rect 35158 21972 35164 21984
rect 35216 21972 35222 22024
rect 35268 22012 35296 22040
rect 35434 22012 35440 22024
rect 35268 21984 35440 22012
rect 35434 21972 35440 21984
rect 35492 21972 35498 22024
rect 35710 21972 35716 22024
rect 35768 21972 35774 22024
rect 36725 22015 36783 22021
rect 35820 21984 36584 22012
rect 35820 21944 35848 21984
rect 34716 21916 35848 21944
rect 36556 21944 36584 21984
rect 36725 21981 36737 22015
rect 36771 22012 36783 22015
rect 36906 22012 36912 22024
rect 36771 21984 36912 22012
rect 36771 21981 36783 21984
rect 36725 21975 36783 21981
rect 36906 21972 36912 21984
rect 36964 21972 36970 22024
rect 37185 22015 37243 22021
rect 37185 21981 37197 22015
rect 37231 22012 37243 22015
rect 37366 22012 37372 22024
rect 37231 21984 37372 22012
rect 37231 21981 37243 21984
rect 37185 21975 37243 21981
rect 37366 21972 37372 21984
rect 37424 21972 37430 22024
rect 37461 22015 37519 22021
rect 37461 21981 37473 22015
rect 37507 21981 37519 22015
rect 37461 21975 37519 21981
rect 37476 21944 37504 21975
rect 37550 21972 37556 22024
rect 37608 22012 37614 22024
rect 38746 22012 38752 22024
rect 37608 21984 38752 22012
rect 37608 21972 37614 21984
rect 38746 21972 38752 21984
rect 38804 21972 38810 22024
rect 39040 22022 39160 22046
rect 39482 22040 39488 22052
rect 39540 22040 39546 22092
rect 42720 22080 42748 22120
rect 42797 22117 42809 22151
rect 42843 22148 42855 22151
rect 42886 22148 42892 22160
rect 42843 22120 42892 22148
rect 42843 22117 42855 22120
rect 42797 22111 42855 22117
rect 42886 22108 42892 22120
rect 42944 22108 42950 22160
rect 39592 22052 39896 22080
rect 38948 22018 39160 22022
rect 38948 21994 39068 22018
rect 38657 21947 38715 21953
rect 38657 21944 38669 21947
rect 36556 21916 37504 21944
rect 38212 21916 38669 21944
rect 26142 21876 26148 21888
rect 25004 21848 26148 21876
rect 25004 21836 25010 21848
rect 26142 21836 26148 21848
rect 26200 21836 26206 21888
rect 27157 21879 27215 21885
rect 27157 21845 27169 21879
rect 27203 21876 27215 21879
rect 27338 21876 27344 21888
rect 27203 21848 27344 21876
rect 27203 21845 27215 21848
rect 27157 21839 27215 21845
rect 27338 21836 27344 21848
rect 27396 21836 27402 21888
rect 27614 21836 27620 21888
rect 27672 21876 27678 21888
rect 28629 21879 28687 21885
rect 28629 21876 28641 21879
rect 27672 21848 28641 21876
rect 27672 21836 27678 21848
rect 28629 21845 28641 21848
rect 28675 21845 28687 21879
rect 28629 21839 28687 21845
rect 28718 21836 28724 21888
rect 28776 21836 28782 21888
rect 30374 21836 30380 21888
rect 30432 21876 30438 21888
rect 31113 21879 31171 21885
rect 31113 21876 31125 21879
rect 30432 21848 31125 21876
rect 30432 21836 30438 21848
rect 31113 21845 31125 21848
rect 31159 21876 31171 21879
rect 31573 21879 31631 21885
rect 31573 21876 31585 21879
rect 31159 21848 31585 21876
rect 31159 21845 31171 21848
rect 31113 21839 31171 21845
rect 31573 21845 31585 21848
rect 31619 21845 31631 21879
rect 31573 21839 31631 21845
rect 33962 21836 33968 21888
rect 34020 21876 34026 21888
rect 35161 21879 35219 21885
rect 35161 21876 35173 21879
rect 34020 21848 35173 21876
rect 34020 21836 34026 21848
rect 35161 21845 35173 21848
rect 35207 21845 35219 21879
rect 35161 21839 35219 21845
rect 35529 21879 35587 21885
rect 35529 21845 35541 21879
rect 35575 21876 35587 21879
rect 36078 21876 36084 21888
rect 35575 21848 36084 21876
rect 35575 21845 35587 21848
rect 35529 21839 35587 21845
rect 36078 21836 36084 21848
rect 36136 21836 36142 21888
rect 36354 21836 36360 21888
rect 36412 21836 36418 21888
rect 36630 21836 36636 21888
rect 36688 21876 36694 21888
rect 38212 21885 38240 21916
rect 38657 21913 38669 21916
rect 38703 21944 38715 21947
rect 38838 21944 38844 21956
rect 38703 21916 38844 21944
rect 38703 21913 38715 21916
rect 38657 21907 38715 21913
rect 38838 21904 38844 21916
rect 38896 21904 38902 21956
rect 38948 21944 38976 21994
rect 39025 21947 39083 21953
rect 39025 21944 39037 21947
rect 38948 21916 39037 21944
rect 39025 21913 39037 21916
rect 39071 21913 39083 21947
rect 39025 21907 39083 21913
rect 36817 21879 36875 21885
rect 36817 21876 36829 21879
rect 36688 21848 36829 21876
rect 36688 21836 36694 21848
rect 36817 21845 36829 21848
rect 36863 21845 36875 21879
rect 36817 21839 36875 21845
rect 38197 21879 38255 21885
rect 38197 21845 38209 21879
rect 38243 21845 38255 21879
rect 38197 21839 38255 21845
rect 38562 21836 38568 21888
rect 38620 21876 38626 21888
rect 39485 21879 39543 21885
rect 39485 21876 39497 21879
rect 38620 21848 39497 21876
rect 38620 21836 38626 21848
rect 39485 21845 39497 21848
rect 39531 21876 39543 21879
rect 39592 21876 39620 22052
rect 39868 22021 39896 22052
rect 42352 22052 43116 22080
rect 39669 22015 39727 22021
rect 39669 21981 39681 22015
rect 39715 21981 39727 22015
rect 39669 21975 39727 21981
rect 39853 22015 39911 22021
rect 39853 21981 39865 22015
rect 39899 21981 39911 22015
rect 39853 21975 39911 21981
rect 39531 21848 39620 21876
rect 39684 21876 39712 21975
rect 40034 21972 40040 22024
rect 40092 22012 40098 22024
rect 42352 22021 42380 22052
rect 40129 22015 40187 22021
rect 40129 22012 40141 22015
rect 40092 21984 40141 22012
rect 40092 21972 40098 21984
rect 40129 21981 40141 21984
rect 40175 21981 40187 22015
rect 40129 21975 40187 21981
rect 42337 22015 42395 22021
rect 42337 21981 42349 22015
rect 42383 21981 42395 22015
rect 42337 21975 42395 21981
rect 42426 21972 42432 22024
rect 42484 21972 42490 22024
rect 42610 21972 42616 22024
rect 42668 21972 42674 22024
rect 42702 21972 42708 22024
rect 42760 21972 42766 22024
rect 42794 21972 42800 22024
rect 42852 22021 42858 22024
rect 43088 22021 43116 22052
rect 42852 22012 42859 22021
rect 43073 22015 43131 22021
rect 42852 21984 42897 22012
rect 42852 21975 42859 21984
rect 43073 21981 43085 22015
rect 43119 21981 43131 22015
rect 43073 21975 43131 21981
rect 42852 21972 42858 21975
rect 39942 21876 39948 21888
rect 39684 21848 39948 21876
rect 39531 21845 39543 21848
rect 39485 21839 39543 21845
rect 39942 21836 39948 21848
rect 40000 21836 40006 21888
rect 40865 21879 40923 21885
rect 40865 21845 40877 21879
rect 40911 21876 40923 21879
rect 41598 21876 41604 21888
rect 40911 21848 41604 21876
rect 40911 21845 40923 21848
rect 40865 21839 40923 21845
rect 41598 21836 41604 21848
rect 41656 21836 41662 21888
rect 42150 21836 42156 21888
rect 42208 21836 42214 21888
rect 42444 21876 42472 21972
rect 42981 21947 43039 21953
rect 42981 21944 42993 21947
rect 42904 21916 42993 21944
rect 42904 21876 42932 21916
rect 42981 21913 42993 21916
rect 43027 21913 43039 21947
rect 42981 21907 43039 21913
rect 42444 21848 42932 21876
rect 1104 21786 47104 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 47104 21786
rect 1104 21712 47104 21734
rect 5810 21632 5816 21684
rect 5868 21672 5874 21684
rect 8573 21675 8631 21681
rect 5868 21644 6914 21672
rect 5868 21632 5874 21644
rect 6886 21604 6914 21644
rect 8573 21641 8585 21675
rect 8619 21672 8631 21675
rect 8846 21672 8852 21684
rect 8619 21644 8852 21672
rect 8619 21641 8631 21644
rect 8573 21635 8631 21641
rect 8846 21632 8852 21644
rect 8904 21632 8910 21684
rect 10321 21675 10379 21681
rect 10321 21641 10333 21675
rect 10367 21641 10379 21675
rect 10321 21635 10379 21641
rect 6886 21576 10180 21604
rect 7190 21496 7196 21548
rect 7248 21496 7254 21548
rect 7466 21545 7472 21548
rect 7460 21499 7472 21545
rect 7466 21496 7472 21499
rect 7524 21496 7530 21548
rect 10152 21468 10180 21576
rect 10229 21539 10287 21545
rect 10229 21505 10241 21539
rect 10275 21536 10287 21539
rect 10336 21536 10364 21635
rect 10778 21632 10784 21684
rect 10836 21632 10842 21684
rect 11330 21632 11336 21684
rect 11388 21672 11394 21684
rect 21545 21675 21603 21681
rect 21545 21672 21557 21675
rect 11388 21644 21557 21672
rect 11388 21632 11394 21644
rect 21545 21641 21557 21644
rect 21591 21641 21603 21675
rect 23842 21672 23848 21684
rect 21545 21635 21603 21641
rect 22066 21644 23848 21672
rect 19242 21564 19248 21616
rect 19300 21564 19306 21616
rect 22066 21604 22094 21644
rect 23842 21632 23848 21644
rect 23900 21632 23906 21684
rect 24489 21675 24547 21681
rect 24489 21641 24501 21675
rect 24535 21672 24547 21675
rect 24578 21672 24584 21684
rect 24535 21644 24584 21672
rect 24535 21641 24547 21644
rect 24489 21635 24547 21641
rect 24578 21632 24584 21644
rect 24636 21632 24642 21684
rect 24762 21632 24768 21684
rect 24820 21672 24826 21684
rect 26605 21675 26663 21681
rect 26605 21672 26617 21675
rect 24820 21644 26617 21672
rect 24820 21632 24826 21644
rect 26605 21641 26617 21644
rect 26651 21641 26663 21675
rect 26605 21635 26663 21641
rect 27338 21632 27344 21684
rect 27396 21632 27402 21684
rect 27798 21632 27804 21684
rect 27856 21632 27862 21684
rect 32398 21672 32404 21684
rect 28276 21644 32404 21672
rect 24213 21607 24271 21613
rect 19352 21576 22094 21604
rect 22388 21576 22692 21604
rect 10275 21508 10364 21536
rect 10275 21505 10287 21508
rect 10229 21499 10287 21505
rect 10686 21496 10692 21548
rect 10744 21496 10750 21548
rect 14550 21536 14556 21548
rect 10796 21508 14556 21536
rect 10796 21468 10824 21508
rect 14550 21496 14556 21508
rect 14608 21496 14614 21548
rect 15841 21539 15899 21545
rect 15841 21505 15853 21539
rect 15887 21536 15899 21539
rect 16114 21536 16120 21548
rect 15887 21508 16120 21536
rect 15887 21505 15899 21508
rect 15841 21499 15899 21505
rect 16114 21496 16120 21508
rect 16172 21536 16178 21548
rect 16172 21508 17448 21536
rect 16172 21496 16178 21508
rect 10152 21440 10824 21468
rect 10873 21471 10931 21477
rect 10873 21437 10885 21471
rect 10919 21437 10931 21471
rect 10873 21431 10931 21437
rect 10410 21360 10416 21412
rect 10468 21400 10474 21412
rect 10888 21400 10916 21431
rect 15746 21428 15752 21480
rect 15804 21468 15810 21480
rect 16025 21471 16083 21477
rect 16025 21468 16037 21471
rect 15804 21440 16037 21468
rect 15804 21428 15810 21440
rect 16025 21437 16037 21440
rect 16071 21437 16083 21471
rect 16025 21431 16083 21437
rect 17126 21428 17132 21480
rect 17184 21428 17190 21480
rect 17218 21428 17224 21480
rect 17276 21468 17282 21480
rect 17313 21471 17371 21477
rect 17313 21468 17325 21471
rect 17276 21440 17325 21468
rect 17276 21428 17282 21440
rect 17313 21437 17325 21440
rect 17359 21437 17371 21471
rect 17420 21468 17448 21508
rect 18046 21496 18052 21548
rect 18104 21496 18110 21548
rect 18138 21496 18144 21548
rect 18196 21545 18202 21548
rect 18196 21539 18224 21545
rect 18212 21505 18224 21539
rect 18196 21499 18224 21505
rect 18196 21496 18202 21499
rect 18322 21496 18328 21548
rect 18380 21496 18386 21548
rect 19058 21496 19064 21548
rect 19116 21536 19122 21548
rect 19352 21536 19380 21576
rect 19116 21508 19380 21536
rect 19116 21496 19122 21508
rect 19886 21496 19892 21548
rect 19944 21536 19950 21548
rect 21361 21539 21419 21545
rect 19944 21508 21312 21536
rect 19944 21496 19950 21508
rect 21284 21468 21312 21508
rect 21361 21505 21373 21539
rect 21407 21536 21419 21539
rect 21450 21536 21456 21548
rect 21407 21508 21456 21536
rect 21407 21505 21419 21508
rect 21361 21499 21419 21505
rect 21450 21496 21456 21508
rect 21508 21496 21514 21548
rect 21634 21496 21640 21548
rect 21692 21536 21698 21548
rect 21818 21536 21824 21548
rect 21692 21508 21824 21536
rect 21692 21496 21698 21508
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 22388 21545 22416 21576
rect 22554 21545 22560 21548
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22525 21539 22560 21545
rect 22525 21505 22537 21539
rect 22525 21499 22560 21505
rect 22554 21496 22560 21499
rect 22612 21496 22618 21548
rect 22094 21468 22100 21480
rect 17420 21440 20944 21468
rect 21284 21440 22100 21468
rect 17313 21431 17371 21437
rect 10468 21372 10916 21400
rect 17773 21403 17831 21409
rect 10468 21360 10474 21372
rect 17773 21369 17785 21403
rect 17819 21400 17831 21403
rect 17862 21400 17868 21412
rect 17819 21372 17868 21400
rect 17819 21369 17831 21372
rect 17773 21363 17831 21369
rect 17862 21360 17868 21372
rect 17920 21360 17926 21412
rect 18969 21403 19027 21409
rect 18969 21369 18981 21403
rect 19015 21400 19027 21403
rect 19521 21403 19579 21409
rect 19521 21400 19533 21403
rect 19015 21372 19533 21400
rect 19015 21369 19027 21372
rect 18969 21363 19027 21369
rect 19521 21369 19533 21372
rect 19567 21369 19579 21403
rect 19521 21363 19579 21369
rect 10045 21335 10103 21341
rect 10045 21301 10057 21335
rect 10091 21332 10103 21335
rect 10134 21332 10140 21344
rect 10091 21304 10140 21332
rect 10091 21301 10103 21304
rect 10045 21295 10103 21301
rect 10134 21292 10140 21304
rect 10192 21292 10198 21344
rect 15838 21292 15844 21344
rect 15896 21332 15902 21344
rect 18138 21332 18144 21344
rect 15896 21304 18144 21332
rect 15896 21292 15902 21304
rect 18138 21292 18144 21304
rect 18196 21292 18202 21344
rect 19705 21335 19763 21341
rect 19705 21301 19717 21335
rect 19751 21332 19763 21335
rect 20806 21332 20812 21344
rect 19751 21304 20812 21332
rect 19751 21301 19763 21304
rect 19705 21295 19763 21301
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 20916 21332 20944 21440
rect 22094 21428 22100 21440
rect 22152 21428 22158 21480
rect 22186 21428 22192 21480
rect 22244 21428 22250 21480
rect 22664 21468 22692 21576
rect 24213 21573 24225 21607
rect 24259 21604 24271 21607
rect 24394 21604 24400 21616
rect 24259 21576 24400 21604
rect 24259 21573 24271 21576
rect 24213 21567 24271 21573
rect 24394 21564 24400 21576
rect 24452 21564 24458 21616
rect 27433 21607 27491 21613
rect 27433 21573 27445 21607
rect 27479 21604 27491 21607
rect 28276 21604 28304 21644
rect 32398 21632 32404 21644
rect 32456 21632 32462 21684
rect 32493 21675 32551 21681
rect 32493 21641 32505 21675
rect 32539 21641 32551 21675
rect 32493 21635 32551 21641
rect 27479 21576 28304 21604
rect 28344 21607 28402 21613
rect 27479 21573 27491 21576
rect 27433 21567 27491 21573
rect 28344 21573 28356 21607
rect 28390 21604 28402 21607
rect 28718 21604 28724 21616
rect 28390 21576 28724 21604
rect 28390 21573 28402 21576
rect 28344 21567 28402 21573
rect 28718 21564 28724 21576
rect 28776 21564 28782 21616
rect 29730 21564 29736 21616
rect 29788 21604 29794 21616
rect 31754 21604 31760 21616
rect 29788 21576 31760 21604
rect 29788 21564 29794 21576
rect 31754 21564 31760 21576
rect 31812 21564 31818 21616
rect 22741 21539 22799 21545
rect 22741 21505 22753 21539
rect 22787 21536 22799 21539
rect 22922 21536 22928 21548
rect 22787 21508 22928 21536
rect 22787 21505 22799 21508
rect 22741 21499 22799 21505
rect 22922 21496 22928 21508
rect 22980 21496 22986 21548
rect 23845 21539 23903 21545
rect 23845 21505 23857 21539
rect 23891 21536 23903 21539
rect 24302 21536 24308 21548
rect 23891 21508 24308 21536
rect 23891 21505 23903 21508
rect 23845 21499 23903 21505
rect 24302 21496 24308 21508
rect 24360 21496 24366 21548
rect 24486 21496 24492 21548
rect 24544 21536 24550 21548
rect 24673 21539 24731 21545
rect 24673 21536 24685 21539
rect 24544 21508 24685 21536
rect 24544 21496 24550 21508
rect 24673 21505 24685 21508
rect 24719 21505 24731 21539
rect 24673 21499 24731 21505
rect 24762 21496 24768 21548
rect 24820 21496 24826 21548
rect 24872 21508 25084 21536
rect 24872 21468 24900 21508
rect 25056 21480 25084 21508
rect 25682 21496 25688 21548
rect 25740 21496 25746 21548
rect 25774 21496 25780 21548
rect 25832 21545 25838 21548
rect 25832 21539 25860 21545
rect 25848 21505 25860 21539
rect 25832 21499 25860 21505
rect 25832 21496 25838 21499
rect 25958 21496 25964 21548
rect 26016 21496 26022 21548
rect 27982 21496 27988 21548
rect 28040 21496 28046 21548
rect 28074 21496 28080 21548
rect 28132 21496 28138 21548
rect 30742 21536 30748 21548
rect 28184 21508 30748 21536
rect 22664 21440 24900 21468
rect 24946 21428 24952 21480
rect 25004 21428 25010 21480
rect 25038 21428 25044 21480
rect 25096 21428 25102 21480
rect 27525 21471 27583 21477
rect 27525 21437 27537 21471
rect 27571 21468 27583 21471
rect 28184 21468 28212 21508
rect 30742 21496 30748 21508
rect 30800 21496 30806 21548
rect 32401 21539 32459 21545
rect 32401 21505 32413 21539
rect 32447 21536 32459 21539
rect 32508 21536 32536 21635
rect 32950 21632 32956 21684
rect 33008 21632 33014 21684
rect 33594 21672 33600 21684
rect 33428 21644 33600 21672
rect 32447 21508 32536 21536
rect 32861 21539 32919 21545
rect 32447 21505 32459 21508
rect 32401 21499 32459 21505
rect 32861 21505 32873 21539
rect 32907 21536 32919 21539
rect 33318 21536 33324 21548
rect 32907 21508 33324 21536
rect 32907 21505 32919 21508
rect 32861 21499 32919 21505
rect 33318 21496 33324 21508
rect 33376 21496 33382 21548
rect 33428 21545 33456 21644
rect 33594 21632 33600 21644
rect 33652 21672 33658 21684
rect 35250 21672 35256 21684
rect 33652 21644 35256 21672
rect 33652 21632 33658 21644
rect 35250 21632 35256 21644
rect 35308 21672 35314 21684
rect 36725 21675 36783 21681
rect 36725 21672 36737 21675
rect 35308 21644 36737 21672
rect 35308 21632 35314 21644
rect 36725 21641 36737 21644
rect 36771 21641 36783 21675
rect 36725 21635 36783 21641
rect 36817 21675 36875 21681
rect 36817 21641 36829 21675
rect 36863 21641 36875 21675
rect 36817 21635 36875 21641
rect 35612 21607 35670 21613
rect 35612 21573 35624 21607
rect 35658 21604 35670 21607
rect 36078 21604 36084 21616
rect 35658 21576 36084 21604
rect 35658 21573 35670 21576
rect 35612 21567 35670 21573
rect 36078 21564 36084 21576
rect 36136 21564 36142 21616
rect 36832 21604 36860 21635
rect 36906 21632 36912 21684
rect 36964 21672 36970 21684
rect 38657 21675 38715 21681
rect 38657 21672 38669 21675
rect 36964 21644 38669 21672
rect 36964 21632 36970 21644
rect 38657 21641 38669 21644
rect 38703 21641 38715 21675
rect 38657 21635 38715 21641
rect 38838 21632 38844 21684
rect 38896 21672 38902 21684
rect 40310 21672 40316 21684
rect 38896 21644 40316 21672
rect 38896 21632 38902 21644
rect 40310 21632 40316 21644
rect 40368 21632 40374 21684
rect 37522 21607 37580 21613
rect 37522 21604 37534 21607
rect 36832 21576 37534 21604
rect 37522 21573 37534 21576
rect 37568 21573 37580 21607
rect 37522 21567 37580 21573
rect 38746 21564 38752 21616
rect 38804 21604 38810 21616
rect 39942 21604 39948 21616
rect 38804 21576 39948 21604
rect 38804 21564 38810 21576
rect 39942 21564 39948 21576
rect 40000 21564 40006 21616
rect 42702 21564 42708 21616
rect 42760 21604 42766 21616
rect 42760 21576 43208 21604
rect 42760 21564 42766 21576
rect 43180 21548 43208 21576
rect 33413 21539 33471 21545
rect 33413 21505 33425 21539
rect 33459 21505 33471 21539
rect 33413 21499 33471 21505
rect 35342 21496 35348 21548
rect 35400 21496 35406 21548
rect 36354 21496 36360 21548
rect 36412 21536 36418 21548
rect 37001 21539 37059 21545
rect 37001 21536 37013 21539
rect 36412 21508 37013 21536
rect 36412 21496 36418 21508
rect 37001 21505 37013 21508
rect 37047 21505 37059 21539
rect 37001 21499 37059 21505
rect 39758 21496 39764 21548
rect 39816 21536 39822 21548
rect 39853 21539 39911 21545
rect 39853 21536 39865 21539
rect 39816 21508 39865 21536
rect 39816 21496 39822 21508
rect 39853 21505 39865 21508
rect 39899 21505 39911 21539
rect 41049 21539 41107 21545
rect 41049 21536 41061 21539
rect 39853 21499 39911 21505
rect 40328 21508 41061 21536
rect 27571 21440 28212 21468
rect 27571 21437 27583 21440
rect 27525 21431 27583 21437
rect 21177 21403 21235 21409
rect 21177 21369 21189 21403
rect 21223 21400 21235 21403
rect 22462 21400 22468 21412
rect 21223 21372 22468 21400
rect 21223 21369 21235 21372
rect 21177 21363 21235 21369
rect 22462 21360 22468 21372
rect 22520 21360 22526 21412
rect 22649 21403 22707 21409
rect 22649 21369 22661 21403
rect 22695 21400 22707 21403
rect 22738 21400 22744 21412
rect 22695 21372 22744 21400
rect 22695 21369 22707 21372
rect 22649 21363 22707 21369
rect 22738 21360 22744 21372
rect 22796 21360 22802 21412
rect 23934 21360 23940 21412
rect 23992 21400 23998 21412
rect 25409 21403 25467 21409
rect 25409 21400 25421 21403
rect 23992 21372 25421 21400
rect 23992 21360 23998 21372
rect 25409 21369 25421 21372
rect 25455 21369 25467 21403
rect 26973 21403 27031 21409
rect 26973 21400 26985 21403
rect 25409 21363 25467 21369
rect 26344 21372 26985 21400
rect 22278 21332 22284 21344
rect 20916 21304 22284 21332
rect 22278 21292 22284 21304
rect 22336 21292 22342 21344
rect 22554 21292 22560 21344
rect 22612 21332 22618 21344
rect 26344 21332 26372 21372
rect 26973 21369 26985 21372
rect 27019 21369 27031 21403
rect 26973 21363 27031 21369
rect 27154 21360 27160 21412
rect 27212 21400 27218 21412
rect 27540 21400 27568 21431
rect 33042 21428 33048 21480
rect 33100 21468 33106 21480
rect 33226 21468 33232 21480
rect 33100 21440 33232 21468
rect 33100 21428 33106 21440
rect 33226 21428 33232 21440
rect 33284 21428 33290 21480
rect 33597 21471 33655 21477
rect 33597 21437 33609 21471
rect 33643 21468 33655 21471
rect 33686 21468 33692 21480
rect 33643 21440 33692 21468
rect 33643 21437 33655 21440
rect 33597 21431 33655 21437
rect 33686 21428 33692 21440
rect 33744 21428 33750 21480
rect 34054 21428 34060 21480
rect 34112 21428 34118 21480
rect 34330 21428 34336 21480
rect 34388 21428 34394 21480
rect 34514 21477 34520 21480
rect 34471 21471 34520 21477
rect 34471 21437 34483 21471
rect 34517 21437 34520 21471
rect 34471 21431 34520 21437
rect 34514 21428 34520 21431
rect 34572 21428 34578 21480
rect 34609 21471 34667 21477
rect 34609 21437 34621 21471
rect 34655 21468 34667 21471
rect 34974 21468 34980 21480
rect 34655 21440 34980 21468
rect 34655 21437 34667 21440
rect 34609 21431 34667 21437
rect 34974 21428 34980 21440
rect 35032 21428 35038 21480
rect 36446 21428 36452 21480
rect 36504 21468 36510 21480
rect 36814 21468 36820 21480
rect 36504 21440 36820 21468
rect 36504 21428 36510 21440
rect 36814 21428 36820 21440
rect 36872 21468 36878 21480
rect 37277 21471 37335 21477
rect 37277 21468 37289 21471
rect 36872 21440 37289 21468
rect 36872 21428 36878 21440
rect 37277 21437 37289 21440
rect 37323 21437 37335 21471
rect 38838 21468 38844 21480
rect 37277 21431 37335 21437
rect 38626 21440 38844 21468
rect 27212 21372 27568 21400
rect 27212 21360 27218 21372
rect 29454 21360 29460 21412
rect 29512 21360 29518 21412
rect 32950 21360 32956 21412
rect 33008 21400 33014 21412
rect 33962 21400 33968 21412
rect 33008 21372 33968 21400
rect 33008 21360 33014 21372
rect 33962 21360 33968 21372
rect 34020 21360 34026 21412
rect 22612 21304 26372 21332
rect 22612 21292 22618 21304
rect 26510 21292 26516 21344
rect 26568 21332 26574 21344
rect 31018 21332 31024 21344
rect 26568 21304 31024 21332
rect 26568 21292 26574 21304
rect 31018 21292 31024 21304
rect 31076 21292 31082 21344
rect 32214 21292 32220 21344
rect 32272 21292 32278 21344
rect 33502 21292 33508 21344
rect 33560 21332 33566 21344
rect 35253 21335 35311 21341
rect 35253 21332 35265 21335
rect 33560 21304 35265 21332
rect 33560 21292 33566 21304
rect 35253 21301 35265 21304
rect 35299 21301 35311 21335
rect 35253 21295 35311 21301
rect 36630 21292 36636 21344
rect 36688 21332 36694 21344
rect 38626 21332 38654 21440
rect 38838 21428 38844 21440
rect 38896 21428 38902 21480
rect 40328 21477 40356 21508
rect 41049 21505 41061 21508
rect 41095 21536 41107 21539
rect 41598 21536 41604 21548
rect 41095 21508 41604 21536
rect 41095 21505 41107 21508
rect 41049 21499 41107 21505
rect 41598 21496 41604 21508
rect 41656 21496 41662 21548
rect 42150 21496 42156 21548
rect 42208 21536 42214 21548
rect 42613 21539 42671 21545
rect 42613 21536 42625 21539
rect 42208 21508 42625 21536
rect 42208 21496 42214 21508
rect 42613 21505 42625 21508
rect 42659 21505 42671 21539
rect 42613 21499 42671 21505
rect 43162 21496 43168 21548
rect 43220 21496 43226 21548
rect 43254 21496 43260 21548
rect 43312 21496 43318 21548
rect 46109 21539 46167 21545
rect 46109 21505 46121 21539
rect 46155 21536 46167 21539
rect 46750 21536 46756 21548
rect 46155 21508 46756 21536
rect 46155 21505 46167 21508
rect 46109 21499 46167 21505
rect 46750 21496 46756 21508
rect 46808 21496 46814 21548
rect 40313 21471 40371 21477
rect 40313 21437 40325 21471
rect 40359 21437 40371 21471
rect 40313 21431 40371 21437
rect 41690 21428 41696 21480
rect 41748 21468 41754 21480
rect 42705 21471 42763 21477
rect 42705 21468 42717 21471
rect 41748 21440 42717 21468
rect 41748 21428 41754 21440
rect 42705 21437 42717 21440
rect 42751 21437 42763 21471
rect 42705 21431 42763 21437
rect 42797 21471 42855 21477
rect 42797 21437 42809 21471
rect 42843 21437 42855 21471
rect 42797 21431 42855 21437
rect 42889 21471 42947 21477
rect 42889 21437 42901 21471
rect 42935 21468 42947 21471
rect 43898 21468 43904 21480
rect 42935 21440 43904 21468
rect 42935 21437 42947 21440
rect 42889 21431 42947 21437
rect 42610 21360 42616 21412
rect 42668 21400 42674 21412
rect 42812 21400 42840 21431
rect 43898 21428 43904 21440
rect 43956 21428 43962 21480
rect 43165 21403 43223 21409
rect 43165 21400 43177 21403
rect 42668 21372 43177 21400
rect 42668 21360 42674 21372
rect 43165 21369 43177 21372
rect 43211 21369 43223 21403
rect 43165 21363 43223 21369
rect 36688 21304 38654 21332
rect 36688 21292 36694 21304
rect 39574 21292 39580 21344
rect 39632 21332 39638 21344
rect 39945 21335 40003 21341
rect 39945 21332 39957 21335
rect 39632 21304 39957 21332
rect 39632 21292 39638 21304
rect 39945 21301 39957 21304
rect 39991 21301 40003 21335
rect 39945 21295 40003 21301
rect 40402 21292 40408 21344
rect 40460 21332 40466 21344
rect 40954 21332 40960 21344
rect 40460 21304 40960 21332
rect 40460 21292 40466 21304
rect 40954 21292 40960 21304
rect 41012 21332 41018 21344
rect 41233 21335 41291 21341
rect 41233 21332 41245 21335
rect 41012 21304 41245 21332
rect 41012 21292 41018 21304
rect 41233 21301 41245 21304
rect 41279 21301 41291 21335
rect 41233 21295 41291 21301
rect 41874 21292 41880 21344
rect 41932 21332 41938 21344
rect 42429 21335 42487 21341
rect 42429 21332 42441 21335
rect 41932 21304 42441 21332
rect 41932 21292 41938 21304
rect 42429 21301 42441 21304
rect 42475 21301 42487 21335
rect 42429 21295 42487 21301
rect 45738 21292 45744 21344
rect 45796 21332 45802 21344
rect 45925 21335 45983 21341
rect 45925 21332 45937 21335
rect 45796 21304 45937 21332
rect 45796 21292 45802 21304
rect 45925 21301 45937 21304
rect 45971 21301 45983 21335
rect 45925 21295 45983 21301
rect 1104 21242 47104 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 47104 21242
rect 1104 21168 47104 21190
rect 7466 21088 7472 21140
rect 7524 21088 7530 21140
rect 10686 21088 10692 21140
rect 10744 21128 10750 21140
rect 11425 21131 11483 21137
rect 11425 21128 11437 21131
rect 10744 21100 11437 21128
rect 10744 21088 10750 21100
rect 11425 21097 11437 21100
rect 11471 21097 11483 21131
rect 11425 21091 11483 21097
rect 13906 21088 13912 21140
rect 13964 21128 13970 21140
rect 18046 21128 18052 21140
rect 13964 21100 18052 21128
rect 13964 21088 13970 21100
rect 18046 21088 18052 21100
rect 18104 21088 18110 21140
rect 20806 21088 20812 21140
rect 20864 21088 20870 21140
rect 20898 21088 20904 21140
rect 20956 21128 20962 21140
rect 21177 21131 21235 21137
rect 21177 21128 21189 21131
rect 20956 21100 21189 21128
rect 20956 21088 20962 21100
rect 21177 21097 21189 21100
rect 21223 21097 21235 21131
rect 21177 21091 21235 21097
rect 22462 21088 22468 21140
rect 22520 21128 22526 21140
rect 22922 21128 22928 21140
rect 22520 21100 22928 21128
rect 22520 21088 22526 21100
rect 22922 21088 22928 21100
rect 22980 21088 22986 21140
rect 23842 21088 23848 21140
rect 23900 21128 23906 21140
rect 25958 21128 25964 21140
rect 23900 21100 25964 21128
rect 23900 21088 23906 21100
rect 25958 21088 25964 21100
rect 26016 21088 26022 21140
rect 26050 21088 26056 21140
rect 26108 21128 26114 21140
rect 33502 21128 33508 21140
rect 26108 21100 33508 21128
rect 26108 21088 26114 21100
rect 33502 21088 33508 21100
rect 33560 21088 33566 21140
rect 33962 21088 33968 21140
rect 34020 21128 34026 21140
rect 34885 21131 34943 21137
rect 34885 21128 34897 21131
rect 34020 21100 34897 21128
rect 34020 21088 34026 21100
rect 34885 21097 34897 21100
rect 34931 21097 34943 21131
rect 34885 21091 34943 21097
rect 35250 21088 35256 21140
rect 35308 21128 35314 21140
rect 35526 21128 35532 21140
rect 35308 21100 35532 21128
rect 35308 21088 35314 21100
rect 35526 21088 35532 21100
rect 35584 21088 35590 21140
rect 38105 21131 38163 21137
rect 38105 21097 38117 21131
rect 38151 21128 38163 21131
rect 39666 21128 39672 21140
rect 38151 21100 39672 21128
rect 38151 21097 38163 21100
rect 38105 21091 38163 21097
rect 39666 21088 39672 21100
rect 39724 21088 39730 21140
rect 43898 21088 43904 21140
rect 43956 21088 43962 21140
rect 46014 21088 46020 21140
rect 46072 21128 46078 21140
rect 46290 21128 46296 21140
rect 46072 21100 46296 21128
rect 46072 21088 46078 21100
rect 46290 21088 46296 21100
rect 46348 21128 46354 21140
rect 46385 21131 46443 21137
rect 46385 21128 46397 21131
rect 46348 21100 46397 21128
rect 46348 21088 46354 21100
rect 46385 21097 46397 21100
rect 46431 21097 46443 21131
rect 46385 21091 46443 21097
rect 46750 21088 46756 21140
rect 46808 21088 46814 21140
rect 11882 21020 11888 21072
rect 11940 21020 11946 21072
rect 18690 21020 18696 21072
rect 18748 21060 18754 21072
rect 23934 21060 23940 21072
rect 18748 21032 23940 21060
rect 18748 21020 18754 21032
rect 23934 21020 23940 21032
rect 23992 21020 23998 21072
rect 26142 21020 26148 21072
rect 26200 21060 26206 21072
rect 29454 21060 29460 21072
rect 26200 21032 29460 21060
rect 26200 21020 26206 21032
rect 29454 21020 29460 21032
rect 29512 21020 29518 21072
rect 33318 21020 33324 21072
rect 33376 21060 33382 21072
rect 34514 21060 34520 21072
rect 33376 21032 34520 21060
rect 33376 21020 33382 21032
rect 34514 21020 34520 21032
rect 34572 21020 34578 21072
rect 45925 21063 45983 21069
rect 45925 21060 45937 21063
rect 43732 21032 45937 21060
rect 3237 20995 3295 21001
rect 3237 20961 3249 20995
rect 3283 20992 3295 20995
rect 3786 20992 3792 21004
rect 3283 20964 3792 20992
rect 3283 20961 3295 20964
rect 3237 20955 3295 20961
rect 3786 20952 3792 20964
rect 3844 20952 3850 21004
rect 7190 20952 7196 21004
rect 7248 20992 7254 21004
rect 10045 20995 10103 21001
rect 10045 20992 10057 20995
rect 7248 20964 10057 20992
rect 7248 20952 7254 20964
rect 10045 20961 10057 20964
rect 10091 20961 10103 20995
rect 10045 20955 10103 20961
rect 11422 20952 11428 21004
rect 11480 20992 11486 21004
rect 12161 20995 12219 21001
rect 12161 20992 12173 20995
rect 11480 20964 12173 20992
rect 11480 20952 11486 20964
rect 12161 20961 12173 20964
rect 12207 20992 12219 20995
rect 12250 20992 12256 21004
rect 12207 20964 12256 20992
rect 12207 20961 12219 20964
rect 12161 20955 12219 20961
rect 12250 20952 12256 20964
rect 12308 20952 12314 21004
rect 17218 20952 17224 21004
rect 17276 20952 17282 21004
rect 17586 20952 17592 21004
rect 17644 20992 17650 21004
rect 17681 20995 17739 21001
rect 17681 20992 17693 20995
rect 17644 20964 17693 20992
rect 17644 20952 17650 20964
rect 17681 20961 17693 20964
rect 17727 20961 17739 20995
rect 17681 20955 17739 20961
rect 18233 20995 18291 21001
rect 18233 20961 18245 20995
rect 18279 20992 18291 20995
rect 18966 20992 18972 21004
rect 18279 20964 18972 20992
rect 18279 20961 18291 20964
rect 18233 20955 18291 20961
rect 18966 20952 18972 20964
rect 19024 20952 19030 21004
rect 20349 20995 20407 21001
rect 20349 20961 20361 20995
rect 20395 20992 20407 20995
rect 20395 20964 31754 20992
rect 20395 20961 20407 20964
rect 20349 20955 20407 20961
rect 2317 20927 2375 20933
rect 2317 20893 2329 20927
rect 2363 20924 2375 20927
rect 2363 20896 2636 20924
rect 2363 20893 2375 20896
rect 2317 20887 2375 20893
rect 2130 20748 2136 20800
rect 2188 20748 2194 20800
rect 2608 20797 2636 20896
rect 4798 20884 4804 20936
rect 4856 20924 4862 20936
rect 4985 20927 5043 20933
rect 4985 20924 4997 20927
rect 4856 20896 4997 20924
rect 4856 20884 4862 20896
rect 4985 20893 4997 20896
rect 5031 20893 5043 20927
rect 4985 20887 5043 20893
rect 7653 20927 7711 20933
rect 7653 20893 7665 20927
rect 7699 20924 7711 20927
rect 8478 20924 8484 20936
rect 7699 20896 8484 20924
rect 7699 20893 7711 20896
rect 7653 20887 7711 20893
rect 8478 20884 8484 20896
rect 8536 20884 8542 20936
rect 10134 20884 10140 20936
rect 10192 20924 10198 20936
rect 10301 20927 10359 20933
rect 10301 20924 10313 20927
rect 10192 20896 10313 20924
rect 10192 20884 10198 20896
rect 10301 20893 10313 20896
rect 10347 20893 10359 20927
rect 10301 20887 10359 20893
rect 10594 20884 10600 20936
rect 10652 20924 10658 20936
rect 11701 20927 11759 20933
rect 11701 20924 11713 20927
rect 10652 20896 11713 20924
rect 10652 20884 10658 20896
rect 10980 20868 11008 20896
rect 11701 20893 11713 20896
rect 11747 20893 11759 20927
rect 11701 20887 11759 20893
rect 5252 20859 5310 20865
rect 5252 20825 5264 20859
rect 5298 20856 5310 20859
rect 5350 20856 5356 20868
rect 5298 20828 5356 20856
rect 5298 20825 5310 20828
rect 5252 20819 5310 20825
rect 5350 20816 5356 20828
rect 5408 20816 5414 20868
rect 10962 20816 10968 20868
rect 11020 20816 11026 20868
rect 2593 20791 2651 20797
rect 2593 20757 2605 20791
rect 2639 20757 2651 20791
rect 2593 20751 2651 20757
rect 2958 20748 2964 20800
rect 3016 20748 3022 20800
rect 3050 20748 3056 20800
rect 3108 20788 3114 20800
rect 3970 20788 3976 20800
rect 3108 20760 3976 20788
rect 3108 20748 3114 20760
rect 3970 20748 3976 20760
rect 4028 20748 4034 20800
rect 6362 20748 6368 20800
rect 6420 20748 6426 20800
rect 11716 20788 11744 20887
rect 11882 20884 11888 20936
rect 11940 20924 11946 20936
rect 11977 20927 12035 20933
rect 11977 20924 11989 20927
rect 11940 20896 11989 20924
rect 11940 20884 11946 20896
rect 11977 20893 11989 20896
rect 12023 20893 12035 20927
rect 11977 20887 12035 20893
rect 12526 20884 12532 20936
rect 12584 20924 12590 20936
rect 14461 20927 14519 20933
rect 14461 20924 14473 20927
rect 12584 20896 14473 20924
rect 12584 20884 12590 20896
rect 14461 20893 14473 20896
rect 14507 20893 14519 20927
rect 15286 20924 15292 20936
rect 14461 20887 14519 20893
rect 14568 20896 15292 20924
rect 12796 20859 12854 20865
rect 12796 20825 12808 20859
rect 12842 20856 12854 20859
rect 12986 20856 12992 20868
rect 12842 20828 12992 20856
rect 12842 20825 12854 20828
rect 12796 20819 12854 20825
rect 12986 20816 12992 20828
rect 13044 20816 13050 20868
rect 14568 20788 14596 20896
rect 15286 20884 15292 20896
rect 15344 20924 15350 20936
rect 15933 20927 15991 20933
rect 15933 20924 15945 20927
rect 15344 20896 15945 20924
rect 15344 20884 15350 20896
rect 15933 20893 15945 20896
rect 15979 20893 15991 20927
rect 15933 20887 15991 20893
rect 17037 20927 17095 20933
rect 17037 20893 17049 20927
rect 17083 20924 17095 20927
rect 17126 20924 17132 20936
rect 17083 20896 17132 20924
rect 17083 20893 17095 20896
rect 17037 20887 17095 20893
rect 17126 20884 17132 20896
rect 17184 20884 17190 20936
rect 14734 20865 14740 20868
rect 14728 20819 14740 20865
rect 14734 20816 14740 20819
rect 14792 20816 14798 20868
rect 11716 20760 14596 20788
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 15746 20788 15752 20800
rect 15252 20760 15752 20788
rect 15252 20748 15258 20760
rect 15746 20748 15752 20760
rect 15804 20748 15810 20800
rect 15838 20748 15844 20800
rect 15896 20748 15902 20800
rect 16114 20748 16120 20800
rect 16172 20748 16178 20800
rect 17236 20788 17264 20952
rect 17954 20884 17960 20936
rect 18012 20884 18018 20936
rect 18138 20933 18144 20936
rect 18095 20927 18144 20933
rect 18095 20893 18107 20927
rect 18141 20893 18144 20927
rect 18095 20887 18144 20893
rect 18138 20884 18144 20887
rect 18196 20884 18202 20936
rect 20533 20927 20591 20933
rect 20533 20893 20545 20927
rect 20579 20893 20591 20927
rect 20533 20887 20591 20893
rect 20625 20927 20683 20933
rect 20625 20893 20637 20927
rect 20671 20893 20683 20927
rect 20625 20887 20683 20893
rect 18506 20788 18512 20800
rect 17236 20760 18512 20788
rect 18506 20748 18512 20760
rect 18564 20748 18570 20800
rect 18877 20791 18935 20797
rect 18877 20757 18889 20791
rect 18923 20788 18935 20791
rect 19242 20788 19248 20800
rect 18923 20760 19248 20788
rect 18923 20757 18935 20760
rect 18877 20751 18935 20757
rect 19242 20748 19248 20760
rect 19300 20748 19306 20800
rect 20548 20788 20576 20887
rect 20640 20856 20668 20887
rect 20714 20884 20720 20936
rect 20772 20924 20778 20936
rect 20901 20927 20959 20933
rect 20901 20924 20913 20927
rect 20772 20896 20913 20924
rect 20772 20884 20778 20896
rect 20901 20893 20913 20896
rect 20947 20893 20959 20927
rect 20901 20887 20959 20893
rect 20990 20884 20996 20936
rect 21048 20884 21054 20936
rect 22278 20884 22284 20936
rect 22336 20924 22342 20936
rect 24302 20924 24308 20936
rect 22336 20896 24308 20924
rect 22336 20884 22342 20896
rect 24302 20884 24308 20896
rect 24360 20884 24366 20936
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 26050 20924 26056 20936
rect 24912 20896 26056 20924
rect 24912 20884 24918 20896
rect 26050 20884 26056 20896
rect 26108 20884 26114 20936
rect 24762 20856 24768 20868
rect 20640 20828 24768 20856
rect 24762 20816 24768 20828
rect 24820 20816 24826 20868
rect 31726 20856 31754 20964
rect 33520 20964 33824 20992
rect 31938 20884 31944 20936
rect 31996 20884 32002 20936
rect 32214 20933 32220 20936
rect 32208 20924 32220 20933
rect 32175 20896 32220 20924
rect 32208 20887 32220 20896
rect 32214 20884 32220 20887
rect 32272 20884 32278 20936
rect 33520 20856 33548 20964
rect 33597 20927 33655 20933
rect 33597 20893 33609 20927
rect 33643 20924 33655 20927
rect 33796 20924 33824 20964
rect 33962 20952 33968 21004
rect 34020 20992 34026 21004
rect 34149 20995 34207 21001
rect 34149 20992 34161 20995
rect 34020 20964 34161 20992
rect 34020 20952 34026 20964
rect 34149 20961 34161 20964
rect 34195 20961 34207 20995
rect 34149 20955 34207 20961
rect 34238 20952 34244 21004
rect 34296 20952 34302 21004
rect 34330 20952 34336 21004
rect 34388 20992 34394 21004
rect 36906 20992 36912 21004
rect 34388 20964 36912 20992
rect 34388 20952 34394 20964
rect 36906 20952 36912 20964
rect 36964 20952 36970 21004
rect 42518 20952 42524 21004
rect 42576 20992 42582 21004
rect 42886 20992 42892 21004
rect 42576 20964 42892 20992
rect 42576 20952 42582 20964
rect 42886 20952 42892 20964
rect 42944 20952 42950 21004
rect 37093 20927 37151 20933
rect 33643 20896 33732 20924
rect 33796 20896 34928 20924
rect 33643 20893 33655 20896
rect 33597 20887 33655 20893
rect 31726 20828 33548 20856
rect 20622 20788 20628 20800
rect 20548 20760 20628 20788
rect 20622 20748 20628 20760
rect 20680 20788 20686 20800
rect 23290 20788 23296 20800
rect 20680 20760 23296 20788
rect 20680 20748 20686 20760
rect 23290 20748 23296 20760
rect 23348 20748 23354 20800
rect 33410 20748 33416 20800
rect 33468 20748 33474 20800
rect 33704 20797 33732 20896
rect 34057 20859 34115 20865
rect 34057 20825 34069 20859
rect 34103 20856 34115 20859
rect 34422 20856 34428 20868
rect 34103 20828 34428 20856
rect 34103 20825 34115 20828
rect 34057 20819 34115 20825
rect 34422 20816 34428 20828
rect 34480 20816 34486 20868
rect 34793 20859 34851 20865
rect 34793 20825 34805 20859
rect 34839 20825 34851 20859
rect 34900 20856 34928 20896
rect 37093 20893 37105 20927
rect 37139 20924 37151 20927
rect 37274 20924 37280 20936
rect 37139 20896 37280 20924
rect 37139 20893 37151 20896
rect 37093 20887 37151 20893
rect 37274 20884 37280 20896
rect 37332 20884 37338 20936
rect 37369 20927 37427 20933
rect 37369 20893 37381 20927
rect 37415 20893 37427 20927
rect 37369 20887 37427 20893
rect 37384 20856 37412 20887
rect 38010 20884 38016 20936
rect 38068 20924 38074 20936
rect 38562 20924 38568 20936
rect 38068 20896 38568 20924
rect 38068 20884 38074 20896
rect 38562 20884 38568 20896
rect 38620 20924 38626 20936
rect 39853 20927 39911 20933
rect 39853 20924 39865 20927
rect 38620 20896 39865 20924
rect 38620 20884 38626 20896
rect 39853 20893 39865 20896
rect 39899 20893 39911 20927
rect 39853 20887 39911 20893
rect 40126 20884 40132 20936
rect 40184 20884 40190 20936
rect 43346 20884 43352 20936
rect 43404 20884 43410 20936
rect 43732 20933 43760 21032
rect 45925 21029 45937 21032
rect 45971 21029 45983 21063
rect 45925 21023 45983 21029
rect 44545 20995 44603 21001
rect 44545 20961 44557 20995
rect 44591 20992 44603 20995
rect 44634 20992 44640 21004
rect 44591 20964 44640 20992
rect 44591 20961 44603 20964
rect 44545 20955 44603 20961
rect 44634 20952 44640 20964
rect 44692 20952 44698 21004
rect 44821 20995 44879 21001
rect 44821 20961 44833 20995
rect 44867 20992 44879 20995
rect 45557 20995 45615 21001
rect 45557 20992 45569 20995
rect 44867 20964 45569 20992
rect 44867 20961 44879 20964
rect 44821 20955 44879 20961
rect 45557 20961 45569 20964
rect 45603 20961 45615 20995
rect 45557 20955 45615 20961
rect 45738 20952 45744 21004
rect 45796 20952 45802 21004
rect 43717 20927 43775 20933
rect 43717 20893 43729 20927
rect 43763 20893 43775 20927
rect 43717 20887 43775 20893
rect 44453 20927 44511 20933
rect 44453 20893 44465 20927
rect 44499 20893 44511 20927
rect 46198 20924 46204 20936
rect 44453 20887 44511 20893
rect 45572 20896 46204 20924
rect 34900 20828 37412 20856
rect 34793 20819 34851 20825
rect 33689 20791 33747 20797
rect 33689 20757 33701 20791
rect 33735 20757 33747 20791
rect 33689 20751 33747 20757
rect 34146 20748 34152 20800
rect 34204 20788 34210 20800
rect 34808 20788 34836 20819
rect 40678 20816 40684 20868
rect 40736 20856 40742 20868
rect 42886 20856 42892 20868
rect 40736 20828 42892 20856
rect 40736 20816 40742 20828
rect 42886 20816 42892 20828
rect 42944 20856 42950 20868
rect 43533 20859 43591 20865
rect 43533 20856 43545 20859
rect 42944 20828 43545 20856
rect 42944 20816 42950 20828
rect 43533 20825 43545 20828
rect 43579 20825 43591 20859
rect 43533 20819 43591 20825
rect 43622 20816 43628 20868
rect 43680 20816 43686 20868
rect 44468 20856 44496 20887
rect 45572 20868 45600 20896
rect 46198 20884 46204 20896
rect 46256 20924 46262 20936
rect 46293 20927 46351 20933
rect 46293 20924 46305 20927
rect 46256 20896 46305 20924
rect 46256 20884 46262 20896
rect 46293 20893 46305 20896
rect 46339 20893 46351 20927
rect 46293 20887 46351 20893
rect 44542 20856 44548 20868
rect 44468 20828 44548 20856
rect 44542 20816 44548 20828
rect 44600 20816 44606 20868
rect 45554 20816 45560 20868
rect 45612 20816 45618 20868
rect 36630 20788 36636 20800
rect 34204 20760 36636 20788
rect 34204 20748 34210 20760
rect 36630 20748 36636 20760
rect 36688 20748 36694 20800
rect 40865 20791 40923 20797
rect 40865 20757 40877 20791
rect 40911 20788 40923 20791
rect 41046 20788 41052 20800
rect 40911 20760 41052 20788
rect 40911 20757 40923 20760
rect 40865 20751 40923 20757
rect 41046 20748 41052 20760
rect 41104 20748 41110 20800
rect 42978 20748 42984 20800
rect 43036 20788 43042 20800
rect 43640 20788 43668 20816
rect 43036 20760 43668 20788
rect 43036 20748 43042 20760
rect 1104 20698 47104 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 47104 20698
rect 1104 20624 47104 20646
rect 2958 20544 2964 20596
rect 3016 20584 3022 20596
rect 3053 20587 3111 20593
rect 3053 20584 3065 20587
rect 3016 20556 3065 20584
rect 3016 20544 3022 20556
rect 3053 20553 3065 20556
rect 3099 20584 3111 20587
rect 3878 20584 3884 20596
rect 3099 20556 3884 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 3878 20544 3884 20556
rect 3936 20544 3942 20596
rect 6914 20584 6920 20596
rect 4448 20556 6920 20584
rect 1940 20519 1998 20525
rect 1940 20485 1952 20519
rect 1986 20516 1998 20519
rect 2130 20516 2136 20528
rect 1986 20488 2136 20516
rect 1986 20485 1998 20488
rect 1940 20479 1998 20485
rect 2130 20476 2136 20488
rect 2188 20476 2194 20528
rect 3970 20476 3976 20528
rect 4028 20516 4034 20528
rect 4448 20516 4476 20556
rect 6914 20544 6920 20556
rect 6972 20584 6978 20596
rect 6972 20556 11836 20584
rect 6972 20544 6978 20556
rect 8294 20525 8300 20528
rect 8288 20516 8300 20525
rect 4028 20488 4476 20516
rect 8255 20488 8300 20516
rect 4028 20476 4034 20488
rect 8288 20479 8300 20488
rect 8294 20476 8300 20479
rect 8352 20476 8358 20528
rect 1581 20451 1639 20457
rect 1581 20417 1593 20451
rect 1627 20448 1639 20451
rect 2498 20448 2504 20460
rect 1627 20420 2504 20448
rect 1627 20417 1639 20420
rect 1581 20411 1639 20417
rect 2498 20408 2504 20420
rect 2556 20408 2562 20460
rect 3881 20451 3939 20457
rect 3881 20417 3893 20451
rect 3927 20448 3939 20451
rect 3927 20420 4292 20448
rect 3927 20417 3939 20420
rect 3881 20411 3939 20417
rect 1670 20340 1676 20392
rect 1728 20340 1734 20392
rect 4062 20340 4068 20392
rect 4120 20340 4126 20392
rect 4264 20380 4292 20420
rect 5534 20408 5540 20460
rect 5592 20408 5598 20460
rect 7650 20408 7656 20460
rect 7708 20448 7714 20460
rect 8110 20448 8116 20460
rect 7708 20420 8116 20448
rect 7708 20408 7714 20420
rect 8110 20408 8116 20420
rect 8168 20408 8174 20460
rect 9769 20451 9827 20457
rect 9769 20417 9781 20451
rect 9815 20448 9827 20451
rect 9858 20448 9864 20460
rect 9815 20420 9864 20448
rect 9815 20417 9827 20420
rect 9769 20411 9827 20417
rect 9858 20408 9864 20420
rect 9916 20408 9922 20460
rect 10321 20451 10379 20457
rect 10321 20417 10333 20451
rect 10367 20417 10379 20451
rect 10321 20411 10379 20417
rect 4341 20383 4399 20389
rect 4341 20380 4353 20383
rect 4264 20352 4353 20380
rect 4341 20349 4353 20352
rect 4387 20380 4399 20383
rect 4430 20380 4436 20392
rect 4387 20352 4436 20380
rect 4387 20349 4399 20352
rect 4341 20343 4399 20349
rect 4430 20340 4436 20352
rect 4488 20340 4494 20392
rect 4525 20383 4583 20389
rect 4525 20349 4537 20383
rect 4571 20349 4583 20383
rect 4525 20343 4583 20349
rect 3326 20272 3332 20324
rect 3384 20312 3390 20324
rect 4154 20312 4160 20324
rect 3384 20284 4160 20312
rect 3384 20272 3390 20284
rect 4154 20272 4160 20284
rect 4212 20272 4218 20324
rect 1397 20247 1455 20253
rect 1397 20213 1409 20247
rect 1443 20244 1455 20247
rect 1946 20244 1952 20256
rect 1443 20216 1952 20244
rect 1443 20213 1455 20216
rect 1397 20207 1455 20213
rect 1946 20204 1952 20216
rect 2004 20204 2010 20256
rect 3510 20204 3516 20256
rect 3568 20204 3574 20256
rect 4540 20244 4568 20343
rect 4706 20340 4712 20392
rect 4764 20380 4770 20392
rect 4764 20352 5028 20380
rect 4764 20340 4770 20352
rect 5000 20321 5028 20352
rect 5258 20340 5264 20392
rect 5316 20340 5322 20392
rect 5442 20389 5448 20392
rect 5399 20383 5448 20389
rect 5399 20349 5411 20383
rect 5445 20349 5448 20383
rect 5399 20343 5448 20349
rect 5442 20340 5448 20343
rect 5500 20340 5506 20392
rect 5718 20340 5724 20392
rect 5776 20380 5782 20392
rect 6365 20383 6423 20389
rect 6365 20380 6377 20383
rect 5776 20352 6377 20380
rect 5776 20340 5782 20352
rect 6365 20349 6377 20352
rect 6411 20349 6423 20383
rect 6365 20343 6423 20349
rect 6641 20383 6699 20389
rect 6641 20349 6653 20383
rect 6687 20349 6699 20383
rect 6641 20343 6699 20349
rect 4985 20315 5043 20321
rect 4985 20281 4997 20315
rect 5031 20281 5043 20315
rect 6656 20312 6684 20343
rect 7190 20340 7196 20392
rect 7248 20380 7254 20392
rect 8021 20383 8079 20389
rect 8021 20380 8033 20383
rect 7248 20352 8033 20380
rect 7248 20340 7254 20352
rect 8021 20349 8033 20352
rect 8067 20349 8079 20383
rect 10336 20380 10364 20411
rect 11146 20408 11152 20460
rect 11204 20448 11210 20460
rect 11609 20451 11667 20457
rect 11609 20448 11621 20451
rect 11204 20420 11621 20448
rect 11204 20408 11210 20420
rect 11609 20417 11621 20420
rect 11655 20417 11667 20451
rect 11808 20448 11836 20556
rect 12066 20544 12072 20596
rect 12124 20584 12130 20596
rect 12161 20587 12219 20593
rect 12161 20584 12173 20587
rect 12124 20556 12173 20584
rect 12124 20544 12130 20556
rect 12161 20553 12173 20556
rect 12207 20553 12219 20587
rect 12161 20547 12219 20553
rect 12986 20544 12992 20596
rect 13044 20544 13050 20596
rect 13265 20587 13323 20593
rect 13265 20553 13277 20587
rect 13311 20553 13323 20587
rect 13265 20547 13323 20553
rect 13633 20587 13691 20593
rect 13633 20553 13645 20587
rect 13679 20584 13691 20587
rect 13906 20584 13912 20596
rect 13679 20556 13912 20584
rect 13679 20553 13691 20556
rect 13633 20547 13691 20553
rect 13173 20451 13231 20457
rect 11808 20420 13124 20448
rect 11609 20411 11667 20417
rect 11882 20380 11888 20392
rect 10336 20352 11888 20380
rect 8021 20343 8079 20349
rect 11882 20340 11888 20352
rect 11940 20340 11946 20392
rect 12526 20340 12532 20392
rect 12584 20340 12590 20392
rect 12618 20340 12624 20392
rect 12676 20340 12682 20392
rect 13096 20380 13124 20420
rect 13173 20417 13185 20451
rect 13219 20448 13231 20451
rect 13280 20448 13308 20547
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 14734 20544 14740 20596
rect 14792 20544 14798 20596
rect 15013 20587 15071 20593
rect 15013 20553 15025 20587
rect 15059 20553 15071 20587
rect 15013 20547 15071 20553
rect 15381 20587 15439 20593
rect 15381 20553 15393 20587
rect 15427 20584 15439 20587
rect 15838 20584 15844 20596
rect 15427 20556 15844 20584
rect 15427 20553 15439 20556
rect 15381 20547 15439 20553
rect 13219 20420 13308 20448
rect 13219 20417 13231 20420
rect 13173 20411 13231 20417
rect 13630 20408 13636 20460
rect 13688 20448 13694 20460
rect 14921 20451 14979 20457
rect 13688 20420 13860 20448
rect 13688 20408 13694 20420
rect 13832 20389 13860 20420
rect 14921 20417 14933 20451
rect 14967 20448 14979 20451
rect 15028 20448 15056 20547
rect 15838 20544 15844 20556
rect 15896 20544 15902 20596
rect 16853 20587 16911 20593
rect 16853 20553 16865 20587
rect 16899 20553 16911 20587
rect 16853 20547 16911 20553
rect 16868 20516 16896 20547
rect 18506 20544 18512 20596
rect 18564 20544 18570 20596
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 31662 20584 31668 20596
rect 19475 20556 30144 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 17374 20519 17432 20525
rect 17374 20516 17386 20519
rect 16868 20488 17386 20516
rect 17374 20485 17386 20488
rect 17420 20485 17432 20519
rect 20254 20516 20260 20528
rect 17374 20479 17432 20485
rect 20180 20488 20260 20516
rect 14967 20420 15056 20448
rect 14967 20417 14979 20420
rect 14921 20411 14979 20417
rect 15930 20408 15936 20460
rect 15988 20408 15994 20460
rect 17034 20408 17040 20460
rect 17092 20408 17098 20460
rect 17129 20451 17187 20457
rect 17129 20417 17141 20451
rect 17175 20448 17187 20451
rect 17678 20448 17684 20460
rect 17175 20420 17684 20448
rect 17175 20417 17187 20420
rect 17129 20411 17187 20417
rect 17678 20408 17684 20420
rect 17736 20408 17742 20460
rect 18969 20451 19027 20457
rect 18969 20417 18981 20451
rect 19015 20448 19027 20451
rect 19978 20448 19984 20460
rect 19015 20420 19984 20448
rect 19015 20417 19027 20420
rect 18969 20411 19027 20417
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 20180 20457 20208 20488
rect 20254 20476 20260 20488
rect 20312 20516 20318 20528
rect 20993 20519 21051 20525
rect 20993 20516 21005 20519
rect 20312 20488 21005 20516
rect 20312 20476 20318 20488
rect 20993 20485 21005 20488
rect 21039 20516 21051 20519
rect 21266 20516 21272 20528
rect 21039 20488 21272 20516
rect 21039 20485 21051 20488
rect 20993 20479 21051 20485
rect 21266 20476 21272 20488
rect 21324 20476 21330 20528
rect 29549 20519 29607 20525
rect 29549 20485 29561 20519
rect 29595 20516 29607 20519
rect 29595 20488 29960 20516
rect 29595 20485 29607 20488
rect 29549 20479 29607 20485
rect 20165 20451 20223 20457
rect 20165 20417 20177 20451
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 13725 20383 13783 20389
rect 13725 20380 13737 20383
rect 13096 20352 13737 20380
rect 13725 20349 13737 20352
rect 13771 20349 13783 20383
rect 13725 20343 13783 20349
rect 13817 20383 13875 20389
rect 13817 20349 13829 20383
rect 13863 20349 13875 20383
rect 13817 20343 13875 20349
rect 15473 20383 15531 20389
rect 15473 20349 15485 20383
rect 15519 20349 15531 20383
rect 15473 20343 15531 20349
rect 15657 20383 15715 20389
rect 15657 20349 15669 20383
rect 15703 20380 15715 20383
rect 16206 20380 16212 20392
rect 15703 20352 16212 20380
rect 15703 20349 15715 20352
rect 15657 20343 15715 20349
rect 4985 20275 5043 20281
rect 5920 20284 6684 20312
rect 4706 20244 4712 20256
rect 4540 20216 4712 20244
rect 4706 20204 4712 20216
rect 4764 20204 4770 20256
rect 4890 20204 4896 20256
rect 4948 20244 4954 20256
rect 5920 20244 5948 20284
rect 9214 20272 9220 20324
rect 9272 20312 9278 20324
rect 10597 20315 10655 20321
rect 10597 20312 10609 20315
rect 9272 20284 10609 20312
rect 9272 20272 9278 20284
rect 10597 20281 10609 20284
rect 10643 20281 10655 20315
rect 13740 20312 13768 20343
rect 15488 20312 15516 20343
rect 16206 20340 16212 20352
rect 16264 20340 16270 20392
rect 19058 20340 19064 20392
rect 19116 20380 19122 20392
rect 20364 20380 20392 20411
rect 20438 20408 20444 20460
rect 20496 20408 20502 20460
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20448 20867 20451
rect 21450 20448 21456 20460
rect 20855 20420 21456 20448
rect 20855 20417 20867 20420
rect 20809 20411 20867 20417
rect 21450 20408 21456 20420
rect 21508 20408 21514 20460
rect 23569 20451 23627 20457
rect 23569 20417 23581 20451
rect 23615 20448 23627 20451
rect 24394 20448 24400 20460
rect 23615 20420 24400 20448
rect 23615 20417 23627 20420
rect 23569 20411 23627 20417
rect 24394 20408 24400 20420
rect 24452 20408 24458 20460
rect 29730 20408 29736 20460
rect 29788 20408 29794 20460
rect 29825 20451 29883 20457
rect 29825 20417 29837 20451
rect 29871 20417 29883 20451
rect 29825 20411 29883 20417
rect 19116 20352 20392 20380
rect 19116 20340 19122 20352
rect 16117 20315 16175 20321
rect 16117 20312 16129 20315
rect 13740 20284 16129 20312
rect 10597 20275 10655 20281
rect 16117 20281 16129 20284
rect 16163 20281 16175 20315
rect 16117 20275 16175 20281
rect 19242 20272 19248 20324
rect 19300 20272 19306 20324
rect 19981 20315 20039 20321
rect 19981 20281 19993 20315
rect 20027 20312 20039 20315
rect 23290 20312 23296 20324
rect 20027 20284 23296 20312
rect 20027 20281 20039 20284
rect 19981 20275 20039 20281
rect 23290 20272 23296 20284
rect 23348 20272 23354 20324
rect 24302 20272 24308 20324
rect 24360 20312 24366 20324
rect 26234 20312 26240 20324
rect 24360 20284 26240 20312
rect 24360 20272 24366 20284
rect 26234 20272 26240 20284
rect 26292 20272 26298 20324
rect 4948 20216 5948 20244
rect 4948 20204 4954 20216
rect 6178 20204 6184 20256
rect 6236 20204 6242 20256
rect 7837 20247 7895 20253
rect 7837 20213 7849 20247
rect 7883 20244 7895 20247
rect 8294 20244 8300 20256
rect 7883 20216 8300 20244
rect 7883 20213 7895 20216
rect 7837 20207 7895 20213
rect 8294 20204 8300 20216
rect 8352 20244 8358 20256
rect 9306 20244 9312 20256
rect 8352 20216 9312 20244
rect 8352 20204 8358 20216
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 9398 20204 9404 20256
rect 9456 20204 9462 20256
rect 9950 20204 9956 20256
rect 10008 20204 10014 20256
rect 10502 20204 10508 20256
rect 10560 20244 10566 20256
rect 11701 20247 11759 20253
rect 11701 20244 11713 20247
rect 10560 20216 11713 20244
rect 10560 20204 10566 20216
rect 11701 20213 11713 20216
rect 11747 20213 11759 20247
rect 11701 20207 11759 20213
rect 12805 20247 12863 20253
rect 12805 20213 12817 20247
rect 12851 20244 12863 20247
rect 20714 20244 20720 20256
rect 12851 20216 20720 20244
rect 12851 20213 12863 20216
rect 12805 20207 12863 20213
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 23382 20204 23388 20256
rect 23440 20204 23446 20256
rect 24670 20204 24676 20256
rect 24728 20244 24734 20256
rect 27890 20244 27896 20256
rect 24728 20216 27896 20244
rect 24728 20204 24734 20216
rect 27890 20204 27896 20216
rect 27948 20204 27954 20256
rect 29840 20244 29868 20411
rect 29932 20312 29960 20488
rect 30116 20457 30144 20556
rect 30576 20556 31668 20584
rect 30576 20457 30604 20556
rect 31662 20544 31668 20556
rect 31720 20544 31726 20596
rect 32125 20587 32183 20593
rect 32125 20553 32137 20587
rect 32171 20553 32183 20587
rect 32125 20547 32183 20553
rect 30828 20519 30886 20525
rect 30828 20485 30840 20519
rect 30874 20516 30886 20519
rect 32140 20516 32168 20547
rect 33686 20544 33692 20596
rect 33744 20584 33750 20596
rect 34330 20584 34336 20596
rect 33744 20556 34336 20584
rect 33744 20544 33750 20556
rect 34330 20544 34336 20556
rect 34388 20544 34394 20596
rect 34698 20544 34704 20596
rect 34756 20584 34762 20596
rect 35345 20587 35403 20593
rect 35345 20584 35357 20587
rect 34756 20556 35357 20584
rect 34756 20544 34762 20556
rect 35345 20553 35357 20556
rect 35391 20553 35403 20587
rect 35345 20547 35403 20553
rect 37458 20544 37464 20596
rect 37516 20584 37522 20596
rect 38378 20584 38384 20596
rect 37516 20556 38384 20584
rect 37516 20544 37522 20556
rect 38378 20544 38384 20556
rect 38436 20544 38442 20596
rect 43438 20584 43444 20596
rect 38672 20556 43444 20584
rect 30874 20488 32168 20516
rect 30874 20485 30886 20488
rect 30828 20479 30886 20485
rect 30101 20451 30159 20457
rect 30101 20417 30113 20451
rect 30147 20417 30159 20451
rect 30101 20411 30159 20417
rect 30561 20451 30619 20457
rect 30561 20417 30573 20451
rect 30607 20417 30619 20451
rect 30561 20411 30619 20417
rect 31386 20408 31392 20460
rect 31444 20448 31450 20460
rect 32309 20451 32367 20457
rect 32309 20448 32321 20451
rect 31444 20420 32321 20448
rect 31444 20408 31450 20420
rect 32309 20417 32321 20420
rect 32355 20417 32367 20451
rect 32309 20411 32367 20417
rect 33505 20451 33563 20457
rect 33505 20417 33517 20451
rect 33551 20448 33563 20451
rect 33594 20448 33600 20460
rect 33551 20420 33600 20448
rect 33551 20417 33563 20420
rect 33505 20411 33563 20417
rect 33594 20408 33600 20420
rect 33652 20408 33658 20460
rect 33704 20457 33732 20544
rect 38672 20525 38700 20556
rect 43438 20544 43444 20556
rect 43496 20544 43502 20596
rect 43533 20587 43591 20593
rect 43533 20553 43545 20587
rect 43579 20584 43591 20587
rect 44542 20584 44548 20596
rect 43579 20556 44548 20584
rect 43579 20553 43591 20556
rect 43533 20547 43591 20553
rect 44542 20544 44548 20556
rect 44600 20544 44606 20596
rect 46658 20544 46664 20596
rect 46716 20544 46722 20596
rect 38657 20519 38715 20525
rect 38657 20485 38669 20519
rect 38703 20485 38715 20519
rect 45925 20519 45983 20525
rect 45925 20516 45937 20519
rect 38657 20479 38715 20485
rect 41156 20488 45937 20516
rect 33689 20451 33747 20457
rect 33689 20417 33701 20451
rect 33735 20417 33747 20451
rect 33689 20411 33747 20417
rect 34514 20408 34520 20460
rect 34572 20457 34578 20460
rect 34572 20451 34600 20457
rect 34588 20417 34600 20451
rect 34572 20411 34600 20417
rect 34572 20408 34578 20411
rect 34698 20408 34704 20460
rect 34756 20408 34762 20460
rect 37458 20408 37464 20460
rect 37516 20448 37522 20460
rect 37918 20448 37924 20460
rect 37516 20420 37924 20448
rect 37516 20408 37522 20420
rect 37918 20408 37924 20420
rect 37976 20448 37982 20460
rect 38381 20451 38439 20457
rect 38381 20448 38393 20451
rect 37976 20420 38393 20448
rect 37976 20408 37982 20420
rect 38381 20417 38393 20420
rect 38427 20417 38439 20451
rect 38381 20411 38439 20417
rect 38565 20451 38623 20457
rect 38565 20417 38577 20451
rect 38611 20417 38623 20451
rect 38565 20411 38623 20417
rect 38754 20451 38812 20457
rect 38754 20417 38766 20451
rect 38800 20417 38812 20451
rect 38754 20411 38812 20417
rect 30006 20340 30012 20392
rect 30064 20340 30070 20392
rect 33134 20340 33140 20392
rect 33192 20380 33198 20392
rect 34149 20383 34207 20389
rect 34149 20380 34161 20383
rect 33192 20352 34161 20380
rect 33192 20340 33198 20352
rect 33980 20324 34008 20352
rect 34149 20349 34161 20352
rect 34195 20349 34207 20383
rect 34149 20343 34207 20349
rect 34422 20340 34428 20392
rect 34480 20340 34486 20392
rect 38580 20380 38608 20411
rect 38654 20380 38660 20392
rect 38580 20352 38660 20380
rect 38654 20340 38660 20352
rect 38712 20340 38718 20392
rect 29932 20284 30604 20312
rect 30466 20244 30472 20256
rect 29840 20216 30472 20244
rect 30466 20204 30472 20216
rect 30524 20204 30530 20256
rect 30576 20244 30604 20284
rect 31726 20284 32076 20312
rect 31726 20244 31754 20284
rect 30576 20216 31754 20244
rect 31846 20204 31852 20256
rect 31904 20244 31910 20256
rect 31941 20247 31999 20253
rect 31941 20244 31953 20247
rect 31904 20216 31953 20244
rect 31904 20204 31910 20216
rect 31941 20213 31953 20216
rect 31987 20213 31999 20247
rect 32048 20244 32076 20284
rect 33962 20272 33968 20324
rect 34020 20272 34026 20324
rect 37918 20272 37924 20324
rect 37976 20312 37982 20324
rect 38764 20312 38792 20411
rect 40678 20408 40684 20460
rect 40736 20448 40742 20460
rect 40954 20448 40960 20460
rect 40736 20420 40960 20448
rect 40736 20408 40742 20420
rect 40954 20408 40960 20420
rect 41012 20448 41018 20460
rect 41156 20457 41184 20488
rect 45925 20485 45937 20488
rect 45971 20485 45983 20519
rect 45925 20479 45983 20485
rect 41049 20451 41107 20457
rect 41049 20448 41061 20451
rect 41012 20420 41061 20448
rect 41012 20408 41018 20420
rect 41049 20417 41061 20420
rect 41095 20417 41107 20451
rect 41049 20411 41107 20417
rect 41141 20451 41199 20457
rect 41141 20417 41153 20451
rect 41187 20417 41199 20451
rect 41141 20411 41199 20417
rect 41322 20408 41328 20460
rect 41380 20408 41386 20460
rect 41414 20408 41420 20460
rect 41472 20408 41478 20460
rect 41598 20408 41604 20460
rect 41656 20448 41662 20460
rect 42153 20451 42211 20457
rect 42153 20448 42165 20451
rect 41656 20420 42165 20448
rect 41656 20408 41662 20420
rect 42153 20417 42165 20420
rect 42199 20417 42211 20451
rect 42153 20411 42211 20417
rect 42334 20408 42340 20460
rect 42392 20448 42398 20460
rect 42429 20451 42487 20457
rect 42429 20448 42441 20451
rect 42392 20420 42441 20448
rect 42392 20408 42398 20420
rect 42429 20417 42441 20420
rect 42475 20417 42487 20451
rect 42429 20411 42487 20417
rect 42613 20451 42671 20457
rect 42613 20417 42625 20451
rect 42659 20417 42671 20451
rect 42613 20411 42671 20417
rect 40218 20340 40224 20392
rect 40276 20380 40282 20392
rect 41340 20380 41368 20408
rect 41877 20383 41935 20389
rect 41877 20380 41889 20383
rect 40276 20352 41368 20380
rect 41616 20352 41889 20380
rect 40276 20340 40282 20352
rect 41616 20324 41644 20352
rect 41877 20349 41889 20352
rect 41923 20349 41935 20383
rect 41877 20343 41935 20349
rect 41969 20383 42027 20389
rect 41969 20349 41981 20383
rect 42015 20349 42027 20383
rect 41969 20343 42027 20349
rect 42061 20383 42119 20389
rect 42061 20349 42073 20383
rect 42107 20380 42119 20383
rect 42628 20380 42656 20411
rect 42702 20408 42708 20460
rect 42760 20408 42766 20460
rect 42978 20408 42984 20460
rect 43036 20448 43042 20460
rect 43349 20451 43407 20457
rect 43349 20448 43361 20451
rect 43036 20420 43361 20448
rect 43036 20408 43042 20420
rect 43349 20417 43361 20420
rect 43395 20417 43407 20451
rect 43349 20411 43407 20417
rect 43530 20408 43536 20460
rect 43588 20408 43594 20460
rect 46198 20408 46204 20460
rect 46256 20408 46262 20460
rect 46474 20408 46480 20460
rect 46532 20408 46538 20460
rect 42107 20352 42656 20380
rect 42107 20349 42119 20352
rect 42061 20343 42119 20349
rect 37976 20284 38792 20312
rect 37976 20272 37982 20284
rect 38838 20272 38844 20324
rect 38896 20312 38902 20324
rect 38933 20315 38991 20321
rect 38933 20312 38945 20315
rect 38896 20284 38945 20312
rect 38896 20272 38902 20284
rect 38933 20281 38945 20284
rect 38979 20281 38991 20315
rect 38933 20275 38991 20281
rect 41598 20272 41604 20324
rect 41656 20272 41662 20324
rect 41984 20312 42012 20343
rect 42334 20312 42340 20324
rect 41984 20284 42340 20312
rect 42334 20272 42340 20284
rect 42392 20272 42398 20324
rect 42628 20312 42656 20352
rect 42797 20383 42855 20389
rect 42797 20349 42809 20383
rect 42843 20380 42855 20383
rect 43548 20380 43576 20408
rect 42843 20352 43576 20380
rect 42843 20349 42855 20352
rect 42797 20343 42855 20349
rect 42812 20312 42840 20343
rect 45278 20340 45284 20392
rect 45336 20340 45342 20392
rect 45465 20383 45523 20389
rect 45465 20349 45477 20383
rect 45511 20349 45523 20383
rect 45465 20343 45523 20349
rect 42628 20284 42840 20312
rect 45480 20312 45508 20343
rect 46017 20315 46075 20321
rect 46017 20312 46029 20315
rect 45480 20284 46029 20312
rect 46017 20281 46029 20284
rect 46063 20281 46075 20315
rect 46017 20275 46075 20281
rect 40034 20244 40040 20256
rect 32048 20216 40040 20244
rect 31941 20207 31999 20213
rect 40034 20204 40040 20216
rect 40092 20204 40098 20256
rect 40862 20204 40868 20256
rect 40920 20204 40926 20256
rect 41506 20204 41512 20256
rect 41564 20244 41570 20256
rect 41693 20247 41751 20253
rect 41693 20244 41705 20247
rect 41564 20216 41705 20244
rect 41564 20204 41570 20216
rect 41693 20213 41705 20216
rect 41739 20213 41751 20247
rect 41693 20207 41751 20213
rect 42426 20204 42432 20256
rect 42484 20204 42490 20256
rect 43162 20204 43168 20256
rect 43220 20204 43226 20256
rect 1104 20154 47104 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 47104 20154
rect 1104 20080 47104 20102
rect 2958 20000 2964 20052
rect 3016 20040 3022 20052
rect 3053 20043 3111 20049
rect 3053 20040 3065 20043
rect 3016 20012 3065 20040
rect 3016 20000 3022 20012
rect 3053 20009 3065 20012
rect 3099 20040 3111 20043
rect 5442 20040 5448 20052
rect 3099 20012 5448 20040
rect 3099 20009 3111 20012
rect 3053 20003 3111 20009
rect 5442 20000 5448 20012
rect 5500 20000 5506 20052
rect 6178 20000 6184 20052
rect 6236 20040 6242 20052
rect 12526 20040 12532 20052
rect 6236 20012 12532 20040
rect 6236 20000 6242 20012
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 17034 20000 17040 20052
rect 17092 20040 17098 20052
rect 17589 20043 17647 20049
rect 17589 20040 17601 20043
rect 17092 20012 17601 20040
rect 17092 20000 17098 20012
rect 17589 20009 17601 20012
rect 17635 20009 17647 20043
rect 17589 20003 17647 20009
rect 18064 20012 24348 20040
rect 4154 19932 4160 19984
rect 4212 19972 4218 19984
rect 4890 19972 4896 19984
rect 4212 19944 4896 19972
rect 4212 19932 4218 19944
rect 4890 19932 4896 19944
rect 4948 19932 4954 19984
rect 5166 19932 5172 19984
rect 5224 19932 5230 19984
rect 6270 19932 6276 19984
rect 6328 19972 6334 19984
rect 8665 19975 8723 19981
rect 8665 19972 8677 19975
rect 6328 19944 8677 19972
rect 6328 19932 6334 19944
rect 3878 19864 3884 19916
rect 3936 19904 3942 19916
rect 5258 19904 5264 19916
rect 3936 19876 5264 19904
rect 3936 19864 3942 19876
rect 5258 19864 5264 19876
rect 5316 19904 5322 19916
rect 5445 19907 5503 19913
rect 5445 19904 5457 19907
rect 5316 19876 5457 19904
rect 5316 19864 5322 19876
rect 5445 19873 5457 19876
rect 5491 19873 5503 19907
rect 5445 19867 5503 19873
rect 5534 19864 5540 19916
rect 5592 19913 5598 19916
rect 5592 19907 5620 19913
rect 5608 19873 5620 19907
rect 5592 19867 5620 19873
rect 5721 19907 5779 19913
rect 5721 19873 5733 19907
rect 5767 19904 5779 19907
rect 6086 19904 6092 19916
rect 5767 19876 6092 19904
rect 5767 19873 5779 19876
rect 5721 19867 5779 19873
rect 5592 19864 5598 19867
rect 6086 19864 6092 19876
rect 6144 19904 6150 19916
rect 6638 19904 6644 19916
rect 6144 19876 6644 19904
rect 6144 19864 6150 19876
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 6914 19864 6920 19916
rect 6972 19864 6978 19916
rect 7116 19913 7144 19944
rect 8665 19941 8677 19944
rect 8711 19972 8723 19975
rect 10410 19972 10416 19984
rect 8711 19944 10416 19972
rect 8711 19941 8723 19944
rect 8665 19935 8723 19941
rect 10410 19932 10416 19944
rect 10468 19932 10474 19984
rect 15930 19932 15936 19984
rect 15988 19972 15994 19984
rect 18064 19972 18092 20012
rect 15988 19944 18092 19972
rect 24320 19972 24348 20012
rect 24394 20000 24400 20052
rect 24452 20000 24458 20052
rect 24762 20000 24768 20052
rect 24820 20040 24826 20052
rect 24820 20012 29684 20040
rect 24820 20000 24826 20012
rect 26142 19972 26148 19984
rect 24320 19944 26148 19972
rect 15988 19932 15994 19944
rect 7101 19907 7159 19913
rect 7101 19873 7113 19907
rect 7147 19904 7159 19907
rect 13814 19904 13820 19916
rect 7147 19876 7181 19904
rect 8496 19876 13820 19904
rect 7147 19873 7159 19876
rect 7101 19867 7159 19873
rect 8496 19848 8524 19876
rect 13814 19864 13820 19876
rect 13872 19904 13878 19916
rect 13998 19904 14004 19916
rect 13872 19876 14004 19904
rect 13872 19864 13878 19876
rect 13998 19864 14004 19876
rect 14056 19864 14062 19916
rect 18064 19913 18092 19944
rect 26142 19932 26148 19944
rect 26200 19932 26206 19984
rect 26234 19932 26240 19984
rect 26292 19932 26298 19984
rect 27525 19975 27583 19981
rect 27525 19941 27537 19975
rect 27571 19972 27583 19975
rect 28902 19972 28908 19984
rect 27571 19944 28908 19972
rect 27571 19941 27583 19944
rect 27525 19935 27583 19941
rect 28902 19932 28908 19944
rect 28960 19932 28966 19984
rect 29362 19972 29368 19984
rect 29012 19944 29368 19972
rect 29012 19916 29040 19944
rect 29362 19932 29368 19944
rect 29420 19932 29426 19984
rect 29656 19972 29684 20012
rect 29730 20000 29736 20052
rect 29788 20040 29794 20052
rect 30929 20043 30987 20049
rect 30929 20040 30941 20043
rect 29788 20012 30941 20040
rect 29788 20000 29794 20012
rect 30929 20009 30941 20012
rect 30975 20009 30987 20043
rect 30929 20003 30987 20009
rect 31386 20000 31392 20052
rect 31444 20000 31450 20052
rect 34422 20000 34428 20052
rect 34480 20040 34486 20052
rect 34517 20043 34575 20049
rect 34517 20040 34529 20043
rect 34480 20012 34529 20040
rect 34480 20000 34486 20012
rect 34517 20009 34529 20012
rect 34563 20009 34575 20043
rect 34517 20003 34575 20009
rect 36906 20000 36912 20052
rect 36964 20040 36970 20052
rect 38562 20040 38568 20052
rect 36964 20012 38568 20040
rect 36964 20000 36970 20012
rect 38562 20000 38568 20012
rect 38620 20040 38626 20052
rect 38749 20043 38807 20049
rect 38749 20040 38761 20043
rect 38620 20012 38761 20040
rect 38620 20000 38626 20012
rect 38749 20009 38761 20012
rect 38795 20009 38807 20043
rect 38749 20003 38807 20009
rect 41414 20000 41420 20052
rect 41472 20040 41478 20052
rect 41509 20043 41567 20049
rect 41509 20040 41521 20043
rect 41472 20012 41521 20040
rect 41472 20000 41478 20012
rect 41509 20009 41521 20012
rect 41555 20009 41567 20043
rect 41509 20003 41567 20009
rect 41598 20000 41604 20052
rect 41656 20040 41662 20052
rect 42610 20040 42616 20052
rect 41656 20012 42616 20040
rect 41656 20000 41662 20012
rect 42610 20000 42616 20012
rect 42668 20000 42674 20052
rect 42978 20000 42984 20052
rect 43036 20040 43042 20052
rect 43165 20043 43223 20049
rect 43165 20040 43177 20043
rect 43036 20012 43177 20040
rect 43036 20000 43042 20012
rect 43165 20009 43177 20012
rect 43211 20009 43223 20043
rect 43165 20003 43223 20009
rect 43349 20043 43407 20049
rect 43349 20009 43361 20043
rect 43395 20040 43407 20043
rect 43530 20040 43536 20052
rect 43395 20012 43536 20040
rect 43395 20009 43407 20012
rect 43349 20003 43407 20009
rect 43530 20000 43536 20012
rect 43588 20000 43594 20052
rect 45922 20000 45928 20052
rect 45980 20000 45986 20052
rect 46198 20000 46204 20052
rect 46256 20000 46262 20052
rect 30837 19975 30895 19981
rect 29656 19944 30788 19972
rect 18049 19907 18107 19913
rect 18049 19873 18061 19907
rect 18095 19873 18107 19907
rect 18049 19867 18107 19873
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19904 18291 19907
rect 18322 19904 18328 19916
rect 18279 19876 18328 19904
rect 18279 19873 18291 19876
rect 18233 19867 18291 19873
rect 18322 19864 18328 19876
rect 18380 19904 18386 19916
rect 18782 19904 18788 19916
rect 18380 19876 18788 19904
rect 18380 19864 18386 19876
rect 18782 19864 18788 19876
rect 18840 19864 18846 19916
rect 19886 19864 19892 19916
rect 19944 19904 19950 19916
rect 20165 19907 20223 19913
rect 20165 19904 20177 19907
rect 19944 19876 20177 19904
rect 19944 19864 19950 19876
rect 20165 19873 20177 19876
rect 20211 19873 20223 19907
rect 20165 19867 20223 19873
rect 21174 19864 21180 19916
rect 21232 19864 21238 19916
rect 22830 19864 22836 19916
rect 22888 19864 22894 19916
rect 24670 19864 24676 19916
rect 24728 19904 24734 19916
rect 24857 19907 24915 19913
rect 24857 19904 24869 19907
rect 24728 19876 24869 19904
rect 24728 19864 24734 19876
rect 24857 19873 24869 19876
rect 24903 19873 24915 19907
rect 24857 19867 24915 19873
rect 24949 19907 25007 19913
rect 24949 19873 24961 19907
rect 24995 19873 25007 19907
rect 24949 19867 25007 19873
rect 1670 19796 1676 19848
rect 1728 19796 1734 19848
rect 1946 19845 1952 19848
rect 1940 19836 1952 19845
rect 1907 19808 1952 19836
rect 1940 19799 1952 19808
rect 1946 19796 1952 19799
rect 2004 19796 2010 19848
rect 3510 19796 3516 19848
rect 3568 19836 3574 19848
rect 4157 19839 4215 19845
rect 4157 19836 4169 19839
rect 3568 19808 4169 19836
rect 3568 19796 3574 19808
rect 4157 19805 4169 19808
rect 4203 19805 4215 19839
rect 4157 19799 4215 19805
rect 4522 19796 4528 19848
rect 4580 19796 4586 19848
rect 4706 19796 4712 19848
rect 4764 19796 4770 19848
rect 6362 19796 6368 19848
rect 6420 19836 6426 19848
rect 6825 19839 6883 19845
rect 6825 19836 6837 19839
rect 6420 19808 6837 19836
rect 6420 19796 6426 19808
rect 6825 19805 6837 19808
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 8478 19796 8484 19848
rect 8536 19796 8542 19848
rect 11606 19796 11612 19848
rect 11664 19836 11670 19848
rect 15289 19839 15347 19845
rect 15289 19836 15301 19839
rect 11664 19808 15301 19836
rect 11664 19796 11670 19808
rect 15289 19805 15301 19808
rect 15335 19836 15347 19839
rect 15654 19836 15660 19848
rect 15335 19808 15660 19836
rect 15335 19805 15347 19808
rect 15289 19799 15347 19805
rect 15654 19796 15660 19808
rect 15712 19796 15718 19848
rect 17221 19839 17279 19845
rect 17221 19805 17233 19839
rect 17267 19836 17279 19839
rect 17310 19836 17316 19848
rect 17267 19808 17316 19836
rect 17267 19805 17279 19808
rect 17221 19799 17279 19805
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 17957 19839 18015 19845
rect 17957 19805 17969 19839
rect 18003 19836 18015 19839
rect 18506 19836 18512 19848
rect 18003 19808 18512 19836
rect 18003 19805 18015 19808
rect 17957 19799 18015 19805
rect 18506 19796 18512 19808
rect 18564 19796 18570 19848
rect 20070 19796 20076 19848
rect 20128 19796 20134 19848
rect 20441 19839 20499 19845
rect 20441 19805 20453 19839
rect 20487 19805 20499 19839
rect 20441 19799 20499 19805
rect 3970 19660 3976 19712
rect 4028 19660 4034 19712
rect 4724 19700 4752 19796
rect 6380 19768 6408 19796
rect 6196 19740 6408 19768
rect 6196 19700 6224 19740
rect 6638 19728 6644 19780
rect 6696 19768 6702 19780
rect 11698 19768 11704 19780
rect 6696 19740 11704 19768
rect 6696 19728 6702 19740
rect 11698 19728 11704 19740
rect 11756 19728 11762 19780
rect 11974 19728 11980 19780
rect 12032 19768 12038 19780
rect 12529 19771 12587 19777
rect 12529 19768 12541 19771
rect 12032 19740 12541 19768
rect 12032 19728 12038 19740
rect 12529 19737 12541 19740
rect 12575 19737 12587 19771
rect 12529 19731 12587 19737
rect 12894 19728 12900 19780
rect 12952 19728 12958 19780
rect 15194 19728 15200 19780
rect 15252 19768 15258 19780
rect 19058 19768 19064 19780
rect 15252 19740 19064 19768
rect 15252 19728 15258 19740
rect 19058 19728 19064 19740
rect 19116 19728 19122 19780
rect 20456 19768 20484 19799
rect 20714 19796 20720 19848
rect 20772 19836 20778 19848
rect 21192 19836 21220 19864
rect 20772 19808 21220 19836
rect 23100 19839 23158 19845
rect 20772 19796 20778 19808
rect 23100 19805 23112 19839
rect 23146 19836 23158 19839
rect 23382 19836 23388 19848
rect 23146 19808 23388 19836
rect 23146 19805 23158 19808
rect 23100 19799 23158 19805
rect 23382 19796 23388 19808
rect 23440 19796 23446 19848
rect 23474 19796 23480 19848
rect 23532 19836 23538 19848
rect 24688 19836 24716 19864
rect 23532 19808 24716 19836
rect 23532 19796 23538 19808
rect 24762 19796 24768 19848
rect 24820 19836 24826 19848
rect 24964 19836 24992 19867
rect 26326 19864 26332 19916
rect 26384 19904 26390 19916
rect 26630 19907 26688 19913
rect 26630 19904 26642 19907
rect 26384 19876 26642 19904
rect 26384 19864 26390 19876
rect 26630 19873 26642 19876
rect 26676 19873 26688 19907
rect 26630 19867 26688 19873
rect 28169 19907 28227 19913
rect 28169 19873 28181 19907
rect 28215 19904 28227 19907
rect 28994 19904 29000 19916
rect 28215 19876 29000 19904
rect 28215 19873 28227 19876
rect 28169 19867 28227 19873
rect 28994 19864 29000 19876
rect 29052 19864 29058 19916
rect 29086 19864 29092 19916
rect 29144 19904 29150 19916
rect 29549 19907 29607 19913
rect 29549 19904 29561 19907
rect 29144 19876 29561 19904
rect 29144 19864 29150 19876
rect 29549 19873 29561 19876
rect 29595 19873 29607 19907
rect 29549 19867 29607 19873
rect 30469 19907 30527 19913
rect 30469 19873 30481 19907
rect 30515 19904 30527 19907
rect 30558 19904 30564 19916
rect 30515 19876 30564 19904
rect 30515 19873 30527 19876
rect 30469 19867 30527 19873
rect 30558 19864 30564 19876
rect 30616 19864 30622 19916
rect 30760 19904 30788 19944
rect 30837 19941 30849 19975
rect 30883 19972 30895 19975
rect 31110 19972 31116 19984
rect 30883 19944 31116 19972
rect 30883 19941 30895 19944
rect 30837 19935 30895 19941
rect 31110 19932 31116 19944
rect 31168 19932 31174 19984
rect 37734 19932 37740 19984
rect 37792 19972 37798 19984
rect 38105 19975 38163 19981
rect 38105 19972 38117 19975
rect 37792 19944 38117 19972
rect 37792 19932 37798 19944
rect 38105 19941 38117 19944
rect 38151 19941 38163 19975
rect 38105 19935 38163 19941
rect 31018 19904 31024 19916
rect 30760 19876 31024 19904
rect 31018 19864 31024 19876
rect 31076 19864 31082 19916
rect 32030 19864 32036 19916
rect 32088 19864 32094 19916
rect 40862 19904 40868 19916
rect 37752 19876 40868 19904
rect 24820 19808 24992 19836
rect 24820 19796 24826 19808
rect 25590 19796 25596 19848
rect 25648 19796 25654 19848
rect 25682 19796 25688 19848
rect 25740 19836 25746 19848
rect 25777 19839 25835 19845
rect 25777 19836 25789 19839
rect 25740 19808 25789 19836
rect 25740 19796 25746 19808
rect 25777 19805 25789 19808
rect 25823 19805 25835 19839
rect 25777 19799 25835 19805
rect 19904 19740 20484 19768
rect 4724 19672 6224 19700
rect 6362 19660 6368 19712
rect 6420 19660 6426 19712
rect 6454 19660 6460 19712
rect 6512 19660 6518 19712
rect 9858 19660 9864 19712
rect 9916 19700 9922 19712
rect 10502 19700 10508 19712
rect 9916 19672 10508 19700
rect 9916 19660 9922 19672
rect 10502 19660 10508 19672
rect 10560 19700 10566 19712
rect 11992 19700 12020 19728
rect 10560 19672 12020 19700
rect 10560 19660 10566 19672
rect 15378 19660 15384 19712
rect 15436 19700 15442 19712
rect 15473 19703 15531 19709
rect 15473 19700 15485 19703
rect 15436 19672 15485 19700
rect 15436 19660 15442 19672
rect 15473 19669 15485 19672
rect 15519 19669 15531 19703
rect 15473 19663 15531 19669
rect 17405 19703 17463 19709
rect 17405 19669 17417 19703
rect 17451 19700 17463 19703
rect 17954 19700 17960 19712
rect 17451 19672 17960 19700
rect 17451 19669 17463 19672
rect 17405 19663 17463 19669
rect 17954 19660 17960 19672
rect 18012 19660 18018 19712
rect 19904 19709 19932 19740
rect 20990 19728 20996 19780
rect 21048 19768 21054 19780
rect 24670 19768 24676 19780
rect 21048 19740 24676 19768
rect 21048 19728 21054 19740
rect 24670 19728 24676 19740
rect 24728 19728 24734 19780
rect 19889 19703 19947 19709
rect 19889 19669 19901 19703
rect 19935 19669 19947 19703
rect 19889 19663 19947 19669
rect 19978 19660 19984 19712
rect 20036 19700 20042 19712
rect 20714 19700 20720 19712
rect 20036 19672 20720 19700
rect 20036 19660 20042 19672
rect 20714 19660 20720 19672
rect 20772 19660 20778 19712
rect 21174 19660 21180 19712
rect 21232 19660 21238 19712
rect 23014 19660 23020 19712
rect 23072 19700 23078 19712
rect 24213 19703 24271 19709
rect 24213 19700 24225 19703
rect 23072 19672 24225 19700
rect 23072 19660 23078 19672
rect 24213 19669 24225 19672
rect 24259 19700 24271 19703
rect 24765 19703 24823 19709
rect 24765 19700 24777 19703
rect 24259 19672 24777 19700
rect 24259 19669 24271 19672
rect 24213 19663 24271 19669
rect 24765 19669 24777 19672
rect 24811 19669 24823 19703
rect 25792 19700 25820 19799
rect 26510 19796 26516 19848
rect 26568 19796 26574 19848
rect 26786 19796 26792 19848
rect 26844 19796 26850 19848
rect 28534 19796 28540 19848
rect 28592 19836 28598 19848
rect 29181 19839 29239 19845
rect 29181 19836 29193 19839
rect 28592 19808 29193 19836
rect 28592 19796 28598 19808
rect 29181 19805 29193 19808
rect 29227 19836 29239 19839
rect 29825 19839 29883 19845
rect 29825 19836 29837 19839
rect 29227 19808 29837 19836
rect 29227 19805 29239 19808
rect 29181 19799 29239 19805
rect 29825 19805 29837 19808
rect 29871 19805 29883 19839
rect 29825 19799 29883 19805
rect 31757 19839 31815 19845
rect 31757 19805 31769 19839
rect 31803 19836 31815 19839
rect 31846 19836 31852 19848
rect 31803 19808 31852 19836
rect 31803 19805 31815 19808
rect 31757 19799 31815 19805
rect 31846 19796 31852 19808
rect 31904 19796 31910 19848
rect 31938 19796 31944 19848
rect 31996 19836 32002 19848
rect 33410 19845 33416 19848
rect 33137 19839 33195 19845
rect 33137 19836 33149 19839
rect 31996 19808 33149 19836
rect 31996 19796 32002 19808
rect 33137 19805 33149 19808
rect 33183 19805 33195 19839
rect 33404 19836 33416 19845
rect 33371 19808 33416 19836
rect 33137 19799 33195 19805
rect 33404 19799 33416 19808
rect 33410 19796 33416 19799
rect 33468 19796 33474 19848
rect 37550 19796 37556 19848
rect 37608 19796 37614 19848
rect 37752 19845 37780 19876
rect 40862 19864 40868 19876
rect 40920 19864 40926 19916
rect 37737 19839 37795 19845
rect 37737 19805 37749 19839
rect 37783 19805 37795 19839
rect 37737 19799 37795 19805
rect 37826 19796 37832 19848
rect 37884 19796 37890 19848
rect 37918 19796 37924 19848
rect 37976 19845 37982 19848
rect 37976 19836 37984 19845
rect 38657 19839 38715 19845
rect 37976 19808 38021 19836
rect 37976 19799 37984 19808
rect 38657 19805 38669 19839
rect 38703 19836 38715 19839
rect 38746 19836 38752 19848
rect 38703 19808 38752 19836
rect 38703 19805 38715 19808
rect 38657 19799 38715 19805
rect 37976 19796 37982 19799
rect 38746 19796 38752 19808
rect 38804 19796 38810 19848
rect 41506 19796 41512 19848
rect 41564 19796 41570 19848
rect 41693 19839 41751 19845
rect 41693 19805 41705 19839
rect 41739 19836 41751 19839
rect 42426 19836 42432 19848
rect 41739 19808 42432 19836
rect 41739 19805 41751 19808
rect 41693 19799 41751 19805
rect 42426 19796 42432 19808
rect 42484 19796 42490 19848
rect 43257 19839 43315 19845
rect 43257 19836 43269 19839
rect 42812 19808 43269 19836
rect 42812 19780 42840 19808
rect 43257 19805 43269 19808
rect 43303 19805 43315 19839
rect 43257 19799 43315 19805
rect 43346 19796 43352 19848
rect 43404 19836 43410 19848
rect 43441 19839 43499 19845
rect 43441 19836 43453 19839
rect 43404 19808 43453 19836
rect 43404 19796 43410 19808
rect 43441 19805 43453 19808
rect 43487 19805 43499 19839
rect 43441 19799 43499 19805
rect 44542 19796 44548 19848
rect 44600 19796 44606 19848
rect 44634 19796 44640 19848
rect 44692 19796 44698 19848
rect 45554 19796 45560 19848
rect 45612 19836 45618 19848
rect 45741 19839 45799 19845
rect 45741 19836 45753 19839
rect 45612 19808 45753 19836
rect 45612 19796 45618 19808
rect 45741 19805 45753 19808
rect 45787 19805 45799 19839
rect 45741 19799 45799 19805
rect 27985 19771 28043 19777
rect 27985 19768 27997 19771
rect 27264 19740 27997 19768
rect 27264 19700 27292 19740
rect 27985 19737 27997 19740
rect 28031 19768 28043 19771
rect 28626 19768 28632 19780
rect 28031 19740 28632 19768
rect 28031 19737 28043 19740
rect 27985 19731 28043 19737
rect 28626 19728 28632 19740
rect 28684 19728 28690 19780
rect 29362 19728 29368 19780
rect 29420 19768 29426 19780
rect 29420 19740 37872 19768
rect 29420 19728 29426 19740
rect 37844 19712 37872 19740
rect 42794 19728 42800 19780
rect 42852 19728 42858 19780
rect 42981 19771 43039 19777
rect 42981 19737 42993 19771
rect 43027 19768 43039 19771
rect 43364 19768 43392 19796
rect 43027 19740 43392 19768
rect 43027 19737 43039 19740
rect 42981 19731 43039 19737
rect 25792 19672 27292 19700
rect 24765 19663 24823 19669
rect 27430 19660 27436 19712
rect 27488 19660 27494 19712
rect 27890 19660 27896 19712
rect 27948 19660 27954 19712
rect 29270 19660 29276 19712
rect 29328 19660 29334 19712
rect 31849 19703 31907 19709
rect 31849 19669 31861 19703
rect 31895 19700 31907 19703
rect 32490 19700 32496 19712
rect 31895 19672 32496 19700
rect 31895 19669 31907 19672
rect 31849 19663 31907 19669
rect 32490 19660 32496 19672
rect 32548 19660 32554 19712
rect 37826 19660 37832 19712
rect 37884 19660 37890 19712
rect 44174 19660 44180 19712
rect 44232 19660 44238 19712
rect 44358 19660 44364 19712
rect 44416 19700 44422 19712
rect 44821 19703 44879 19709
rect 44821 19700 44833 19703
rect 44416 19672 44833 19700
rect 44416 19660 44422 19672
rect 44821 19669 44833 19672
rect 44867 19669 44879 19703
rect 44821 19663 44879 19669
rect 1104 19610 47104 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 47104 19610
rect 1104 19536 47104 19558
rect 1302 19456 1308 19508
rect 1360 19496 1366 19508
rect 1581 19499 1639 19505
rect 1581 19496 1593 19499
rect 1360 19468 1593 19496
rect 1360 19456 1366 19468
rect 1581 19465 1593 19468
rect 1627 19465 1639 19499
rect 1581 19459 1639 19465
rect 2498 19456 2504 19508
rect 2556 19496 2562 19508
rect 2593 19499 2651 19505
rect 2593 19496 2605 19499
rect 2556 19468 2605 19496
rect 2556 19456 2562 19468
rect 2593 19465 2605 19468
rect 2639 19465 2651 19499
rect 2593 19459 2651 19465
rect 2958 19456 2964 19508
rect 3016 19456 3022 19508
rect 3050 19456 3056 19508
rect 3108 19456 3114 19508
rect 4522 19456 4528 19508
rect 4580 19496 4586 19508
rect 4893 19499 4951 19505
rect 4893 19496 4905 19499
rect 4580 19468 4905 19496
rect 4580 19456 4586 19468
rect 4893 19465 4905 19468
rect 4939 19465 4951 19499
rect 4893 19459 4951 19465
rect 5350 19456 5356 19508
rect 5408 19456 5414 19508
rect 8294 19496 8300 19508
rect 5460 19468 8300 19496
rect 3326 19428 3332 19440
rect 1412 19400 3332 19428
rect 1412 19369 1440 19400
rect 3326 19388 3332 19400
rect 3384 19388 3390 19440
rect 3780 19431 3838 19437
rect 3780 19397 3792 19431
rect 3826 19428 3838 19431
rect 3970 19428 3976 19440
rect 3826 19400 3976 19428
rect 3826 19397 3838 19400
rect 3780 19391 3838 19397
rect 3970 19388 3976 19400
rect 4028 19388 4034 19440
rect 4062 19388 4068 19440
rect 4120 19428 4126 19440
rect 5460 19428 5488 19468
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 10502 19456 10508 19508
rect 10560 19456 10566 19508
rect 11698 19456 11704 19508
rect 11756 19456 11762 19508
rect 15381 19499 15439 19505
rect 15381 19465 15393 19499
rect 15427 19465 15439 19499
rect 15381 19459 15439 19465
rect 4120 19400 5488 19428
rect 4120 19388 4126 19400
rect 6362 19388 6368 19440
rect 6420 19428 6426 19440
rect 15194 19428 15200 19440
rect 6420 19400 15200 19428
rect 6420 19388 6426 19400
rect 15194 19388 15200 19400
rect 15252 19388 15258 19440
rect 15396 19428 15424 19459
rect 17678 19456 17684 19508
rect 17736 19496 17742 19508
rect 18141 19499 18199 19505
rect 18141 19496 18153 19499
rect 17736 19468 18153 19496
rect 17736 19456 17742 19468
rect 18141 19465 18153 19468
rect 18187 19465 18199 19499
rect 18141 19459 18199 19465
rect 20070 19456 20076 19508
rect 20128 19496 20134 19508
rect 20165 19499 20223 19505
rect 20165 19496 20177 19499
rect 20128 19468 20177 19496
rect 20128 19456 20134 19468
rect 20165 19465 20177 19468
rect 20211 19465 20223 19499
rect 20165 19459 20223 19465
rect 22649 19499 22707 19505
rect 22649 19465 22661 19499
rect 22695 19496 22707 19499
rect 24118 19496 24124 19508
rect 22695 19468 24124 19496
rect 22695 19465 22707 19468
rect 22649 19459 22707 19465
rect 24118 19456 24124 19468
rect 24176 19456 24182 19508
rect 26973 19499 27031 19505
rect 26973 19465 26985 19499
rect 27019 19465 27031 19499
rect 29270 19496 29276 19508
rect 26973 19459 27031 19465
rect 27264 19468 29276 19496
rect 20625 19431 20683 19437
rect 20625 19428 20637 19431
rect 15396 19400 20637 19428
rect 20625 19397 20637 19400
rect 20671 19397 20683 19431
rect 20625 19391 20683 19397
rect 22741 19431 22799 19437
rect 22741 19397 22753 19431
rect 22787 19428 22799 19431
rect 23290 19428 23296 19440
rect 22787 19400 23296 19428
rect 22787 19397 22799 19400
rect 22741 19391 22799 19397
rect 23290 19388 23296 19400
rect 23348 19388 23354 19440
rect 25676 19431 25734 19437
rect 25676 19397 25688 19431
rect 25722 19428 25734 19431
rect 26988 19428 27016 19459
rect 27264 19428 27292 19468
rect 25722 19400 27016 19428
rect 27080 19400 27292 19428
rect 25722 19397 25734 19400
rect 25676 19391 25734 19397
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19329 1455 19363
rect 1397 19323 1455 19329
rect 1670 19320 1676 19372
rect 1728 19360 1734 19372
rect 3513 19363 3571 19369
rect 3513 19360 3525 19363
rect 1728 19332 3525 19360
rect 1728 19320 1734 19332
rect 3513 19329 3525 19332
rect 3559 19360 3571 19363
rect 4154 19360 4160 19372
rect 3559 19332 4160 19360
rect 3559 19329 3571 19332
rect 3513 19323 3571 19329
rect 4154 19320 4160 19332
rect 4212 19320 4218 19372
rect 4798 19320 4804 19372
rect 4856 19360 4862 19372
rect 5350 19360 5356 19372
rect 4856 19332 5356 19360
rect 4856 19320 4862 19332
rect 5350 19320 5356 19332
rect 5408 19320 5414 19372
rect 5537 19363 5595 19369
rect 5537 19329 5549 19363
rect 5583 19360 5595 19363
rect 6454 19360 6460 19372
rect 5583 19332 6460 19360
rect 5583 19329 5595 19332
rect 5537 19323 5595 19329
rect 6454 19320 6460 19332
rect 6512 19320 6518 19372
rect 9398 19320 9404 19372
rect 9456 19360 9462 19372
rect 10413 19363 10471 19369
rect 10413 19360 10425 19363
rect 9456 19332 10425 19360
rect 9456 19320 9462 19332
rect 10413 19329 10425 19332
rect 10459 19360 10471 19363
rect 11422 19360 11428 19372
rect 10459 19332 11428 19360
rect 10459 19329 10471 19332
rect 10413 19323 10471 19329
rect 11422 19320 11428 19332
rect 11480 19320 11486 19372
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19360 11575 19363
rect 11563 19332 11744 19360
rect 11563 19329 11575 19332
rect 11517 19323 11575 19329
rect 3234 19252 3240 19304
rect 3292 19252 3298 19304
rect 11716 19236 11744 19332
rect 13078 19320 13084 19372
rect 13136 19320 13142 19372
rect 15746 19320 15752 19372
rect 15804 19320 15810 19372
rect 15838 19320 15844 19372
rect 15896 19320 15902 19372
rect 15948 19332 16160 19360
rect 15562 19252 15568 19304
rect 15620 19292 15626 19304
rect 15948 19301 15976 19332
rect 15933 19295 15991 19301
rect 15933 19292 15945 19295
rect 15620 19264 15945 19292
rect 15620 19252 15626 19264
rect 15933 19261 15945 19264
rect 15979 19261 15991 19295
rect 16132 19292 16160 19332
rect 18230 19320 18236 19372
rect 18288 19360 18294 19372
rect 18325 19363 18383 19369
rect 18325 19360 18337 19363
rect 18288 19332 18337 19360
rect 18288 19320 18294 19332
rect 18325 19329 18337 19332
rect 18371 19329 18383 19363
rect 18325 19323 18383 19329
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19360 20591 19363
rect 23474 19360 23480 19372
rect 20579 19332 23480 19360
rect 20579 19329 20591 19332
rect 20533 19323 20591 19329
rect 23474 19320 23480 19332
rect 23532 19320 23538 19372
rect 25409 19363 25467 19369
rect 25409 19329 25421 19363
rect 25455 19360 25467 19363
rect 26786 19360 26792 19372
rect 25455 19332 26792 19360
rect 25455 19329 25467 19332
rect 25409 19323 25467 19329
rect 26786 19320 26792 19332
rect 26844 19360 26850 19372
rect 27080 19360 27108 19400
rect 26844 19332 27108 19360
rect 26844 19320 26850 19332
rect 27154 19320 27160 19372
rect 27212 19320 27218 19372
rect 27264 19369 27292 19400
rect 27516 19431 27574 19437
rect 27516 19397 27528 19431
rect 27562 19428 27574 19431
rect 27562 19400 28764 19428
rect 27562 19397 27574 19400
rect 27516 19391 27574 19397
rect 27249 19363 27307 19369
rect 27249 19329 27261 19363
rect 27295 19329 27307 19363
rect 27249 19323 27307 19329
rect 19978 19292 19984 19304
rect 16132 19264 19984 19292
rect 15933 19255 15991 19261
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 20809 19295 20867 19301
rect 20809 19261 20821 19295
rect 20855 19261 20867 19295
rect 20809 19255 20867 19261
rect 11698 19184 11704 19236
rect 11756 19224 11762 19236
rect 11756 19196 14780 19224
rect 11756 19184 11762 19196
rect 12802 19116 12808 19168
rect 12860 19156 12866 19168
rect 12897 19159 12955 19165
rect 12897 19156 12909 19159
rect 12860 19128 12909 19156
rect 12860 19116 12866 19128
rect 12897 19125 12909 19128
rect 12943 19125 12955 19159
rect 14752 19156 14780 19196
rect 14826 19184 14832 19236
rect 14884 19224 14890 19236
rect 19058 19224 19064 19236
rect 14884 19196 19064 19224
rect 14884 19184 14890 19196
rect 19058 19184 19064 19196
rect 19116 19184 19122 19236
rect 20824 19224 20852 19255
rect 22922 19252 22928 19304
rect 22980 19252 22986 19304
rect 23014 19252 23020 19304
rect 23072 19292 23078 19304
rect 23109 19295 23167 19301
rect 23109 19292 23121 19295
rect 23072 19264 23121 19292
rect 23072 19252 23078 19264
rect 23109 19261 23121 19264
rect 23155 19261 23167 19295
rect 23109 19255 23167 19261
rect 23290 19252 23296 19304
rect 23348 19292 23354 19304
rect 23348 19264 23888 19292
rect 23348 19252 23354 19264
rect 23198 19224 23204 19236
rect 20824 19196 23204 19224
rect 23198 19184 23204 19196
rect 23256 19184 23262 19236
rect 23658 19184 23664 19236
rect 23716 19224 23722 19236
rect 23753 19227 23811 19233
rect 23753 19224 23765 19227
rect 23716 19196 23765 19224
rect 23716 19184 23722 19196
rect 23753 19193 23765 19196
rect 23799 19193 23811 19227
rect 23753 19187 23811 19193
rect 16022 19156 16028 19168
rect 14752 19128 16028 19156
rect 12897 19119 12955 19125
rect 16022 19116 16028 19128
rect 16080 19116 16086 19168
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 21450 19156 21456 19168
rect 21232 19128 21456 19156
rect 21232 19116 21238 19128
rect 21450 19116 21456 19128
rect 21508 19116 21514 19168
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22281 19159 22339 19165
rect 22281 19156 22293 19159
rect 22152 19128 22293 19156
rect 22152 19116 22158 19128
rect 22281 19125 22293 19128
rect 22327 19125 22339 19159
rect 23860 19156 23888 19264
rect 24026 19252 24032 19304
rect 24084 19252 24090 19304
rect 24118 19252 24124 19304
rect 24176 19301 24182 19304
rect 24176 19295 24204 19301
rect 24192 19261 24204 19295
rect 24176 19255 24204 19261
rect 24305 19295 24363 19301
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 24670 19292 24676 19304
rect 24351 19264 24676 19292
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 24176 19252 24182 19255
rect 24670 19252 24676 19264
rect 24728 19252 24734 19304
rect 28626 19184 28632 19236
rect 28684 19184 28690 19236
rect 28736 19233 28764 19400
rect 28902 19320 28908 19372
rect 28960 19320 28966 19372
rect 29012 19369 29040 19468
rect 29270 19456 29276 19468
rect 29328 19456 29334 19508
rect 30837 19499 30895 19505
rect 30837 19465 30849 19499
rect 30883 19496 30895 19499
rect 34054 19496 34060 19508
rect 30883 19468 34060 19496
rect 30883 19465 30895 19468
rect 30837 19459 30895 19465
rect 34054 19456 34060 19468
rect 34112 19456 34118 19508
rect 35986 19456 35992 19508
rect 36044 19496 36050 19508
rect 36354 19496 36360 19508
rect 36044 19468 36360 19496
rect 36044 19456 36050 19468
rect 36354 19456 36360 19468
rect 36412 19456 36418 19508
rect 37550 19456 37556 19508
rect 37608 19496 37614 19508
rect 37921 19499 37979 19505
rect 37921 19496 37933 19499
rect 37608 19468 37933 19496
rect 37608 19456 37614 19468
rect 37921 19465 37933 19468
rect 37967 19465 37979 19499
rect 37921 19459 37979 19465
rect 38746 19456 38752 19508
rect 38804 19496 38810 19508
rect 39577 19499 39635 19505
rect 38804 19468 39528 19496
rect 38804 19456 38810 19468
rect 31481 19431 31539 19437
rect 31481 19397 31493 19431
rect 31527 19428 31539 19431
rect 31527 19400 33640 19428
rect 31527 19397 31539 19400
rect 31481 19391 31539 19397
rect 29270 19369 29276 19372
rect 28997 19363 29055 19369
rect 28997 19329 29009 19363
rect 29043 19329 29055 19363
rect 28997 19323 29055 19329
rect 29264 19323 29276 19369
rect 29270 19320 29276 19323
rect 29328 19320 29334 19372
rect 30190 19320 30196 19372
rect 30248 19360 30254 19372
rect 30653 19363 30711 19369
rect 30653 19360 30665 19363
rect 30248 19332 30665 19360
rect 30248 19320 30254 19332
rect 30653 19329 30665 19332
rect 30699 19329 30711 19363
rect 30653 19323 30711 19329
rect 30834 19320 30840 19372
rect 30892 19360 30898 19372
rect 30929 19363 30987 19369
rect 30929 19360 30941 19363
rect 30892 19332 30941 19360
rect 30892 19320 30898 19332
rect 30929 19329 30941 19332
rect 30975 19360 30987 19363
rect 31294 19360 31300 19372
rect 30975 19332 31300 19360
rect 30975 19329 30987 19332
rect 30929 19323 30987 19329
rect 31294 19320 31300 19332
rect 31352 19320 31358 19372
rect 31389 19363 31447 19369
rect 31389 19329 31401 19363
rect 31435 19360 31447 19363
rect 31662 19360 31668 19372
rect 31435 19332 31668 19360
rect 31435 19329 31447 19332
rect 31389 19323 31447 19329
rect 31662 19320 31668 19332
rect 31720 19320 31726 19372
rect 30466 19252 30472 19304
rect 30524 19252 30530 19304
rect 31570 19292 31576 19304
rect 31531 19264 31576 19292
rect 31570 19252 31576 19264
rect 31628 19292 31634 19304
rect 31846 19292 31852 19304
rect 31628 19264 31852 19292
rect 31628 19252 31634 19264
rect 31846 19252 31852 19264
rect 31904 19252 31910 19304
rect 33502 19252 33508 19304
rect 33560 19252 33566 19304
rect 28721 19227 28779 19233
rect 28721 19193 28733 19227
rect 28767 19193 28779 19227
rect 28721 19187 28779 19193
rect 31018 19184 31024 19236
rect 31076 19184 31082 19236
rect 24210 19156 24216 19168
rect 23860 19128 24216 19156
rect 22281 19119 22339 19125
rect 24210 19116 24216 19128
rect 24268 19116 24274 19168
rect 24854 19116 24860 19168
rect 24912 19156 24918 19168
rect 24949 19159 25007 19165
rect 24949 19156 24961 19159
rect 24912 19128 24961 19156
rect 24912 19116 24918 19128
rect 24949 19125 24961 19128
rect 24995 19125 25007 19159
rect 24949 19119 25007 19125
rect 25590 19116 25596 19168
rect 25648 19156 25654 19168
rect 26789 19159 26847 19165
rect 26789 19156 26801 19159
rect 25648 19128 26801 19156
rect 25648 19116 25654 19128
rect 26789 19125 26801 19128
rect 26835 19156 26847 19159
rect 27614 19156 27620 19168
rect 26835 19128 27620 19156
rect 26835 19125 26847 19128
rect 26789 19119 26847 19125
rect 27614 19116 27620 19128
rect 27672 19116 27678 19168
rect 28166 19116 28172 19168
rect 28224 19156 28230 19168
rect 29638 19156 29644 19168
rect 28224 19128 29644 19156
rect 28224 19116 28230 19128
rect 29638 19116 29644 19128
rect 29696 19116 29702 19168
rect 30377 19159 30435 19165
rect 30377 19125 30389 19159
rect 30423 19156 30435 19159
rect 30558 19156 30564 19168
rect 30423 19128 30564 19156
rect 30423 19125 30435 19128
rect 30377 19119 30435 19125
rect 30558 19116 30564 19128
rect 30616 19116 30622 19168
rect 33612 19156 33640 19400
rect 37660 19400 38884 19428
rect 35897 19363 35955 19369
rect 35897 19329 35909 19363
rect 35943 19360 35955 19363
rect 35986 19360 35992 19372
rect 35943 19332 35992 19360
rect 35943 19329 35955 19332
rect 35897 19323 35955 19329
rect 35986 19320 35992 19332
rect 36044 19320 36050 19372
rect 33686 19252 33692 19304
rect 33744 19252 33750 19304
rect 33870 19252 33876 19304
rect 33928 19292 33934 19304
rect 34149 19295 34207 19301
rect 34149 19292 34161 19295
rect 33928 19264 34161 19292
rect 33928 19252 33934 19264
rect 34149 19261 34161 19264
rect 34195 19261 34207 19295
rect 34149 19255 34207 19261
rect 34238 19252 34244 19304
rect 34296 19292 34302 19304
rect 34425 19295 34483 19301
rect 34425 19292 34437 19295
rect 34296 19264 34437 19292
rect 34296 19252 34302 19264
rect 34425 19261 34437 19264
rect 34471 19261 34483 19295
rect 34425 19255 34483 19261
rect 34514 19252 34520 19304
rect 34572 19301 34578 19304
rect 34572 19295 34600 19301
rect 34588 19261 34600 19295
rect 34572 19255 34600 19261
rect 34701 19295 34759 19301
rect 34701 19261 34713 19295
rect 34747 19292 34759 19295
rect 34882 19292 34888 19304
rect 34747 19264 34888 19292
rect 34747 19261 34759 19264
rect 34701 19255 34759 19261
rect 34572 19252 34578 19255
rect 34882 19252 34888 19264
rect 34940 19252 34946 19304
rect 37660 19233 37688 19400
rect 37826 19320 37832 19372
rect 37884 19320 37890 19372
rect 38105 19363 38163 19369
rect 38105 19329 38117 19363
rect 38151 19360 38163 19363
rect 38151 19332 38332 19360
rect 38151 19329 38163 19332
rect 38105 19323 38163 19329
rect 38304 19292 38332 19332
rect 38378 19320 38384 19372
rect 38436 19320 38442 19372
rect 38746 19360 38752 19372
rect 38488 19332 38752 19360
rect 38488 19292 38516 19332
rect 38746 19320 38752 19332
rect 38804 19320 38810 19372
rect 38856 19369 38884 19400
rect 38841 19363 38899 19369
rect 38841 19329 38853 19363
rect 38887 19329 38899 19363
rect 39500 19360 39528 19468
rect 39577 19465 39589 19499
rect 39623 19465 39635 19499
rect 39577 19459 39635 19465
rect 43533 19499 43591 19505
rect 43533 19465 43545 19499
rect 43579 19496 43591 19499
rect 43806 19496 43812 19508
rect 43579 19468 43812 19496
rect 43579 19465 43591 19468
rect 43533 19459 43591 19465
rect 39592 19428 39620 19459
rect 43806 19456 43812 19468
rect 43864 19496 43870 19508
rect 44174 19496 44180 19508
rect 43864 19468 44180 19496
rect 43864 19456 43870 19468
rect 44174 19456 44180 19468
rect 44232 19456 44238 19508
rect 42794 19428 42800 19440
rect 39592 19400 42800 19428
rect 40221 19363 40279 19369
rect 40221 19360 40233 19363
rect 39500 19332 40233 19360
rect 38841 19323 38899 19329
rect 40221 19329 40233 19332
rect 40267 19329 40279 19363
rect 40221 19323 40279 19329
rect 38304 19264 38516 19292
rect 38562 19252 38568 19304
rect 38620 19252 38626 19304
rect 40236 19292 40264 19323
rect 40494 19320 40500 19372
rect 40552 19320 40558 19372
rect 40586 19320 40592 19372
rect 40644 19360 40650 19372
rect 40880 19369 40908 19400
rect 42794 19388 42800 19400
rect 42852 19388 42858 19440
rect 40681 19363 40739 19369
rect 40681 19360 40693 19363
rect 40644 19332 40693 19360
rect 40644 19320 40650 19332
rect 40681 19329 40693 19332
rect 40727 19329 40739 19363
rect 40681 19323 40739 19329
rect 40865 19363 40923 19369
rect 40865 19329 40877 19363
rect 40911 19329 40923 19363
rect 40865 19323 40923 19329
rect 41417 19363 41475 19369
rect 41417 19329 41429 19363
rect 41463 19329 41475 19363
rect 41417 19323 41475 19329
rect 43073 19363 43131 19369
rect 43073 19329 43085 19363
rect 43119 19360 43131 19363
rect 43346 19360 43352 19372
rect 43119 19332 43352 19360
rect 43119 19329 43131 19332
rect 43073 19323 43131 19329
rect 41322 19292 41328 19304
rect 40236 19264 41328 19292
rect 41322 19252 41328 19264
rect 41380 19292 41386 19304
rect 41432 19292 41460 19323
rect 43346 19320 43352 19332
rect 43404 19320 43410 19372
rect 44266 19320 44272 19372
rect 44324 19320 44330 19372
rect 41380 19264 41460 19292
rect 41509 19295 41567 19301
rect 41380 19252 41386 19264
rect 41509 19261 41521 19295
rect 41555 19261 41567 19295
rect 41509 19255 41567 19261
rect 42245 19295 42303 19301
rect 42245 19261 42257 19295
rect 42291 19292 42303 19295
rect 42334 19292 42340 19304
rect 42291 19264 42340 19292
rect 42291 19261 42303 19264
rect 42245 19255 42303 19261
rect 37645 19227 37703 19233
rect 37645 19193 37657 19227
rect 37691 19193 37703 19227
rect 37645 19187 37703 19193
rect 37826 19184 37832 19236
rect 37884 19224 37890 19236
rect 38197 19227 38255 19233
rect 38197 19224 38209 19227
rect 37884 19196 38209 19224
rect 37884 19184 37890 19196
rect 38197 19193 38209 19196
rect 38243 19193 38255 19227
rect 38197 19187 38255 19193
rect 38289 19227 38347 19233
rect 38289 19193 38301 19227
rect 38335 19193 38347 19227
rect 38289 19187 38347 19193
rect 35345 19159 35403 19165
rect 35345 19156 35357 19159
rect 33612 19128 35357 19156
rect 35345 19125 35357 19128
rect 35391 19125 35403 19159
rect 35345 19119 35403 19125
rect 35710 19116 35716 19168
rect 35768 19116 35774 19168
rect 38304 19156 38332 19187
rect 40586 19184 40592 19236
rect 40644 19184 40650 19236
rect 41414 19184 41420 19236
rect 41472 19224 41478 19236
rect 41524 19224 41552 19255
rect 42334 19252 42340 19264
rect 42392 19292 42398 19304
rect 44284 19292 44312 19320
rect 42392 19264 44312 19292
rect 42392 19252 42398 19264
rect 44358 19252 44364 19304
rect 44416 19252 44422 19304
rect 44637 19295 44695 19301
rect 44637 19261 44649 19295
rect 44683 19292 44695 19295
rect 45278 19292 45284 19304
rect 44683 19264 45284 19292
rect 44683 19261 44695 19264
rect 44637 19255 44695 19261
rect 45278 19252 45284 19264
rect 45336 19252 45342 19304
rect 41472 19196 41552 19224
rect 41472 19184 41478 19196
rect 39206 19156 39212 19168
rect 38304 19128 39212 19156
rect 39206 19116 39212 19128
rect 39264 19116 39270 19168
rect 42794 19116 42800 19168
rect 42852 19156 42858 19168
rect 43165 19159 43223 19165
rect 43165 19156 43177 19159
rect 42852 19128 43177 19156
rect 42852 19116 42858 19128
rect 43165 19125 43177 19128
rect 43211 19125 43223 19159
rect 43165 19119 43223 19125
rect 1104 19066 47104 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 47104 19066
rect 1104 18992 47104 19014
rect 3234 18912 3240 18964
rect 3292 18952 3298 18964
rect 3970 18952 3976 18964
rect 3292 18924 3976 18952
rect 3292 18912 3298 18924
rect 3970 18912 3976 18924
rect 4028 18912 4034 18964
rect 16669 18955 16727 18961
rect 11164 18924 16620 18952
rect 11164 18896 11192 18924
rect 10318 18844 10324 18896
rect 10376 18844 10382 18896
rect 11146 18844 11152 18896
rect 11204 18844 11210 18896
rect 15488 18893 15516 18924
rect 15473 18887 15531 18893
rect 15473 18853 15485 18887
rect 15519 18853 15531 18887
rect 15473 18847 15531 18853
rect 11238 18776 11244 18828
rect 11296 18816 11302 18828
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 11296 18788 11437 18816
rect 11296 18776 11302 18788
rect 11425 18785 11437 18788
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 11698 18776 11704 18828
rect 11756 18776 11762 18828
rect 14458 18776 14464 18828
rect 14516 18816 14522 18828
rect 14826 18816 14832 18828
rect 14516 18788 14832 18816
rect 14516 18776 14522 18788
rect 14826 18776 14832 18788
rect 14884 18776 14890 18828
rect 15102 18776 15108 18828
rect 15160 18816 15166 18828
rect 15160 18788 15792 18816
rect 15160 18776 15166 18788
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 8202 18748 8208 18760
rect 6972 18720 8208 18748
rect 6972 18708 6978 18720
rect 8202 18708 8208 18720
rect 8260 18748 8266 18760
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8260 18720 8953 18748
rect 8260 18708 8266 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 10318 18708 10324 18760
rect 10376 18748 10382 18760
rect 10505 18751 10563 18757
rect 10505 18748 10517 18751
rect 10376 18720 10517 18748
rect 10376 18708 10382 18720
rect 10505 18717 10517 18720
rect 10551 18717 10563 18751
rect 10505 18711 10563 18717
rect 10686 18708 10692 18760
rect 10744 18708 10750 18760
rect 11514 18708 11520 18760
rect 11572 18757 11578 18760
rect 11572 18751 11600 18757
rect 11588 18717 11600 18751
rect 11572 18711 11600 18717
rect 11572 18708 11578 18711
rect 12526 18708 12532 18760
rect 12584 18708 12590 18760
rect 12802 18757 12808 18760
rect 12796 18748 12808 18757
rect 12763 18720 12808 18748
rect 12796 18711 12808 18720
rect 12802 18708 12808 18711
rect 12860 18708 12866 18760
rect 14274 18708 14280 18760
rect 14332 18708 14338 18760
rect 14734 18708 14740 18760
rect 14792 18748 14798 18760
rect 15764 18757 15792 18788
rect 15930 18757 15936 18760
rect 15013 18751 15071 18757
rect 15013 18748 15025 18751
rect 14792 18720 15025 18748
rect 14792 18708 14798 18720
rect 15013 18717 15025 18720
rect 15059 18717 15071 18751
rect 15013 18711 15071 18717
rect 15749 18751 15807 18757
rect 15749 18717 15761 18751
rect 15795 18717 15807 18751
rect 15749 18711 15807 18717
rect 15887 18751 15936 18757
rect 15887 18717 15899 18751
rect 15933 18717 15936 18751
rect 15887 18711 15936 18717
rect 15930 18708 15936 18711
rect 15988 18708 15994 18760
rect 16022 18708 16028 18760
rect 16080 18708 16086 18760
rect 16592 18748 16620 18924
rect 16669 18921 16681 18955
rect 16715 18952 16727 18955
rect 16715 18924 19932 18952
rect 16715 18921 16727 18924
rect 16669 18915 16727 18921
rect 16758 18844 16764 18896
rect 16816 18884 16822 18896
rect 17310 18884 17316 18896
rect 16816 18856 17316 18884
rect 16816 18844 16822 18856
rect 17310 18844 17316 18856
rect 17368 18844 17374 18896
rect 19058 18844 19064 18896
rect 19116 18884 19122 18896
rect 19116 18856 19656 18884
rect 19116 18844 19122 18856
rect 16666 18776 16672 18828
rect 16724 18816 16730 18828
rect 17678 18816 17684 18828
rect 16724 18788 17684 18816
rect 16724 18776 16730 18788
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 17497 18751 17555 18757
rect 16592 18720 17448 18748
rect 6638 18640 6644 18692
rect 6696 18680 6702 18692
rect 7162 18683 7220 18689
rect 7162 18680 7174 18683
rect 6696 18652 7174 18680
rect 6696 18640 6702 18652
rect 7162 18649 7174 18652
rect 7208 18649 7220 18683
rect 7162 18643 7220 18649
rect 8570 18640 8576 18692
rect 8628 18680 8634 18692
rect 9186 18683 9244 18689
rect 9186 18680 9198 18683
rect 8628 18652 9198 18680
rect 8628 18640 8634 18652
rect 9186 18649 9198 18652
rect 9232 18649 9244 18683
rect 9186 18643 9244 18649
rect 12345 18683 12403 18689
rect 12345 18649 12357 18683
rect 12391 18680 12403 18683
rect 12391 18652 15056 18680
rect 12391 18649 12403 18652
rect 12345 18643 12403 18649
rect 8297 18615 8355 18621
rect 8297 18581 8309 18615
rect 8343 18612 8355 18615
rect 8386 18612 8392 18624
rect 8343 18584 8392 18612
rect 8343 18581 8355 18584
rect 8297 18575 8355 18581
rect 8386 18572 8392 18584
rect 8444 18612 8450 18624
rect 11330 18612 11336 18624
rect 8444 18584 11336 18612
rect 8444 18572 8450 18584
rect 11330 18572 11336 18584
rect 11388 18572 11394 18624
rect 13906 18572 13912 18624
rect 13964 18572 13970 18624
rect 14090 18572 14096 18624
rect 14148 18572 14154 18624
rect 15028 18612 15056 18652
rect 17310 18640 17316 18692
rect 17368 18640 17374 18692
rect 17420 18680 17448 18720
rect 17497 18717 17509 18751
rect 17543 18748 17555 18751
rect 19058 18748 19064 18760
rect 17543 18720 19064 18748
rect 17543 18717 17555 18720
rect 17497 18711 17555 18717
rect 19058 18708 19064 18720
rect 19116 18708 19122 18760
rect 19628 18757 19656 18856
rect 19794 18776 19800 18828
rect 19852 18776 19858 18828
rect 19904 18816 19932 18924
rect 20346 18912 20352 18964
rect 20404 18952 20410 18964
rect 24029 18955 24087 18961
rect 20404 18924 21496 18952
rect 20404 18912 20410 18924
rect 20073 18887 20131 18893
rect 20073 18853 20085 18887
rect 20119 18884 20131 18887
rect 21082 18884 21088 18896
rect 20119 18856 21088 18884
rect 20119 18853 20131 18856
rect 20073 18847 20131 18853
rect 21082 18844 21088 18856
rect 21140 18844 21146 18896
rect 21174 18844 21180 18896
rect 21232 18884 21238 18896
rect 21361 18887 21419 18893
rect 21361 18884 21373 18887
rect 21232 18856 21373 18884
rect 21232 18844 21238 18856
rect 21361 18853 21373 18856
rect 21407 18853 21419 18887
rect 21361 18847 21419 18853
rect 20717 18819 20775 18825
rect 19904 18788 20668 18816
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 20254 18708 20260 18760
rect 20312 18708 20318 18760
rect 20438 18708 20444 18760
rect 20496 18748 20502 18760
rect 20533 18751 20591 18757
rect 20533 18748 20545 18751
rect 20496 18720 20545 18748
rect 20496 18708 20502 18720
rect 20533 18717 20545 18720
rect 20579 18717 20591 18751
rect 20640 18748 20668 18788
rect 20717 18785 20729 18819
rect 20763 18816 20775 18819
rect 20990 18816 20996 18828
rect 20763 18788 20996 18816
rect 20763 18785 20775 18788
rect 20717 18779 20775 18785
rect 20990 18776 20996 18788
rect 21048 18776 21054 18828
rect 21468 18816 21496 18924
rect 24029 18921 24041 18955
rect 24075 18952 24087 18955
rect 24118 18952 24124 18964
rect 24075 18924 24124 18952
rect 24075 18921 24087 18924
rect 24029 18915 24087 18921
rect 24118 18912 24124 18924
rect 24176 18912 24182 18964
rect 24210 18912 24216 18964
rect 24268 18952 24274 18964
rect 24268 18924 27108 18952
rect 24268 18912 24274 18924
rect 27080 18884 27108 18924
rect 27154 18912 27160 18964
rect 27212 18952 27218 18964
rect 27433 18955 27491 18961
rect 27433 18952 27445 18955
rect 27212 18924 27445 18952
rect 27212 18912 27218 18924
rect 27433 18921 27445 18924
rect 27479 18921 27491 18955
rect 27433 18915 27491 18921
rect 29181 18955 29239 18961
rect 29181 18921 29193 18955
rect 29227 18952 29239 18955
rect 29270 18952 29276 18964
rect 29227 18924 29276 18952
rect 29227 18921 29239 18924
rect 29181 18915 29239 18921
rect 29270 18912 29276 18924
rect 29328 18912 29334 18964
rect 30098 18912 30104 18964
rect 30156 18952 30162 18964
rect 30282 18952 30288 18964
rect 30156 18924 30288 18952
rect 30156 18912 30162 18924
rect 30282 18912 30288 18924
rect 30340 18912 30346 18964
rect 37642 18952 37648 18964
rect 31772 18924 37648 18952
rect 31772 18884 31800 18924
rect 37642 18912 37648 18924
rect 37700 18952 37706 18964
rect 38289 18955 38347 18961
rect 38289 18952 38301 18955
rect 37700 18924 38301 18952
rect 37700 18912 37706 18924
rect 38289 18921 38301 18924
rect 38335 18921 38347 18955
rect 38289 18915 38347 18921
rect 38654 18912 38660 18964
rect 38712 18952 38718 18964
rect 40405 18955 40463 18961
rect 40405 18952 40417 18955
rect 38712 18924 40417 18952
rect 38712 18912 38718 18924
rect 40405 18921 40417 18924
rect 40451 18921 40463 18955
rect 40405 18915 40463 18921
rect 41322 18912 41328 18964
rect 41380 18912 41386 18964
rect 27080 18856 31800 18884
rect 38746 18844 38752 18896
rect 38804 18884 38810 18896
rect 38933 18887 38991 18893
rect 38933 18884 38945 18887
rect 38804 18856 38945 18884
rect 38804 18844 38810 18856
rect 38933 18853 38945 18856
rect 38979 18853 38991 18887
rect 38933 18847 38991 18853
rect 40313 18887 40371 18893
rect 40313 18853 40325 18887
rect 40359 18884 40371 18887
rect 41509 18887 41567 18893
rect 41509 18884 41521 18887
rect 40359 18856 41521 18884
rect 40359 18853 40371 18856
rect 40313 18847 40371 18853
rect 41509 18853 41521 18856
rect 41555 18853 41567 18887
rect 41509 18847 41567 18853
rect 21754 18819 21812 18825
rect 21754 18816 21766 18819
rect 21468 18788 21766 18816
rect 21754 18785 21766 18788
rect 21800 18785 21812 18819
rect 21754 18779 21812 18785
rect 21910 18776 21916 18828
rect 21968 18776 21974 18828
rect 23658 18776 23664 18828
rect 23716 18816 23722 18828
rect 24302 18816 24308 18828
rect 23716 18788 24308 18816
rect 23716 18776 23722 18788
rect 24302 18776 24308 18788
rect 24360 18776 24366 18828
rect 24854 18776 24860 18828
rect 24912 18776 24918 18828
rect 24949 18819 25007 18825
rect 24949 18785 24961 18819
rect 24995 18785 25007 18819
rect 24949 18779 25007 18785
rect 25501 18819 25559 18825
rect 25501 18785 25513 18819
rect 25547 18816 25559 18819
rect 25590 18816 25596 18828
rect 25547 18788 25596 18816
rect 25547 18785 25559 18788
rect 25501 18779 25559 18785
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20640 18720 20913 18748
rect 20533 18711 20591 18717
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 21634 18708 21640 18760
rect 21692 18708 21698 18760
rect 22554 18708 22560 18760
rect 22612 18748 22618 18760
rect 22649 18751 22707 18757
rect 22649 18748 22661 18751
rect 22612 18720 22661 18748
rect 22612 18708 22618 18720
rect 22649 18717 22661 18720
rect 22695 18717 22707 18751
rect 22649 18711 22707 18717
rect 22738 18708 22744 18760
rect 22796 18748 22802 18760
rect 24964 18748 24992 18779
rect 25590 18776 25596 18788
rect 25648 18776 25654 18828
rect 25682 18776 25688 18828
rect 25740 18776 25746 18828
rect 25866 18776 25872 18828
rect 25924 18816 25930 18828
rect 26145 18819 26203 18825
rect 26145 18816 26157 18819
rect 25924 18788 26157 18816
rect 25924 18776 25930 18788
rect 26145 18785 26157 18788
rect 26191 18785 26203 18819
rect 26145 18779 26203 18785
rect 26418 18776 26424 18828
rect 26476 18776 26482 18828
rect 27338 18776 27344 18828
rect 27396 18776 27402 18828
rect 27890 18776 27896 18828
rect 27948 18776 27954 18828
rect 28077 18819 28135 18825
rect 28077 18785 28089 18819
rect 28123 18816 28135 18819
rect 28166 18816 28172 18828
rect 28123 18788 28172 18816
rect 28123 18785 28135 18788
rect 28077 18779 28135 18785
rect 28166 18776 28172 18788
rect 28224 18776 28230 18828
rect 30101 18819 30159 18825
rect 30101 18816 30113 18819
rect 28460 18788 30113 18816
rect 26602 18757 26608 18760
rect 22796 18720 24992 18748
rect 26559 18751 26608 18757
rect 22796 18708 22802 18720
rect 26559 18717 26571 18751
rect 26605 18717 26608 18751
rect 26559 18711 26608 18717
rect 26602 18708 26608 18711
rect 26660 18708 26666 18760
rect 26694 18708 26700 18760
rect 26752 18708 26758 18760
rect 27614 18708 27620 18760
rect 27672 18748 27678 18760
rect 27801 18751 27859 18757
rect 27801 18748 27813 18751
rect 27672 18720 27813 18748
rect 27672 18708 27678 18720
rect 27801 18717 27813 18720
rect 27847 18717 27859 18751
rect 27801 18711 27859 18717
rect 28460 18692 28488 18788
rect 30101 18785 30113 18788
rect 30147 18785 30159 18819
rect 30101 18779 30159 18785
rect 31570 18776 31576 18828
rect 31628 18816 31634 18828
rect 31849 18819 31907 18825
rect 31849 18816 31861 18819
rect 31628 18788 31861 18816
rect 31628 18776 31634 18788
rect 31849 18785 31861 18788
rect 31895 18785 31907 18819
rect 31849 18779 31907 18785
rect 40402 18776 40408 18828
rect 40460 18816 40466 18828
rect 41414 18816 41420 18828
rect 40460 18788 41420 18816
rect 40460 18776 40466 18788
rect 41414 18776 41420 18788
rect 41472 18816 41478 18828
rect 41782 18816 41788 18828
rect 41472 18788 41788 18816
rect 41472 18776 41478 18788
rect 41782 18776 41788 18788
rect 41840 18776 41846 18828
rect 44085 18819 44143 18825
rect 44085 18785 44097 18819
rect 44131 18816 44143 18819
rect 44266 18816 44272 18828
rect 44131 18788 44272 18816
rect 44131 18785 44143 18788
rect 44085 18779 44143 18785
rect 44266 18776 44272 18788
rect 44324 18776 44330 18828
rect 29365 18751 29423 18757
rect 29365 18717 29377 18751
rect 29411 18748 29423 18751
rect 29411 18720 29592 18748
rect 29411 18717 29423 18720
rect 29365 18711 29423 18717
rect 17678 18680 17684 18692
rect 17420 18652 17684 18680
rect 17678 18640 17684 18652
rect 17736 18640 17742 18692
rect 17948 18683 18006 18689
rect 17948 18649 17960 18683
rect 17994 18680 18006 18683
rect 18690 18680 18696 18692
rect 17994 18652 18696 18680
rect 17994 18649 18006 18652
rect 17948 18643 18006 18649
rect 18690 18640 18696 18652
rect 18748 18640 18754 18692
rect 20346 18680 20352 18692
rect 18800 18652 20352 18680
rect 18800 18612 18828 18652
rect 20346 18640 20352 18652
rect 20404 18640 20410 18692
rect 22462 18640 22468 18692
rect 22520 18680 22526 18692
rect 22894 18683 22952 18689
rect 22894 18680 22906 18683
rect 22520 18652 22906 18680
rect 22520 18640 22526 18652
rect 22894 18649 22906 18652
rect 22940 18649 22952 18683
rect 24946 18680 24952 18692
rect 22894 18643 22952 18649
rect 23400 18652 24952 18680
rect 15028 18584 18828 18612
rect 19242 18572 19248 18624
rect 19300 18572 19306 18624
rect 19702 18572 19708 18624
rect 19760 18572 19766 18624
rect 20438 18572 20444 18624
rect 20496 18572 20502 18624
rect 22557 18615 22615 18621
rect 22557 18581 22569 18615
rect 22603 18612 22615 18615
rect 23400 18612 23428 18652
rect 24946 18640 24952 18652
rect 25004 18640 25010 18692
rect 27522 18640 27528 18692
rect 27580 18680 27586 18692
rect 28442 18680 28448 18692
rect 27580 18652 28448 18680
rect 27580 18640 27586 18652
rect 28442 18640 28448 18652
rect 28500 18640 28506 18692
rect 22603 18584 23428 18612
rect 22603 18581 22615 18584
rect 22557 18575 22615 18581
rect 23474 18572 23480 18624
rect 23532 18612 23538 18624
rect 24397 18615 24455 18621
rect 24397 18612 24409 18615
rect 23532 18584 24409 18612
rect 23532 18572 23538 18584
rect 24397 18581 24409 18584
rect 24443 18581 24455 18615
rect 24397 18575 24455 18581
rect 24765 18615 24823 18621
rect 24765 18581 24777 18615
rect 24811 18612 24823 18615
rect 27430 18612 27436 18624
rect 24811 18584 27436 18612
rect 24811 18581 24823 18584
rect 24765 18575 24823 18581
rect 27430 18572 27436 18584
rect 27488 18572 27494 18624
rect 29564 18621 29592 18720
rect 29730 18708 29736 18760
rect 29788 18748 29794 18760
rect 30006 18748 30012 18760
rect 29788 18720 30012 18748
rect 29788 18708 29794 18720
rect 30006 18708 30012 18720
rect 30064 18708 30070 18760
rect 31754 18708 31760 18760
rect 31812 18708 31818 18760
rect 33689 18751 33747 18757
rect 33689 18717 33701 18751
rect 33735 18748 33747 18751
rect 33778 18748 33784 18760
rect 33735 18720 33784 18748
rect 33735 18717 33747 18720
rect 33689 18711 33747 18717
rect 33778 18708 33784 18720
rect 33836 18708 33842 18760
rect 33965 18751 34023 18757
rect 33965 18717 33977 18751
rect 34011 18748 34023 18751
rect 34146 18748 34152 18760
rect 34011 18720 34152 18748
rect 34011 18717 34023 18720
rect 33965 18711 34023 18717
rect 29917 18683 29975 18689
rect 29917 18649 29929 18683
rect 29963 18680 29975 18683
rect 30558 18680 30564 18692
rect 29963 18652 30564 18680
rect 29963 18649 29975 18652
rect 29917 18643 29975 18649
rect 30558 18640 30564 18652
rect 30616 18640 30622 18692
rect 32094 18683 32152 18689
rect 32094 18649 32106 18683
rect 32140 18649 32152 18683
rect 32094 18643 32152 18649
rect 29549 18615 29607 18621
rect 29549 18581 29561 18615
rect 29595 18581 29607 18615
rect 29549 18575 29607 18581
rect 31573 18615 31631 18621
rect 31573 18581 31585 18615
rect 31619 18612 31631 18615
rect 32109 18612 32137 18643
rect 32490 18640 32496 18692
rect 32548 18680 32554 18692
rect 33980 18680 34008 18711
rect 34146 18708 34152 18720
rect 34204 18708 34210 18760
rect 34330 18708 34336 18760
rect 34388 18748 34394 18760
rect 35710 18757 35716 18760
rect 35437 18751 35495 18757
rect 35437 18748 35449 18751
rect 34388 18720 35449 18748
rect 34388 18708 34394 18720
rect 35437 18717 35449 18720
rect 35483 18717 35495 18751
rect 35704 18748 35716 18757
rect 35671 18720 35716 18748
rect 35437 18711 35495 18717
rect 35704 18711 35716 18720
rect 32548 18652 34008 18680
rect 35452 18680 35480 18711
rect 35710 18708 35716 18711
rect 35768 18708 35774 18760
rect 36814 18748 36820 18760
rect 35912 18720 36820 18748
rect 35912 18680 35940 18720
rect 36814 18708 36820 18720
rect 36872 18748 36878 18760
rect 36909 18751 36967 18757
rect 36909 18748 36921 18751
rect 36872 18720 36921 18748
rect 36872 18708 36878 18720
rect 36909 18717 36921 18720
rect 36955 18717 36967 18751
rect 36909 18711 36967 18717
rect 38102 18708 38108 18760
rect 38160 18748 38166 18760
rect 38378 18748 38384 18760
rect 38160 18720 38384 18748
rect 38160 18708 38166 18720
rect 38378 18708 38384 18720
rect 38436 18708 38442 18760
rect 38654 18708 38660 18760
rect 38712 18748 38718 18760
rect 38749 18751 38807 18757
rect 38749 18748 38761 18751
rect 38712 18720 38761 18748
rect 38712 18708 38718 18720
rect 38749 18717 38761 18720
rect 38795 18717 38807 18751
rect 38749 18711 38807 18717
rect 40034 18708 40040 18760
rect 40092 18708 40098 18760
rect 40175 18751 40233 18757
rect 40175 18717 40187 18751
rect 40221 18748 40233 18751
rect 40221 18720 40448 18748
rect 40221 18717 40233 18720
rect 40175 18711 40233 18717
rect 35452 18652 35940 18680
rect 32548 18640 32554 18652
rect 36630 18640 36636 18692
rect 36688 18680 36694 18692
rect 37154 18683 37212 18689
rect 37154 18680 37166 18683
rect 36688 18652 37166 18680
rect 36688 18640 36694 18652
rect 37154 18649 37166 18652
rect 37200 18649 37212 18683
rect 37154 18643 37212 18649
rect 37826 18640 37832 18692
rect 37884 18680 37890 18692
rect 39114 18680 39120 18692
rect 37884 18652 39120 18680
rect 37884 18640 37890 18652
rect 39114 18640 39120 18652
rect 39172 18640 39178 18692
rect 40420 18680 40448 18720
rect 40494 18708 40500 18760
rect 40552 18708 40558 18760
rect 40586 18708 40592 18760
rect 40644 18748 40650 18760
rect 40898 18751 40956 18757
rect 40898 18748 40910 18751
rect 40644 18720 40910 18748
rect 40644 18708 40650 18720
rect 40898 18717 40910 18720
rect 40944 18748 40956 18751
rect 41138 18748 41144 18760
rect 40944 18720 41144 18748
rect 40944 18717 40956 18720
rect 40898 18711 40956 18717
rect 41138 18708 41144 18720
rect 41196 18708 41202 18760
rect 41509 18751 41567 18757
rect 41509 18748 41521 18751
rect 41386 18720 41521 18748
rect 41386 18680 41414 18720
rect 41509 18717 41521 18720
rect 41555 18717 41567 18751
rect 41509 18711 41567 18717
rect 41693 18751 41751 18757
rect 41693 18717 41705 18751
rect 41739 18748 41751 18751
rect 42058 18748 42064 18760
rect 41739 18720 42064 18748
rect 41739 18717 41751 18720
rect 41693 18711 41751 18717
rect 42058 18708 42064 18720
rect 42116 18708 42122 18760
rect 44177 18751 44235 18757
rect 44177 18717 44189 18751
rect 44223 18748 44235 18751
rect 44223 18720 44312 18748
rect 44223 18717 44235 18720
rect 44177 18711 44235 18717
rect 44284 18692 44312 18720
rect 44542 18708 44548 18760
rect 44600 18708 44606 18760
rect 44726 18708 44732 18760
rect 44784 18708 44790 18760
rect 46106 18708 46112 18760
rect 46164 18708 46170 18760
rect 40420 18652 40632 18680
rect 40604 18624 40632 18652
rect 40788 18652 41414 18680
rect 31619 18584 32137 18612
rect 31619 18581 31631 18584
rect 31573 18575 31631 18581
rect 32582 18572 32588 18624
rect 32640 18612 32646 18624
rect 33229 18615 33287 18621
rect 33229 18612 33241 18615
rect 32640 18584 33241 18612
rect 32640 18572 32646 18584
rect 33229 18581 33241 18584
rect 33275 18581 33287 18615
rect 33229 18575 33287 18581
rect 36078 18572 36084 18624
rect 36136 18612 36142 18624
rect 36817 18615 36875 18621
rect 36817 18612 36829 18615
rect 36136 18584 36829 18612
rect 36136 18572 36142 18584
rect 36817 18581 36829 18584
rect 36863 18581 36875 18615
rect 36817 18575 36875 18581
rect 37918 18572 37924 18624
rect 37976 18612 37982 18624
rect 38565 18615 38623 18621
rect 38565 18612 38577 18615
rect 37976 18584 38577 18612
rect 37976 18572 37982 18584
rect 38565 18581 38577 18584
rect 38611 18581 38623 18615
rect 38565 18575 38623 18581
rect 40586 18572 40592 18624
rect 40644 18572 40650 18624
rect 40788 18621 40816 18652
rect 44266 18640 44272 18692
rect 44324 18680 44330 18692
rect 44634 18680 44640 18692
rect 44324 18652 44640 18680
rect 44324 18640 44330 18652
rect 44634 18640 44640 18652
rect 44692 18640 44698 18692
rect 40773 18615 40831 18621
rect 40773 18581 40785 18615
rect 40819 18581 40831 18615
rect 40773 18575 40831 18581
rect 40957 18615 41015 18621
rect 40957 18581 40969 18615
rect 41003 18612 41015 18615
rect 41506 18612 41512 18624
rect 41003 18584 41512 18612
rect 41003 18581 41015 18584
rect 40957 18575 41015 18581
rect 41506 18572 41512 18584
rect 41564 18572 41570 18624
rect 44818 18572 44824 18624
rect 44876 18572 44882 18624
rect 45830 18572 45836 18624
rect 45888 18612 45894 18624
rect 45925 18615 45983 18621
rect 45925 18612 45937 18615
rect 45888 18584 45937 18612
rect 45888 18572 45894 18584
rect 45925 18581 45937 18584
rect 45971 18581 45983 18615
rect 45925 18575 45983 18581
rect 1104 18522 47104 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 47104 18522
rect 1104 18448 47104 18470
rect 6365 18411 6423 18417
rect 6365 18377 6377 18411
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 2685 18343 2743 18349
rect 2685 18309 2697 18343
rect 2731 18340 2743 18343
rect 2958 18340 2964 18352
rect 2731 18312 2964 18340
rect 2731 18309 2743 18312
rect 2685 18303 2743 18309
rect 2958 18300 2964 18312
rect 3016 18340 3022 18352
rect 3418 18340 3424 18352
rect 3016 18312 3424 18340
rect 3016 18300 3022 18312
rect 3418 18300 3424 18312
rect 3476 18300 3482 18352
rect 6380 18340 6408 18371
rect 6638 18368 6644 18420
rect 6696 18368 6702 18420
rect 8294 18368 8300 18420
rect 8352 18408 8358 18420
rect 11238 18408 11244 18420
rect 8352 18380 11244 18408
rect 8352 18368 8358 18380
rect 11238 18368 11244 18380
rect 11296 18368 11302 18420
rect 14461 18411 14519 18417
rect 14461 18377 14473 18411
rect 14507 18408 14519 18411
rect 14550 18408 14556 18420
rect 14507 18380 14556 18408
rect 14507 18377 14519 18380
rect 14461 18371 14519 18377
rect 14550 18368 14556 18380
rect 14608 18408 14614 18420
rect 15562 18408 15568 18420
rect 14608 18380 15568 18408
rect 14608 18368 14614 18380
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 15746 18368 15752 18420
rect 15804 18408 15810 18420
rect 16393 18411 16451 18417
rect 16393 18408 16405 18411
rect 15804 18380 16405 18408
rect 15804 18368 15810 18380
rect 16393 18377 16405 18380
rect 16439 18377 16451 18411
rect 16393 18371 16451 18377
rect 18322 18368 18328 18420
rect 18380 18368 18386 18420
rect 18690 18368 18696 18420
rect 18748 18368 18754 18420
rect 20254 18417 20260 18420
rect 20211 18411 20260 18417
rect 20211 18377 20223 18411
rect 20257 18377 20260 18411
rect 20211 18371 20260 18377
rect 20254 18368 20260 18371
rect 20312 18368 20318 18420
rect 21913 18411 21971 18417
rect 21913 18377 21925 18411
rect 21959 18408 21971 18411
rect 22462 18408 22468 18420
rect 21959 18380 22468 18408
rect 21959 18377 21971 18380
rect 21913 18371 21971 18377
rect 22462 18368 22468 18380
rect 22520 18368 22526 18420
rect 24857 18411 24915 18417
rect 24857 18408 24869 18411
rect 23216 18380 24869 18408
rect 7162 18343 7220 18349
rect 7162 18340 7174 18343
rect 6380 18312 7174 18340
rect 7162 18309 7174 18312
rect 7208 18309 7220 18343
rect 7162 18303 7220 18309
rect 9674 18300 9680 18352
rect 9732 18340 9738 18352
rect 10198 18343 10256 18349
rect 10198 18340 10210 18343
rect 9732 18312 10210 18340
rect 9732 18300 9738 18312
rect 10198 18309 10210 18312
rect 10244 18309 10256 18343
rect 10198 18303 10256 18309
rect 10410 18300 10416 18352
rect 10468 18340 10474 18352
rect 13348 18343 13406 18349
rect 10468 18312 12020 18340
rect 10468 18300 10474 18312
rect 1394 18232 1400 18284
rect 1452 18272 1458 18284
rect 2133 18275 2191 18281
rect 2133 18272 2145 18275
rect 1452 18244 2145 18272
rect 1452 18232 1458 18244
rect 2133 18241 2145 18244
rect 2179 18272 2191 18275
rect 3050 18272 3056 18284
rect 2179 18244 3056 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 3878 18232 3884 18284
rect 3936 18272 3942 18284
rect 4689 18275 4747 18281
rect 4689 18272 4701 18275
rect 3936 18244 4701 18272
rect 3936 18232 3942 18244
rect 4689 18241 4701 18244
rect 4735 18241 4747 18275
rect 4689 18235 4747 18241
rect 6549 18275 6607 18281
rect 6549 18241 6561 18275
rect 6595 18241 6607 18275
rect 6549 18235 6607 18241
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18272 6883 18275
rect 7558 18272 7564 18284
rect 6871 18244 7564 18272
rect 6871 18241 6883 18244
rect 6825 18235 6883 18241
rect 2222 18164 2228 18216
rect 2280 18164 2286 18216
rect 2409 18207 2467 18213
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 3602 18204 3608 18216
rect 2455 18176 3608 18204
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 3602 18164 3608 18176
rect 3660 18164 3666 18216
rect 4430 18164 4436 18216
rect 4488 18164 4494 18216
rect 1765 18139 1823 18145
rect 1765 18105 1777 18139
rect 1811 18136 1823 18139
rect 3326 18136 3332 18148
rect 1811 18108 3332 18136
rect 1811 18105 1823 18108
rect 1765 18099 1823 18105
rect 3326 18096 3332 18108
rect 3384 18096 3390 18148
rect 6564 18136 6592 18235
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 8202 18232 8208 18284
rect 8260 18272 8266 18284
rect 8849 18275 8907 18281
rect 8849 18272 8861 18275
rect 8260 18244 8861 18272
rect 8260 18232 8266 18244
rect 8849 18241 8861 18244
rect 8895 18241 8907 18275
rect 8849 18235 8907 18241
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18272 9919 18275
rect 11885 18275 11943 18281
rect 9907 18244 11560 18272
rect 9907 18241 9919 18244
rect 9861 18235 9919 18241
rect 6914 18164 6920 18216
rect 6972 18164 6978 18216
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 9398 18204 9404 18216
rect 8619 18176 9404 18204
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 9398 18164 9404 18176
rect 9456 18204 9462 18216
rect 9766 18204 9772 18216
rect 9456 18176 9772 18204
rect 9456 18164 9462 18176
rect 9766 18164 9772 18176
rect 9824 18204 9830 18216
rect 9953 18207 10011 18213
rect 9953 18204 9965 18207
rect 9824 18176 9965 18204
rect 9824 18164 9830 18176
rect 9953 18173 9965 18176
rect 9999 18173 10011 18207
rect 9953 18167 10011 18173
rect 6564 18108 6914 18136
rect 4614 18028 4620 18080
rect 4672 18068 4678 18080
rect 5442 18068 5448 18080
rect 4672 18040 5448 18068
rect 4672 18028 4678 18040
rect 5442 18028 5448 18040
rect 5500 18068 5506 18080
rect 5813 18071 5871 18077
rect 5813 18068 5825 18071
rect 5500 18040 5825 18068
rect 5500 18028 5506 18040
rect 5813 18037 5825 18040
rect 5859 18037 5871 18071
rect 6886 18068 6914 18108
rect 9674 18096 9680 18148
rect 9732 18096 9738 18148
rect 11532 18145 11560 18244
rect 11885 18241 11897 18275
rect 11931 18241 11943 18275
rect 11992 18272 12020 18312
rect 13348 18309 13360 18343
rect 13394 18340 13406 18343
rect 14090 18340 14096 18352
rect 13394 18312 14096 18340
rect 13394 18309 13406 18312
rect 13348 18303 13406 18309
rect 14090 18300 14096 18312
rect 14148 18300 14154 18352
rect 16316 18312 19380 18340
rect 11992 18244 12112 18272
rect 11885 18235 11943 18241
rect 11517 18139 11575 18145
rect 11517 18105 11529 18139
rect 11563 18105 11575 18139
rect 11517 18099 11575 18105
rect 7282 18068 7288 18080
rect 6886 18040 7288 18068
rect 5813 18031 5871 18037
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 10686 18028 10692 18080
rect 10744 18068 10750 18080
rect 11333 18071 11391 18077
rect 11333 18068 11345 18071
rect 10744 18040 11345 18068
rect 10744 18028 10750 18040
rect 11333 18037 11345 18040
rect 11379 18068 11391 18071
rect 11900 18068 11928 18235
rect 11974 18164 11980 18216
rect 12032 18164 12038 18216
rect 12084 18213 12112 18244
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 13081 18275 13139 18281
rect 13081 18272 13093 18275
rect 12584 18244 13093 18272
rect 12584 18232 12590 18244
rect 13081 18241 13093 18244
rect 13127 18272 13139 18275
rect 13814 18272 13820 18284
rect 13127 18244 13820 18272
rect 13127 18241 13139 18244
rect 13081 18235 13139 18241
rect 13814 18232 13820 18244
rect 13872 18232 13878 18284
rect 13906 18232 13912 18284
rect 13964 18272 13970 18284
rect 13964 18244 14872 18272
rect 13964 18232 13970 18244
rect 12069 18207 12127 18213
rect 12069 18173 12081 18207
rect 12115 18173 12127 18207
rect 12069 18167 12127 18173
rect 14458 18164 14464 18216
rect 14516 18204 14522 18216
rect 14553 18207 14611 18213
rect 14553 18204 14565 18207
rect 14516 18176 14565 18204
rect 14516 18164 14522 18176
rect 14553 18173 14565 18176
rect 14599 18173 14611 18207
rect 14553 18167 14611 18173
rect 14734 18164 14740 18216
rect 14792 18164 14798 18216
rect 14844 18204 14872 18244
rect 15746 18232 15752 18284
rect 15804 18232 15810 18284
rect 15102 18204 15108 18216
rect 14844 18176 15108 18204
rect 15102 18164 15108 18176
rect 15160 18204 15166 18216
rect 15473 18207 15531 18213
rect 15473 18204 15485 18207
rect 15160 18176 15485 18204
rect 15160 18164 15166 18176
rect 15473 18173 15485 18176
rect 15519 18173 15531 18207
rect 15473 18167 15531 18173
rect 15562 18164 15568 18216
rect 15620 18213 15626 18216
rect 15620 18207 15669 18213
rect 15620 18173 15623 18207
rect 15657 18204 15669 18207
rect 15930 18204 15936 18216
rect 15657 18176 15936 18204
rect 15657 18173 15669 18176
rect 15620 18167 15669 18173
rect 15620 18164 15626 18167
rect 15930 18164 15936 18176
rect 15988 18164 15994 18216
rect 16114 18164 16120 18216
rect 16172 18204 16178 18216
rect 16316 18204 16344 18312
rect 16925 18275 16983 18281
rect 16925 18272 16937 18275
rect 16172 18176 16344 18204
rect 16408 18244 16937 18272
rect 16172 18164 16178 18176
rect 11379 18040 11928 18068
rect 14752 18068 14780 18164
rect 15197 18139 15255 18145
rect 15197 18105 15209 18139
rect 15243 18136 15255 18139
rect 15286 18136 15292 18148
rect 15243 18108 15292 18136
rect 15243 18105 15255 18108
rect 15197 18099 15255 18105
rect 15286 18096 15292 18108
rect 15344 18096 15350 18148
rect 16298 18096 16304 18148
rect 16356 18136 16362 18148
rect 16408 18136 16436 18244
rect 16925 18241 16937 18244
rect 16971 18241 16983 18275
rect 16925 18235 16983 18241
rect 18141 18275 18199 18281
rect 18141 18241 18153 18275
rect 18187 18241 18199 18275
rect 18141 18235 18199 18241
rect 18877 18275 18935 18281
rect 18877 18241 18889 18275
rect 18923 18272 18935 18275
rect 19242 18272 19248 18284
rect 18923 18244 19248 18272
rect 18923 18241 18935 18244
rect 18877 18235 18935 18241
rect 16666 18164 16672 18216
rect 16724 18164 16730 18216
rect 18156 18204 18184 18235
rect 19242 18232 19248 18244
rect 19300 18232 19306 18284
rect 19352 18272 19380 18312
rect 21634 18300 21640 18352
rect 21692 18340 21698 18352
rect 23216 18340 23244 18380
rect 24857 18377 24869 18380
rect 24903 18377 24915 18411
rect 24857 18371 24915 18377
rect 24946 18368 24952 18420
rect 25004 18408 25010 18420
rect 29362 18408 29368 18420
rect 25004 18380 29368 18408
rect 25004 18368 25010 18380
rect 29362 18368 29368 18380
rect 29420 18368 29426 18420
rect 30006 18408 30012 18420
rect 29472 18380 30012 18408
rect 21692 18312 23244 18340
rect 21692 18300 21698 18312
rect 22002 18272 22008 18284
rect 19352 18244 22008 18272
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 22094 18232 22100 18284
rect 22152 18232 22158 18284
rect 23014 18232 23020 18284
rect 23072 18232 23078 18284
rect 23934 18232 23940 18284
rect 23992 18232 23998 18284
rect 24118 18281 24124 18284
rect 24075 18275 24124 18281
rect 24075 18241 24087 18275
rect 24121 18241 24124 18275
rect 24075 18235 24124 18241
rect 24118 18232 24124 18235
rect 24176 18232 24182 18284
rect 29472 18281 29500 18380
rect 30006 18368 30012 18380
rect 30064 18408 30070 18420
rect 30064 18380 30972 18408
rect 30064 18368 30070 18380
rect 30944 18340 30972 18380
rect 31110 18368 31116 18420
rect 31168 18368 31174 18420
rect 31754 18368 31760 18420
rect 31812 18408 31818 18420
rect 32125 18411 32183 18417
rect 32125 18408 32137 18411
rect 31812 18380 32137 18408
rect 31812 18368 31818 18380
rect 32125 18377 32137 18380
rect 32171 18377 32183 18411
rect 32125 18371 32183 18377
rect 32490 18368 32496 18420
rect 32548 18368 32554 18420
rect 32582 18368 32588 18420
rect 32640 18368 32646 18420
rect 33686 18368 33692 18420
rect 33744 18408 33750 18420
rect 33744 18380 35204 18408
rect 33744 18368 33750 18380
rect 32600 18340 32628 18368
rect 30944 18312 32628 18340
rect 35176 18340 35204 18380
rect 35250 18368 35256 18420
rect 35308 18408 35314 18420
rect 35526 18408 35532 18420
rect 35308 18380 35532 18408
rect 35308 18368 35314 18380
rect 35526 18368 35532 18380
rect 35584 18368 35590 18420
rect 35713 18411 35771 18417
rect 35713 18377 35725 18411
rect 35759 18408 35771 18411
rect 35986 18408 35992 18420
rect 35759 18380 35992 18408
rect 35759 18377 35771 18380
rect 35713 18371 35771 18377
rect 35986 18368 35992 18380
rect 36044 18368 36050 18420
rect 36170 18368 36176 18420
rect 36228 18368 36234 18420
rect 36630 18368 36636 18420
rect 36688 18368 36694 18420
rect 37277 18411 37335 18417
rect 37277 18377 37289 18411
rect 37323 18377 37335 18411
rect 37277 18371 37335 18377
rect 36078 18340 36084 18352
rect 35176 18312 36084 18340
rect 36078 18300 36084 18312
rect 36136 18300 36142 18352
rect 29457 18275 29515 18281
rect 29457 18241 29469 18275
rect 29503 18241 29515 18275
rect 29457 18235 29515 18241
rect 30466 18232 30472 18284
rect 30524 18232 30530 18284
rect 33686 18232 33692 18284
rect 33744 18232 33750 18284
rect 34514 18232 34520 18284
rect 34572 18281 34578 18284
rect 34572 18275 34600 18281
rect 34588 18241 34600 18275
rect 34572 18235 34600 18241
rect 36817 18275 36875 18281
rect 36817 18241 36829 18275
rect 36863 18272 36875 18275
rect 37292 18272 37320 18371
rect 37642 18368 37648 18420
rect 37700 18368 37706 18420
rect 40034 18368 40040 18420
rect 40092 18408 40098 18420
rect 40770 18408 40776 18420
rect 40092 18380 40776 18408
rect 40092 18368 40098 18380
rect 40770 18368 40776 18380
rect 40828 18408 40834 18420
rect 41325 18411 41383 18417
rect 41325 18408 41337 18411
rect 40828 18380 41337 18408
rect 40828 18368 40834 18380
rect 41325 18377 41337 18380
rect 41371 18377 41383 18411
rect 41325 18371 41383 18377
rect 44085 18411 44143 18417
rect 44085 18377 44097 18411
rect 44131 18408 44143 18411
rect 44726 18408 44732 18420
rect 44131 18380 44732 18408
rect 44131 18377 44143 18380
rect 44085 18371 44143 18377
rect 44726 18368 44732 18380
rect 44784 18368 44790 18420
rect 40310 18300 40316 18352
rect 40368 18340 40374 18352
rect 40589 18343 40647 18349
rect 40589 18340 40601 18343
rect 40368 18312 40601 18340
rect 40368 18300 40374 18312
rect 40589 18309 40601 18312
rect 40635 18309 40647 18343
rect 40865 18343 40923 18349
rect 40865 18340 40877 18343
rect 40589 18303 40647 18309
rect 40696 18312 40877 18340
rect 36863 18244 37320 18272
rect 36863 18241 36875 18244
rect 36817 18235 36875 18241
rect 34572 18232 34578 18235
rect 39114 18232 39120 18284
rect 39172 18272 39178 18284
rect 40126 18272 40132 18284
rect 39172 18244 40132 18272
rect 39172 18232 39178 18244
rect 40126 18232 40132 18244
rect 40184 18272 40190 18284
rect 40696 18272 40724 18312
rect 40865 18309 40877 18312
rect 40911 18309 40923 18343
rect 46293 18343 46351 18349
rect 46293 18340 46305 18343
rect 40865 18303 40923 18309
rect 41156 18312 46305 18340
rect 40184 18244 40724 18272
rect 40773 18275 40831 18281
rect 40184 18232 40190 18244
rect 40773 18241 40785 18275
rect 40819 18241 40831 18275
rect 40773 18235 40831 18241
rect 40993 18275 41051 18281
rect 40993 18241 41005 18275
rect 41039 18272 41051 18275
rect 41156 18272 41184 18312
rect 46293 18309 46305 18312
rect 46339 18309 46351 18343
rect 46293 18303 46351 18309
rect 41039 18244 41184 18272
rect 41325 18275 41383 18281
rect 41039 18241 41051 18244
rect 40993 18235 41051 18241
rect 41325 18241 41337 18275
rect 41371 18241 41383 18275
rect 41325 18235 41383 18241
rect 19150 18204 19156 18216
rect 18156 18176 19156 18204
rect 18892 18148 18920 18176
rect 19150 18164 19156 18176
rect 19208 18164 19214 18216
rect 19978 18164 19984 18216
rect 20036 18204 20042 18216
rect 22738 18204 22744 18216
rect 20036 18176 22744 18204
rect 20036 18164 20042 18176
rect 22738 18164 22744 18176
rect 22796 18164 22802 18216
rect 23201 18207 23259 18213
rect 23201 18173 23213 18207
rect 23247 18204 23259 18207
rect 23290 18204 23296 18216
rect 23247 18176 23296 18204
rect 23247 18173 23259 18176
rect 23201 18167 23259 18173
rect 23290 18164 23296 18176
rect 23348 18164 23354 18216
rect 24213 18207 24271 18213
rect 24213 18204 24225 18207
rect 23584 18176 24225 18204
rect 16356 18108 16436 18136
rect 16356 18096 16362 18108
rect 17678 18096 17684 18148
rect 17736 18136 17742 18148
rect 17736 18108 18184 18136
rect 17736 18096 17742 18108
rect 17310 18068 17316 18080
rect 14752 18040 17316 18068
rect 11379 18037 11391 18040
rect 11333 18031 11391 18037
rect 17310 18028 17316 18040
rect 17368 18068 17374 18080
rect 18049 18071 18107 18077
rect 18049 18068 18061 18071
rect 17368 18040 18061 18068
rect 17368 18028 17374 18040
rect 18049 18037 18061 18040
rect 18095 18037 18107 18071
rect 18156 18068 18184 18108
rect 18874 18096 18880 18148
rect 18932 18096 18938 18148
rect 19794 18096 19800 18148
rect 19852 18136 19858 18148
rect 22278 18136 22284 18148
rect 19852 18108 22284 18136
rect 19852 18096 19858 18108
rect 22278 18096 22284 18108
rect 22336 18096 22342 18148
rect 22462 18096 22468 18148
rect 22520 18136 22526 18148
rect 23584 18136 23612 18176
rect 24213 18173 24225 18176
rect 24259 18204 24271 18207
rect 25498 18204 25504 18216
rect 24259 18176 25504 18204
rect 24259 18173 24271 18176
rect 24213 18167 24271 18173
rect 25498 18164 25504 18176
rect 25556 18204 25562 18216
rect 26694 18204 26700 18216
rect 25556 18176 26700 18204
rect 25556 18164 25562 18176
rect 26694 18164 26700 18176
rect 26752 18164 26758 18216
rect 29273 18207 29331 18213
rect 29273 18173 29285 18207
rect 29319 18204 29331 18207
rect 29822 18204 29828 18216
rect 29319 18176 29828 18204
rect 29319 18173 29331 18176
rect 29273 18167 29331 18173
rect 29822 18164 29828 18176
rect 29880 18164 29886 18216
rect 30193 18207 30251 18213
rect 30193 18204 30205 18207
rect 30024 18176 30205 18204
rect 22520 18108 23612 18136
rect 23661 18139 23719 18145
rect 22520 18096 22526 18108
rect 23661 18105 23673 18139
rect 23707 18105 23719 18139
rect 23661 18099 23719 18105
rect 23676 18068 23704 18099
rect 24670 18096 24676 18148
rect 24728 18136 24734 18148
rect 26234 18136 26240 18148
rect 24728 18108 26240 18136
rect 24728 18096 24734 18108
rect 26234 18096 26240 18108
rect 26292 18136 26298 18148
rect 26878 18136 26884 18148
rect 26292 18108 26884 18136
rect 26292 18096 26298 18108
rect 26878 18096 26884 18108
rect 26936 18096 26942 18148
rect 29454 18096 29460 18148
rect 29512 18136 29518 18148
rect 29917 18139 29975 18145
rect 29917 18136 29929 18139
rect 29512 18108 29929 18136
rect 29512 18096 29518 18108
rect 29917 18105 29929 18108
rect 29963 18105 29975 18139
rect 29917 18099 29975 18105
rect 25866 18068 25872 18080
rect 18156 18040 25872 18068
rect 18049 18031 18107 18037
rect 25866 18028 25872 18040
rect 25924 18028 25930 18080
rect 26142 18028 26148 18080
rect 26200 18068 26206 18080
rect 29086 18068 29092 18080
rect 26200 18040 29092 18068
rect 26200 18028 26206 18040
rect 29086 18028 29092 18040
rect 29144 18068 29150 18080
rect 29730 18068 29736 18080
rect 29144 18040 29736 18068
rect 29144 18028 29150 18040
rect 29730 18028 29736 18040
rect 29788 18028 29794 18080
rect 30024 18068 30052 18176
rect 30193 18173 30205 18176
rect 30239 18173 30251 18207
rect 30193 18167 30251 18173
rect 30282 18164 30288 18216
rect 30340 18213 30346 18216
rect 30340 18207 30368 18213
rect 30356 18173 30368 18207
rect 30340 18167 30368 18173
rect 32677 18207 32735 18213
rect 32677 18173 32689 18207
rect 32723 18173 32735 18207
rect 32677 18167 32735 18173
rect 30340 18164 30346 18167
rect 32692 18136 32720 18167
rect 33502 18164 33508 18216
rect 33560 18204 33566 18216
rect 33870 18204 33876 18216
rect 33560 18176 33876 18204
rect 33560 18164 33566 18176
rect 33870 18164 33876 18176
rect 33928 18164 33934 18216
rect 34238 18164 34244 18216
rect 34296 18204 34302 18216
rect 34425 18207 34483 18213
rect 34425 18204 34437 18207
rect 34296 18176 34437 18204
rect 34296 18164 34302 18176
rect 34425 18173 34437 18176
rect 34471 18173 34483 18207
rect 34425 18167 34483 18173
rect 34701 18207 34759 18213
rect 34701 18173 34713 18207
rect 34747 18204 34759 18207
rect 35434 18204 35440 18216
rect 34747 18176 35440 18204
rect 34747 18173 34759 18176
rect 34701 18167 34759 18173
rect 35434 18164 35440 18176
rect 35492 18204 35498 18216
rect 36170 18204 36176 18216
rect 35492 18176 36176 18204
rect 35492 18164 35498 18176
rect 36170 18164 36176 18176
rect 36228 18164 36234 18216
rect 36262 18164 36268 18216
rect 36320 18164 36326 18216
rect 37734 18164 37740 18216
rect 37792 18164 37798 18216
rect 37829 18207 37887 18213
rect 37829 18173 37841 18207
rect 37875 18173 37887 18207
rect 37829 18167 37887 18173
rect 31726 18108 32720 18136
rect 30558 18068 30564 18080
rect 30024 18040 30564 18068
rect 30558 18028 30564 18040
rect 30616 18028 30622 18080
rect 30650 18028 30656 18080
rect 30708 18068 30714 18080
rect 31726 18068 31754 18108
rect 33134 18096 33140 18148
rect 33192 18136 33198 18148
rect 33318 18136 33324 18148
rect 33192 18108 33324 18136
rect 33192 18096 33198 18108
rect 33318 18096 33324 18108
rect 33376 18136 33382 18148
rect 34149 18139 34207 18145
rect 34149 18136 34161 18139
rect 33376 18108 34161 18136
rect 33376 18096 33382 18108
rect 34149 18105 34161 18108
rect 34195 18105 34207 18139
rect 36280 18136 36308 18164
rect 37844 18136 37872 18167
rect 40494 18164 40500 18216
rect 40552 18204 40558 18216
rect 40681 18207 40739 18213
rect 40681 18204 40693 18207
rect 40552 18176 40693 18204
rect 40552 18164 40558 18176
rect 40681 18173 40693 18176
rect 40727 18173 40739 18207
rect 40681 18167 40739 18173
rect 36280 18108 37872 18136
rect 34149 18099 34207 18105
rect 30708 18040 31754 18068
rect 30708 18028 30714 18040
rect 34054 18028 34060 18080
rect 34112 18068 34118 18080
rect 35345 18071 35403 18077
rect 35345 18068 35357 18071
rect 34112 18040 35357 18068
rect 34112 18028 34118 18040
rect 35345 18037 35357 18040
rect 35391 18037 35403 18071
rect 40788 18068 40816 18235
rect 41138 18164 41144 18216
rect 41196 18164 41202 18216
rect 41340 18204 41368 18235
rect 41414 18232 41420 18284
rect 41472 18272 41478 18284
rect 41785 18275 41843 18281
rect 41785 18272 41797 18275
rect 41472 18244 41797 18272
rect 41472 18232 41478 18244
rect 41785 18241 41797 18244
rect 41831 18272 41843 18275
rect 42429 18275 42487 18281
rect 42429 18272 42441 18275
rect 41831 18244 42441 18272
rect 41831 18241 41843 18244
rect 41785 18235 41843 18241
rect 42429 18241 42441 18244
rect 42475 18241 42487 18275
rect 42429 18235 42487 18241
rect 43806 18232 43812 18284
rect 43864 18272 43870 18284
rect 44174 18272 44180 18284
rect 43864 18244 44180 18272
rect 43864 18232 43870 18244
rect 44174 18232 44180 18244
rect 44232 18232 44238 18284
rect 45002 18232 45008 18284
rect 45060 18232 45066 18284
rect 45830 18232 45836 18284
rect 45888 18232 45894 18284
rect 41506 18204 41512 18216
rect 41340 18176 41512 18204
rect 41506 18164 41512 18176
rect 41564 18164 41570 18216
rect 41690 18164 41696 18216
rect 41748 18164 41754 18216
rect 42058 18164 42064 18216
rect 42116 18164 42122 18216
rect 42889 18207 42947 18213
rect 42889 18173 42901 18207
rect 42935 18204 42947 18207
rect 44085 18207 44143 18213
rect 44085 18204 44097 18207
rect 42935 18176 44097 18204
rect 42935 18173 42947 18176
rect 42889 18167 42947 18173
rect 44085 18173 44097 18176
rect 44131 18204 44143 18207
rect 44358 18204 44364 18216
rect 44131 18176 44364 18204
rect 44131 18173 44143 18176
rect 44085 18167 44143 18173
rect 44358 18164 44364 18176
rect 44416 18164 44422 18216
rect 44818 18164 44824 18216
rect 44876 18204 44882 18216
rect 44913 18207 44971 18213
rect 44913 18204 44925 18207
rect 44876 18176 44925 18204
rect 44876 18164 44882 18176
rect 44913 18173 44925 18176
rect 44959 18173 44971 18207
rect 44913 18167 44971 18173
rect 45373 18207 45431 18213
rect 45373 18173 45385 18207
rect 45419 18204 45431 18207
rect 45649 18207 45707 18213
rect 45649 18204 45661 18207
rect 45419 18176 45661 18204
rect 45419 18173 45431 18176
rect 45373 18167 45431 18173
rect 45649 18173 45661 18176
rect 45695 18173 45707 18207
rect 45649 18167 45707 18173
rect 41782 18096 41788 18148
rect 41840 18136 41846 18148
rect 41877 18139 41935 18145
rect 41877 18136 41889 18139
rect 41840 18108 41889 18136
rect 41840 18096 41846 18108
rect 41877 18105 41889 18108
rect 41923 18136 41935 18139
rect 41923 18108 42564 18136
rect 41923 18105 41935 18108
rect 41877 18099 41935 18105
rect 41230 18068 41236 18080
rect 40788 18040 41236 18068
rect 35345 18031 35403 18037
rect 41230 18028 41236 18040
rect 41288 18028 41294 18080
rect 41690 18028 41696 18080
rect 41748 18068 41754 18080
rect 42536 18077 42564 18108
rect 41969 18071 42027 18077
rect 41969 18068 41981 18071
rect 41748 18040 41981 18068
rect 41748 18028 41754 18040
rect 41969 18037 41981 18040
rect 42015 18037 42027 18071
rect 41969 18031 42027 18037
rect 42521 18071 42579 18077
rect 42521 18037 42533 18071
rect 42567 18037 42579 18071
rect 42521 18031 42579 18037
rect 43806 18028 43812 18080
rect 43864 18068 43870 18080
rect 43901 18071 43959 18077
rect 43901 18068 43913 18071
rect 43864 18040 43913 18068
rect 43864 18028 43870 18040
rect 43901 18037 43913 18040
rect 43947 18037 43959 18071
rect 43901 18031 43959 18037
rect 1104 17978 47104 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 47104 17978
rect 1104 17904 47104 17926
rect 2958 17824 2964 17876
rect 3016 17824 3022 17876
rect 3878 17824 3884 17876
rect 3936 17824 3942 17876
rect 4706 17824 4712 17876
rect 4764 17864 4770 17876
rect 5810 17864 5816 17876
rect 4764 17836 5816 17864
rect 4764 17824 4770 17836
rect 5810 17824 5816 17836
rect 5868 17864 5874 17876
rect 6273 17867 6331 17873
rect 6273 17864 6285 17867
rect 5868 17836 6285 17864
rect 5868 17824 5874 17836
rect 6273 17833 6285 17836
rect 6319 17833 6331 17867
rect 6273 17827 6331 17833
rect 7558 17824 7564 17876
rect 7616 17824 7622 17876
rect 8570 17824 8576 17876
rect 8628 17824 8634 17876
rect 8754 17824 8760 17876
rect 8812 17864 8818 17876
rect 8941 17867 8999 17873
rect 8941 17864 8953 17867
rect 8812 17836 8953 17864
rect 8812 17824 8818 17836
rect 8941 17833 8953 17836
rect 8987 17833 8999 17867
rect 8941 17827 8999 17833
rect 13078 17824 13084 17876
rect 13136 17824 13142 17876
rect 16298 17824 16304 17876
rect 16356 17824 16362 17876
rect 16577 17867 16635 17873
rect 16577 17864 16589 17867
rect 16500 17836 16589 17864
rect 5997 17799 6055 17805
rect 4724 17768 4936 17796
rect 4724 17740 4752 17768
rect 4246 17728 4252 17740
rect 3252 17700 4252 17728
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17660 1639 17663
rect 3252 17660 3280 17700
rect 4246 17688 4252 17700
rect 4304 17688 4310 17740
rect 4341 17731 4399 17737
rect 4341 17697 4353 17731
rect 4387 17728 4399 17731
rect 4522 17728 4528 17740
rect 4387 17700 4528 17728
rect 4387 17697 4399 17700
rect 4341 17691 4399 17697
rect 4522 17688 4528 17700
rect 4580 17688 4586 17740
rect 4706 17688 4712 17740
rect 4764 17688 4770 17740
rect 4798 17688 4804 17740
rect 4856 17688 4862 17740
rect 4908 17728 4936 17768
rect 5736 17768 5948 17796
rect 5736 17728 5764 17768
rect 4908 17700 5120 17728
rect 1627 17632 3280 17660
rect 1627 17629 1639 17632
rect 1581 17623 1639 17629
rect 3326 17620 3332 17672
rect 3384 17620 3390 17672
rect 4065 17663 4123 17669
rect 4065 17629 4077 17663
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 1848 17595 1906 17601
rect 1848 17561 1860 17595
rect 1894 17592 1906 17595
rect 1894 17564 3188 17592
rect 1894 17561 1906 17564
rect 1848 17555 1906 17561
rect 3160 17533 3188 17564
rect 3145 17527 3203 17533
rect 3145 17493 3157 17527
rect 3191 17493 3203 17527
rect 4080 17524 4108 17623
rect 4154 17620 4160 17672
rect 4212 17620 4218 17672
rect 5092 17669 5120 17700
rect 5368 17700 5764 17728
rect 5258 17669 5264 17672
rect 5077 17663 5135 17669
rect 5077 17629 5089 17663
rect 5123 17629 5135 17663
rect 5077 17623 5135 17629
rect 5215 17663 5264 17669
rect 5215 17629 5227 17663
rect 5261 17629 5264 17663
rect 5215 17623 5264 17629
rect 5258 17620 5264 17623
rect 5316 17620 5322 17672
rect 5368 17669 5396 17700
rect 5353 17663 5411 17669
rect 5353 17629 5365 17663
rect 5399 17629 5411 17663
rect 5920 17660 5948 17768
rect 5997 17765 6009 17799
rect 6043 17796 6055 17799
rect 11054 17796 11060 17808
rect 6043 17768 11060 17796
rect 6043 17765 6055 17768
rect 5997 17759 6055 17765
rect 11054 17756 11060 17768
rect 11112 17756 11118 17808
rect 15838 17796 15844 17808
rect 13372 17768 15844 17796
rect 7190 17688 7196 17740
rect 7248 17728 7254 17740
rect 8113 17731 8171 17737
rect 8113 17728 8125 17731
rect 7248 17700 8125 17728
rect 7248 17688 7254 17700
rect 8113 17697 8125 17700
rect 8159 17697 8171 17731
rect 8113 17691 8171 17697
rect 8570 17688 8576 17740
rect 8628 17728 8634 17740
rect 9490 17728 9496 17740
rect 8628 17700 9496 17728
rect 8628 17688 8634 17700
rect 9490 17688 9496 17700
rect 9548 17688 9554 17740
rect 10505 17731 10563 17737
rect 10505 17697 10517 17731
rect 10551 17728 10563 17731
rect 10686 17728 10692 17740
rect 10551 17700 10692 17728
rect 10551 17697 10563 17700
rect 10505 17691 10563 17697
rect 10686 17688 10692 17700
rect 10744 17688 10750 17740
rect 10962 17688 10968 17740
rect 11020 17688 11026 17740
rect 6086 17660 6092 17672
rect 5920 17632 6092 17660
rect 5353 17623 5411 17629
rect 6086 17620 6092 17632
rect 6144 17620 6150 17672
rect 6181 17663 6239 17669
rect 6181 17629 6193 17663
rect 6227 17629 6239 17663
rect 6181 17623 6239 17629
rect 6196 17592 6224 17623
rect 7006 17620 7012 17672
rect 7064 17660 7070 17672
rect 7466 17660 7472 17672
rect 7064 17632 7472 17660
rect 7064 17620 7070 17632
rect 7466 17620 7472 17632
rect 7524 17620 7530 17672
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17660 7987 17663
rect 8386 17660 8392 17672
rect 7975 17632 8392 17660
rect 7975 17629 7987 17632
rect 7929 17623 7987 17629
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 8754 17620 8760 17672
rect 8812 17620 8818 17672
rect 9309 17663 9367 17669
rect 9309 17629 9321 17663
rect 9355 17660 9367 17663
rect 10318 17660 10324 17672
rect 9355 17632 10324 17660
rect 9355 17629 9367 17632
rect 9309 17623 9367 17629
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 11238 17620 11244 17672
rect 11296 17620 11302 17672
rect 11330 17620 11336 17672
rect 11388 17669 11394 17672
rect 11388 17663 11416 17669
rect 11404 17629 11416 17663
rect 11388 17623 11416 17629
rect 11388 17620 11394 17623
rect 11514 17620 11520 17672
rect 11572 17620 11578 17672
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17660 12219 17663
rect 13372 17660 13400 17768
rect 15838 17756 15844 17768
rect 15896 17756 15902 17808
rect 13630 17688 13636 17740
rect 13688 17688 13694 17740
rect 13814 17688 13820 17740
rect 13872 17728 13878 17740
rect 14369 17731 14427 17737
rect 14369 17728 14381 17731
rect 13872 17700 14381 17728
rect 13872 17688 13878 17700
rect 14369 17697 14381 17700
rect 14415 17728 14427 17731
rect 14458 17728 14464 17740
rect 14415 17700 14464 17728
rect 14415 17697 14427 17700
rect 14369 17691 14427 17697
rect 14458 17688 14464 17700
rect 14516 17688 14522 17740
rect 14642 17688 14648 17740
rect 14700 17728 14706 17740
rect 15102 17728 15108 17740
rect 14700 17700 15108 17728
rect 14700 17688 14706 17700
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 12207 17632 13400 17660
rect 13449 17663 13507 17669
rect 12207 17629 12219 17632
rect 12161 17623 12219 17629
rect 13449 17629 13461 17663
rect 13495 17660 13507 17663
rect 13906 17660 13912 17672
rect 13495 17632 13912 17660
rect 13495 17629 13507 17632
rect 13449 17623 13507 17629
rect 13906 17620 13912 17632
rect 13964 17620 13970 17672
rect 14090 17620 14096 17672
rect 14148 17620 14154 17672
rect 15381 17663 15439 17669
rect 15381 17629 15393 17663
rect 15427 17660 15439 17663
rect 15470 17660 15476 17672
rect 15427 17632 15476 17660
rect 15427 17629 15439 17632
rect 15381 17623 15439 17629
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 15654 17620 15660 17672
rect 15712 17620 15718 17672
rect 16500 17669 16528 17836
rect 16577 17833 16589 17836
rect 16623 17833 16635 17867
rect 16577 17827 16635 17833
rect 19702 17824 19708 17876
rect 19760 17864 19766 17876
rect 20533 17867 20591 17873
rect 20533 17864 20545 17867
rect 19760 17836 20545 17864
rect 19760 17824 19766 17836
rect 20533 17833 20545 17836
rect 20579 17833 20591 17867
rect 20533 17827 20591 17833
rect 17034 17756 17040 17808
rect 17092 17796 17098 17808
rect 20438 17796 20444 17808
rect 17092 17768 20444 17796
rect 17092 17756 17098 17768
rect 20438 17756 20444 17768
rect 20496 17756 20502 17808
rect 20548 17796 20576 17827
rect 21266 17824 21272 17876
rect 21324 17864 21330 17876
rect 21324 17836 38516 17864
rect 21324 17824 21330 17836
rect 23566 17796 23572 17808
rect 20548 17768 23572 17796
rect 23566 17756 23572 17768
rect 23624 17756 23630 17808
rect 28629 17799 28687 17805
rect 28629 17765 28641 17799
rect 28675 17796 28687 17799
rect 28675 17768 29776 17796
rect 28675 17765 28687 17768
rect 28629 17759 28687 17765
rect 17221 17731 17279 17737
rect 17221 17697 17233 17731
rect 17267 17728 17279 17731
rect 17770 17728 17776 17740
rect 17267 17700 17776 17728
rect 17267 17697 17279 17700
rect 17221 17691 17279 17697
rect 17770 17688 17776 17700
rect 17828 17728 17834 17740
rect 18322 17728 18328 17740
rect 17828 17700 18328 17728
rect 17828 17688 17834 17700
rect 18322 17688 18328 17700
rect 18380 17688 18386 17740
rect 25406 17688 25412 17740
rect 25464 17728 25470 17740
rect 28258 17728 28264 17740
rect 25464 17700 28264 17728
rect 25464 17688 25470 17700
rect 28258 17688 28264 17700
rect 28316 17688 28322 17740
rect 29086 17688 29092 17740
rect 29144 17688 29150 17740
rect 29178 17688 29184 17740
rect 29236 17688 29242 17740
rect 16485 17663 16543 17669
rect 16485 17629 16497 17663
rect 16531 17629 16543 17663
rect 16485 17623 16543 17629
rect 16945 17663 17003 17669
rect 16945 17629 16957 17663
rect 16991 17660 17003 17663
rect 17310 17660 17316 17672
rect 16991 17632 17316 17660
rect 16991 17629 17003 17632
rect 16945 17623 17003 17629
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 23198 17620 23204 17672
rect 23256 17620 23262 17672
rect 26602 17620 26608 17672
rect 26660 17620 26666 17672
rect 29748 17669 29776 17768
rect 30098 17756 30104 17808
rect 30156 17796 30162 17808
rect 30469 17799 30527 17805
rect 30469 17796 30481 17799
rect 30156 17768 30481 17796
rect 30156 17756 30162 17768
rect 30469 17765 30481 17768
rect 30515 17765 30527 17799
rect 30469 17759 30527 17765
rect 31662 17756 31668 17808
rect 31720 17756 31726 17808
rect 37734 17796 37740 17808
rect 35176 17768 37740 17796
rect 29822 17688 29828 17740
rect 29880 17688 29886 17740
rect 30006 17688 30012 17740
rect 30064 17688 30070 17740
rect 30558 17688 30564 17740
rect 30616 17728 30622 17740
rect 30745 17731 30803 17737
rect 30745 17728 30757 17731
rect 30616 17700 30757 17728
rect 30616 17688 30622 17700
rect 30745 17697 30757 17700
rect 30791 17697 30803 17731
rect 30745 17691 30803 17697
rect 31386 17688 31392 17740
rect 31444 17728 31450 17740
rect 35176 17728 35204 17768
rect 37734 17756 37740 17768
rect 37792 17796 37798 17808
rect 38381 17799 38439 17805
rect 38381 17796 38393 17799
rect 37792 17768 38393 17796
rect 37792 17756 37798 17768
rect 38381 17765 38393 17768
rect 38427 17765 38439 17799
rect 38381 17759 38439 17765
rect 31444 17700 35204 17728
rect 35253 17731 35311 17737
rect 31444 17688 31450 17700
rect 35253 17697 35265 17731
rect 35299 17728 35311 17731
rect 35526 17728 35532 17740
rect 35299 17700 35532 17728
rect 35299 17697 35311 17700
rect 35253 17691 35311 17697
rect 29733 17663 29791 17669
rect 29733 17629 29745 17663
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 30834 17620 30840 17672
rect 30892 17669 30898 17672
rect 30892 17663 30920 17669
rect 30908 17629 30920 17663
rect 30892 17623 30920 17629
rect 30892 17620 30898 17623
rect 31018 17620 31024 17672
rect 31076 17620 31082 17672
rect 34514 17620 34520 17672
rect 34572 17660 34578 17672
rect 34698 17660 34704 17672
rect 34572 17632 34704 17660
rect 34572 17620 34578 17632
rect 34698 17620 34704 17632
rect 34756 17620 34762 17672
rect 34974 17620 34980 17672
rect 35032 17660 35038 17672
rect 35268 17660 35296 17691
rect 35526 17688 35532 17700
rect 35584 17688 35590 17740
rect 35032 17632 35296 17660
rect 35032 17620 35038 17632
rect 37458 17620 37464 17672
rect 37516 17660 37522 17672
rect 37829 17663 37887 17669
rect 37829 17660 37841 17663
rect 37516 17632 37841 17660
rect 37516 17620 37522 17632
rect 37829 17629 37841 17632
rect 37875 17629 37887 17663
rect 37829 17623 37887 17629
rect 37918 17620 37924 17672
rect 37976 17660 37982 17672
rect 38202 17663 38260 17669
rect 38202 17660 38214 17663
rect 37976 17632 38214 17660
rect 37976 17620 37982 17632
rect 38202 17629 38214 17632
rect 38248 17629 38260 17663
rect 38488 17660 38516 17836
rect 41230 17824 41236 17876
rect 41288 17864 41294 17876
rect 42886 17864 42892 17876
rect 41288 17836 42892 17864
rect 41288 17824 41294 17836
rect 42886 17824 42892 17836
rect 42944 17824 42950 17876
rect 45830 17824 45836 17876
rect 45888 17824 45894 17876
rect 46106 17824 46112 17876
rect 46164 17864 46170 17876
rect 46201 17867 46259 17873
rect 46201 17864 46213 17867
rect 46164 17836 46213 17864
rect 46164 17824 46170 17836
rect 46201 17833 46213 17836
rect 46247 17833 46259 17867
rect 46201 17827 46259 17833
rect 41046 17756 41052 17808
rect 41104 17796 41110 17808
rect 44082 17796 44088 17808
rect 41104 17768 44088 17796
rect 41104 17756 41110 17768
rect 44082 17756 44088 17768
rect 44140 17756 44146 17808
rect 40402 17728 40408 17740
rect 38856 17700 40408 17728
rect 38856 17672 38884 17700
rect 40402 17688 40408 17700
rect 40460 17688 40466 17740
rect 38654 17660 38660 17672
rect 38488 17632 38660 17660
rect 38202 17623 38260 17629
rect 38654 17620 38660 17632
rect 38712 17620 38718 17672
rect 38838 17620 38844 17672
rect 38896 17620 38902 17672
rect 39942 17620 39948 17672
rect 40000 17660 40006 17672
rect 41322 17660 41328 17672
rect 40000 17632 41328 17660
rect 40000 17620 40006 17632
rect 41322 17620 41328 17632
rect 41380 17620 41386 17672
rect 44174 17620 44180 17672
rect 44232 17620 44238 17672
rect 44269 17663 44327 17669
rect 44269 17629 44281 17663
rect 44315 17629 44327 17663
rect 44269 17623 44327 17629
rect 6914 17592 6920 17604
rect 6196 17564 6920 17592
rect 4798 17524 4804 17536
rect 4080 17496 4804 17524
rect 3145 17487 3203 17493
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 5166 17484 5172 17536
rect 5224 17524 5230 17536
rect 6196 17524 6224 17564
rect 6914 17552 6920 17564
rect 6972 17552 6978 17604
rect 12406 17564 13584 17592
rect 5224 17496 6224 17524
rect 5224 17484 5230 17496
rect 7190 17484 7196 17536
rect 7248 17484 7254 17536
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 7984 17496 8033 17524
rect 7984 17484 7990 17496
rect 8021 17493 8033 17496
rect 8067 17524 8079 17527
rect 9401 17527 9459 17533
rect 9401 17524 9413 17527
rect 8067 17496 9413 17524
rect 8067 17493 8079 17496
rect 8021 17487 8079 17493
rect 9401 17493 9413 17496
rect 9447 17524 9459 17527
rect 11974 17524 11980 17536
rect 9447 17496 11980 17524
rect 9447 17493 9459 17496
rect 9401 17487 9459 17493
rect 11974 17484 11980 17496
rect 12032 17524 12038 17536
rect 12406 17524 12434 17564
rect 13556 17533 13584 17564
rect 17034 17552 17040 17604
rect 17092 17592 17098 17604
rect 20441 17595 20499 17601
rect 20441 17592 20453 17595
rect 17092 17564 20453 17592
rect 17092 17552 17098 17564
rect 20441 17561 20453 17564
rect 20487 17592 20499 17595
rect 26878 17592 26884 17604
rect 20487 17564 26884 17592
rect 20487 17561 20499 17564
rect 20441 17555 20499 17561
rect 26878 17552 26884 17564
rect 26936 17552 26942 17604
rect 33870 17552 33876 17604
rect 33928 17592 33934 17604
rect 35069 17595 35127 17601
rect 35069 17592 35081 17595
rect 33928 17564 35081 17592
rect 33928 17552 33934 17564
rect 35069 17561 35081 17564
rect 35115 17592 35127 17595
rect 35342 17592 35348 17604
rect 35115 17564 35348 17592
rect 35115 17561 35127 17564
rect 35069 17555 35127 17561
rect 35342 17552 35348 17564
rect 35400 17552 35406 17604
rect 38013 17595 38071 17601
rect 38013 17561 38025 17595
rect 38059 17561 38071 17595
rect 38013 17555 38071 17561
rect 12032 17496 12434 17524
rect 13541 17527 13599 17533
rect 12032 17484 12038 17496
rect 13541 17493 13553 17527
rect 13587 17524 13599 17527
rect 15654 17524 15660 17536
rect 13587 17496 15660 17524
rect 13587 17493 13599 17496
rect 13541 17487 13599 17493
rect 15654 17484 15660 17496
rect 15712 17484 15718 17536
rect 23014 17484 23020 17536
rect 23072 17484 23078 17536
rect 26418 17484 26424 17536
rect 26476 17484 26482 17536
rect 26694 17484 26700 17536
rect 26752 17524 26758 17536
rect 26970 17524 26976 17536
rect 26752 17496 26976 17524
rect 26752 17484 26758 17496
rect 26970 17484 26976 17496
rect 27028 17484 27034 17536
rect 28994 17484 29000 17536
rect 29052 17484 29058 17536
rect 29546 17484 29552 17536
rect 29604 17484 29610 17536
rect 30282 17484 30288 17536
rect 30340 17524 30346 17536
rect 30834 17524 30840 17536
rect 30340 17496 30840 17524
rect 30340 17484 30346 17496
rect 30834 17484 30840 17496
rect 30892 17484 30898 17536
rect 34698 17484 34704 17536
rect 34756 17484 34762 17536
rect 35158 17484 35164 17536
rect 35216 17524 35222 17536
rect 35986 17524 35992 17536
rect 35216 17496 35992 17524
rect 35216 17484 35222 17496
rect 35986 17484 35992 17496
rect 36044 17484 36050 17536
rect 38028 17524 38056 17555
rect 38102 17552 38108 17604
rect 38160 17552 38166 17604
rect 39669 17595 39727 17601
rect 39669 17561 39681 17595
rect 39715 17592 39727 17595
rect 42794 17592 42800 17604
rect 39715 17564 42800 17592
rect 39715 17561 39727 17564
rect 39669 17555 39727 17561
rect 42794 17552 42800 17564
rect 42852 17592 42858 17604
rect 43806 17592 43812 17604
rect 42852 17564 43812 17592
rect 42852 17552 42858 17564
rect 43806 17552 43812 17564
rect 43864 17592 43870 17604
rect 44284 17592 44312 17623
rect 44358 17620 44364 17672
rect 44416 17620 44422 17672
rect 44542 17620 44548 17672
rect 44600 17620 44606 17672
rect 45554 17620 45560 17672
rect 45612 17660 45618 17672
rect 45741 17663 45799 17669
rect 45741 17660 45753 17663
rect 45612 17632 45753 17660
rect 45612 17620 45618 17632
rect 45741 17629 45753 17632
rect 45787 17629 45799 17663
rect 45741 17623 45799 17629
rect 46382 17620 46388 17672
rect 46440 17620 46446 17672
rect 46750 17620 46756 17672
rect 46808 17620 46814 17672
rect 43864 17564 44312 17592
rect 43864 17552 43870 17564
rect 41874 17524 41880 17536
rect 38028 17496 41880 17524
rect 41874 17484 41880 17496
rect 41932 17484 41938 17536
rect 43901 17527 43959 17533
rect 43901 17493 43913 17527
rect 43947 17524 43959 17527
rect 45002 17524 45008 17536
rect 43947 17496 45008 17524
rect 43947 17493 43959 17496
rect 43901 17487 43959 17493
rect 45002 17484 45008 17496
rect 45060 17484 45066 17536
rect 1104 17434 47104 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 47104 17434
rect 1104 17360 47104 17382
rect 1397 17323 1455 17329
rect 1397 17289 1409 17323
rect 1443 17320 1455 17323
rect 2222 17320 2228 17332
rect 1443 17292 2228 17320
rect 1443 17289 1455 17292
rect 1397 17283 1455 17289
rect 2222 17280 2228 17292
rect 2280 17280 2286 17332
rect 3786 17280 3792 17332
rect 3844 17320 3850 17332
rect 6638 17320 6644 17332
rect 3844 17292 6644 17320
rect 3844 17280 3850 17292
rect 6638 17280 6644 17292
rect 6696 17320 6702 17332
rect 6733 17323 6791 17329
rect 6733 17320 6745 17323
rect 6696 17292 6745 17320
rect 6696 17280 6702 17292
rect 6733 17289 6745 17292
rect 6779 17289 6791 17323
rect 6733 17283 6791 17289
rect 7282 17280 7288 17332
rect 7340 17320 7346 17332
rect 7469 17323 7527 17329
rect 7469 17320 7481 17323
rect 7340 17292 7481 17320
rect 7340 17280 7346 17292
rect 7469 17289 7481 17292
rect 7515 17289 7527 17323
rect 7469 17283 7527 17289
rect 7837 17323 7895 17329
rect 7837 17289 7849 17323
rect 7883 17320 7895 17323
rect 8294 17320 8300 17332
rect 7883 17292 8300 17320
rect 7883 17289 7895 17292
rect 7837 17283 7895 17289
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 14185 17323 14243 17329
rect 14185 17289 14197 17323
rect 14231 17320 14243 17323
rect 14274 17320 14280 17332
rect 14231 17292 14280 17320
rect 14231 17289 14243 17292
rect 14185 17283 14243 17289
rect 14274 17280 14280 17292
rect 14332 17280 14338 17332
rect 14550 17280 14556 17332
rect 14608 17280 14614 17332
rect 14645 17323 14703 17329
rect 14645 17289 14657 17323
rect 14691 17320 14703 17323
rect 15654 17320 15660 17332
rect 14691 17292 15660 17320
rect 14691 17289 14703 17292
rect 14645 17283 14703 17289
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 21266 17320 21272 17332
rect 18248 17292 21272 17320
rect 6822 17212 6828 17264
rect 6880 17252 6886 17264
rect 18248 17252 18276 17292
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 22646 17320 22652 17332
rect 21560 17292 22652 17320
rect 6880 17224 18276 17252
rect 6880 17212 6886 17224
rect 20346 17212 20352 17264
rect 20404 17252 20410 17264
rect 20404 17224 20576 17252
rect 20404 17212 20410 17224
rect 934 17144 940 17196
rect 992 17184 998 17196
rect 2314 17193 2320 17196
rect 1581 17187 1639 17193
rect 1581 17184 1593 17187
rect 992 17156 1593 17184
rect 992 17144 998 17156
rect 1581 17153 1593 17156
rect 1627 17153 1639 17187
rect 1581 17147 1639 17153
rect 2308 17147 2320 17193
rect 2314 17144 2320 17147
rect 2372 17144 2378 17196
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17184 4399 17187
rect 4522 17184 4528 17196
rect 4387 17156 4528 17184
rect 4387 17153 4399 17156
rect 4341 17147 4399 17153
rect 4522 17144 4528 17156
rect 4580 17144 4586 17196
rect 6546 17144 6552 17196
rect 6604 17144 6610 17196
rect 7926 17144 7932 17196
rect 7984 17144 7990 17196
rect 14182 17144 14188 17196
rect 14240 17184 14246 17196
rect 14826 17184 14832 17196
rect 14240 17156 14832 17184
rect 14240 17144 14246 17156
rect 14826 17144 14832 17156
rect 14884 17144 14890 17196
rect 19242 17144 19248 17196
rect 19300 17144 19306 17196
rect 20548 17193 20576 17224
rect 21560 17193 21588 17292
rect 22646 17280 22652 17292
rect 22704 17320 22710 17332
rect 23474 17320 23480 17332
rect 22704 17292 23480 17320
rect 22704 17280 22710 17292
rect 23474 17280 23480 17292
rect 23532 17280 23538 17332
rect 24026 17280 24032 17332
rect 24084 17280 24090 17332
rect 25869 17323 25927 17329
rect 25869 17289 25881 17323
rect 25915 17320 25927 17323
rect 26326 17320 26332 17332
rect 25915 17292 26332 17320
rect 25915 17289 25927 17292
rect 25869 17283 25927 17289
rect 26326 17280 26332 17292
rect 26384 17280 26390 17332
rect 26510 17280 26516 17332
rect 26568 17320 26574 17332
rect 28353 17323 28411 17329
rect 28353 17320 28365 17323
rect 26568 17292 28365 17320
rect 26568 17280 26574 17292
rect 28353 17289 28365 17292
rect 28399 17289 28411 17323
rect 28353 17283 28411 17289
rect 28994 17280 29000 17332
rect 29052 17320 29058 17332
rect 29917 17323 29975 17329
rect 29917 17320 29929 17323
rect 29052 17292 29929 17320
rect 29052 17280 29058 17292
rect 29917 17289 29929 17292
rect 29963 17320 29975 17323
rect 30282 17320 30288 17332
rect 29963 17292 30288 17320
rect 29963 17289 29975 17292
rect 29917 17283 29975 17289
rect 30282 17280 30288 17292
rect 30340 17280 30346 17332
rect 33413 17323 33471 17329
rect 33413 17289 33425 17323
rect 33459 17320 33471 17323
rect 34422 17320 34428 17332
rect 33459 17292 34428 17320
rect 33459 17289 33471 17292
rect 33413 17283 33471 17289
rect 34422 17280 34428 17292
rect 34480 17280 34486 17332
rect 38289 17323 38347 17329
rect 38289 17289 38301 17323
rect 38335 17320 38347 17323
rect 38838 17320 38844 17332
rect 38335 17292 38844 17320
rect 38335 17289 38347 17292
rect 38289 17283 38347 17289
rect 38838 17280 38844 17292
rect 38896 17280 38902 17332
rect 39942 17280 39948 17332
rect 40000 17320 40006 17332
rect 40129 17323 40187 17329
rect 40129 17320 40141 17323
rect 40000 17292 40141 17320
rect 40000 17280 40006 17292
rect 40129 17289 40141 17292
rect 40175 17289 40187 17323
rect 40129 17283 40187 17289
rect 40310 17280 40316 17332
rect 40368 17320 40374 17332
rect 41230 17320 41236 17332
rect 40368 17292 41236 17320
rect 40368 17280 40374 17292
rect 41230 17280 41236 17292
rect 41288 17280 41294 17332
rect 41322 17280 41328 17332
rect 41380 17320 41386 17332
rect 42150 17320 42156 17332
rect 41380 17292 42156 17320
rect 41380 17280 41386 17292
rect 42150 17280 42156 17292
rect 42208 17280 42214 17332
rect 42242 17280 42248 17332
rect 42300 17320 42306 17332
rect 42521 17323 42579 17329
rect 42521 17320 42533 17323
rect 42300 17292 42533 17320
rect 42300 17280 42306 17292
rect 42521 17289 42533 17292
rect 42567 17289 42579 17323
rect 42521 17283 42579 17289
rect 42613 17323 42671 17329
rect 42613 17289 42625 17323
rect 42659 17320 42671 17323
rect 42794 17320 42800 17332
rect 42659 17292 42800 17320
rect 42659 17289 42671 17292
rect 42613 17283 42671 17289
rect 42794 17280 42800 17292
rect 42852 17280 42858 17332
rect 44542 17280 44548 17332
rect 44600 17280 44606 17332
rect 22916 17255 22974 17261
rect 22916 17221 22928 17255
rect 22962 17252 22974 17255
rect 23014 17252 23020 17264
rect 22962 17224 23020 17252
rect 22962 17221 22974 17224
rect 22916 17215 22974 17221
rect 23014 17212 23020 17224
rect 23072 17212 23078 17264
rect 24756 17255 24814 17261
rect 24756 17221 24768 17255
rect 24802 17252 24814 17255
rect 24854 17252 24860 17264
rect 24802 17224 24860 17252
rect 24802 17221 24814 17224
rect 24756 17215 24814 17221
rect 24854 17212 24860 17224
rect 24912 17212 24918 17264
rect 26418 17212 26424 17264
rect 26476 17252 26482 17264
rect 27218 17255 27276 17261
rect 27218 17252 27230 17255
rect 26476 17224 27230 17252
rect 26476 17212 26482 17224
rect 27218 17221 27230 17224
rect 27264 17221 27276 17255
rect 27218 17215 27276 17221
rect 28804 17255 28862 17261
rect 28804 17221 28816 17255
rect 28850 17252 28862 17255
rect 29546 17252 29552 17264
rect 28850 17224 29552 17252
rect 28850 17221 28862 17224
rect 28804 17215 28862 17221
rect 29546 17212 29552 17224
rect 29604 17212 29610 17264
rect 29822 17212 29828 17264
rect 29880 17252 29886 17264
rect 31573 17255 31631 17261
rect 31573 17252 31585 17255
rect 29880 17224 31585 17252
rect 29880 17212 29886 17224
rect 31573 17221 31585 17224
rect 31619 17252 31631 17255
rect 32122 17252 32128 17264
rect 31619 17224 32128 17252
rect 31619 17221 31631 17224
rect 31573 17215 31631 17221
rect 32122 17212 32128 17224
rect 32180 17212 32186 17264
rect 38378 17212 38384 17264
rect 38436 17252 38442 17264
rect 40589 17255 40647 17261
rect 38436 17224 38976 17252
rect 38436 17212 38442 17224
rect 20533 17187 20591 17193
rect 20533 17153 20545 17187
rect 20579 17153 20591 17187
rect 20533 17147 20591 17153
rect 21545 17187 21603 17193
rect 21545 17153 21557 17187
rect 21591 17153 21603 17187
rect 21545 17147 21603 17153
rect 22554 17144 22560 17196
rect 22612 17184 22618 17196
rect 22649 17187 22707 17193
rect 22649 17184 22661 17187
rect 22612 17156 22661 17184
rect 22612 17144 22618 17156
rect 22649 17153 22661 17156
rect 22695 17184 22707 17187
rect 24489 17187 24547 17193
rect 24489 17184 24501 17187
rect 22695 17156 24501 17184
rect 22695 17153 22707 17156
rect 22649 17147 22707 17153
rect 24489 17153 24501 17156
rect 24535 17184 24547 17187
rect 26878 17184 26884 17196
rect 24535 17156 26280 17184
rect 24535 17153 24547 17156
rect 24489 17147 24547 17153
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 2056 16980 2084 17079
rect 4154 17076 4160 17128
rect 4212 17076 4218 17128
rect 4706 17076 4712 17128
rect 4764 17116 4770 17128
rect 5258 17125 5264 17128
rect 5077 17119 5135 17125
rect 5077 17116 5089 17119
rect 4764 17088 5089 17116
rect 4764 17076 4770 17088
rect 5077 17085 5089 17088
rect 5123 17085 5135 17119
rect 5077 17079 5135 17085
rect 5215 17119 5264 17125
rect 5215 17085 5227 17119
rect 5261 17085 5264 17119
rect 5215 17079 5264 17085
rect 5258 17076 5264 17079
rect 5316 17076 5322 17128
rect 5353 17119 5411 17125
rect 5353 17085 5365 17119
rect 5399 17116 5411 17119
rect 5534 17116 5540 17128
rect 5399 17088 5540 17116
rect 5399 17085 5411 17088
rect 5353 17079 5411 17085
rect 5534 17076 5540 17088
rect 5592 17116 5598 17128
rect 6730 17116 6736 17128
rect 5592 17088 6736 17116
rect 5592 17076 5598 17088
rect 6730 17076 6736 17088
rect 6788 17076 6794 17128
rect 7834 17076 7840 17128
rect 7892 17116 7898 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7892 17088 8033 17116
rect 7892 17076 7898 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 14737 17119 14795 17125
rect 14737 17085 14749 17119
rect 14783 17116 14795 17119
rect 16206 17116 16212 17128
rect 14783 17088 16212 17116
rect 14783 17085 14795 17088
rect 14737 17079 14795 17085
rect 16206 17076 16212 17088
rect 16264 17076 16270 17128
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17116 18107 17119
rect 18138 17116 18144 17128
rect 18095 17088 18144 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18138 17076 18144 17088
rect 18196 17076 18202 17128
rect 18230 17076 18236 17128
rect 18288 17076 18294 17128
rect 18782 17076 18788 17128
rect 18840 17116 18846 17128
rect 19150 17125 19156 17128
rect 18969 17119 19027 17125
rect 18969 17116 18981 17119
rect 18840 17088 18981 17116
rect 18840 17076 18846 17088
rect 18969 17085 18981 17088
rect 19015 17085 19027 17119
rect 18969 17079 19027 17085
rect 19107 17119 19156 17125
rect 19107 17085 19119 17119
rect 19153 17085 19156 17119
rect 19107 17079 19156 17085
rect 19150 17076 19156 17079
rect 19208 17076 19214 17128
rect 19886 17076 19892 17128
rect 19944 17116 19950 17128
rect 20257 17119 20315 17125
rect 20257 17116 20269 17119
rect 19944 17088 20269 17116
rect 19944 17076 19950 17088
rect 20257 17085 20269 17088
rect 20303 17085 20315 17119
rect 20257 17079 20315 17085
rect 4172 17048 4200 17076
rect 4614 17048 4620 17060
rect 4172 17020 4620 17048
rect 4614 17008 4620 17020
rect 4672 17008 4678 17060
rect 2406 16980 2412 16992
rect 2056 16952 2412 16980
rect 2406 16940 2412 16952
rect 2464 16940 2470 16992
rect 3421 16983 3479 16989
rect 3421 16949 3433 16983
rect 3467 16980 3479 16983
rect 4724 16980 4752 17076
rect 4801 17051 4859 17057
rect 4801 17017 4813 17051
rect 4847 17017 4859 17051
rect 4801 17011 4859 17017
rect 5997 17051 6055 17057
rect 5997 17017 6009 17051
rect 6043 17048 6055 17051
rect 12342 17048 12348 17060
rect 6043 17020 12348 17048
rect 6043 17017 6055 17020
rect 5997 17011 6055 17017
rect 3467 16952 4752 16980
rect 4816 16980 4844 17011
rect 12342 17008 12348 17020
rect 12400 17008 12406 17060
rect 17954 17008 17960 17060
rect 18012 17048 18018 17060
rect 18690 17048 18696 17060
rect 18012 17020 18696 17048
rect 18012 17008 18018 17020
rect 18690 17008 18696 17020
rect 18748 17008 18754 17060
rect 19812 17020 20392 17048
rect 5350 16980 5356 16992
rect 4816 16952 5356 16980
rect 3467 16949 3479 16952
rect 3421 16943 3479 16949
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 6638 16940 6644 16992
rect 6696 16980 6702 16992
rect 7190 16980 7196 16992
rect 6696 16952 7196 16980
rect 6696 16940 6702 16952
rect 7190 16940 7196 16952
rect 7248 16980 7254 16992
rect 7834 16980 7840 16992
rect 7248 16952 7840 16980
rect 7248 16940 7254 16952
rect 7834 16940 7840 16952
rect 7892 16940 7898 16992
rect 11054 16940 11060 16992
rect 11112 16980 11118 16992
rect 13078 16980 13084 16992
rect 11112 16952 13084 16980
rect 11112 16940 11118 16952
rect 13078 16940 13084 16952
rect 13136 16940 13142 16992
rect 16942 16940 16948 16992
rect 17000 16980 17006 16992
rect 19812 16980 19840 17020
rect 17000 16952 19840 16980
rect 19889 16983 19947 16989
rect 17000 16940 17006 16952
rect 19889 16949 19901 16983
rect 19935 16980 19947 16983
rect 20070 16980 20076 16992
rect 19935 16952 20076 16980
rect 19935 16949 19947 16952
rect 19889 16943 19947 16949
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 20364 16980 20392 17020
rect 20990 16980 20996 16992
rect 20364 16952 20996 16980
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 21174 16940 21180 16992
rect 21232 16980 21238 16992
rect 21545 16983 21603 16989
rect 21545 16980 21557 16983
rect 21232 16952 21557 16980
rect 21232 16940 21238 16952
rect 21545 16949 21557 16952
rect 21591 16980 21603 16983
rect 21634 16980 21640 16992
rect 21591 16952 21640 16980
rect 21591 16949 21603 16952
rect 21545 16943 21603 16949
rect 21634 16940 21640 16952
rect 21692 16940 21698 16992
rect 25958 16940 25964 16992
rect 26016 16940 26022 16992
rect 26252 16980 26280 17156
rect 26436 17156 26884 17184
rect 26436 17125 26464 17156
rect 26878 17144 26884 17156
rect 26936 17184 26942 17196
rect 31386 17184 31392 17196
rect 26936 17156 31392 17184
rect 26936 17144 26942 17156
rect 31386 17144 31392 17156
rect 31444 17144 31450 17196
rect 31665 17187 31723 17193
rect 31665 17153 31677 17187
rect 31711 17184 31723 17187
rect 31711 17156 33180 17184
rect 31711 17153 31723 17156
rect 31665 17147 31723 17153
rect 26421 17119 26479 17125
rect 26421 17085 26433 17119
rect 26467 17085 26479 17119
rect 26421 17079 26479 17085
rect 26605 17119 26663 17125
rect 26605 17085 26617 17119
rect 26651 17116 26663 17119
rect 26694 17116 26700 17128
rect 26651 17088 26700 17116
rect 26651 17085 26663 17088
rect 26605 17079 26663 17085
rect 26694 17076 26700 17088
rect 26752 17076 26758 17128
rect 26786 17076 26792 17128
rect 26844 17116 26850 17128
rect 26973 17119 27031 17125
rect 26973 17116 26985 17119
rect 26844 17088 26985 17116
rect 26844 17076 26850 17088
rect 26973 17085 26985 17088
rect 27019 17085 27031 17119
rect 26973 17079 27031 17085
rect 28534 17076 28540 17128
rect 28592 17076 28598 17128
rect 29914 17076 29920 17128
rect 29972 17116 29978 17128
rect 31018 17116 31024 17128
rect 29972 17088 31024 17116
rect 29972 17076 29978 17088
rect 31018 17076 31024 17088
rect 31076 17076 31082 17128
rect 31849 17119 31907 17125
rect 31849 17085 31861 17119
rect 31895 17085 31907 17119
rect 33152 17116 33180 17156
rect 33226 17144 33232 17196
rect 33284 17184 33290 17196
rect 33284 17156 33640 17184
rect 33284 17144 33290 17156
rect 33612 17128 33640 17156
rect 34330 17144 34336 17196
rect 34388 17144 34394 17196
rect 34698 17144 34704 17196
rect 34756 17184 34762 17196
rect 35437 17187 35495 17193
rect 35437 17184 35449 17187
rect 34756 17156 35449 17184
rect 34756 17144 34762 17156
rect 35437 17153 35449 17156
rect 35483 17153 35495 17187
rect 35437 17147 35495 17153
rect 36078 17144 36084 17196
rect 36136 17184 36142 17196
rect 37553 17187 37611 17193
rect 37553 17184 37565 17187
rect 36136 17156 37565 17184
rect 36136 17144 36142 17156
rect 37553 17153 37565 17156
rect 37599 17153 37611 17187
rect 37553 17147 37611 17153
rect 38565 17187 38623 17193
rect 38565 17153 38577 17187
rect 38611 17153 38623 17187
rect 38565 17147 38623 17153
rect 38657 17187 38715 17193
rect 38657 17153 38669 17187
rect 38703 17153 38715 17187
rect 38657 17147 38715 17153
rect 33505 17119 33563 17125
rect 33505 17116 33517 17119
rect 33152 17088 33517 17116
rect 31849 17079 31907 17085
rect 33505 17085 33517 17088
rect 33551 17085 33563 17119
rect 33505 17079 33563 17085
rect 28552 16980 28580 17076
rect 29638 17008 29644 17060
rect 29696 17048 29702 17060
rect 30466 17048 30472 17060
rect 29696 17020 30472 17048
rect 29696 17008 29702 17020
rect 30466 17008 30472 17020
rect 30524 17048 30530 17060
rect 31864 17048 31892 17079
rect 30524 17020 31892 17048
rect 33520 17048 33548 17079
rect 33594 17076 33600 17128
rect 33652 17076 33658 17128
rect 34146 17116 34152 17128
rect 33704 17088 34152 17116
rect 33704 17048 33732 17088
rect 34146 17076 34152 17088
rect 34204 17116 34210 17128
rect 35158 17116 35164 17128
rect 34204 17088 35164 17116
rect 34204 17076 34210 17088
rect 35158 17076 35164 17088
rect 35216 17076 35222 17128
rect 37277 17119 37335 17125
rect 37277 17085 37289 17119
rect 37323 17085 37335 17119
rect 37277 17079 37335 17085
rect 33520 17020 33732 17048
rect 30524 17008 30530 17020
rect 34330 17008 34336 17060
rect 34388 17048 34394 17060
rect 34563 17051 34621 17057
rect 34563 17048 34575 17051
rect 34388 17020 34575 17048
rect 34388 17008 34394 17020
rect 34563 17017 34575 17020
rect 34609 17017 34621 17051
rect 34563 17011 34621 17017
rect 26252 16952 28580 16980
rect 31205 16983 31263 16989
rect 31205 16949 31217 16983
rect 31251 16980 31263 16983
rect 31294 16980 31300 16992
rect 31251 16952 31300 16980
rect 31251 16949 31263 16952
rect 31205 16943 31263 16949
rect 31294 16940 31300 16952
rect 31352 16940 31358 16992
rect 32858 16940 32864 16992
rect 32916 16980 32922 16992
rect 33045 16983 33103 16989
rect 33045 16980 33057 16983
rect 32916 16952 33057 16980
rect 32916 16940 32922 16952
rect 33045 16949 33057 16952
rect 33091 16949 33103 16983
rect 33045 16943 33103 16949
rect 34146 16940 34152 16992
rect 34204 16980 34210 16992
rect 34974 16980 34980 16992
rect 34204 16952 34980 16980
rect 34204 16940 34210 16952
rect 34974 16940 34980 16952
rect 35032 16940 35038 16992
rect 35253 16983 35311 16989
rect 35253 16949 35265 16983
rect 35299 16980 35311 16983
rect 35526 16980 35532 16992
rect 35299 16952 35532 16980
rect 35299 16949 35311 16952
rect 35253 16943 35311 16949
rect 35526 16940 35532 16952
rect 35584 16940 35590 16992
rect 37292 16980 37320 17079
rect 38010 16980 38016 16992
rect 37292 16952 38016 16980
rect 38010 16940 38016 16952
rect 38068 16940 38074 16992
rect 38381 16983 38439 16989
rect 38381 16949 38393 16983
rect 38427 16980 38439 16983
rect 38470 16980 38476 16992
rect 38427 16952 38476 16980
rect 38427 16949 38439 16952
rect 38381 16943 38439 16949
rect 38470 16940 38476 16952
rect 38528 16940 38534 16992
rect 38580 16980 38608 17147
rect 38672 17116 38700 17147
rect 38838 17144 38844 17196
rect 38896 17144 38902 17196
rect 38948 17193 38976 17224
rect 40589 17221 40601 17255
rect 40635 17252 40647 17255
rect 42058 17252 42064 17264
rect 40635 17224 42064 17252
rect 40635 17221 40647 17224
rect 40589 17215 40647 17221
rect 42058 17212 42064 17224
rect 42116 17212 42122 17264
rect 42260 17224 44128 17252
rect 38933 17187 38991 17193
rect 38933 17153 38945 17187
rect 38979 17153 38991 17187
rect 38933 17147 38991 17153
rect 39945 17187 40003 17193
rect 39945 17153 39957 17187
rect 39991 17184 40003 17187
rect 40034 17184 40040 17196
rect 39991 17156 40040 17184
rect 39991 17153 40003 17156
rect 39945 17147 40003 17153
rect 40034 17144 40040 17156
rect 40092 17144 40098 17196
rect 40221 17187 40279 17193
rect 40221 17153 40233 17187
rect 40267 17153 40279 17187
rect 40221 17147 40279 17153
rect 40773 17187 40831 17193
rect 40773 17153 40785 17187
rect 40819 17153 40831 17187
rect 40773 17147 40831 17153
rect 40957 17187 41015 17193
rect 40957 17153 40969 17187
rect 41003 17184 41015 17187
rect 41690 17184 41696 17196
rect 41003 17156 41696 17184
rect 41003 17153 41015 17156
rect 40957 17147 41015 17153
rect 38672 17088 38976 17116
rect 38948 17060 38976 17088
rect 39850 17076 39856 17128
rect 39908 17116 39914 17128
rect 40236 17116 40264 17147
rect 39908 17088 40264 17116
rect 39908 17076 39914 17088
rect 38930 17008 38936 17060
rect 38988 17008 38994 17060
rect 39945 17051 40003 17057
rect 39945 17017 39957 17051
rect 39991 17048 40003 17051
rect 40788 17048 40816 17147
rect 41690 17144 41696 17156
rect 41748 17144 41754 17196
rect 42260 17174 42288 17224
rect 42076 17146 42288 17174
rect 42429 17187 42487 17193
rect 42429 17153 42441 17187
rect 42475 17184 42487 17187
rect 43070 17184 43076 17196
rect 42475 17182 42656 17184
rect 42720 17182 43076 17184
rect 42475 17156 43076 17182
rect 42475 17153 42487 17156
rect 42628 17154 42748 17156
rect 42429 17147 42487 17153
rect 41049 17119 41107 17125
rect 41049 17085 41061 17119
rect 41095 17116 41107 17119
rect 41138 17116 41144 17128
rect 41095 17088 41144 17116
rect 41095 17085 41107 17088
rect 41049 17079 41107 17085
rect 41138 17076 41144 17088
rect 41196 17076 41202 17128
rect 41230 17076 41236 17128
rect 41288 17116 41294 17128
rect 42076 17116 42104 17146
rect 42444 17116 42472 17147
rect 43070 17144 43076 17156
rect 43128 17144 43134 17196
rect 44100 17193 44128 17224
rect 44085 17187 44143 17193
rect 44085 17153 44097 17187
rect 44131 17184 44143 17187
rect 44358 17184 44364 17196
rect 44131 17156 44364 17184
rect 44131 17153 44143 17156
rect 44085 17147 44143 17153
rect 44358 17144 44364 17156
rect 44416 17144 44422 17196
rect 41288 17088 42104 17116
rect 42168 17088 42472 17116
rect 42797 17119 42855 17125
rect 41288 17076 41294 17088
rect 39991 17020 40816 17048
rect 39991 17017 40003 17020
rect 39945 17011 40003 17017
rect 40862 17008 40868 17060
rect 40920 17048 40926 17060
rect 42168 17048 42196 17088
rect 42797 17085 42809 17119
rect 42843 17116 42855 17119
rect 43162 17116 43168 17128
rect 42843 17088 43168 17116
rect 42843 17085 42855 17088
rect 42797 17079 42855 17085
rect 43162 17076 43168 17088
rect 43220 17116 43226 17128
rect 43530 17116 43536 17128
rect 43220 17088 43536 17116
rect 43220 17076 43226 17088
rect 43530 17076 43536 17088
rect 43588 17076 43594 17128
rect 44560 17116 44588 17280
rect 44818 17212 44824 17264
rect 44876 17252 44882 17264
rect 44876 17224 45416 17252
rect 44876 17212 44882 17224
rect 44726 17144 44732 17196
rect 44784 17184 44790 17196
rect 45388 17193 45416 17224
rect 45281 17187 45339 17193
rect 45281 17184 45293 17187
rect 44784 17156 45293 17184
rect 44784 17144 44790 17156
rect 45281 17153 45293 17156
rect 45327 17153 45339 17187
rect 45281 17147 45339 17153
rect 45373 17187 45431 17193
rect 45373 17153 45385 17187
rect 45419 17153 45431 17187
rect 45373 17147 45431 17153
rect 45005 17119 45063 17125
rect 45005 17116 45017 17119
rect 44560 17088 45017 17116
rect 45005 17085 45017 17088
rect 45051 17116 45063 17119
rect 45557 17119 45615 17125
rect 45557 17116 45569 17119
rect 45051 17088 45569 17116
rect 45051 17085 45063 17088
rect 45005 17079 45063 17085
rect 45557 17085 45569 17088
rect 45603 17085 45615 17119
rect 45557 17079 45615 17085
rect 40920 17020 42196 17048
rect 40920 17008 40926 17020
rect 42242 17008 42248 17060
rect 42300 17048 42306 17060
rect 43346 17048 43352 17060
rect 42300 17020 43352 17048
rect 42300 17008 42306 17020
rect 43346 17008 43352 17020
rect 43404 17048 43410 17060
rect 44910 17048 44916 17060
rect 43404 17020 44916 17048
rect 43404 17008 43410 17020
rect 44910 17008 44916 17020
rect 44968 17008 44974 17060
rect 40218 16980 40224 16992
rect 38580 16952 40224 16980
rect 40218 16940 40224 16952
rect 40276 16940 40282 16992
rect 42334 16940 42340 16992
rect 42392 16980 42398 16992
rect 42521 16983 42579 16989
rect 42521 16980 42533 16983
rect 42392 16952 42533 16980
rect 42392 16940 42398 16952
rect 42521 16949 42533 16952
rect 42567 16949 42579 16983
rect 42521 16943 42579 16949
rect 44082 16940 44088 16992
rect 44140 16980 44146 16992
rect 44177 16983 44235 16989
rect 44177 16980 44189 16983
rect 44140 16952 44189 16980
rect 44140 16940 44146 16952
rect 44177 16949 44189 16952
rect 44223 16949 44235 16983
rect 44177 16943 44235 16949
rect 45094 16940 45100 16992
rect 45152 16980 45158 16992
rect 45465 16983 45523 16989
rect 45465 16980 45477 16983
rect 45152 16952 45477 16980
rect 45152 16940 45158 16952
rect 45465 16949 45477 16952
rect 45511 16949 45523 16983
rect 45465 16943 45523 16949
rect 1104 16890 47104 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 47104 16890
rect 1104 16816 47104 16838
rect 2314 16736 2320 16788
rect 2372 16776 2378 16788
rect 2501 16779 2559 16785
rect 2501 16776 2513 16779
rect 2372 16748 2513 16776
rect 2372 16736 2378 16748
rect 2501 16745 2513 16748
rect 2547 16745 2559 16779
rect 2501 16739 2559 16745
rect 4798 16736 4804 16788
rect 4856 16776 4862 16788
rect 5077 16779 5135 16785
rect 5077 16776 5089 16779
rect 4856 16748 5089 16776
rect 4856 16736 4862 16748
rect 5077 16745 5089 16748
rect 5123 16745 5135 16779
rect 5077 16739 5135 16745
rect 12621 16779 12679 16785
rect 12621 16745 12633 16779
rect 12667 16776 12679 16779
rect 12667 16748 18184 16776
rect 12667 16745 12679 16748
rect 12621 16739 12679 16745
rect 2130 16668 2136 16720
rect 2188 16708 2194 16720
rect 6822 16708 6828 16720
rect 2188 16680 6828 16708
rect 2188 16668 2194 16680
rect 6822 16668 6828 16680
rect 6880 16668 6886 16720
rect 13357 16711 13415 16717
rect 12636 16680 13216 16708
rect 12636 16652 12664 16680
rect 3786 16600 3792 16652
rect 3844 16640 3850 16652
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 3844 16612 4353 16640
rect 3844 16600 3850 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 5350 16600 5356 16652
rect 5408 16640 5414 16652
rect 5721 16643 5779 16649
rect 5408 16612 5580 16640
rect 5408 16600 5414 16612
rect 2685 16575 2743 16581
rect 2685 16541 2697 16575
rect 2731 16541 2743 16575
rect 2685 16535 2743 16541
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16572 4215 16575
rect 4706 16572 4712 16584
rect 4203 16544 4712 16572
rect 4203 16541 4215 16544
rect 4157 16535 4215 16541
rect 2700 16436 2728 16535
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 5442 16532 5448 16584
rect 5500 16532 5506 16584
rect 5552 16572 5580 16612
rect 5721 16609 5733 16643
rect 5767 16640 5779 16643
rect 6270 16640 6276 16652
rect 5767 16612 6276 16640
rect 5767 16609 5779 16612
rect 5721 16603 5779 16609
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 9398 16600 9404 16652
rect 9456 16600 9462 16652
rect 12342 16600 12348 16652
rect 12400 16600 12406 16652
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16640 12495 16643
rect 12618 16640 12624 16652
rect 12483 16612 12624 16640
rect 12483 16609 12495 16612
rect 12437 16603 12495 16609
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 13078 16600 13084 16652
rect 13136 16600 13142 16652
rect 13188 16649 13216 16680
rect 13357 16677 13369 16711
rect 13403 16708 13415 16711
rect 16942 16708 16948 16720
rect 13403 16680 16948 16708
rect 13403 16677 13415 16680
rect 13357 16671 13415 16677
rect 16942 16668 16948 16680
rect 17000 16668 17006 16720
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 15565 16643 15623 16649
rect 15565 16609 15577 16643
rect 15611 16640 15623 16643
rect 15930 16640 15936 16652
rect 15611 16612 15936 16640
rect 15611 16609 15623 16612
rect 15565 16603 15623 16609
rect 15930 16600 15936 16612
rect 15988 16640 15994 16652
rect 16206 16640 16212 16652
rect 15988 16612 16212 16640
rect 15988 16600 15994 16612
rect 16206 16600 16212 16612
rect 16264 16600 16270 16652
rect 16666 16600 16672 16652
rect 16724 16640 16730 16652
rect 18156 16640 18184 16748
rect 18230 16736 18236 16788
rect 18288 16776 18294 16788
rect 18325 16779 18383 16785
rect 18325 16776 18337 16779
rect 18288 16748 18337 16776
rect 18288 16736 18294 16748
rect 18325 16745 18337 16748
rect 18371 16745 18383 16779
rect 18325 16739 18383 16745
rect 20346 16736 20352 16788
rect 20404 16736 20410 16788
rect 20809 16779 20867 16785
rect 20809 16776 20821 16779
rect 20548 16748 20821 16776
rect 20070 16668 20076 16720
rect 20128 16668 20134 16720
rect 20257 16711 20315 16717
rect 20257 16677 20269 16711
rect 20303 16708 20315 16711
rect 20548 16708 20576 16748
rect 20809 16745 20821 16748
rect 20855 16745 20867 16779
rect 20809 16739 20867 16745
rect 23198 16736 23204 16788
rect 23256 16736 23262 16788
rect 23492 16748 24808 16776
rect 23492 16708 23520 16748
rect 20303 16680 20576 16708
rect 20640 16680 23520 16708
rect 20303 16677 20315 16680
rect 20257 16671 20315 16677
rect 16724 16612 16988 16640
rect 18156 16612 20392 16640
rect 16724 16600 16730 16612
rect 16960 16584 16988 16612
rect 8294 16572 8300 16584
rect 5552 16544 8300 16572
rect 8294 16532 8300 16544
rect 8352 16572 8358 16584
rect 9214 16572 9220 16584
rect 8352 16544 9220 16572
rect 8352 16532 8358 16544
rect 9214 16532 9220 16544
rect 9272 16532 9278 16584
rect 14829 16575 14887 16581
rect 14829 16541 14841 16575
rect 14875 16572 14887 16575
rect 14875 16544 14964 16572
rect 14875 16541 14887 16544
rect 14829 16535 14887 16541
rect 9668 16507 9726 16513
rect 9668 16473 9680 16507
rect 9714 16504 9726 16507
rect 10686 16504 10692 16516
rect 9714 16476 10692 16504
rect 9714 16473 9726 16476
rect 9668 16467 9726 16473
rect 10686 16464 10692 16476
rect 10744 16464 10750 16516
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 2700 16408 3801 16436
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 4246 16396 4252 16448
rect 4304 16436 4310 16448
rect 5537 16439 5595 16445
rect 5537 16436 5549 16439
rect 4304 16408 5549 16436
rect 4304 16396 4310 16408
rect 5537 16405 5549 16408
rect 5583 16405 5595 16439
rect 5537 16399 5595 16405
rect 10134 16396 10140 16448
rect 10192 16436 10198 16448
rect 10781 16439 10839 16445
rect 10781 16436 10793 16439
rect 10192 16408 10793 16436
rect 10192 16396 10198 16408
rect 10781 16405 10793 16408
rect 10827 16405 10839 16439
rect 10781 16399 10839 16405
rect 11977 16439 12035 16445
rect 11977 16405 11989 16439
rect 12023 16436 12035 16439
rect 12066 16436 12072 16448
rect 12023 16408 12072 16436
rect 12023 16405 12035 16408
rect 11977 16399 12035 16405
rect 12066 16396 12072 16408
rect 12124 16436 12130 16448
rect 12434 16436 12440 16448
rect 12124 16408 12440 16436
rect 12124 16396 12130 16408
rect 12434 16396 12440 16408
rect 12492 16436 12498 16448
rect 12713 16439 12771 16445
rect 12713 16436 12725 16439
rect 12492 16408 12725 16436
rect 12492 16396 12498 16408
rect 12713 16405 12725 16408
rect 12759 16405 12771 16439
rect 12713 16399 12771 16405
rect 13630 16396 13636 16448
rect 13688 16436 13694 16448
rect 14090 16436 14096 16448
rect 13688 16408 14096 16436
rect 13688 16396 13694 16408
rect 14090 16396 14096 16408
rect 14148 16396 14154 16448
rect 14645 16439 14703 16445
rect 14645 16405 14657 16439
rect 14691 16436 14703 16439
rect 14734 16436 14740 16448
rect 14691 16408 14740 16436
rect 14691 16405 14703 16408
rect 14645 16399 14703 16405
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 14936 16445 14964 16544
rect 16942 16532 16948 16584
rect 17000 16532 17006 16584
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16572 19855 16575
rect 20254 16572 20260 16584
rect 19843 16544 20260 16572
rect 19843 16541 19855 16544
rect 19797 16535 19855 16541
rect 20254 16532 20260 16544
rect 20312 16532 20318 16584
rect 17218 16513 17224 16516
rect 17212 16467 17224 16513
rect 17218 16464 17224 16467
rect 17276 16464 17282 16516
rect 20364 16504 20392 16612
rect 20530 16532 20536 16584
rect 20588 16532 20594 16584
rect 20640 16581 20668 16680
rect 23566 16668 23572 16720
rect 23624 16708 23630 16720
rect 24780 16708 24808 16748
rect 24854 16736 24860 16788
rect 24912 16736 24918 16788
rect 26421 16779 26479 16785
rect 26421 16745 26433 16779
rect 26467 16776 26479 16779
rect 26602 16776 26608 16788
rect 26467 16748 26608 16776
rect 26467 16745 26479 16748
rect 26421 16739 26479 16745
rect 26602 16736 26608 16748
rect 26660 16736 26666 16788
rect 32122 16736 32128 16788
rect 32180 16736 32186 16788
rect 34333 16779 34391 16785
rect 34333 16745 34345 16779
rect 34379 16776 34391 16779
rect 34422 16776 34428 16788
rect 34379 16748 34428 16776
rect 34379 16745 34391 16748
rect 34333 16739 34391 16745
rect 34422 16736 34428 16748
rect 34480 16736 34486 16788
rect 39850 16736 39856 16788
rect 39908 16776 39914 16788
rect 39908 16748 41414 16776
rect 39908 16736 39914 16748
rect 30650 16708 30656 16720
rect 23624 16680 23704 16708
rect 24780 16680 30656 16708
rect 23624 16668 23630 16680
rect 23676 16649 23704 16680
rect 30650 16668 30656 16680
rect 30708 16668 30714 16720
rect 40678 16708 40684 16720
rect 40052 16680 40684 16708
rect 23661 16643 23719 16649
rect 23661 16609 23673 16643
rect 23707 16609 23719 16643
rect 23661 16603 23719 16609
rect 23842 16600 23848 16652
rect 23900 16600 23906 16652
rect 26878 16600 26884 16652
rect 26936 16600 26942 16652
rect 27065 16643 27123 16649
rect 27065 16609 27077 16643
rect 27111 16640 27123 16643
rect 28442 16640 28448 16652
rect 27111 16612 28448 16640
rect 27111 16609 27123 16612
rect 27065 16603 27123 16609
rect 28442 16600 28448 16612
rect 28500 16600 28506 16652
rect 32953 16643 33011 16649
rect 32953 16640 32965 16643
rect 32784 16612 32965 16640
rect 20625 16575 20683 16581
rect 20625 16541 20637 16575
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 20901 16575 20959 16581
rect 20901 16541 20913 16575
rect 20947 16572 20959 16575
rect 20990 16572 20996 16584
rect 20947 16544 20996 16572
rect 20947 16541 20959 16544
rect 20901 16535 20959 16541
rect 20990 16532 20996 16544
rect 21048 16532 21054 16584
rect 23569 16575 23627 16581
rect 23569 16541 23581 16575
rect 23615 16572 23627 16575
rect 24026 16572 24032 16584
rect 23615 16544 24032 16572
rect 23615 16541 23627 16544
rect 23569 16535 23627 16541
rect 24026 16532 24032 16544
rect 24084 16532 24090 16584
rect 25041 16575 25099 16581
rect 25041 16541 25053 16575
rect 25087 16572 25099 16575
rect 25958 16572 25964 16584
rect 25087 16544 25964 16572
rect 25087 16541 25099 16544
rect 25041 16535 25099 16541
rect 25958 16532 25964 16544
rect 26016 16532 26022 16584
rect 26510 16532 26516 16584
rect 26568 16572 26574 16584
rect 26789 16575 26847 16581
rect 26789 16572 26801 16575
rect 26568 16544 26801 16572
rect 26568 16532 26574 16544
rect 26789 16541 26801 16544
rect 26835 16541 26847 16575
rect 26789 16535 26847 16541
rect 29086 16532 29092 16584
rect 29144 16572 29150 16584
rect 29638 16572 29644 16584
rect 29144 16544 29644 16572
rect 29144 16532 29150 16544
rect 29638 16532 29644 16544
rect 29696 16572 29702 16584
rect 30282 16572 30288 16584
rect 29696 16544 30288 16572
rect 29696 16532 29702 16544
rect 30282 16532 30288 16544
rect 30340 16532 30346 16584
rect 30745 16575 30803 16581
rect 30745 16541 30757 16575
rect 30791 16572 30803 16575
rect 31570 16572 31576 16584
rect 30791 16544 31576 16572
rect 30791 16541 30803 16544
rect 30745 16535 30803 16541
rect 31570 16532 31576 16544
rect 31628 16572 31634 16584
rect 32784 16572 32812 16612
rect 32953 16609 32965 16612
rect 32999 16609 33011 16643
rect 34701 16643 34759 16649
rect 34701 16640 34713 16643
rect 32953 16603 33011 16609
rect 34348 16612 34713 16640
rect 31628 16544 32812 16572
rect 31628 16532 31634 16544
rect 32858 16532 32864 16584
rect 32916 16532 32922 16584
rect 32968 16572 32996 16603
rect 34348 16584 34376 16612
rect 34701 16609 34713 16612
rect 34747 16609 34759 16643
rect 34701 16603 34759 16609
rect 38010 16600 38016 16652
rect 38068 16600 38074 16652
rect 34330 16572 34336 16584
rect 32968 16544 34336 16572
rect 34330 16532 34336 16544
rect 34388 16532 34394 16584
rect 34606 16532 34612 16584
rect 34664 16572 34670 16584
rect 35526 16572 35532 16584
rect 34664 16544 35532 16572
rect 34664 16532 34670 16544
rect 35526 16532 35532 16544
rect 35584 16532 35590 16584
rect 37093 16575 37151 16581
rect 37093 16541 37105 16575
rect 37139 16541 37151 16575
rect 37093 16535 37151 16541
rect 21266 16504 21272 16516
rect 20364 16476 21272 16504
rect 21266 16464 21272 16476
rect 21324 16464 21330 16516
rect 21818 16464 21824 16516
rect 21876 16504 21882 16516
rect 23934 16504 23940 16516
rect 21876 16476 23940 16504
rect 21876 16464 21882 16476
rect 23934 16464 23940 16476
rect 23992 16464 23998 16516
rect 25130 16504 25136 16516
rect 24228 16476 25136 16504
rect 14921 16439 14979 16445
rect 14921 16405 14933 16439
rect 14967 16405 14979 16439
rect 14921 16399 14979 16405
rect 15286 16396 15292 16448
rect 15344 16396 15350 16448
rect 15381 16439 15439 16445
rect 15381 16405 15393 16439
rect 15427 16436 15439 16439
rect 15838 16436 15844 16448
rect 15427 16408 15844 16436
rect 15427 16405 15439 16408
rect 15381 16399 15439 16405
rect 15838 16396 15844 16408
rect 15896 16396 15902 16448
rect 17954 16396 17960 16448
rect 18012 16436 18018 16448
rect 19150 16436 19156 16448
rect 18012 16408 19156 16436
rect 18012 16396 18018 16408
rect 19150 16396 19156 16408
rect 19208 16396 19214 16448
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 19794 16436 19800 16448
rect 19392 16408 19800 16436
rect 19392 16396 19398 16408
rect 19794 16396 19800 16408
rect 19852 16396 19858 16448
rect 21174 16396 21180 16448
rect 21232 16436 21238 16448
rect 24228 16436 24256 16476
rect 25130 16464 25136 16476
rect 25188 16464 25194 16516
rect 31012 16507 31070 16513
rect 31012 16473 31024 16507
rect 31058 16504 31070 16507
rect 31110 16504 31116 16516
rect 31058 16476 31116 16504
rect 31058 16473 31070 16476
rect 31012 16467 31070 16473
rect 31110 16464 31116 16476
rect 31168 16464 31174 16516
rect 33198 16507 33256 16513
rect 33198 16504 33210 16507
rect 32692 16476 33210 16504
rect 21232 16408 24256 16436
rect 21232 16396 21238 16408
rect 24302 16396 24308 16448
rect 24360 16436 24366 16448
rect 27062 16436 27068 16448
rect 24360 16408 27068 16436
rect 24360 16396 24366 16408
rect 27062 16396 27068 16408
rect 27120 16396 27126 16448
rect 32692 16445 32720 16476
rect 33198 16473 33210 16476
rect 33244 16473 33256 16507
rect 33198 16467 33256 16473
rect 34054 16464 34060 16516
rect 34112 16504 34118 16516
rect 34946 16507 35004 16513
rect 34946 16504 34958 16507
rect 34112 16476 34958 16504
rect 34112 16464 34118 16476
rect 34946 16473 34958 16476
rect 34992 16473 35004 16507
rect 37108 16504 37136 16535
rect 37274 16532 37280 16584
rect 37332 16532 37338 16584
rect 38286 16532 38292 16584
rect 38344 16532 38350 16584
rect 38470 16532 38476 16584
rect 38528 16532 38534 16584
rect 38838 16532 38844 16584
rect 38896 16572 38902 16584
rect 39942 16572 39948 16584
rect 38896 16544 39948 16572
rect 38896 16532 38902 16544
rect 39942 16532 39948 16544
rect 40000 16532 40006 16584
rect 40052 16581 40080 16680
rect 40678 16668 40684 16680
rect 40736 16668 40742 16720
rect 40773 16711 40831 16717
rect 40773 16677 40785 16711
rect 40819 16708 40831 16711
rect 40862 16708 40868 16720
rect 40819 16680 40868 16708
rect 40819 16677 40831 16680
rect 40773 16671 40831 16677
rect 40788 16640 40816 16671
rect 40862 16668 40868 16680
rect 40920 16668 40926 16720
rect 41386 16708 41414 16748
rect 42058 16736 42064 16788
rect 42116 16776 42122 16788
rect 42702 16776 42708 16788
rect 42116 16748 42708 16776
rect 42116 16736 42122 16748
rect 42702 16736 42708 16748
rect 42760 16736 42766 16788
rect 42794 16736 42800 16788
rect 42852 16776 42858 16788
rect 43441 16779 43499 16785
rect 43441 16776 43453 16779
rect 42852 16748 43453 16776
rect 42852 16736 42858 16748
rect 43441 16745 43453 16748
rect 43487 16745 43499 16779
rect 43441 16739 43499 16745
rect 44726 16736 44732 16788
rect 44784 16736 44790 16788
rect 44818 16736 44824 16788
rect 44876 16776 44882 16788
rect 45005 16779 45063 16785
rect 45005 16776 45017 16779
rect 44876 16748 45017 16776
rect 44876 16736 44882 16748
rect 45005 16745 45017 16748
rect 45051 16745 45063 16779
rect 45005 16739 45063 16745
rect 41969 16711 42027 16717
rect 41386 16680 41920 16708
rect 40420 16612 40816 16640
rect 40420 16581 40448 16612
rect 41046 16600 41052 16652
rect 41104 16640 41110 16652
rect 41104 16612 41368 16640
rect 41104 16600 41110 16612
rect 40037 16575 40095 16581
rect 40037 16541 40049 16575
rect 40083 16541 40095 16575
rect 40037 16535 40095 16541
rect 40221 16575 40279 16581
rect 40221 16541 40233 16575
rect 40267 16541 40279 16575
rect 40221 16535 40279 16541
rect 40405 16575 40463 16581
rect 40405 16541 40417 16575
rect 40451 16541 40463 16575
rect 40405 16535 40463 16541
rect 40681 16575 40739 16581
rect 40681 16541 40693 16575
rect 40727 16541 40739 16575
rect 40681 16535 40739 16541
rect 37918 16504 37924 16516
rect 37108 16476 37924 16504
rect 34946 16467 35004 16473
rect 37918 16464 37924 16476
rect 37976 16464 37982 16516
rect 32677 16439 32735 16445
rect 32677 16405 32689 16439
rect 32723 16405 32735 16439
rect 32677 16399 32735 16405
rect 34238 16396 34244 16448
rect 34296 16436 34302 16448
rect 34422 16436 34428 16448
rect 34296 16408 34428 16436
rect 34296 16396 34302 16408
rect 34422 16396 34428 16408
rect 34480 16436 34486 16448
rect 36081 16439 36139 16445
rect 36081 16436 36093 16439
rect 34480 16408 36093 16436
rect 34480 16396 34486 16408
rect 36081 16405 36093 16408
rect 36127 16405 36139 16439
rect 36081 16399 36139 16405
rect 38930 16396 38936 16448
rect 38988 16396 38994 16448
rect 40034 16396 40040 16448
rect 40092 16436 40098 16448
rect 40236 16436 40264 16535
rect 40310 16464 40316 16516
rect 40368 16464 40374 16516
rect 40696 16504 40724 16535
rect 40770 16532 40776 16584
rect 40828 16572 40834 16584
rect 40865 16575 40923 16581
rect 40865 16572 40877 16575
rect 40828 16544 40877 16572
rect 40828 16532 40834 16544
rect 40865 16541 40877 16544
rect 40911 16541 40923 16575
rect 40865 16535 40923 16541
rect 40954 16532 40960 16584
rect 41012 16532 41018 16584
rect 41230 16532 41236 16584
rect 41288 16532 41294 16584
rect 41340 16581 41368 16612
rect 41325 16575 41383 16581
rect 41325 16541 41337 16575
rect 41371 16541 41383 16575
rect 41892 16572 41920 16680
rect 41969 16677 41981 16711
rect 42015 16708 42027 16711
rect 42015 16680 43576 16708
rect 42015 16677 42027 16680
rect 41969 16671 42027 16677
rect 42610 16600 42616 16652
rect 42668 16600 42674 16652
rect 41969 16575 42027 16581
rect 41969 16572 41981 16575
rect 41892 16544 41981 16572
rect 41325 16535 41383 16541
rect 41969 16541 41981 16544
rect 42015 16541 42027 16575
rect 41969 16535 42027 16541
rect 41509 16507 41567 16513
rect 41509 16504 41521 16507
rect 40420 16476 41521 16504
rect 40420 16436 40448 16476
rect 41509 16473 41521 16476
rect 41555 16473 41567 16507
rect 41509 16467 41567 16473
rect 40092 16408 40448 16436
rect 40497 16439 40555 16445
rect 40092 16396 40098 16408
rect 40497 16405 40509 16439
rect 40543 16436 40555 16439
rect 40770 16436 40776 16448
rect 40543 16408 40776 16436
rect 40543 16405 40555 16408
rect 40497 16399 40555 16405
rect 40770 16396 40776 16408
rect 40828 16396 40834 16448
rect 40954 16396 40960 16448
rect 41012 16436 41018 16448
rect 41322 16436 41328 16448
rect 41012 16408 41328 16436
rect 41012 16396 41018 16408
rect 41322 16396 41328 16408
rect 41380 16436 41386 16448
rect 41598 16436 41604 16448
rect 41380 16408 41604 16436
rect 41380 16396 41386 16408
rect 41598 16396 41604 16408
rect 41656 16396 41662 16448
rect 41984 16436 42012 16535
rect 42150 16532 42156 16584
rect 42208 16532 42214 16584
rect 42334 16532 42340 16584
rect 42392 16532 42398 16584
rect 42518 16532 42524 16584
rect 42576 16532 42582 16584
rect 42702 16532 42708 16584
rect 42760 16572 42766 16584
rect 42996 16581 43024 16680
rect 43346 16600 43352 16652
rect 43404 16600 43410 16652
rect 42797 16575 42855 16581
rect 42797 16572 42809 16575
rect 42760 16544 42809 16572
rect 42760 16532 42766 16544
rect 42797 16541 42809 16544
rect 42843 16541 42855 16575
rect 42797 16535 42855 16541
rect 42981 16575 43039 16581
rect 42981 16541 42993 16575
rect 43027 16541 43039 16575
rect 42981 16535 43039 16541
rect 43070 16532 43076 16584
rect 43128 16572 43134 16584
rect 43165 16575 43223 16581
rect 43165 16572 43177 16575
rect 43128 16544 43177 16572
rect 43128 16532 43134 16544
rect 43165 16541 43177 16544
rect 43211 16541 43223 16575
rect 43548 16572 43576 16680
rect 44082 16668 44088 16720
rect 44140 16708 44146 16720
rect 44545 16711 44603 16717
rect 44545 16708 44557 16711
rect 44140 16680 44557 16708
rect 44140 16668 44146 16680
rect 44545 16677 44557 16680
rect 44591 16677 44603 16711
rect 44545 16671 44603 16677
rect 44744 16640 44772 16736
rect 44910 16668 44916 16720
rect 44968 16708 44974 16720
rect 44968 16680 45968 16708
rect 44968 16668 44974 16680
rect 45097 16643 45155 16649
rect 45097 16640 45109 16643
rect 44744 16612 45109 16640
rect 45097 16609 45109 16612
rect 45143 16609 45155 16643
rect 45097 16603 45155 16609
rect 45370 16600 45376 16652
rect 45428 16640 45434 16652
rect 45940 16649 45968 16680
rect 45649 16643 45707 16649
rect 45649 16640 45661 16643
rect 45428 16612 45661 16640
rect 45428 16600 45434 16612
rect 45649 16609 45661 16612
rect 45695 16609 45707 16643
rect 45649 16603 45707 16609
rect 45925 16643 45983 16649
rect 45925 16609 45937 16643
rect 45971 16609 45983 16643
rect 45925 16603 45983 16609
rect 43625 16575 43683 16581
rect 43625 16572 43637 16575
rect 43548 16544 43637 16572
rect 43165 16535 43223 16541
rect 43625 16541 43637 16544
rect 43671 16541 43683 16575
rect 43625 16535 43683 16541
rect 43180 16504 43208 16535
rect 43806 16532 43812 16584
rect 43864 16532 43870 16584
rect 45002 16532 45008 16584
rect 45060 16532 45066 16584
rect 43180 16476 43484 16504
rect 42702 16436 42708 16448
rect 41984 16408 42708 16436
rect 42702 16396 42708 16408
rect 42760 16396 42766 16448
rect 43254 16396 43260 16448
rect 43312 16396 43318 16448
rect 43456 16436 43484 16476
rect 43530 16464 43536 16516
rect 43588 16464 43594 16516
rect 44269 16507 44327 16513
rect 44269 16473 44281 16507
rect 44315 16504 44327 16507
rect 44358 16504 44364 16516
rect 44315 16476 44364 16504
rect 44315 16473 44327 16476
rect 44269 16467 44327 16473
rect 44358 16464 44364 16476
rect 44416 16464 44422 16516
rect 45738 16464 45744 16516
rect 45796 16464 45802 16516
rect 43717 16439 43775 16445
rect 43717 16436 43729 16439
rect 43456 16408 43729 16436
rect 43717 16405 43729 16408
rect 43763 16436 43775 16439
rect 44726 16436 44732 16448
rect 43763 16408 44732 16436
rect 43763 16405 43775 16408
rect 43717 16399 43775 16405
rect 44726 16396 44732 16408
rect 44784 16396 44790 16448
rect 44818 16396 44824 16448
rect 44876 16436 44882 16448
rect 45373 16439 45431 16445
rect 45373 16436 45385 16439
rect 44876 16408 45385 16436
rect 44876 16396 44882 16408
rect 45373 16405 45385 16408
rect 45419 16405 45431 16439
rect 45373 16399 45431 16405
rect 1104 16346 47104 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 47104 16346
rect 1104 16272 47104 16294
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 4157 16235 4215 16241
rect 4157 16232 4169 16235
rect 3743 16204 4169 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 4157 16201 4169 16204
rect 4203 16232 4215 16235
rect 5258 16232 5264 16244
rect 4203 16204 5264 16232
rect 4203 16201 4215 16204
rect 4157 16195 4215 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 7282 16232 7288 16244
rect 6972 16204 7288 16232
rect 6972 16192 6978 16204
rect 7282 16192 7288 16204
rect 7340 16192 7346 16244
rect 9490 16192 9496 16244
rect 9548 16232 9554 16244
rect 10042 16232 10048 16244
rect 9548 16204 10048 16232
rect 9548 16192 9554 16204
rect 10042 16192 10048 16204
rect 10100 16192 10106 16244
rect 10686 16192 10692 16244
rect 10744 16192 10750 16244
rect 11793 16235 11851 16241
rect 11793 16201 11805 16235
rect 11839 16201 11851 16235
rect 13541 16235 13599 16241
rect 13541 16232 13553 16235
rect 11793 16195 11851 16201
rect 12406 16204 13553 16232
rect 7009 16167 7067 16173
rect 7009 16133 7021 16167
rect 7055 16164 7067 16167
rect 7098 16164 7104 16176
rect 7055 16136 7104 16164
rect 7055 16133 7067 16136
rect 7009 16127 7067 16133
rect 7098 16124 7104 16136
rect 7156 16124 7162 16176
rect 10597 16167 10655 16173
rect 10597 16133 10609 16167
rect 10643 16164 10655 16167
rect 11054 16164 11060 16176
rect 10643 16136 11060 16164
rect 10643 16133 10655 16136
rect 10597 16127 10655 16133
rect 11054 16124 11060 16136
rect 11112 16124 11118 16176
rect 11808 16164 11836 16195
rect 12314 16167 12372 16173
rect 12314 16164 12326 16167
rect 11808 16136 12326 16164
rect 12314 16133 12326 16136
rect 12360 16133 12372 16167
rect 12314 16127 12372 16133
rect 2317 16099 2375 16105
rect 2317 16065 2329 16099
rect 2363 16096 2375 16099
rect 2406 16096 2412 16108
rect 2363 16068 2412 16096
rect 2363 16065 2375 16068
rect 2317 16059 2375 16065
rect 2406 16056 2412 16068
rect 2464 16056 2470 16108
rect 2590 16105 2596 16108
rect 2584 16059 2596 16105
rect 2590 16056 2596 16059
rect 2648 16056 2654 16108
rect 4246 16056 4252 16108
rect 4304 16096 4310 16108
rect 4706 16096 4712 16108
rect 4304 16068 4712 16096
rect 4304 16056 4310 16068
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 7116 16096 7144 16124
rect 7116 16068 9076 16096
rect 3970 15988 3976 16040
rect 4028 16028 4034 16040
rect 4433 16031 4491 16037
rect 4433 16028 4445 16031
rect 4028 16000 4445 16028
rect 4028 15988 4034 16000
rect 4433 15997 4445 16000
rect 4479 16028 4491 16031
rect 6914 16028 6920 16040
rect 4479 16000 6920 16028
rect 4479 15997 4491 16000
rect 4433 15991 4491 15997
rect 6914 15988 6920 16000
rect 6972 15988 6978 16040
rect 7101 16031 7159 16037
rect 7101 15997 7113 16031
rect 7147 15997 7159 16031
rect 7101 15991 7159 15997
rect 5718 15920 5724 15972
rect 5776 15960 5782 15972
rect 6641 15963 6699 15969
rect 6641 15960 6653 15963
rect 5776 15932 6653 15960
rect 5776 15920 5782 15932
rect 6641 15929 6653 15932
rect 6687 15929 6699 15963
rect 7116 15960 7144 15991
rect 7190 15988 7196 16040
rect 7248 15988 7254 16040
rect 8754 15988 8760 16040
rect 8812 15988 8818 16040
rect 8938 15988 8944 16040
rect 8996 15988 9002 16040
rect 9048 16028 9076 16068
rect 9950 16056 9956 16108
rect 10008 16056 10014 16108
rect 10686 16056 10692 16108
rect 10744 16096 10750 16108
rect 10873 16099 10931 16105
rect 10873 16096 10885 16099
rect 10744 16068 10885 16096
rect 10744 16056 10750 16068
rect 10873 16065 10885 16068
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16096 12035 16099
rect 12406 16096 12434 16204
rect 13541 16201 13553 16204
rect 13587 16201 13599 16235
rect 13541 16195 13599 16201
rect 13909 16235 13967 16241
rect 13909 16201 13921 16235
rect 13955 16232 13967 16235
rect 16666 16232 16672 16244
rect 13955 16204 16672 16232
rect 13955 16201 13967 16204
rect 13909 16195 13967 16201
rect 12023 16068 12434 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 9674 16028 9680 16040
rect 9048 16000 9680 16028
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 9766 15988 9772 16040
rect 9824 16037 9830 16040
rect 9824 16031 9852 16037
rect 9840 15997 9852 16031
rect 9824 15991 9852 15997
rect 9824 15988 9830 15991
rect 12066 15988 12072 16040
rect 12124 15988 12130 16040
rect 7116 15932 7236 15960
rect 6641 15923 6699 15929
rect 7208 15904 7236 15932
rect 9214 15920 9220 15972
rect 9272 15960 9278 15972
rect 9401 15963 9459 15969
rect 9401 15960 9413 15963
rect 9272 15932 9413 15960
rect 9272 15920 9278 15932
rect 9401 15929 9413 15932
rect 9447 15929 9459 15963
rect 9401 15923 9459 15929
rect 13449 15963 13507 15969
rect 13449 15929 13461 15963
rect 13495 15960 13507 15963
rect 13924 15960 13952 16195
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 17218 16192 17224 16244
rect 17276 16192 17282 16244
rect 17497 16235 17555 16241
rect 17497 16201 17509 16235
rect 17543 16201 17555 16235
rect 17957 16235 18015 16241
rect 17957 16232 17969 16235
rect 17497 16195 17555 16201
rect 17604 16204 17969 16232
rect 14001 16167 14059 16173
rect 14001 16133 14013 16167
rect 14047 16164 14059 16167
rect 15838 16164 15844 16176
rect 14047 16136 15844 16164
rect 14047 16133 14059 16136
rect 14001 16127 14059 16133
rect 13495 15932 13952 15960
rect 13495 15929 13507 15932
rect 13449 15923 13507 15929
rect 3786 15852 3792 15904
rect 3844 15852 3850 15904
rect 6362 15852 6368 15904
rect 6420 15852 6426 15904
rect 7190 15852 7196 15904
rect 7248 15852 7254 15904
rect 10318 15852 10324 15904
rect 10376 15892 10382 15904
rect 14016 15892 14044 16127
rect 15838 16124 15844 16136
rect 15896 16124 15902 16176
rect 14458 16056 14464 16108
rect 14516 16056 14522 16108
rect 14734 16105 14740 16108
rect 14728 16096 14740 16105
rect 14695 16068 14740 16096
rect 14728 16059 14740 16068
rect 14734 16056 14740 16059
rect 14792 16056 14798 16108
rect 15286 16056 15292 16108
rect 15344 16096 15350 16108
rect 16209 16099 16267 16105
rect 15344 16068 15884 16096
rect 15344 16056 15350 16068
rect 14090 15988 14096 16040
rect 14148 15988 14154 16040
rect 10376 15864 14044 15892
rect 14476 15892 14504 16056
rect 15856 15969 15884 16068
rect 16209 16065 16221 16099
rect 16255 16096 16267 16099
rect 17310 16096 17316 16108
rect 16255 16068 17316 16096
rect 16255 16065 16267 16068
rect 16209 16059 16267 16065
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16096 17463 16099
rect 17512 16096 17540 16195
rect 17451 16068 17540 16096
rect 17451 16065 17463 16068
rect 17405 16059 17463 16065
rect 17126 15988 17132 16040
rect 17184 16028 17190 16040
rect 17604 16028 17632 16204
rect 17957 16201 17969 16204
rect 18003 16232 18015 16235
rect 20990 16232 20996 16244
rect 18003 16204 20996 16232
rect 18003 16201 18015 16204
rect 17957 16195 18015 16201
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 21174 16192 21180 16244
rect 21232 16192 21238 16244
rect 21266 16192 21272 16244
rect 21324 16232 21330 16244
rect 21324 16204 23612 16232
rect 21324 16192 21330 16204
rect 21082 16124 21088 16176
rect 21140 16164 21146 16176
rect 23477 16167 23535 16173
rect 23477 16164 23489 16167
rect 21140 16136 22094 16164
rect 21140 16124 21146 16136
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16096 17923 16099
rect 18230 16096 18236 16108
rect 17911 16068 18236 16096
rect 17911 16065 17923 16068
rect 17865 16059 17923 16065
rect 18230 16056 18236 16068
rect 18288 16096 18294 16108
rect 18509 16099 18567 16105
rect 18509 16096 18521 16099
rect 18288 16068 18521 16096
rect 18288 16056 18294 16068
rect 18509 16065 18521 16068
rect 18555 16065 18567 16099
rect 18509 16059 18567 16065
rect 19334 16056 19340 16108
rect 19392 16105 19398 16108
rect 19392 16099 19420 16105
rect 19408 16065 19420 16099
rect 19392 16059 19420 16065
rect 19392 16056 19398 16059
rect 20162 16056 20168 16108
rect 20220 16096 20226 16108
rect 21266 16096 21272 16108
rect 20220 16068 21272 16096
rect 20220 16056 20226 16068
rect 21266 16056 21272 16068
rect 21324 16056 21330 16108
rect 21358 16056 21364 16108
rect 21416 16056 21422 16108
rect 21450 16056 21456 16108
rect 21508 16096 21514 16108
rect 21545 16099 21603 16105
rect 21545 16096 21557 16099
rect 21508 16068 21557 16096
rect 21508 16056 21514 16068
rect 21545 16065 21557 16068
rect 21591 16065 21603 16099
rect 21545 16059 21603 16065
rect 21637 16099 21695 16105
rect 21637 16065 21649 16099
rect 21683 16096 21695 16099
rect 21818 16096 21824 16108
rect 21683 16068 21824 16096
rect 21683 16065 21695 16068
rect 21637 16059 21695 16065
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 22066 16096 22094 16136
rect 22756 16136 23489 16164
rect 22373 16099 22431 16105
rect 22373 16096 22385 16099
rect 22066 16068 22385 16096
rect 22373 16065 22385 16068
rect 22419 16065 22431 16099
rect 22373 16059 22431 16065
rect 22462 16056 22468 16108
rect 22520 16056 22526 16108
rect 22756 16105 22784 16136
rect 23477 16133 23489 16136
rect 23523 16133 23535 16167
rect 23477 16127 23535 16133
rect 22741 16099 22799 16105
rect 22741 16065 22753 16099
rect 22787 16065 22799 16099
rect 22741 16059 22799 16065
rect 23017 16099 23075 16105
rect 23017 16065 23029 16099
rect 23063 16065 23075 16099
rect 23017 16059 23075 16065
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16065 23167 16099
rect 23109 16059 23167 16065
rect 23385 16099 23443 16105
rect 23385 16065 23397 16099
rect 23431 16096 23443 16099
rect 23584 16096 23612 16204
rect 26694 16192 26700 16244
rect 26752 16232 26758 16244
rect 28077 16235 28135 16241
rect 28077 16232 28089 16235
rect 26752 16204 28089 16232
rect 26752 16192 26758 16204
rect 28077 16201 28089 16204
rect 28123 16232 28135 16235
rect 29178 16232 29184 16244
rect 28123 16204 29184 16232
rect 28123 16201 28135 16204
rect 28077 16195 28135 16201
rect 29178 16192 29184 16204
rect 29236 16192 29242 16244
rect 31110 16192 31116 16244
rect 31168 16192 31174 16244
rect 33505 16235 33563 16241
rect 33505 16201 33517 16235
rect 33551 16201 33563 16235
rect 33505 16195 33563 16201
rect 23845 16167 23903 16173
rect 23845 16133 23857 16167
rect 23891 16164 23903 16167
rect 24210 16164 24216 16176
rect 23891 16136 24216 16164
rect 23891 16133 23903 16136
rect 23845 16127 23903 16133
rect 24210 16124 24216 16136
rect 24268 16124 24274 16176
rect 28902 16164 28908 16176
rect 24964 16136 28908 16164
rect 23431 16068 23612 16096
rect 23431 16065 23443 16068
rect 23385 16059 23443 16065
rect 17184 16000 17632 16028
rect 17184 15988 17190 16000
rect 17770 15988 17776 16040
rect 17828 16028 17834 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17828 16000 18061 16028
rect 17828 15988 17834 16000
rect 18049 15997 18061 16000
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 18322 15988 18328 16040
rect 18380 15988 18386 16040
rect 19245 16031 19303 16037
rect 19245 16028 19257 16031
rect 18800 16000 19257 16028
rect 18800 15972 18828 16000
rect 19245 15997 19257 16000
rect 19291 15997 19303 16031
rect 19245 15991 19303 15997
rect 19521 16031 19579 16037
rect 19521 15997 19533 16031
rect 19567 16028 19579 16031
rect 19567 16000 20116 16028
rect 19567 15997 19579 16000
rect 19521 15991 19579 15997
rect 15841 15963 15899 15969
rect 15841 15929 15853 15963
rect 15887 15960 15899 15963
rect 17954 15960 17960 15972
rect 15887 15932 17960 15960
rect 15887 15929 15899 15932
rect 15841 15923 15899 15929
rect 17954 15920 17960 15932
rect 18012 15920 18018 15972
rect 18782 15920 18788 15972
rect 18840 15920 18846 15972
rect 18969 15963 19027 15969
rect 18969 15929 18981 15963
rect 19015 15960 19027 15963
rect 19015 15932 19104 15960
rect 19015 15929 19027 15932
rect 18969 15923 19027 15929
rect 14642 15892 14648 15904
rect 14476 15864 14648 15892
rect 10376 15852 10382 15864
rect 14642 15852 14648 15864
rect 14700 15852 14706 15904
rect 16298 15852 16304 15904
rect 16356 15852 16362 15904
rect 16666 15852 16672 15904
rect 16724 15892 16730 15904
rect 18800 15892 18828 15920
rect 16724 15864 18828 15892
rect 19076 15892 19104 15932
rect 19978 15892 19984 15904
rect 19076 15864 19984 15892
rect 16724 15852 16730 15864
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 20088 15892 20116 16000
rect 20530 15988 20536 16040
rect 20588 16028 20594 16040
rect 23032 16028 23060 16059
rect 20588 16000 23060 16028
rect 23124 16028 23152 16059
rect 23658 16056 23664 16108
rect 23716 16056 23722 16108
rect 23934 16056 23940 16108
rect 23992 16056 23998 16108
rect 24854 16056 24860 16108
rect 24912 16056 24918 16108
rect 24964 16105 24992 16136
rect 28902 16124 28908 16136
rect 28960 16124 28966 16176
rect 29086 16124 29092 16176
rect 29144 16164 29150 16176
rect 31938 16164 31944 16176
rect 29144 16136 31944 16164
rect 29144 16124 29150 16136
rect 31938 16124 31944 16136
rect 31996 16164 32002 16176
rect 33520 16164 33548 16195
rect 34054 16192 34060 16244
rect 34112 16192 34118 16244
rect 35342 16192 35348 16244
rect 35400 16232 35406 16244
rect 35713 16235 35771 16241
rect 35713 16232 35725 16235
rect 35400 16204 35725 16232
rect 35400 16192 35406 16204
rect 35713 16201 35725 16204
rect 35759 16201 35771 16235
rect 35713 16195 35771 16201
rect 38286 16192 38292 16244
rect 38344 16232 38350 16244
rect 40037 16235 40095 16241
rect 40037 16232 40049 16235
rect 38344 16204 40049 16232
rect 38344 16192 38350 16204
rect 40037 16201 40049 16204
rect 40083 16201 40095 16235
rect 40037 16195 40095 16201
rect 42889 16235 42947 16241
rect 42889 16201 42901 16235
rect 42935 16232 42947 16235
rect 43806 16232 43812 16244
rect 42935 16204 43812 16232
rect 42935 16201 42947 16204
rect 42889 16195 42947 16201
rect 43806 16192 43812 16204
rect 43864 16192 43870 16244
rect 45370 16192 45376 16244
rect 45428 16192 45434 16244
rect 34606 16173 34612 16176
rect 34600 16164 34612 16173
rect 31996 16136 33548 16164
rect 34567 16136 34612 16164
rect 31996 16124 32002 16136
rect 34600 16127 34612 16136
rect 34606 16124 34612 16127
rect 34664 16124 34670 16176
rect 38930 16124 38936 16176
rect 38988 16164 38994 16176
rect 38988 16136 43024 16164
rect 38988 16124 38994 16136
rect 24949 16099 25007 16105
rect 24949 16065 24961 16099
rect 24995 16065 25007 16099
rect 24949 16059 25007 16065
rect 25130 16056 25136 16108
rect 25188 16096 25194 16108
rect 25225 16099 25283 16105
rect 25225 16096 25237 16099
rect 25188 16068 25237 16096
rect 25188 16056 25194 16068
rect 25225 16065 25237 16068
rect 25271 16065 25283 16099
rect 25225 16059 25283 16065
rect 26510 16056 26516 16108
rect 26568 16056 26574 16108
rect 27062 16056 27068 16108
rect 27120 16056 27126 16108
rect 27706 16056 27712 16108
rect 27764 16096 27770 16108
rect 27890 16096 27896 16108
rect 27764 16068 27896 16096
rect 27764 16056 27770 16068
rect 27890 16056 27896 16068
rect 27948 16056 27954 16108
rect 28258 16056 28264 16108
rect 28316 16056 28322 16108
rect 28994 16056 29000 16108
rect 29052 16056 29058 16108
rect 31294 16056 31300 16108
rect 31352 16056 31358 16108
rect 31570 16056 31576 16108
rect 31628 16096 31634 16108
rect 32398 16105 32404 16108
rect 32125 16099 32183 16105
rect 32125 16096 32137 16099
rect 31628 16068 32137 16096
rect 31628 16056 31634 16068
rect 32125 16065 32137 16068
rect 32171 16065 32183 16099
rect 32125 16059 32183 16065
rect 32392 16059 32404 16105
rect 32398 16056 32404 16059
rect 32456 16056 32462 16108
rect 34238 16056 34244 16108
rect 34296 16056 34302 16108
rect 34330 16056 34336 16108
rect 34388 16056 34394 16108
rect 37550 16056 37556 16108
rect 37608 16056 37614 16108
rect 39390 16056 39396 16108
rect 39448 16096 39454 16108
rect 39577 16099 39635 16105
rect 39577 16096 39589 16099
rect 39448 16068 39589 16096
rect 39448 16056 39454 16068
rect 39577 16065 39589 16068
rect 39623 16065 39635 16099
rect 39577 16059 39635 16065
rect 40129 16099 40187 16105
rect 40129 16065 40141 16099
rect 40175 16096 40187 16099
rect 40218 16096 40224 16108
rect 40175 16068 40224 16096
rect 40175 16065 40187 16068
rect 40129 16059 40187 16065
rect 40218 16056 40224 16068
rect 40276 16056 40282 16108
rect 40770 16056 40776 16108
rect 40828 16056 40834 16108
rect 41233 16099 41291 16105
rect 41233 16065 41245 16099
rect 41279 16065 41291 16099
rect 41233 16059 41291 16065
rect 24026 16028 24032 16040
rect 23124 16000 24032 16028
rect 20588 15988 20594 16000
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 24121 16031 24179 16037
rect 24121 15997 24133 16031
rect 24167 16028 24179 16031
rect 24673 16031 24731 16037
rect 24167 16000 24532 16028
rect 24167 15997 24179 16000
rect 24121 15991 24179 15997
rect 20165 15963 20223 15969
rect 20165 15929 20177 15963
rect 20211 15960 20223 15963
rect 24397 15963 24455 15969
rect 24397 15960 24409 15963
rect 20211 15932 24409 15960
rect 20211 15929 20223 15932
rect 20165 15923 20223 15929
rect 24397 15929 24409 15932
rect 24443 15929 24455 15963
rect 24397 15923 24455 15929
rect 20806 15892 20812 15904
rect 20088 15864 20812 15892
rect 20806 15852 20812 15864
rect 20864 15892 20870 15904
rect 22002 15892 22008 15904
rect 20864 15864 22008 15892
rect 20864 15852 20870 15864
rect 22002 15852 22008 15864
rect 22060 15852 22066 15904
rect 22189 15895 22247 15901
rect 22189 15861 22201 15895
rect 22235 15892 22247 15895
rect 22554 15892 22560 15904
rect 22235 15864 22560 15892
rect 22235 15861 22247 15864
rect 22189 15855 22247 15861
rect 22554 15852 22560 15864
rect 22612 15852 22618 15904
rect 22646 15852 22652 15904
rect 22704 15852 22710 15904
rect 22830 15852 22836 15904
rect 22888 15852 22894 15904
rect 23290 15852 23296 15904
rect 23348 15852 23354 15904
rect 24504 15892 24532 16000
rect 24673 15997 24685 16031
rect 24719 16028 24731 16031
rect 24719 16000 32168 16028
rect 24719 15997 24731 16000
rect 24673 15991 24731 15997
rect 24581 15963 24639 15969
rect 24581 15929 24593 15963
rect 24627 15960 24639 15963
rect 25133 15963 25191 15969
rect 25133 15960 25145 15963
rect 24627 15932 25145 15960
rect 24627 15929 24639 15932
rect 24581 15923 24639 15929
rect 25133 15929 25145 15932
rect 25179 15929 25191 15963
rect 25133 15923 25191 15929
rect 27341 15963 27399 15969
rect 27341 15929 27353 15963
rect 27387 15960 27399 15963
rect 27706 15960 27712 15972
rect 27387 15932 27712 15960
rect 27387 15929 27399 15932
rect 27341 15923 27399 15929
rect 27706 15920 27712 15932
rect 27764 15960 27770 15972
rect 30098 15960 30104 15972
rect 27764 15932 30104 15960
rect 27764 15920 27770 15932
rect 30098 15920 30104 15932
rect 30156 15960 30162 15972
rect 30282 15960 30288 15972
rect 30156 15932 30288 15960
rect 30156 15920 30162 15932
rect 30282 15920 30288 15932
rect 30340 15920 30346 15972
rect 25314 15892 25320 15904
rect 24504 15864 25320 15892
rect 25314 15852 25320 15864
rect 25372 15892 25378 15904
rect 26050 15892 26056 15904
rect 25372 15864 26056 15892
rect 25372 15852 25378 15864
rect 26050 15852 26056 15864
rect 26108 15852 26114 15904
rect 26697 15895 26755 15901
rect 26697 15861 26709 15895
rect 26743 15892 26755 15895
rect 28166 15892 28172 15904
rect 26743 15864 28172 15892
rect 26743 15861 26755 15864
rect 26697 15855 26755 15861
rect 28166 15852 28172 15864
rect 28224 15852 28230 15904
rect 28442 15852 28448 15904
rect 28500 15852 28506 15904
rect 29181 15895 29239 15901
rect 29181 15861 29193 15895
rect 29227 15892 29239 15895
rect 29638 15892 29644 15904
rect 29227 15864 29644 15892
rect 29227 15861 29239 15864
rect 29181 15855 29239 15861
rect 29638 15852 29644 15864
rect 29696 15852 29702 15904
rect 32140 15892 32168 16000
rect 37274 15988 37280 16040
rect 37332 15988 37338 16040
rect 40310 15988 40316 16040
rect 40368 16028 40374 16040
rect 40681 16031 40739 16037
rect 40681 16028 40693 16031
rect 40368 16000 40693 16028
rect 40368 15988 40374 16000
rect 40681 15997 40693 16000
rect 40727 15997 40739 16031
rect 40681 15991 40739 15997
rect 38289 15963 38347 15969
rect 38289 15929 38301 15963
rect 38335 15960 38347 15963
rect 38838 15960 38844 15972
rect 38335 15932 38844 15960
rect 38335 15929 38347 15932
rect 38289 15923 38347 15929
rect 38838 15920 38844 15932
rect 38896 15920 38902 15972
rect 39022 15920 39028 15972
rect 39080 15960 39086 15972
rect 39761 15963 39819 15969
rect 39761 15960 39773 15963
rect 39080 15932 39773 15960
rect 39080 15920 39086 15932
rect 39761 15929 39773 15932
rect 39807 15960 39819 15963
rect 41248 15960 41276 16059
rect 42150 16056 42156 16108
rect 42208 16096 42214 16108
rect 42521 16099 42579 16105
rect 42521 16096 42533 16099
rect 42208 16068 42533 16096
rect 42208 16056 42214 16068
rect 42521 16065 42533 16068
rect 42567 16065 42579 16099
rect 42521 16059 42579 16065
rect 42702 16056 42708 16108
rect 42760 16056 42766 16108
rect 42996 16105 43024 16136
rect 42981 16099 43039 16105
rect 42981 16065 42993 16099
rect 43027 16065 43039 16099
rect 42981 16059 43039 16065
rect 44726 16056 44732 16108
rect 44784 16096 44790 16108
rect 45005 16099 45063 16105
rect 45005 16096 45017 16099
rect 44784 16068 45017 16096
rect 44784 16056 44790 16068
rect 45005 16065 45017 16068
rect 45051 16065 45063 16099
rect 45005 16059 45063 16065
rect 45741 16099 45799 16105
rect 45741 16065 45753 16099
rect 45787 16096 45799 16099
rect 45830 16096 45836 16108
rect 45787 16068 45836 16096
rect 45787 16065 45799 16068
rect 45741 16059 45799 16065
rect 45830 16056 45836 16068
rect 45888 16056 45894 16108
rect 46474 16056 46480 16108
rect 46532 16056 46538 16108
rect 41325 16031 41383 16037
rect 41325 15997 41337 16031
rect 41371 16028 41383 16031
rect 42720 16028 42748 16056
rect 43073 16031 43131 16037
rect 43073 16028 43085 16031
rect 41371 16000 42656 16028
rect 42720 16000 43085 16028
rect 41371 15997 41383 16000
rect 41325 15991 41383 15997
rect 42518 15960 42524 15972
rect 39807 15932 42524 15960
rect 39807 15929 39819 15932
rect 39761 15923 39819 15929
rect 42518 15920 42524 15932
rect 42576 15920 42582 15972
rect 42628 15960 42656 16000
rect 43073 15997 43085 16000
rect 43119 15997 43131 16031
rect 43073 15991 43131 15997
rect 43257 16031 43315 16037
rect 43257 15997 43269 16031
rect 43303 16028 43315 16031
rect 44818 16028 44824 16040
rect 43303 16000 44824 16028
rect 43303 15997 43315 16000
rect 43257 15991 43315 15997
rect 44818 15988 44824 16000
rect 44876 15988 44882 16040
rect 45094 15988 45100 16040
rect 45152 15988 45158 16040
rect 45462 15988 45468 16040
rect 45520 15988 45526 16040
rect 44910 15960 44916 15972
rect 42628 15932 44916 15960
rect 44910 15920 44916 15932
rect 44968 15920 44974 15972
rect 36078 15892 36084 15904
rect 32140 15864 36084 15892
rect 36078 15852 36084 15864
rect 36136 15852 36142 15904
rect 43165 15895 43223 15901
rect 43165 15861 43177 15895
rect 43211 15892 43223 15895
rect 43714 15892 43720 15904
rect 43211 15864 43720 15892
rect 43211 15861 43223 15864
rect 43165 15855 43223 15861
rect 43714 15852 43720 15864
rect 43772 15852 43778 15904
rect 46658 15852 46664 15904
rect 46716 15852 46722 15904
rect 1104 15802 47104 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 47104 15802
rect 1104 15728 47104 15750
rect 2590 15648 2596 15700
rect 2648 15688 2654 15700
rect 2777 15691 2835 15697
rect 2777 15688 2789 15691
rect 2648 15660 2789 15688
rect 2648 15648 2654 15660
rect 2777 15657 2789 15660
rect 2823 15657 2835 15691
rect 8570 15688 8576 15700
rect 2777 15651 2835 15657
rect 5828 15660 8576 15688
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 5828 15552 5856 15660
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 8938 15648 8944 15700
rect 8996 15688 9002 15700
rect 10134 15688 10140 15700
rect 8996 15660 10140 15688
rect 8996 15648 9002 15660
rect 7098 15580 7104 15632
rect 7156 15620 7162 15632
rect 7193 15623 7251 15629
rect 7193 15620 7205 15623
rect 7156 15592 7205 15620
rect 7156 15580 7162 15592
rect 7193 15589 7205 15592
rect 7239 15589 7251 15623
rect 7193 15583 7251 15589
rect 8021 15623 8079 15629
rect 8021 15589 8033 15623
rect 8067 15589 8079 15623
rect 8021 15583 8079 15589
rect 4847 15524 5856 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 3786 15484 3792 15496
rect 3007 15456 3792 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 4525 15487 4583 15493
rect 4525 15453 4537 15487
rect 4571 15484 4583 15487
rect 4614 15484 4620 15496
rect 4571 15456 4620 15484
rect 4571 15453 4583 15456
rect 4525 15447 4583 15453
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 5718 15444 5724 15496
rect 5776 15444 5782 15496
rect 5810 15444 5816 15496
rect 5868 15444 5874 15496
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8036 15484 8064 15583
rect 8570 15512 8576 15564
rect 8628 15512 8634 15564
rect 9140 15561 9168 15660
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 10781 15691 10839 15697
rect 10781 15657 10793 15691
rect 10827 15688 10839 15691
rect 21450 15688 21456 15700
rect 10827 15660 21456 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 22097 15691 22155 15697
rect 22097 15657 22109 15691
rect 22143 15688 22155 15691
rect 22462 15688 22468 15700
rect 22143 15660 22468 15688
rect 22143 15657 22155 15660
rect 22097 15651 22155 15657
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 22554 15648 22560 15700
rect 22612 15688 22618 15700
rect 22612 15660 30604 15688
rect 22612 15648 22618 15660
rect 14553 15623 14611 15629
rect 14553 15589 14565 15623
rect 14599 15589 14611 15623
rect 14553 15583 14611 15589
rect 9125 15555 9183 15561
rect 9125 15521 9137 15555
rect 9171 15521 9183 15555
rect 9125 15515 9183 15521
rect 9490 15512 9496 15564
rect 9548 15552 9554 15564
rect 9585 15555 9643 15561
rect 9585 15552 9597 15555
rect 9548 15524 9597 15552
rect 9548 15512 9554 15524
rect 9585 15521 9597 15524
rect 9631 15521 9643 15555
rect 9585 15515 9643 15521
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 9861 15555 9919 15561
rect 9861 15552 9873 15555
rect 9732 15524 9873 15552
rect 9732 15512 9738 15524
rect 9861 15521 9873 15524
rect 9907 15521 9919 15555
rect 9861 15515 9919 15521
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15552 10195 15555
rect 10502 15552 10508 15564
rect 10183 15524 10508 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 10502 15512 10508 15524
rect 10560 15512 10566 15564
rect 12066 15512 12072 15564
rect 12124 15552 12130 15564
rect 12161 15555 12219 15561
rect 12161 15552 12173 15555
rect 12124 15524 12173 15552
rect 12124 15512 12130 15524
rect 12161 15521 12173 15524
rect 12207 15521 12219 15555
rect 14568 15552 14596 15583
rect 14642 15580 14648 15632
rect 14700 15620 14706 15632
rect 14700 15592 14872 15620
rect 14700 15580 14706 15592
rect 14844 15561 14872 15592
rect 15838 15580 15844 15632
rect 15896 15620 15902 15632
rect 17129 15623 17187 15629
rect 17129 15620 17141 15623
rect 15896 15592 17141 15620
rect 15896 15580 15902 15592
rect 17129 15589 17141 15592
rect 17175 15589 17187 15623
rect 17129 15583 17187 15589
rect 17497 15623 17555 15629
rect 17497 15589 17509 15623
rect 17543 15589 17555 15623
rect 17497 15583 17555 15589
rect 17604 15592 20116 15620
rect 14829 15555 14887 15561
rect 14568 15524 14688 15552
rect 12161 15515 12219 15521
rect 7975 15456 8064 15484
rect 8389 15487 8447 15493
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 8754 15484 8760 15496
rect 8435 15456 8760 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 8754 15444 8760 15456
rect 8812 15484 8818 15496
rect 8938 15484 8944 15496
rect 8812 15456 8944 15484
rect 8812 15444 8818 15456
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 9950 15444 9956 15496
rect 10008 15493 10014 15496
rect 10008 15487 10036 15493
rect 10024 15453 10036 15487
rect 10008 15447 10036 15453
rect 10008 15444 10014 15447
rect 6058 15419 6116 15425
rect 6058 15416 6070 15419
rect 5552 15388 6070 15416
rect 4154 15308 4160 15360
rect 4212 15308 4218 15360
rect 4617 15351 4675 15357
rect 4617 15317 4629 15351
rect 4663 15348 4675 15351
rect 4706 15348 4712 15360
rect 4663 15320 4712 15348
rect 4663 15317 4675 15320
rect 4617 15311 4675 15317
rect 4706 15308 4712 15320
rect 4764 15348 4770 15360
rect 5258 15348 5264 15360
rect 4764 15320 5264 15348
rect 4764 15308 4770 15320
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 5552 15357 5580 15388
rect 6058 15385 6070 15388
rect 6104 15385 6116 15419
rect 6058 15379 6116 15385
rect 7190 15376 7196 15428
rect 7248 15416 7254 15428
rect 8481 15419 8539 15425
rect 8481 15416 8493 15419
rect 7248 15388 8493 15416
rect 7248 15376 7254 15388
rect 8481 15385 8493 15388
rect 8527 15385 8539 15419
rect 8481 15379 8539 15385
rect 12428 15419 12486 15425
rect 12428 15385 12440 15419
rect 12474 15416 12486 15419
rect 12526 15416 12532 15428
rect 12474 15388 12532 15416
rect 12474 15385 12486 15388
rect 12428 15379 12486 15385
rect 5537 15351 5595 15357
rect 5537 15317 5549 15351
rect 5583 15317 5595 15351
rect 5537 15311 5595 15317
rect 7742 15308 7748 15360
rect 7800 15308 7806 15360
rect 8496 15348 8524 15379
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 14660 15416 14688 15524
rect 14829 15521 14841 15555
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 17405 15487 17463 15493
rect 14783 15456 15240 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 15074 15419 15132 15425
rect 15074 15416 15086 15419
rect 14660 15388 15086 15416
rect 15074 15385 15086 15388
rect 15120 15385 15132 15419
rect 15212 15416 15240 15456
rect 15396 15456 17080 15484
rect 15286 15416 15292 15428
rect 15212 15388 15292 15416
rect 15074 15379 15132 15385
rect 15286 15376 15292 15388
rect 15344 15376 15350 15428
rect 10226 15348 10232 15360
rect 8496 15320 10232 15348
rect 10226 15308 10232 15320
rect 10284 15308 10290 15360
rect 13170 15308 13176 15360
rect 13228 15348 13234 15360
rect 13541 15351 13599 15357
rect 13541 15348 13553 15351
rect 13228 15320 13553 15348
rect 13228 15308 13234 15320
rect 13541 15317 13553 15320
rect 13587 15348 13599 15351
rect 15396 15348 15424 15456
rect 16945 15419 17003 15425
rect 16945 15385 16957 15419
rect 16991 15385 17003 15419
rect 17052 15416 17080 15456
rect 17405 15453 17417 15487
rect 17451 15484 17463 15487
rect 17512 15484 17540 15583
rect 17451 15456 17540 15484
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 17604 15416 17632 15592
rect 20088 15564 20116 15592
rect 20346 15580 20352 15632
rect 20404 15580 20410 15632
rect 21545 15623 21603 15629
rect 21545 15589 21557 15623
rect 21591 15620 21603 15623
rect 21913 15623 21971 15629
rect 21913 15620 21925 15623
rect 21591 15592 21925 15620
rect 21591 15589 21603 15592
rect 21545 15583 21603 15589
rect 21913 15589 21925 15592
rect 21959 15589 21971 15623
rect 21913 15583 21971 15589
rect 22002 15580 22008 15632
rect 22060 15620 22066 15632
rect 25130 15620 25136 15632
rect 22060 15592 25136 15620
rect 22060 15580 22066 15592
rect 25130 15580 25136 15592
rect 25188 15580 25194 15632
rect 17770 15512 17776 15564
rect 17828 15552 17834 15564
rect 18049 15555 18107 15561
rect 18049 15552 18061 15555
rect 17828 15524 18061 15552
rect 17828 15512 17834 15524
rect 18049 15521 18061 15524
rect 18095 15521 18107 15555
rect 18049 15515 18107 15521
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 19889 15555 19947 15561
rect 19889 15552 19901 15555
rect 19392 15524 19901 15552
rect 19392 15512 19398 15524
rect 19889 15521 19901 15524
rect 19935 15521 19947 15555
rect 19889 15515 19947 15521
rect 20070 15512 20076 15564
rect 20128 15552 20134 15564
rect 20625 15555 20683 15561
rect 20625 15552 20637 15555
rect 20128 15524 20637 15552
rect 20128 15512 20134 15524
rect 20625 15521 20637 15524
rect 20671 15521 20683 15555
rect 20625 15515 20683 15521
rect 20898 15512 20904 15564
rect 20956 15512 20962 15564
rect 21266 15512 21272 15564
rect 21324 15552 21330 15564
rect 24118 15552 24124 15564
rect 21324 15524 24124 15552
rect 21324 15512 21330 15524
rect 24118 15512 24124 15524
rect 24176 15512 24182 15564
rect 29549 15555 29607 15561
rect 29549 15552 29561 15555
rect 29012 15524 29561 15552
rect 17957 15487 18015 15493
rect 17957 15484 17969 15487
rect 17052 15388 17632 15416
rect 17696 15456 17969 15484
rect 16945 15379 17003 15385
rect 13587 15320 15424 15348
rect 13587 15317 13599 15320
rect 13541 15311 13599 15317
rect 16206 15308 16212 15360
rect 16264 15308 16270 15360
rect 16960 15348 16988 15379
rect 17126 15348 17132 15360
rect 16960 15320 17132 15348
rect 17126 15308 17132 15320
rect 17184 15308 17190 15360
rect 17218 15308 17224 15360
rect 17276 15308 17282 15360
rect 17310 15308 17316 15360
rect 17368 15348 17374 15360
rect 17696 15348 17724 15456
rect 17957 15453 17969 15456
rect 18003 15484 18015 15487
rect 19518 15484 19524 15496
rect 18003 15456 19524 15484
rect 18003 15453 18015 15456
rect 17957 15447 18015 15453
rect 19518 15444 19524 15456
rect 19576 15444 19582 15496
rect 19702 15444 19708 15496
rect 19760 15444 19766 15496
rect 20714 15444 20720 15496
rect 20772 15493 20778 15496
rect 20772 15487 20800 15493
rect 20788 15453 20800 15487
rect 20772 15447 20800 15453
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15484 21695 15487
rect 21910 15484 21916 15496
rect 21683 15456 21916 15484
rect 21683 15453 21695 15456
rect 21637 15447 21695 15453
rect 20772 15444 20778 15447
rect 21910 15444 21916 15456
rect 21968 15444 21974 15496
rect 23474 15444 23480 15496
rect 23532 15484 23538 15496
rect 24854 15484 24860 15496
rect 23532 15456 24860 15484
rect 23532 15444 23538 15456
rect 24854 15444 24860 15456
rect 24912 15444 24918 15496
rect 26053 15487 26111 15493
rect 26053 15453 26065 15487
rect 26099 15484 26111 15487
rect 26786 15484 26792 15496
rect 26099 15456 26792 15484
rect 26099 15453 26111 15456
rect 26053 15447 26111 15453
rect 26786 15444 26792 15456
rect 26844 15484 26850 15496
rect 29012 15484 29040 15524
rect 29549 15521 29561 15524
rect 29595 15521 29607 15555
rect 29549 15515 29607 15521
rect 26844 15456 29040 15484
rect 26844 15444 26850 15456
rect 29362 15444 29368 15496
rect 29420 15444 29426 15496
rect 17865 15419 17923 15425
rect 17865 15385 17877 15419
rect 17911 15416 17923 15419
rect 18322 15416 18328 15428
rect 17911 15388 18328 15416
rect 17911 15385 17923 15388
rect 17865 15379 17923 15385
rect 18322 15376 18328 15388
rect 18380 15376 18386 15428
rect 26326 15425 26332 15428
rect 26320 15379 26332 15425
rect 26326 15376 26332 15379
rect 26384 15376 26390 15428
rect 29086 15416 29092 15428
rect 26896 15388 29092 15416
rect 17368 15320 17724 15348
rect 17368 15308 17374 15320
rect 18230 15308 18236 15360
rect 18288 15348 18294 15360
rect 26896 15348 26924 15388
rect 29086 15376 29092 15388
rect 29144 15376 29150 15428
rect 29794 15419 29852 15425
rect 29794 15416 29806 15419
rect 29196 15388 29806 15416
rect 18288 15320 26924 15348
rect 18288 15308 18294 15320
rect 27338 15308 27344 15360
rect 27396 15348 27402 15360
rect 29196 15357 29224 15388
rect 29794 15385 29806 15388
rect 29840 15385 29852 15419
rect 30576 15416 30604 15660
rect 32398 15648 32404 15700
rect 32456 15648 32462 15700
rect 34238 15648 34244 15700
rect 34296 15688 34302 15700
rect 34701 15691 34759 15697
rect 34701 15688 34713 15691
rect 34296 15660 34713 15688
rect 34296 15648 34302 15660
rect 34701 15657 34713 15660
rect 34747 15657 34759 15691
rect 34701 15651 34759 15657
rect 36262 15648 36268 15700
rect 36320 15688 36326 15700
rect 36357 15691 36415 15697
rect 36357 15688 36369 15691
rect 36320 15660 36369 15688
rect 36320 15648 36326 15660
rect 36357 15657 36369 15660
rect 36403 15688 36415 15691
rect 36998 15688 37004 15700
rect 36403 15660 37004 15688
rect 36403 15657 36415 15660
rect 36357 15651 36415 15657
rect 36998 15648 37004 15660
rect 37056 15648 37062 15700
rect 37921 15691 37979 15697
rect 37921 15657 37933 15691
rect 37967 15688 37979 15691
rect 39850 15688 39856 15700
rect 37967 15660 39856 15688
rect 37967 15657 37979 15660
rect 37921 15651 37979 15657
rect 39850 15648 39856 15660
rect 39908 15648 39914 15700
rect 45738 15648 45744 15700
rect 45796 15688 45802 15700
rect 46201 15691 46259 15697
rect 46201 15688 46213 15691
rect 45796 15660 46213 15688
rect 45796 15648 45802 15660
rect 46201 15657 46213 15660
rect 46247 15657 46259 15691
rect 46201 15651 46259 15657
rect 31573 15623 31631 15629
rect 31573 15589 31585 15623
rect 31619 15620 31631 15623
rect 31619 15592 31754 15620
rect 31619 15589 31631 15592
rect 31573 15583 31631 15589
rect 31726 15484 31754 15592
rect 38102 15580 38108 15632
rect 38160 15620 38166 15632
rect 46474 15620 46480 15632
rect 38160 15592 46480 15620
rect 38160 15580 38166 15592
rect 46474 15580 46480 15592
rect 46532 15580 46538 15632
rect 32030 15512 32036 15564
rect 32088 15552 32094 15564
rect 32125 15555 32183 15561
rect 32125 15552 32137 15555
rect 32088 15524 32137 15552
rect 32088 15512 32094 15524
rect 32125 15521 32137 15524
rect 32171 15521 32183 15555
rect 32125 15515 32183 15521
rect 33686 15512 33692 15564
rect 33744 15552 33750 15564
rect 35253 15555 35311 15561
rect 35253 15552 35265 15555
rect 33744 15524 35265 15552
rect 33744 15512 33750 15524
rect 35253 15521 35265 15524
rect 35299 15521 35311 15555
rect 35253 15515 35311 15521
rect 39206 15512 39212 15564
rect 39264 15552 39270 15564
rect 39577 15555 39635 15561
rect 39577 15552 39589 15555
rect 39264 15524 39589 15552
rect 39264 15512 39270 15524
rect 39577 15521 39589 15524
rect 39623 15552 39635 15555
rect 40037 15555 40095 15561
rect 40037 15552 40049 15555
rect 39623 15524 40049 15552
rect 39623 15521 39635 15524
rect 39577 15515 39635 15521
rect 40037 15521 40049 15524
rect 40083 15521 40095 15555
rect 40037 15515 40095 15521
rect 45554 15512 45560 15564
rect 45612 15512 45618 15564
rect 32585 15487 32643 15493
rect 32585 15484 32597 15487
rect 31726 15456 32597 15484
rect 32585 15453 32597 15456
rect 32631 15453 32643 15487
rect 32585 15447 32643 15453
rect 34422 15444 34428 15496
rect 34480 15484 34486 15496
rect 35069 15487 35127 15493
rect 35069 15484 35081 15487
rect 34480 15456 35081 15484
rect 34480 15444 34486 15456
rect 35069 15453 35081 15456
rect 35115 15453 35127 15487
rect 35069 15447 35127 15453
rect 35161 15487 35219 15493
rect 35161 15453 35173 15487
rect 35207 15484 35219 15487
rect 35986 15484 35992 15496
rect 35207 15456 35992 15484
rect 35207 15453 35219 15456
rect 35161 15447 35219 15453
rect 35986 15444 35992 15456
rect 36044 15444 36050 15496
rect 36173 15487 36231 15493
rect 36173 15453 36185 15487
rect 36219 15484 36231 15487
rect 36538 15484 36544 15496
rect 36219 15456 36544 15484
rect 36219 15453 36231 15456
rect 36173 15447 36231 15453
rect 36538 15444 36544 15456
rect 36596 15444 36602 15496
rect 36906 15444 36912 15496
rect 36964 15444 36970 15496
rect 37185 15487 37243 15493
rect 37185 15453 37197 15487
rect 37231 15453 37243 15487
rect 37185 15447 37243 15453
rect 40313 15487 40371 15493
rect 40313 15453 40325 15487
rect 40359 15484 40371 15487
rect 41230 15484 41236 15496
rect 40359 15456 41236 15484
rect 40359 15453 40371 15456
rect 40313 15447 40371 15453
rect 37200 15416 37228 15447
rect 41230 15444 41236 15456
rect 41288 15444 41294 15496
rect 45186 15444 45192 15496
rect 45244 15484 45250 15496
rect 45281 15487 45339 15493
rect 45281 15484 45293 15487
rect 45244 15456 45293 15484
rect 45244 15444 45250 15456
rect 45281 15453 45293 15456
rect 45327 15453 45339 15487
rect 45281 15447 45339 15453
rect 46382 15444 46388 15496
rect 46440 15444 46446 15496
rect 30576 15388 37228 15416
rect 39393 15419 39451 15425
rect 29794 15379 29852 15385
rect 39393 15385 39405 15419
rect 39439 15416 39451 15419
rect 39758 15416 39764 15428
rect 39439 15388 39764 15416
rect 39439 15385 39451 15388
rect 39393 15379 39451 15385
rect 39758 15376 39764 15388
rect 39816 15376 39822 15428
rect 27433 15351 27491 15357
rect 27433 15348 27445 15351
rect 27396 15320 27445 15348
rect 27396 15308 27402 15320
rect 27433 15317 27445 15320
rect 27479 15317 27491 15351
rect 27433 15311 27491 15317
rect 29181 15351 29239 15357
rect 29181 15317 29193 15351
rect 29227 15317 29239 15351
rect 29181 15311 29239 15317
rect 30926 15308 30932 15360
rect 30984 15308 30990 15360
rect 31938 15308 31944 15360
rect 31996 15308 32002 15360
rect 32033 15351 32091 15357
rect 32033 15317 32045 15351
rect 32079 15348 32091 15351
rect 32490 15348 32496 15360
rect 32079 15320 32496 15348
rect 32079 15317 32091 15320
rect 32033 15311 32091 15317
rect 32490 15308 32496 15320
rect 32548 15308 32554 15360
rect 1104 15258 47104 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 47104 15258
rect 1104 15184 47104 15206
rect 4614 15104 4620 15156
rect 4672 15144 4678 15156
rect 4801 15147 4859 15153
rect 4801 15144 4813 15147
rect 4672 15116 4813 15144
rect 4672 15104 4678 15116
rect 4801 15113 4813 15116
rect 4847 15113 4859 15147
rect 4801 15107 4859 15113
rect 5258 15104 5264 15156
rect 5316 15144 5322 15156
rect 5316 15116 8892 15144
rect 5316 15104 5322 15116
rect 5810 15076 5816 15088
rect 3436 15048 5816 15076
rect 2406 14968 2412 15020
rect 2464 15008 2470 15020
rect 3436 15017 3464 15048
rect 5810 15036 5816 15048
rect 5868 15036 5874 15088
rect 6362 15036 6368 15088
rect 6420 15076 6426 15088
rect 6610 15079 6668 15085
rect 6610 15076 6622 15079
rect 6420 15048 6622 15076
rect 6420 15036 6426 15048
rect 6610 15045 6622 15048
rect 6656 15045 6668 15079
rect 6610 15039 6668 15045
rect 7742 15036 7748 15088
rect 7800 15076 7806 15088
rect 8174 15079 8232 15085
rect 8174 15076 8186 15079
rect 7800 15048 8186 15076
rect 7800 15036 7806 15048
rect 8174 15045 8186 15048
rect 8220 15045 8232 15079
rect 8174 15039 8232 15045
rect 3694 15017 3700 15020
rect 3421 15011 3479 15017
rect 3421 15008 3433 15011
rect 2464 14980 3433 15008
rect 2464 14968 2470 14980
rect 3421 14977 3433 14980
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3688 14971 3700 15017
rect 3694 14968 3700 14971
rect 3752 14968 3758 15020
rect 5828 14940 5856 15036
rect 7006 14968 7012 15020
rect 7064 15008 7070 15020
rect 7929 15011 7987 15017
rect 7929 15008 7941 15011
rect 7064 14980 7941 15008
rect 7064 14968 7070 14980
rect 7929 14977 7941 14980
rect 7975 14977 7987 15011
rect 8864 15008 8892 15116
rect 8938 15104 8944 15156
rect 8996 15144 9002 15156
rect 9309 15147 9367 15153
rect 9309 15144 9321 15147
rect 8996 15116 9321 15144
rect 8996 15104 9002 15116
rect 9309 15113 9321 15116
rect 9355 15113 9367 15147
rect 9309 15107 9367 15113
rect 9769 15147 9827 15153
rect 9769 15113 9781 15147
rect 9815 15144 9827 15147
rect 10686 15144 10692 15156
rect 9815 15116 10692 15144
rect 9815 15113 9827 15116
rect 9769 15107 9827 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 12526 15104 12532 15156
rect 12584 15104 12590 15156
rect 12805 15147 12863 15153
rect 12805 15113 12817 15147
rect 12851 15113 12863 15147
rect 12805 15107 12863 15113
rect 10134 15036 10140 15088
rect 10192 15036 10198 15088
rect 10226 15036 10232 15088
rect 10284 15036 10290 15088
rect 12713 15011 12771 15017
rect 8864 14980 12434 15008
rect 7929 14971 7987 14977
rect 6365 14943 6423 14949
rect 6365 14940 6377 14943
rect 5828 14912 6377 14940
rect 6365 14909 6377 14912
rect 6411 14909 6423 14943
rect 6365 14903 6423 14909
rect 10410 14900 10416 14952
rect 10468 14900 10474 14952
rect 12406 14940 12434 14980
rect 12713 14977 12725 15011
rect 12759 15008 12771 15011
rect 12820 15008 12848 15107
rect 13170 15104 13176 15156
rect 13228 15104 13234 15156
rect 15286 15104 15292 15156
rect 15344 15104 15350 15156
rect 15657 15147 15715 15153
rect 15657 15113 15669 15147
rect 15703 15144 15715 15147
rect 16206 15144 16212 15156
rect 15703 15116 16212 15144
rect 15703 15113 15715 15116
rect 15657 15107 15715 15113
rect 16206 15104 16212 15116
rect 16264 15104 16270 15156
rect 18322 15104 18328 15156
rect 18380 15144 18386 15156
rect 19334 15144 19340 15156
rect 18380 15116 19340 15144
rect 18380 15104 18386 15116
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 20254 15104 20260 15156
rect 20312 15144 20318 15156
rect 21545 15147 21603 15153
rect 20312 15116 21128 15144
rect 20312 15104 20318 15116
rect 13265 15079 13323 15085
rect 13265 15045 13277 15079
rect 13311 15076 13323 15079
rect 15749 15079 15807 15085
rect 15749 15076 15761 15079
rect 13311 15048 15761 15076
rect 13311 15045 13323 15048
rect 13265 15039 13323 15045
rect 15749 15045 15761 15048
rect 15795 15076 15807 15079
rect 16298 15076 16304 15088
rect 15795 15048 16304 15076
rect 15795 15045 15807 15048
rect 15749 15039 15807 15045
rect 12759 14980 12848 15008
rect 12759 14977 12771 14980
rect 12713 14971 12771 14977
rect 13280 14940 13308 15039
rect 16298 15036 16304 15048
rect 16356 15036 16362 15088
rect 17218 15085 17224 15088
rect 17212 15076 17224 15085
rect 17179 15048 17224 15076
rect 17212 15039 17224 15048
rect 17218 15036 17224 15039
rect 17276 15036 17282 15088
rect 21100 15085 21128 15116
rect 21545 15113 21557 15147
rect 21591 15144 21603 15147
rect 21591 15116 22094 15144
rect 21591 15113 21603 15116
rect 21545 15107 21603 15113
rect 21085 15079 21143 15085
rect 21085 15045 21097 15079
rect 21131 15045 21143 15079
rect 22066 15076 22094 15116
rect 22646 15104 22652 15156
rect 22704 15144 22710 15156
rect 23109 15147 23167 15153
rect 23109 15144 23121 15147
rect 22704 15116 23121 15144
rect 22704 15104 22710 15116
rect 23109 15113 23121 15116
rect 23155 15113 23167 15147
rect 23109 15107 23167 15113
rect 26326 15104 26332 15156
rect 26384 15104 26390 15156
rect 26973 15147 27031 15153
rect 26973 15113 26985 15147
rect 27019 15113 27031 15147
rect 26973 15107 27031 15113
rect 29273 15147 29331 15153
rect 29273 15113 29285 15147
rect 29319 15144 29331 15147
rect 29362 15144 29368 15156
rect 29319 15116 29368 15144
rect 29319 15113 29331 15116
rect 29273 15107 29331 15113
rect 23290 15076 23296 15088
rect 22066 15048 23296 15076
rect 21085 15039 21143 15045
rect 23290 15036 23296 15048
rect 23348 15036 23354 15088
rect 16942 14968 16948 15020
rect 17000 14968 17006 15020
rect 19334 14968 19340 15020
rect 19392 14968 19398 15020
rect 20070 14968 20076 15020
rect 20128 14968 20134 15020
rect 20346 14968 20352 15020
rect 20404 14968 20410 15020
rect 20990 14968 20996 15020
rect 21048 15008 21054 15020
rect 26418 15008 26424 15020
rect 21048 14980 26424 15008
rect 21048 14968 21054 14980
rect 26418 14968 26424 14980
rect 26476 14968 26482 15020
rect 26513 15011 26571 15017
rect 26513 14977 26525 15011
rect 26559 15008 26571 15011
rect 26988 15008 27016 15107
rect 29362 15104 29368 15116
rect 29420 15104 29426 15156
rect 29641 15147 29699 15153
rect 29641 15113 29653 15147
rect 29687 15144 29699 15147
rect 30650 15144 30656 15156
rect 29687 15116 30656 15144
rect 29687 15113 29699 15116
rect 29641 15107 29699 15113
rect 30650 15104 30656 15116
rect 30708 15144 30714 15156
rect 30926 15144 30932 15156
rect 30708 15116 30932 15144
rect 30708 15104 30714 15116
rect 30926 15104 30932 15116
rect 30984 15104 30990 15156
rect 42521 15147 42579 15153
rect 42521 15113 42533 15147
rect 42567 15144 42579 15147
rect 45186 15144 45192 15156
rect 42567 15116 45192 15144
rect 42567 15113 42579 15116
rect 42521 15107 42579 15113
rect 45186 15104 45192 15116
rect 45244 15104 45250 15156
rect 45649 15147 45707 15153
rect 45649 15113 45661 15147
rect 45695 15144 45707 15147
rect 46382 15144 46388 15156
rect 45695 15116 46388 15144
rect 45695 15113 45707 15116
rect 45649 15107 45707 15113
rect 46382 15104 46388 15116
rect 46440 15104 46446 15156
rect 28166 15036 28172 15088
rect 28224 15076 28230 15088
rect 29914 15076 29920 15088
rect 28224 15048 29920 15076
rect 28224 15036 28230 15048
rect 29914 15036 29920 15048
rect 29972 15076 29978 15088
rect 31294 15076 31300 15088
rect 29972 15048 31300 15076
rect 29972 15036 29978 15048
rect 31294 15036 31300 15048
rect 31352 15036 31358 15088
rect 40126 15076 40132 15088
rect 38948 15048 40132 15076
rect 26559 14980 27016 15008
rect 26559 14977 26571 14980
rect 26513 14971 26571 14977
rect 27338 14968 27344 15020
rect 27396 14968 27402 15020
rect 28626 14968 28632 15020
rect 28684 15008 28690 15020
rect 29181 15011 29239 15017
rect 29181 15008 29193 15011
rect 28684 14980 29193 15008
rect 28684 14968 28690 14980
rect 29181 14977 29193 14980
rect 29227 14977 29239 15011
rect 29181 14971 29239 14977
rect 33778 14968 33784 15020
rect 33836 14968 33842 15020
rect 35342 14968 35348 15020
rect 35400 15008 35406 15020
rect 35529 15011 35587 15017
rect 35529 15008 35541 15011
rect 35400 14980 35541 15008
rect 35400 14968 35406 14980
rect 35529 14977 35541 14980
rect 35575 15008 35587 15011
rect 37090 15008 37096 15020
rect 35575 14980 37096 15008
rect 35575 14977 35587 14980
rect 35529 14971 35587 14977
rect 37090 14968 37096 14980
rect 37148 14968 37154 15020
rect 38470 14968 38476 15020
rect 38528 15008 38534 15020
rect 38948 15017 38976 15048
rect 40126 15036 40132 15048
rect 40184 15036 40190 15088
rect 44266 15076 44272 15088
rect 43364 15048 44272 15076
rect 38841 15011 38899 15017
rect 38841 15008 38853 15011
rect 38528 14980 38853 15008
rect 38528 14968 38534 14980
rect 38841 14977 38853 14980
rect 38887 14977 38899 15011
rect 38841 14971 38899 14977
rect 38933 15011 38991 15017
rect 38933 14977 38945 15011
rect 38979 14977 38991 15011
rect 38933 14971 38991 14977
rect 39117 15011 39175 15017
rect 39117 14977 39129 15011
rect 39163 14977 39175 15011
rect 39117 14971 39175 14977
rect 12406 14912 13308 14940
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14940 13507 14943
rect 13630 14940 13636 14952
rect 13495 14912 13636 14940
rect 13495 14909 13507 14912
rect 13449 14903 13507 14909
rect 13630 14900 13636 14912
rect 13688 14900 13694 14952
rect 15930 14900 15936 14952
rect 15988 14900 15994 14952
rect 19153 14943 19211 14949
rect 19153 14909 19165 14943
rect 19199 14940 19211 14943
rect 19702 14940 19708 14952
rect 19199 14912 19708 14940
rect 19199 14909 19211 14912
rect 19153 14903 19211 14909
rect 19702 14900 19708 14912
rect 19760 14900 19766 14952
rect 20211 14943 20269 14949
rect 20211 14909 20223 14943
rect 20257 14940 20269 14943
rect 20714 14940 20720 14952
rect 20257 14912 20720 14940
rect 20257 14909 20269 14912
rect 20211 14903 20269 14909
rect 20714 14900 20720 14912
rect 20772 14900 20778 14952
rect 21726 14900 21732 14952
rect 21784 14940 21790 14952
rect 22649 14943 22707 14949
rect 22649 14940 22661 14943
rect 21784 14912 22661 14940
rect 21784 14900 21790 14912
rect 22649 14909 22661 14912
rect 22695 14909 22707 14943
rect 22649 14903 22707 14909
rect 26878 14900 26884 14952
rect 26936 14940 26942 14952
rect 27356 14940 27384 14968
rect 26936 14912 27384 14940
rect 26936 14900 26942 14912
rect 27430 14900 27436 14952
rect 27488 14900 27494 14952
rect 27525 14943 27583 14949
rect 27525 14909 27537 14943
rect 27571 14940 27583 14943
rect 28442 14940 28448 14952
rect 27571 14912 28448 14940
rect 27571 14909 27583 14912
rect 27525 14903 27583 14909
rect 28442 14900 28448 14912
rect 28500 14900 28506 14952
rect 29730 14900 29736 14952
rect 29788 14900 29794 14952
rect 29825 14943 29883 14949
rect 29825 14909 29837 14943
rect 29871 14909 29883 14943
rect 29825 14903 29883 14909
rect 35805 14943 35863 14949
rect 35805 14909 35817 14943
rect 35851 14940 35863 14943
rect 35894 14940 35900 14952
rect 35851 14912 35900 14940
rect 35851 14909 35863 14912
rect 35805 14903 35863 14909
rect 18690 14832 18696 14884
rect 18748 14872 18754 14884
rect 19797 14875 19855 14881
rect 19797 14872 19809 14875
rect 18748 14844 19809 14872
rect 18748 14832 18754 14844
rect 19797 14841 19809 14844
rect 19843 14841 19855 14875
rect 19797 14835 19855 14841
rect 7742 14764 7748 14816
rect 7800 14804 7806 14816
rect 9582 14804 9588 14816
rect 7800 14776 9588 14804
rect 7800 14764 7806 14776
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 20732 14804 20760 14900
rect 20993 14875 21051 14881
rect 20993 14841 21005 14875
rect 21039 14872 21051 14875
rect 21361 14875 21419 14881
rect 21361 14872 21373 14875
rect 21039 14844 21373 14872
rect 21039 14841 21051 14844
rect 20993 14835 21051 14841
rect 21361 14841 21373 14844
rect 21407 14841 21419 14875
rect 21361 14835 21419 14841
rect 23017 14875 23075 14881
rect 23017 14841 23029 14875
rect 23063 14872 23075 14875
rect 27798 14872 27804 14884
rect 23063 14844 27804 14872
rect 23063 14841 23075 14844
rect 23017 14835 23075 14841
rect 27798 14832 27804 14844
rect 27856 14832 27862 14884
rect 28460 14872 28488 14900
rect 29840 14872 29868 14903
rect 35894 14900 35900 14912
rect 35952 14900 35958 14952
rect 39132 14940 39160 14971
rect 39298 14968 39304 15020
rect 39356 14968 39362 15020
rect 39390 14968 39396 15020
rect 39448 14968 39454 15020
rect 41325 15011 41383 15017
rect 41325 14977 41337 15011
rect 41371 15008 41383 15011
rect 42150 15008 42156 15020
rect 41371 14980 42156 15008
rect 41371 14977 41383 14980
rect 41325 14971 41383 14977
rect 42150 14968 42156 14980
rect 42208 14968 42214 15020
rect 42518 14968 42524 15020
rect 42576 15008 42582 15020
rect 42705 15011 42763 15017
rect 42705 15008 42717 15011
rect 42576 14980 42717 15008
rect 42576 14968 42582 14980
rect 42705 14977 42717 14980
rect 42751 14977 42763 15011
rect 42705 14971 42763 14977
rect 43165 15011 43223 15017
rect 43165 14977 43177 15011
rect 43211 15008 43223 15011
rect 43254 15008 43260 15020
rect 43211 14980 43260 15008
rect 43211 14977 43223 14980
rect 43165 14971 43223 14977
rect 43254 14968 43260 14980
rect 43312 14968 43318 15020
rect 43364 15017 43392 15048
rect 43349 15011 43407 15017
rect 43349 14977 43361 15011
rect 43395 14977 43407 15011
rect 43349 14971 43407 14977
rect 43714 14968 43720 15020
rect 43772 14968 43778 15020
rect 44008 15017 44036 15048
rect 44266 15036 44272 15048
rect 44324 15036 44330 15088
rect 43809 15011 43867 15017
rect 43809 14977 43821 15011
rect 43855 14977 43867 15011
rect 43809 14971 43867 14977
rect 43993 15011 44051 15017
rect 43993 14977 44005 15011
rect 44039 14977 44051 15011
rect 43993 14971 44051 14977
rect 39853 14943 39911 14949
rect 39853 14940 39865 14943
rect 39132 14912 39865 14940
rect 39853 14909 39865 14912
rect 39899 14909 39911 14943
rect 43272 14940 43300 14968
rect 43824 14940 43852 14971
rect 45186 14968 45192 15020
rect 45244 14968 45250 15020
rect 43272 14912 43852 14940
rect 39853 14903 39911 14909
rect 28460 14844 29868 14872
rect 39025 14875 39083 14881
rect 39025 14841 39037 14875
rect 39071 14872 39083 14875
rect 39206 14872 39212 14884
rect 39071 14844 39212 14872
rect 39071 14841 39083 14844
rect 39025 14835 39083 14841
rect 39206 14832 39212 14844
rect 39264 14832 39270 14884
rect 43622 14832 43628 14884
rect 43680 14832 43686 14884
rect 16264 14776 20760 14804
rect 16264 14764 16270 14776
rect 23382 14764 23388 14816
rect 23440 14804 23446 14816
rect 26510 14804 26516 14816
rect 23440 14776 26516 14804
rect 23440 14764 23446 14776
rect 26510 14764 26516 14776
rect 26568 14764 26574 14816
rect 28997 14807 29055 14813
rect 28997 14773 29009 14807
rect 29043 14804 29055 14807
rect 29086 14804 29092 14816
rect 29043 14776 29092 14804
rect 29043 14773 29055 14776
rect 28997 14767 29055 14773
rect 29086 14764 29092 14776
rect 29144 14764 29150 14816
rect 33965 14807 34023 14813
rect 33965 14773 33977 14807
rect 34011 14804 34023 14807
rect 34146 14804 34152 14816
rect 34011 14776 34152 14804
rect 34011 14773 34023 14776
rect 33965 14767 34023 14773
rect 34146 14764 34152 14776
rect 34204 14804 34210 14816
rect 34330 14804 34336 14816
rect 34204 14776 34336 14804
rect 34204 14764 34210 14776
rect 34330 14764 34336 14776
rect 34388 14764 34394 14816
rect 38654 14764 38660 14816
rect 38712 14764 38718 14816
rect 39666 14764 39672 14816
rect 39724 14764 39730 14816
rect 41138 14764 41144 14816
rect 41196 14764 41202 14816
rect 42978 14764 42984 14816
rect 43036 14804 43042 14816
rect 43901 14807 43959 14813
rect 43901 14804 43913 14807
rect 43036 14776 43913 14804
rect 43036 14764 43042 14776
rect 43901 14773 43913 14776
rect 43947 14773 43959 14807
rect 43901 14767 43959 14773
rect 45462 14764 45468 14816
rect 45520 14764 45526 14816
rect 1104 14714 47104 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 47104 14714
rect 1104 14640 47104 14662
rect 3694 14560 3700 14612
rect 3752 14600 3758 14612
rect 3881 14603 3939 14609
rect 3881 14600 3893 14603
rect 3752 14572 3893 14600
rect 3752 14560 3758 14572
rect 3881 14569 3893 14572
rect 3927 14569 3939 14603
rect 3881 14563 3939 14569
rect 6546 14560 6552 14612
rect 6604 14560 6610 14612
rect 10226 14560 10232 14612
rect 10284 14600 10290 14612
rect 10284 14572 12434 14600
rect 10284 14560 10290 14572
rect 6914 14424 6920 14476
rect 6972 14464 6978 14476
rect 7101 14467 7159 14473
rect 7101 14464 7113 14467
rect 6972 14436 7113 14464
rect 6972 14424 6978 14436
rect 7101 14433 7113 14436
rect 7147 14433 7159 14467
rect 12406 14464 12434 14572
rect 18322 14560 18328 14612
rect 18380 14600 18386 14612
rect 19058 14600 19064 14612
rect 18380 14572 19064 14600
rect 18380 14560 18386 14572
rect 19058 14560 19064 14572
rect 19116 14600 19122 14612
rect 20346 14600 20352 14612
rect 19116 14572 20352 14600
rect 19116 14560 19122 14572
rect 20346 14560 20352 14572
rect 20404 14560 20410 14612
rect 24026 14560 24032 14612
rect 24084 14600 24090 14612
rect 24397 14603 24455 14609
rect 24397 14600 24409 14603
rect 24084 14572 24409 14600
rect 24084 14560 24090 14572
rect 24397 14569 24409 14572
rect 24443 14569 24455 14603
rect 24397 14563 24455 14569
rect 26418 14560 26424 14612
rect 26476 14600 26482 14612
rect 26476 14572 27752 14600
rect 26476 14560 26482 14572
rect 19794 14492 19800 14544
rect 19852 14532 19858 14544
rect 20530 14532 20536 14544
rect 19852 14504 20536 14532
rect 19852 14492 19858 14504
rect 20530 14492 20536 14504
rect 20588 14492 20594 14544
rect 27724 14532 27752 14572
rect 27798 14560 27804 14612
rect 27856 14560 27862 14612
rect 28626 14560 28632 14612
rect 28684 14560 28690 14612
rect 28902 14560 28908 14612
rect 28960 14600 28966 14612
rect 30653 14603 30711 14609
rect 30653 14600 30665 14603
rect 28960 14572 30665 14600
rect 28960 14560 28966 14572
rect 30653 14569 30665 14572
rect 30699 14569 30711 14603
rect 30653 14563 30711 14569
rect 30742 14560 30748 14612
rect 30800 14600 30806 14612
rect 31481 14603 31539 14609
rect 31481 14600 31493 14603
rect 30800 14572 31493 14600
rect 30800 14560 30806 14572
rect 31481 14569 31493 14572
rect 31527 14569 31539 14603
rect 31481 14563 31539 14569
rect 33502 14560 33508 14612
rect 33560 14600 33566 14612
rect 37185 14603 37243 14609
rect 37185 14600 37197 14603
rect 33560 14572 37197 14600
rect 33560 14560 33566 14572
rect 37185 14569 37197 14572
rect 37231 14600 37243 14603
rect 37642 14600 37648 14612
rect 37231 14572 37648 14600
rect 37231 14569 37243 14572
rect 37185 14563 37243 14569
rect 37642 14560 37648 14572
rect 37700 14560 37706 14612
rect 38013 14603 38071 14609
rect 38013 14569 38025 14603
rect 38059 14600 38071 14603
rect 38194 14600 38200 14612
rect 38059 14572 38200 14600
rect 38059 14569 38071 14572
rect 38013 14563 38071 14569
rect 38194 14560 38200 14572
rect 38252 14560 38258 14612
rect 39666 14560 39672 14612
rect 39724 14600 39730 14612
rect 40221 14603 40279 14609
rect 40221 14600 40233 14603
rect 39724 14572 40233 14600
rect 39724 14560 39730 14572
rect 40221 14569 40233 14572
rect 40267 14569 40279 14603
rect 40221 14563 40279 14569
rect 40310 14560 40316 14612
rect 40368 14560 40374 14612
rect 41230 14560 41236 14612
rect 41288 14600 41294 14612
rect 41969 14603 42027 14609
rect 41969 14600 41981 14603
rect 41288 14572 41981 14600
rect 41288 14560 41294 14572
rect 41969 14569 41981 14572
rect 42015 14569 42027 14603
rect 41969 14563 42027 14569
rect 29730 14532 29736 14544
rect 27724 14504 29736 14532
rect 18509 14467 18567 14473
rect 18509 14464 18521 14467
rect 12406 14436 18521 14464
rect 7101 14427 7159 14433
rect 18509 14433 18521 14436
rect 18555 14464 18567 14467
rect 19889 14467 19947 14473
rect 19889 14464 19901 14467
rect 18555 14436 19901 14464
rect 18555 14433 18567 14436
rect 18509 14427 18567 14433
rect 19889 14433 19901 14436
rect 19935 14433 19947 14467
rect 19889 14427 19947 14433
rect 22278 14424 22284 14476
rect 22336 14424 22342 14476
rect 25041 14467 25099 14473
rect 25041 14433 25053 14467
rect 25087 14464 25099 14467
rect 25222 14464 25228 14476
rect 25087 14436 25228 14464
rect 25087 14433 25099 14436
rect 25041 14427 25099 14433
rect 25222 14424 25228 14436
rect 25280 14424 25286 14476
rect 26602 14424 26608 14476
rect 26660 14424 26666 14476
rect 26970 14424 26976 14476
rect 27028 14473 27034 14476
rect 27028 14467 27056 14473
rect 27044 14433 27056 14467
rect 27028 14427 27056 14433
rect 27028 14424 27034 14427
rect 27522 14424 27528 14476
rect 27580 14464 27586 14476
rect 29104 14473 29132 14504
rect 29730 14492 29736 14504
rect 29788 14532 29794 14544
rect 40328 14532 40356 14560
rect 41984 14532 42012 14563
rect 42150 14560 42156 14612
rect 42208 14560 42214 14612
rect 43809 14603 43867 14609
rect 43809 14569 43821 14603
rect 43855 14600 43867 14603
rect 45370 14600 45376 14612
rect 43855 14572 45376 14600
rect 43855 14569 43867 14572
rect 43809 14563 43867 14569
rect 43824 14532 43852 14563
rect 45370 14560 45376 14572
rect 45428 14560 45434 14612
rect 29788 14504 31754 14532
rect 40328 14504 41092 14532
rect 41984 14504 43852 14532
rect 29788 14492 29794 14504
rect 28537 14467 28595 14473
rect 28537 14464 28549 14467
rect 27580 14436 28549 14464
rect 27580 14424 27586 14436
rect 28537 14433 28549 14436
rect 28583 14433 28595 14467
rect 28537 14427 28595 14433
rect 29089 14467 29147 14473
rect 29089 14433 29101 14467
rect 29135 14433 29147 14467
rect 29089 14427 29147 14433
rect 29178 14424 29184 14476
rect 29236 14424 29242 14476
rect 30558 14424 30564 14476
rect 30616 14464 30622 14476
rect 30834 14464 30840 14476
rect 30616 14436 30840 14464
rect 30616 14424 30622 14436
rect 30834 14424 30840 14436
rect 30892 14464 30898 14476
rect 31205 14467 31263 14473
rect 31205 14464 31217 14467
rect 30892 14436 31217 14464
rect 30892 14424 30898 14436
rect 31205 14433 31217 14436
rect 31251 14433 31263 14467
rect 31205 14427 31263 14433
rect 1394 14356 1400 14408
rect 1452 14356 1458 14408
rect 4062 14356 4068 14408
rect 4120 14356 4126 14408
rect 7009 14399 7067 14405
rect 7009 14365 7021 14399
rect 7055 14396 7067 14399
rect 7190 14396 7196 14408
rect 7055 14368 7196 14396
rect 7055 14365 7067 14368
rect 7009 14359 7067 14365
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 12158 14356 12164 14408
rect 12216 14396 12222 14408
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 12216 14368 12265 14396
rect 12216 14356 12222 14368
rect 12253 14365 12265 14368
rect 12299 14396 12311 14399
rect 13630 14396 13636 14408
rect 12299 14368 13636 14396
rect 12299 14365 12311 14368
rect 12253 14359 12311 14365
rect 13630 14356 13636 14368
rect 13688 14356 13694 14408
rect 15378 14356 15384 14408
rect 15436 14396 15442 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15436 14368 15853 14396
rect 15436 14356 15442 14368
rect 15841 14365 15853 14368
rect 15887 14396 15899 14399
rect 18233 14399 18291 14405
rect 15887 14368 17816 14396
rect 15887 14365 15899 14368
rect 15841 14359 15899 14365
rect 6917 14331 6975 14337
rect 6917 14297 6929 14331
rect 6963 14328 6975 14331
rect 7742 14328 7748 14340
rect 6963 14300 7748 14328
rect 6963 14297 6975 14300
rect 6917 14291 6975 14297
rect 7742 14288 7748 14300
rect 7800 14288 7806 14340
rect 12434 14288 12440 14340
rect 12492 14288 12498 14340
rect 15930 14288 15936 14340
rect 15988 14328 15994 14340
rect 16114 14328 16120 14340
rect 15988 14300 16120 14328
rect 15988 14288 15994 14300
rect 16114 14288 16120 14300
rect 16172 14288 16178 14340
rect 17788 14328 17816 14368
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 18598 14396 18604 14408
rect 18279 14368 18604 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 20070 14356 20076 14408
rect 20128 14396 20134 14408
rect 20165 14399 20223 14405
rect 20165 14396 20177 14399
rect 20128 14368 20177 14396
rect 20128 14356 20134 14368
rect 20165 14365 20177 14368
rect 20211 14396 20223 14399
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20211 14368 20913 14396
rect 20211 14365 20223 14368
rect 20165 14359 20223 14365
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 22066 14368 24072 14396
rect 20438 14328 20444 14340
rect 17788 14300 20444 14328
rect 20438 14288 20444 14300
rect 20496 14288 20502 14340
rect 20806 14288 20812 14340
rect 20864 14328 20870 14340
rect 22066 14328 22094 14368
rect 20864 14300 22094 14328
rect 23293 14331 23351 14337
rect 20864 14288 20870 14300
rect 23293 14297 23305 14331
rect 23339 14297 23351 14331
rect 23293 14291 23351 14297
rect 934 14220 940 14272
rect 992 14260 998 14272
rect 1581 14263 1639 14269
rect 1581 14260 1593 14263
rect 992 14232 1593 14260
rect 992 14220 998 14232
rect 1581 14229 1593 14232
rect 1627 14229 1639 14263
rect 1581 14223 1639 14229
rect 19794 14220 19800 14272
rect 19852 14260 19858 14272
rect 20993 14263 21051 14269
rect 20993 14260 21005 14263
rect 19852 14232 21005 14260
rect 19852 14220 19858 14232
rect 20993 14229 21005 14232
rect 21039 14229 21051 14263
rect 20993 14223 21051 14229
rect 21726 14220 21732 14272
rect 21784 14220 21790 14272
rect 22094 14220 22100 14272
rect 22152 14220 22158 14272
rect 22189 14263 22247 14269
rect 22189 14229 22201 14263
rect 22235 14260 22247 14263
rect 22738 14260 22744 14272
rect 22235 14232 22744 14260
rect 22235 14229 22247 14232
rect 22189 14223 22247 14229
rect 22738 14220 22744 14232
rect 22796 14220 22802 14272
rect 23308 14260 23336 14291
rect 23658 14288 23664 14340
rect 23716 14288 23722 14340
rect 24044 14328 24072 14368
rect 25590 14356 25596 14408
rect 25648 14356 25654 14408
rect 25961 14399 26019 14405
rect 25961 14365 25973 14399
rect 26007 14365 26019 14399
rect 25961 14359 26019 14365
rect 25866 14328 25872 14340
rect 24044 14300 25872 14328
rect 25866 14288 25872 14300
rect 25924 14288 25930 14340
rect 24302 14260 24308 14272
rect 23308 14232 24308 14260
rect 24302 14220 24308 14232
rect 24360 14220 24366 14272
rect 24762 14220 24768 14272
rect 24820 14220 24826 14272
rect 24854 14220 24860 14272
rect 24912 14220 24918 14272
rect 25406 14220 25412 14272
rect 25464 14220 25470 14272
rect 25976 14260 26004 14359
rect 26142 14356 26148 14408
rect 26200 14356 26206 14408
rect 26878 14356 26884 14408
rect 26936 14356 26942 14408
rect 27154 14356 27160 14408
rect 27212 14356 27218 14408
rect 28353 14399 28411 14405
rect 28353 14365 28365 14399
rect 28399 14396 28411 14399
rect 29546 14396 29552 14408
rect 28399 14368 29552 14396
rect 28399 14365 28411 14368
rect 28353 14359 28411 14365
rect 29546 14356 29552 14368
rect 29604 14356 29610 14408
rect 31726 14396 31754 14504
rect 31846 14424 31852 14476
rect 31904 14464 31910 14476
rect 32030 14464 32036 14476
rect 31904 14436 32036 14464
rect 31904 14424 31910 14436
rect 32030 14424 32036 14436
rect 32088 14424 32094 14476
rect 32490 14424 32496 14476
rect 32548 14464 32554 14476
rect 33873 14467 33931 14473
rect 33873 14464 33885 14467
rect 32548 14436 33885 14464
rect 32548 14424 32554 14436
rect 33873 14433 33885 14436
rect 33919 14464 33931 14467
rect 34238 14464 34244 14476
rect 33919 14436 34244 14464
rect 33919 14433 33931 14436
rect 33873 14427 33931 14433
rect 34238 14424 34244 14436
rect 34296 14424 34302 14476
rect 37734 14424 37740 14476
rect 37792 14464 37798 14476
rect 38197 14467 38255 14473
rect 38197 14464 38209 14467
rect 37792 14436 38209 14464
rect 37792 14424 37798 14436
rect 38197 14433 38209 14436
rect 38243 14464 38255 14467
rect 38470 14464 38476 14476
rect 38243 14436 38476 14464
rect 38243 14433 38255 14436
rect 38197 14427 38255 14433
rect 38470 14424 38476 14436
rect 38528 14424 38534 14476
rect 40586 14424 40592 14476
rect 40644 14424 40650 14476
rect 33597 14399 33655 14405
rect 33597 14396 33609 14399
rect 31726 14368 33609 14396
rect 33597 14365 33609 14368
rect 33643 14396 33655 14399
rect 35805 14399 35863 14405
rect 33643 14368 35388 14396
rect 33643 14365 33655 14368
rect 33597 14359 33655 14365
rect 28997 14331 29055 14337
rect 28997 14297 29009 14331
rect 29043 14328 29055 14331
rect 30742 14328 30748 14340
rect 29043 14300 30748 14328
rect 29043 14297 29055 14300
rect 28997 14291 29055 14297
rect 30742 14288 30748 14300
rect 30800 14288 30806 14340
rect 31113 14331 31171 14337
rect 31113 14297 31125 14331
rect 31159 14328 31171 14331
rect 35250 14328 35256 14340
rect 31159 14300 35256 14328
rect 31159 14297 31171 14300
rect 31113 14291 31171 14297
rect 35250 14288 35256 14300
rect 35308 14288 35314 14340
rect 26970 14260 26976 14272
rect 25976 14232 26976 14260
rect 26970 14220 26976 14232
rect 27028 14220 27034 14272
rect 27154 14220 27160 14272
rect 27212 14260 27218 14272
rect 28626 14260 28632 14272
rect 27212 14232 28632 14260
rect 27212 14220 27218 14232
rect 28626 14220 28632 14232
rect 28684 14260 28690 14272
rect 29779 14263 29837 14269
rect 29779 14260 29791 14263
rect 28684 14232 29791 14260
rect 28684 14220 28690 14232
rect 29779 14229 29791 14232
rect 29825 14229 29837 14263
rect 29779 14223 29837 14229
rect 31018 14220 31024 14272
rect 31076 14220 31082 14272
rect 31846 14220 31852 14272
rect 31904 14220 31910 14272
rect 31941 14263 31999 14269
rect 31941 14229 31953 14263
rect 31987 14260 31999 14263
rect 34514 14260 34520 14272
rect 31987 14232 34520 14260
rect 31987 14229 31999 14232
rect 31941 14223 31999 14229
rect 34514 14220 34520 14232
rect 34572 14220 34578 14272
rect 35360 14260 35388 14368
rect 35805 14365 35817 14399
rect 35851 14396 35863 14399
rect 35894 14396 35900 14408
rect 35851 14368 35900 14396
rect 35851 14365 35863 14368
rect 35805 14359 35863 14365
rect 35894 14356 35900 14368
rect 35952 14356 35958 14408
rect 38289 14399 38347 14405
rect 38289 14365 38301 14399
rect 38335 14396 38347 14399
rect 38562 14396 38568 14408
rect 38335 14368 38568 14396
rect 38335 14365 38347 14368
rect 38289 14359 38347 14365
rect 38562 14356 38568 14368
rect 38620 14356 38626 14408
rect 39850 14356 39856 14408
rect 39908 14356 39914 14408
rect 40037 14399 40095 14405
rect 40037 14365 40049 14399
rect 40083 14396 40095 14399
rect 40126 14396 40132 14408
rect 40083 14368 40132 14396
rect 40083 14365 40095 14368
rect 40037 14359 40095 14365
rect 40126 14356 40132 14368
rect 40184 14356 40190 14408
rect 40218 14356 40224 14408
rect 40276 14396 40282 14408
rect 40865 14399 40923 14405
rect 40865 14396 40877 14399
rect 40276 14368 40877 14396
rect 40276 14356 40282 14368
rect 40865 14365 40877 14368
rect 40911 14365 40923 14399
rect 40865 14359 40923 14365
rect 40954 14356 40960 14408
rect 41012 14405 41018 14408
rect 41012 14359 41020 14405
rect 41012 14356 41018 14359
rect 36078 14337 36084 14340
rect 36072 14291 36084 14337
rect 36078 14288 36084 14291
rect 36136 14288 36142 14340
rect 38013 14331 38071 14337
rect 38013 14297 38025 14331
rect 38059 14297 38071 14331
rect 38013 14291 38071 14297
rect 37826 14260 37832 14272
rect 35360 14232 37832 14260
rect 37826 14220 37832 14232
rect 37884 14220 37890 14272
rect 38028 14260 38056 14291
rect 38102 14288 38108 14340
rect 38160 14328 38166 14340
rect 38381 14331 38439 14337
rect 38381 14328 38393 14331
rect 38160 14300 38393 14328
rect 38160 14288 38166 14300
rect 38381 14297 38393 14300
rect 38427 14297 38439 14331
rect 38381 14291 38439 14297
rect 40589 14331 40647 14337
rect 40589 14297 40601 14331
rect 40635 14297 40647 14331
rect 40589 14291 40647 14297
rect 40773 14331 40831 14337
rect 40773 14297 40785 14331
rect 40819 14328 40831 14331
rect 41064 14328 41092 14504
rect 43714 14464 43720 14476
rect 43180 14436 43720 14464
rect 43180 14405 43208 14436
rect 43714 14424 43720 14436
rect 43772 14424 43778 14476
rect 41141 14399 41199 14405
rect 41141 14365 41153 14399
rect 41187 14396 41199 14399
rect 41693 14399 41751 14405
rect 41693 14396 41705 14399
rect 41187 14368 41705 14396
rect 41187 14365 41199 14368
rect 41141 14359 41199 14365
rect 41693 14365 41705 14368
rect 41739 14365 41751 14399
rect 41693 14359 41751 14365
rect 43165 14399 43223 14405
rect 43165 14365 43177 14399
rect 43211 14365 43223 14399
rect 43165 14359 43223 14365
rect 43533 14399 43591 14405
rect 43533 14365 43545 14399
rect 43579 14396 43591 14399
rect 45186 14396 45192 14408
rect 43579 14368 45192 14396
rect 43579 14365 43591 14368
rect 43533 14359 43591 14365
rect 40819 14300 41092 14328
rect 41708 14328 41736 14359
rect 43548 14328 43576 14359
rect 45186 14356 45192 14368
rect 45244 14356 45250 14408
rect 41708 14300 43576 14328
rect 40819 14297 40831 14300
rect 40773 14291 40831 14297
rect 38470 14260 38476 14272
rect 38028 14232 38476 14260
rect 38470 14220 38476 14232
rect 38528 14260 38534 14272
rect 40494 14260 40500 14272
rect 38528 14232 40500 14260
rect 38528 14220 38534 14232
rect 40494 14220 40500 14232
rect 40552 14260 40558 14272
rect 40604 14260 40632 14291
rect 40552 14232 40632 14260
rect 40552 14220 40558 14232
rect 40678 14220 40684 14272
rect 40736 14260 40742 14272
rect 41601 14263 41659 14269
rect 41601 14260 41613 14263
rect 40736 14232 41613 14260
rect 40736 14220 40742 14232
rect 41601 14229 41613 14232
rect 41647 14229 41659 14263
rect 41601 14223 41659 14229
rect 43070 14220 43076 14272
rect 43128 14260 43134 14272
rect 43257 14263 43315 14269
rect 43257 14260 43269 14263
rect 43128 14232 43269 14260
rect 43128 14220 43134 14232
rect 43257 14229 43269 14232
rect 43303 14229 43315 14263
rect 43257 14223 43315 14229
rect 43993 14263 44051 14269
rect 43993 14229 44005 14263
rect 44039 14260 44051 14263
rect 44174 14260 44180 14272
rect 44039 14232 44180 14260
rect 44039 14229 44051 14232
rect 43993 14223 44051 14229
rect 44174 14220 44180 14232
rect 44232 14220 44238 14272
rect 1104 14170 47104 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 47104 14170
rect 1104 14096 47104 14118
rect 19702 14016 19708 14068
rect 19760 14056 19766 14068
rect 21085 14059 21143 14065
rect 21085 14056 21097 14059
rect 19760 14028 21097 14056
rect 19760 14016 19766 14028
rect 21085 14025 21097 14028
rect 21131 14056 21143 14059
rect 22094 14056 22100 14068
rect 21131 14028 22100 14056
rect 21131 14025 21143 14028
rect 21085 14019 21143 14025
rect 22094 14016 22100 14028
rect 22152 14016 22158 14068
rect 23382 14056 23388 14068
rect 22480 14028 23388 14056
rect 10226 13948 10232 14000
rect 10284 13948 10290 14000
rect 13265 13991 13323 13997
rect 13265 13957 13277 13991
rect 13311 13988 13323 13991
rect 13354 13988 13360 14000
rect 13311 13960 13360 13988
rect 13311 13957 13323 13960
rect 13265 13951 13323 13957
rect 13354 13948 13360 13960
rect 13412 13948 13418 14000
rect 14642 13948 14648 14000
rect 14700 13988 14706 14000
rect 14700 13960 15516 13988
rect 14700 13948 14706 13960
rect 7098 13880 7104 13932
rect 7156 13880 7162 13932
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13920 9551 13923
rect 9674 13920 9680 13932
rect 9539 13892 9680 13920
rect 9539 13889 9551 13892
rect 9493 13883 9551 13889
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 11054 13880 11060 13932
rect 11112 13920 11118 13932
rect 12529 13923 12587 13929
rect 12529 13920 12541 13923
rect 11112 13892 12541 13920
rect 11112 13880 11118 13892
rect 12529 13889 12541 13892
rect 12575 13889 12587 13923
rect 12529 13883 12587 13889
rect 12618 13880 12624 13932
rect 12676 13920 12682 13932
rect 13449 13923 13507 13929
rect 13449 13920 13461 13923
rect 12676 13892 13461 13920
rect 12676 13880 12682 13892
rect 13449 13889 13461 13892
rect 13495 13889 13507 13923
rect 13449 13883 13507 13889
rect 15286 13880 15292 13932
rect 15344 13880 15350 13932
rect 15488 13920 15516 13960
rect 19518 13948 19524 14000
rect 19576 13988 19582 14000
rect 19576 13960 20392 13988
rect 19576 13948 19582 13960
rect 19705 13923 19763 13929
rect 19705 13920 19717 13923
rect 15488 13892 19717 13920
rect 19705 13889 19717 13892
rect 19751 13920 19763 13923
rect 19794 13920 19800 13932
rect 19751 13892 19800 13920
rect 19751 13889 19763 13892
rect 19705 13883 19763 13889
rect 19794 13880 19800 13892
rect 19852 13880 19858 13932
rect 19972 13923 20030 13929
rect 19972 13889 19984 13923
rect 20018 13920 20030 13923
rect 20254 13920 20260 13932
rect 20018 13892 20260 13920
rect 20018 13889 20030 13892
rect 19972 13883 20030 13889
rect 20254 13880 20260 13892
rect 20312 13880 20318 13932
rect 20364 13920 20392 13960
rect 20438 13948 20444 14000
rect 20496 13988 20502 14000
rect 22480 13988 22508 14028
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 24762 14016 24768 14068
rect 24820 14056 24826 14068
rect 28813 14059 28871 14065
rect 28813 14056 28825 14059
rect 24820 14028 28825 14056
rect 24820 14016 24826 14028
rect 28813 14025 28825 14028
rect 28859 14025 28871 14059
rect 28813 14019 28871 14025
rect 31018 14016 31024 14068
rect 31076 14056 31082 14068
rect 31573 14059 31631 14065
rect 31573 14056 31585 14059
rect 31076 14028 31585 14056
rect 31076 14016 31082 14028
rect 31573 14025 31585 14028
rect 31619 14025 31631 14059
rect 31573 14019 31631 14025
rect 32125 14059 32183 14065
rect 32125 14025 32137 14059
rect 32171 14025 32183 14059
rect 32125 14019 32183 14025
rect 20496 13960 22508 13988
rect 22557 13991 22615 13997
rect 20496 13948 20502 13960
rect 22557 13957 22569 13991
rect 22603 13988 22615 13991
rect 22603 13960 23336 13988
rect 22603 13957 22615 13960
rect 22557 13951 22615 13957
rect 22572 13920 22600 13951
rect 20364 13892 22600 13920
rect 12161 13855 12219 13861
rect 12161 13821 12173 13855
rect 12207 13852 12219 13855
rect 12434 13852 12440 13864
rect 12207 13824 12440 13852
rect 12207 13821 12219 13824
rect 12161 13815 12219 13821
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12805 13855 12863 13861
rect 12805 13821 12817 13855
rect 12851 13852 12863 13855
rect 19242 13852 19248 13864
rect 12851 13824 19248 13852
rect 12851 13821 12863 13824
rect 12805 13815 12863 13821
rect 19242 13812 19248 13824
rect 19300 13812 19306 13864
rect 23308 13852 23336 13960
rect 23400 13929 23428 14016
rect 25406 13997 25412 14000
rect 25400 13988 25412 13997
rect 25367 13960 25412 13988
rect 25400 13951 25412 13960
rect 25406 13948 25412 13951
rect 25464 13948 25470 14000
rect 27154 13988 27160 14000
rect 26804 13960 27160 13988
rect 23385 13923 23443 13929
rect 23385 13889 23397 13923
rect 23431 13889 23443 13923
rect 23385 13883 23443 13889
rect 25133 13923 25191 13929
rect 25133 13889 25145 13923
rect 25179 13920 25191 13923
rect 26804 13920 26832 13960
rect 27154 13948 27160 13960
rect 27212 13948 27218 14000
rect 25179 13892 26832 13920
rect 25179 13889 25191 13892
rect 25133 13883 25191 13889
rect 26878 13880 26884 13932
rect 26936 13920 26942 13932
rect 26936 13892 27292 13920
rect 26936 13880 26942 13892
rect 25038 13852 25044 13864
rect 23308 13824 25044 13852
rect 25038 13812 25044 13824
rect 25096 13812 25102 13864
rect 26142 13812 26148 13864
rect 26200 13852 26206 13864
rect 26200 13824 26924 13852
rect 26200 13812 26206 13824
rect 7742 13744 7748 13796
rect 7800 13784 7806 13796
rect 8018 13784 8024 13796
rect 7800 13756 8024 13784
rect 7800 13744 7806 13756
rect 8018 13744 8024 13756
rect 8076 13784 8082 13796
rect 12710 13784 12716 13796
rect 8076 13756 12716 13784
rect 8076 13744 8082 13756
rect 12710 13744 12716 13756
rect 12768 13744 12774 13796
rect 22738 13744 22744 13796
rect 22796 13744 22802 13796
rect 26896 13784 26924 13824
rect 26970 13812 26976 13864
rect 27028 13812 27034 13864
rect 27154 13852 27160 13864
rect 27080 13824 27160 13852
rect 27080 13784 27108 13824
rect 27154 13812 27160 13824
rect 27212 13812 27218 13864
rect 27264 13852 27292 13892
rect 28166 13880 28172 13932
rect 28224 13880 28230 13932
rect 29270 13880 29276 13932
rect 29328 13880 29334 13932
rect 30650 13880 30656 13932
rect 30708 13880 30714 13932
rect 30742 13880 30748 13932
rect 30800 13929 30806 13932
rect 30800 13923 30828 13929
rect 30816 13889 30828 13923
rect 30800 13883 30828 13889
rect 30929 13923 30987 13929
rect 30929 13889 30941 13923
rect 30975 13889 30987 13923
rect 30929 13883 30987 13889
rect 31941 13923 31999 13929
rect 31941 13889 31953 13923
rect 31987 13920 31999 13923
rect 32140 13920 32168 14019
rect 32490 14016 32496 14068
rect 32548 14016 32554 14068
rect 35250 14016 35256 14068
rect 35308 14016 35314 14068
rect 35437 14059 35495 14065
rect 35437 14025 35449 14059
rect 35483 14025 35495 14059
rect 35437 14019 35495 14025
rect 35452 13988 35480 14019
rect 37642 14016 37648 14068
rect 37700 14016 37706 14068
rect 37737 14059 37795 14065
rect 37737 14025 37749 14059
rect 37783 14056 37795 14059
rect 37826 14056 37832 14068
rect 37783 14028 37832 14056
rect 37783 14025 37795 14028
rect 37737 14019 37795 14025
rect 37826 14016 37832 14028
rect 37884 14016 37890 14068
rect 40126 14016 40132 14068
rect 40184 14016 40190 14068
rect 40954 14016 40960 14068
rect 41012 14056 41018 14068
rect 41601 14059 41659 14065
rect 41601 14056 41613 14059
rect 41012 14028 41613 14056
rect 41012 14016 41018 14028
rect 41601 14025 41613 14028
rect 41647 14025 41659 14059
rect 41601 14019 41659 14025
rect 42978 14016 42984 14068
rect 43036 14016 43042 14068
rect 43993 14059 44051 14065
rect 43993 14025 44005 14059
rect 44039 14025 44051 14059
rect 43993 14019 44051 14025
rect 35958 13991 36016 13997
rect 35958 13988 35970 13991
rect 35452 13960 35970 13988
rect 35958 13957 35970 13960
rect 36004 13957 36016 13991
rect 35958 13951 36016 13957
rect 40494 13948 40500 14000
rect 40552 13988 40558 14000
rect 40552 13960 43392 13988
rect 40552 13948 40558 13960
rect 31987 13892 32168 13920
rect 32585 13923 32643 13929
rect 31987 13889 31999 13892
rect 31941 13883 31999 13889
rect 32585 13889 32597 13923
rect 32631 13920 32643 13923
rect 33226 13920 33232 13932
rect 32631 13892 33232 13920
rect 32631 13889 32643 13892
rect 32585 13883 32643 13889
rect 30800 13880 30806 13883
rect 27893 13855 27951 13861
rect 27893 13852 27905 13855
rect 27264 13824 27905 13852
rect 27893 13821 27905 13824
rect 27939 13821 27951 13855
rect 27893 13815 27951 13821
rect 27982 13812 27988 13864
rect 28040 13861 28046 13864
rect 28040 13855 28068 13861
rect 28056 13821 28068 13855
rect 28040 13815 28068 13821
rect 28040 13812 28046 13815
rect 28718 13812 28724 13864
rect 28776 13852 28782 13864
rect 29365 13855 29423 13861
rect 29365 13852 29377 13855
rect 28776 13824 29377 13852
rect 28776 13812 28782 13824
rect 29365 13821 29377 13824
rect 29411 13821 29423 13855
rect 29365 13815 29423 13821
rect 29549 13855 29607 13861
rect 29549 13821 29561 13855
rect 29595 13821 29607 13855
rect 29549 13815 29607 13821
rect 29733 13855 29791 13861
rect 29733 13821 29745 13855
rect 29779 13821 29791 13855
rect 29733 13815 29791 13821
rect 29917 13855 29975 13861
rect 29917 13821 29929 13855
rect 29963 13852 29975 13855
rect 30098 13852 30104 13864
rect 29963 13824 30104 13852
rect 29963 13821 29975 13824
rect 29917 13815 29975 13821
rect 26896 13756 27108 13784
rect 27617 13787 27675 13793
rect 27617 13753 27629 13787
rect 27663 13784 27675 13787
rect 27706 13784 27712 13796
rect 27663 13756 27712 13784
rect 27663 13753 27675 13756
rect 27617 13747 27675 13753
rect 27706 13744 27712 13756
rect 27764 13744 27770 13796
rect 29564 13784 29592 13815
rect 29638 13784 29644 13796
rect 29564 13756 29644 13784
rect 29638 13744 29644 13756
rect 29696 13744 29702 13796
rect 29748 13784 29776 13815
rect 30098 13812 30104 13824
rect 30156 13852 30162 13864
rect 30944 13852 30972 13883
rect 31110 13852 31116 13864
rect 30156 13824 30512 13852
rect 30944 13824 31116 13852
rect 30156 13812 30162 13824
rect 30006 13784 30012 13796
rect 29748 13756 30012 13784
rect 30006 13744 30012 13756
rect 30064 13744 30070 13796
rect 30374 13744 30380 13796
rect 30432 13744 30438 13796
rect 6914 13676 6920 13728
rect 6972 13676 6978 13728
rect 9306 13676 9312 13728
rect 9364 13676 9370 13728
rect 10318 13676 10324 13728
rect 10376 13676 10382 13728
rect 15010 13676 15016 13728
rect 15068 13716 15074 13728
rect 15105 13719 15163 13725
rect 15105 13716 15117 13719
rect 15068 13688 15117 13716
rect 15068 13676 15074 13688
rect 15105 13685 15117 13688
rect 15151 13685 15163 13719
rect 15105 13679 15163 13685
rect 23569 13719 23627 13725
rect 23569 13685 23581 13719
rect 23615 13716 23627 13719
rect 24578 13716 24584 13728
rect 23615 13688 24584 13716
rect 23615 13685 23627 13688
rect 23569 13679 23627 13685
rect 24578 13676 24584 13688
rect 24636 13676 24642 13728
rect 26510 13676 26516 13728
rect 26568 13716 26574 13728
rect 27062 13716 27068 13728
rect 26568 13688 27068 13716
rect 26568 13676 26574 13688
rect 27062 13676 27068 13688
rect 27120 13716 27126 13728
rect 27982 13716 27988 13728
rect 27120 13688 27988 13716
rect 27120 13676 27126 13688
rect 27982 13676 27988 13688
rect 28040 13676 28046 13728
rect 28902 13676 28908 13728
rect 28960 13676 28966 13728
rect 30484 13716 30512 13824
rect 31110 13812 31116 13824
rect 31168 13812 31174 13864
rect 32600 13852 32628 13883
rect 33226 13880 33232 13892
rect 33284 13880 33290 13932
rect 33318 13880 33324 13932
rect 33376 13920 33382 13932
rect 33376 13892 33732 13920
rect 33376 13880 33382 13892
rect 31312 13824 32628 13852
rect 31312 13716 31340 13824
rect 32674 13812 32680 13864
rect 32732 13812 32738 13864
rect 33413 13855 33471 13861
rect 33413 13821 33425 13855
rect 33459 13821 33471 13855
rect 33413 13815 33471 13821
rect 33428 13784 33456 13815
rect 33502 13812 33508 13864
rect 33560 13852 33566 13864
rect 33597 13855 33655 13861
rect 33597 13852 33609 13855
rect 33560 13824 33609 13852
rect 33560 13812 33566 13824
rect 33597 13821 33609 13824
rect 33643 13821 33655 13855
rect 33704 13852 33732 13892
rect 34606 13880 34612 13932
rect 34664 13880 34670 13932
rect 35621 13923 35679 13929
rect 35621 13889 35633 13923
rect 35667 13920 35679 13923
rect 36262 13920 36268 13932
rect 35667 13892 36268 13920
rect 35667 13889 35679 13892
rect 35621 13883 35679 13889
rect 36262 13880 36268 13892
rect 36320 13880 36326 13932
rect 40313 13923 40371 13929
rect 40313 13889 40325 13923
rect 40359 13920 40371 13923
rect 40678 13920 40684 13932
rect 40359 13892 40684 13920
rect 40359 13889 40371 13892
rect 40313 13883 40371 13889
rect 40678 13880 40684 13892
rect 40736 13880 40742 13932
rect 41138 13880 41144 13932
rect 41196 13880 41202 13932
rect 42242 13880 42248 13932
rect 42300 13920 42306 13932
rect 42797 13923 42855 13929
rect 42797 13920 42809 13923
rect 42300 13892 42809 13920
rect 42300 13880 42306 13892
rect 42797 13889 42809 13892
rect 42843 13889 42855 13923
rect 42797 13883 42855 13889
rect 43070 13880 43076 13932
rect 43128 13880 43134 13932
rect 33962 13852 33968 13864
rect 33704 13824 33968 13852
rect 33597 13815 33655 13821
rect 33962 13812 33968 13824
rect 34020 13852 34026 13864
rect 34057 13855 34115 13861
rect 34057 13852 34069 13855
rect 34020 13824 34069 13852
rect 34020 13812 34026 13824
rect 34057 13821 34069 13824
rect 34103 13821 34115 13855
rect 34057 13815 34115 13821
rect 34146 13812 34152 13864
rect 34204 13852 34210 13864
rect 34333 13855 34391 13861
rect 34333 13852 34345 13855
rect 34204 13824 34345 13852
rect 34204 13812 34210 13824
rect 34333 13821 34345 13824
rect 34379 13821 34391 13855
rect 34333 13815 34391 13821
rect 34422 13812 34428 13864
rect 34480 13861 34486 13864
rect 34480 13855 34508 13861
rect 34496 13821 34508 13855
rect 34480 13815 34508 13821
rect 34480 13812 34486 13815
rect 35710 13812 35716 13864
rect 35768 13812 35774 13864
rect 37829 13855 37887 13861
rect 37829 13821 37841 13855
rect 37875 13821 37887 13855
rect 37829 13815 37887 13821
rect 33870 13784 33876 13796
rect 33428 13756 33876 13784
rect 33870 13744 33876 13756
rect 33928 13744 33934 13796
rect 36998 13744 37004 13796
rect 37056 13784 37062 13796
rect 37844 13784 37872 13815
rect 40954 13812 40960 13864
rect 41012 13812 41018 13864
rect 43162 13812 43168 13864
rect 43220 13852 43226 13864
rect 43257 13855 43315 13861
rect 43257 13852 43269 13855
rect 43220 13824 43269 13852
rect 43220 13812 43226 13824
rect 43257 13821 43269 13824
rect 43303 13821 43315 13855
rect 43364 13852 43392 13960
rect 43441 13923 43499 13929
rect 43441 13889 43453 13923
rect 43487 13920 43499 13923
rect 44008 13920 44036 14019
rect 43487 13892 44036 13920
rect 43487 13889 43499 13892
rect 43441 13883 43499 13889
rect 44174 13880 44180 13932
rect 44232 13880 44238 13932
rect 45005 13923 45063 13929
rect 45005 13889 45017 13923
rect 45051 13920 45063 13923
rect 45186 13920 45192 13932
rect 45051 13892 45192 13920
rect 45051 13889 45063 13892
rect 45005 13883 45063 13889
rect 45186 13880 45192 13892
rect 45244 13880 45250 13932
rect 46842 13852 46848 13864
rect 43364 13824 46848 13852
rect 43257 13815 43315 13821
rect 46842 13812 46848 13824
rect 46900 13812 46906 13864
rect 37056 13756 37872 13784
rect 37056 13744 37062 13756
rect 30484 13688 31340 13716
rect 31757 13719 31815 13725
rect 31757 13685 31769 13719
rect 31803 13716 31815 13719
rect 31938 13716 31944 13728
rect 31803 13688 31944 13716
rect 31803 13685 31815 13688
rect 31757 13679 31815 13685
rect 31938 13676 31944 13688
rect 31996 13676 32002 13728
rect 33410 13676 33416 13728
rect 33468 13716 33474 13728
rect 35342 13716 35348 13728
rect 33468 13688 35348 13716
rect 33468 13676 33474 13688
rect 35342 13676 35348 13688
rect 35400 13676 35406 13728
rect 37090 13676 37096 13728
rect 37148 13676 37154 13728
rect 37274 13676 37280 13728
rect 37332 13676 37338 13728
rect 42794 13676 42800 13728
rect 42852 13676 42858 13728
rect 43254 13676 43260 13728
rect 43312 13716 43318 13728
rect 43625 13719 43683 13725
rect 43625 13716 43637 13719
rect 43312 13688 43637 13716
rect 43312 13676 43318 13688
rect 43625 13685 43637 13688
rect 43671 13685 43683 13719
rect 43625 13679 43683 13685
rect 45281 13719 45339 13725
rect 45281 13685 45293 13719
rect 45327 13716 45339 13719
rect 45370 13716 45376 13728
rect 45327 13688 45376 13716
rect 45327 13685 45339 13688
rect 45281 13679 45339 13685
rect 45370 13676 45376 13688
rect 45428 13676 45434 13728
rect 45462 13676 45468 13728
rect 45520 13676 45526 13728
rect 1104 13626 47104 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 47104 13626
rect 1104 13552 47104 13574
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 6472 13484 9045 13512
rect 6472 13385 6500 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 9033 13475 9091 13481
rect 6457 13379 6515 13385
rect 6457 13345 6469 13379
rect 6503 13345 6515 13379
rect 6457 13339 6515 13345
rect 8938 13336 8944 13388
rect 8996 13376 9002 13388
rect 9048 13376 9076 13475
rect 17770 13472 17776 13524
rect 17828 13512 17834 13524
rect 18690 13512 18696 13524
rect 17828 13484 18696 13512
rect 17828 13472 17834 13484
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 20254 13472 20260 13524
rect 20312 13472 20318 13524
rect 20898 13472 20904 13524
rect 20956 13512 20962 13524
rect 21358 13512 21364 13524
rect 20956 13484 21364 13512
rect 20956 13472 20962 13484
rect 21358 13472 21364 13484
rect 21416 13512 21422 13524
rect 21453 13515 21511 13521
rect 21453 13512 21465 13515
rect 21416 13484 21465 13512
rect 21416 13472 21422 13484
rect 21453 13481 21465 13484
rect 21499 13481 21511 13515
rect 21453 13475 21511 13481
rect 22066 13484 23980 13512
rect 14642 13404 14648 13456
rect 14700 13404 14706 13456
rect 20717 13447 20775 13453
rect 20717 13413 20729 13447
rect 20763 13444 20775 13447
rect 22066 13444 22094 13484
rect 20763 13416 22094 13444
rect 23952 13444 23980 13484
rect 24210 13472 24216 13524
rect 24268 13472 24274 13524
rect 25501 13515 25559 13521
rect 25501 13481 25513 13515
rect 25547 13512 25559 13515
rect 25590 13512 25596 13524
rect 25547 13484 25596 13512
rect 25547 13481 25559 13484
rect 25501 13475 25559 13481
rect 25590 13472 25596 13484
rect 25648 13472 25654 13524
rect 27154 13472 27160 13524
rect 27212 13512 27218 13524
rect 28718 13512 28724 13524
rect 27212 13484 28724 13512
rect 27212 13472 27218 13484
rect 28718 13472 28724 13484
rect 28776 13512 28782 13524
rect 28813 13515 28871 13521
rect 28813 13512 28825 13515
rect 28776 13484 28825 13512
rect 28776 13472 28782 13484
rect 28813 13481 28825 13484
rect 28859 13481 28871 13515
rect 28813 13475 28871 13481
rect 29638 13472 29644 13524
rect 29696 13512 29702 13524
rect 31018 13512 31024 13524
rect 29696 13484 31024 13512
rect 29696 13472 29702 13484
rect 31018 13472 31024 13484
rect 31076 13472 31082 13524
rect 31757 13515 31815 13521
rect 31757 13481 31769 13515
rect 31803 13512 31815 13515
rect 31846 13512 31852 13524
rect 31803 13484 31852 13512
rect 31803 13481 31815 13484
rect 31757 13475 31815 13481
rect 31846 13472 31852 13484
rect 31904 13472 31910 13524
rect 33226 13472 33232 13524
rect 33284 13472 33290 13524
rect 36173 13515 36231 13521
rect 33428 13484 35756 13512
rect 26326 13444 26332 13456
rect 23952 13416 26332 13444
rect 20763 13413 20775 13416
rect 20717 13407 20775 13413
rect 26326 13404 26332 13416
rect 26384 13404 26390 13456
rect 27430 13444 27436 13456
rect 27356 13416 27436 13444
rect 9309 13379 9367 13385
rect 9309 13376 9321 13379
rect 8996 13348 9321 13376
rect 8996 13336 9002 13348
rect 9309 13345 9321 13348
rect 9355 13345 9367 13379
rect 9309 13339 9367 13345
rect 14274 13336 14280 13388
rect 14332 13376 14338 13388
rect 14660 13376 14688 13404
rect 14737 13379 14795 13385
rect 14737 13376 14749 13379
rect 14332 13348 14749 13376
rect 14332 13336 14338 13348
rect 14737 13345 14749 13348
rect 14783 13345 14795 13379
rect 21726 13376 21732 13388
rect 14737 13339 14795 13345
rect 20456 13348 21732 13376
rect 4430 13268 4436 13320
rect 4488 13268 4494 13320
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 10318 13308 10324 13320
rect 9263 13280 10324 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 10965 13311 11023 13317
rect 10965 13308 10977 13311
rect 10468 13280 10977 13308
rect 10468 13268 10474 13280
rect 10965 13277 10977 13280
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 11698 13268 11704 13320
rect 11756 13268 11762 13320
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13308 11851 13311
rect 14292 13308 14320 13336
rect 11839 13280 14320 13308
rect 11839 13277 11851 13280
rect 11793 13271 11851 13277
rect 14642 13268 14648 13320
rect 14700 13268 14706 13320
rect 15010 13317 15016 13320
rect 15004 13308 15016 13317
rect 14971 13280 15016 13308
rect 15004 13271 15016 13280
rect 15010 13268 15016 13271
rect 15068 13268 15074 13320
rect 16666 13268 16672 13320
rect 16724 13308 16730 13320
rect 16853 13311 16911 13317
rect 16853 13308 16865 13311
rect 16724 13280 16865 13308
rect 16724 13268 16730 13280
rect 16853 13277 16865 13280
rect 16899 13308 16911 13311
rect 20070 13308 20076 13320
rect 16899 13280 20076 13308
rect 16899 13277 16911 13280
rect 16853 13271 16911 13277
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 20456 13317 20484 13348
rect 21726 13336 21732 13348
rect 21784 13336 21790 13388
rect 23017 13379 23075 13385
rect 23017 13376 23029 13379
rect 22066 13348 23029 13376
rect 20441 13311 20499 13317
rect 20441 13277 20453 13311
rect 20487 13277 20499 13311
rect 20441 13271 20499 13277
rect 20898 13268 20904 13320
rect 20956 13268 20962 13320
rect 21174 13268 21180 13320
rect 21232 13308 21238 13320
rect 21910 13308 21916 13320
rect 21232 13280 21916 13308
rect 21232 13268 21238 13280
rect 21910 13268 21916 13280
rect 21968 13268 21974 13320
rect 6724 13243 6782 13249
rect 6724 13209 6736 13243
rect 6770 13240 6782 13243
rect 6914 13240 6920 13252
rect 6770 13212 6920 13240
rect 6770 13209 6782 13212
rect 6724 13203 6782 13209
rect 6914 13200 6920 13212
rect 6972 13200 6978 13252
rect 9576 13243 9634 13249
rect 9576 13209 9588 13243
rect 9622 13240 9634 13243
rect 12038 13243 12096 13249
rect 12038 13240 12050 13243
rect 9622 13212 10824 13240
rect 9622 13209 9634 13212
rect 9576 13203 9634 13209
rect 4246 13132 4252 13184
rect 4304 13132 4310 13184
rect 6546 13132 6552 13184
rect 6604 13172 6610 13184
rect 7834 13172 7840 13184
rect 6604 13144 7840 13172
rect 6604 13132 6610 13144
rect 7834 13132 7840 13144
rect 7892 13132 7898 13184
rect 10686 13132 10692 13184
rect 10744 13132 10750 13184
rect 10796 13181 10824 13212
rect 11532 13212 12050 13240
rect 11532 13181 11560 13212
rect 12038 13209 12050 13212
rect 12084 13209 12096 13243
rect 12038 13203 12096 13209
rect 16942 13200 16948 13252
rect 17000 13240 17006 13252
rect 17098 13243 17156 13249
rect 17098 13240 17110 13243
rect 17000 13212 17110 13240
rect 17000 13200 17006 13212
rect 17098 13209 17110 13212
rect 17144 13209 17156 13243
rect 18138 13240 18144 13252
rect 17098 13203 17156 13209
rect 17236 13212 18144 13240
rect 10781 13175 10839 13181
rect 10781 13141 10793 13175
rect 10827 13141 10839 13175
rect 10781 13135 10839 13141
rect 11517 13175 11575 13181
rect 11517 13141 11529 13175
rect 11563 13141 11575 13175
rect 11517 13135 11575 13141
rect 11882 13132 11888 13184
rect 11940 13172 11946 13184
rect 13173 13175 13231 13181
rect 13173 13172 13185 13175
rect 11940 13144 13185 13172
rect 11940 13132 11946 13144
rect 13173 13141 13185 13144
rect 13219 13172 13231 13175
rect 13814 13172 13820 13184
rect 13219 13144 13820 13172
rect 13219 13141 13231 13144
rect 13173 13135 13231 13141
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 14461 13175 14519 13181
rect 14461 13141 14473 13175
rect 14507 13172 14519 13175
rect 14550 13172 14556 13184
rect 14507 13144 14556 13172
rect 14507 13141 14519 13144
rect 14461 13135 14519 13141
rect 14550 13132 14556 13144
rect 14608 13132 14614 13184
rect 16114 13132 16120 13184
rect 16172 13172 16178 13184
rect 17236 13172 17264 13212
rect 18138 13200 18144 13212
rect 18196 13200 18202 13252
rect 20622 13200 20628 13252
rect 20680 13240 20686 13252
rect 21361 13243 21419 13249
rect 20680 13212 21220 13240
rect 20680 13200 20686 13212
rect 16172 13144 17264 13172
rect 16172 13132 16178 13144
rect 17310 13132 17316 13184
rect 17368 13172 17374 13184
rect 18233 13175 18291 13181
rect 18233 13172 18245 13175
rect 17368 13144 18245 13172
rect 17368 13132 17374 13144
rect 18233 13141 18245 13144
rect 18279 13172 18291 13175
rect 19150 13172 19156 13184
rect 18279 13144 19156 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 19150 13132 19156 13144
rect 19208 13132 19214 13184
rect 21082 13132 21088 13184
rect 21140 13132 21146 13184
rect 21192 13172 21220 13212
rect 21361 13209 21373 13243
rect 21407 13240 21419 13243
rect 21634 13240 21640 13252
rect 21407 13212 21640 13240
rect 21407 13209 21419 13212
rect 21361 13203 21419 13209
rect 21634 13200 21640 13212
rect 21692 13200 21698 13252
rect 22066 13172 22094 13348
rect 23017 13345 23029 13348
rect 23063 13345 23075 13379
rect 23017 13339 23075 13345
rect 23566 13336 23572 13388
rect 23624 13336 23630 13388
rect 24670 13336 24676 13388
rect 24728 13376 24734 13388
rect 25041 13379 25099 13385
rect 25041 13376 25053 13379
rect 24728 13348 25053 13376
rect 24728 13336 24734 13348
rect 25041 13345 25053 13348
rect 25087 13376 25099 13379
rect 25958 13376 25964 13388
rect 25087 13348 25964 13376
rect 25087 13345 25099 13348
rect 25041 13339 25099 13345
rect 25958 13336 25964 13348
rect 26016 13336 26022 13388
rect 26145 13379 26203 13385
rect 26145 13345 26157 13379
rect 26191 13376 26203 13379
rect 26694 13376 26700 13388
rect 26191 13348 26700 13376
rect 26191 13345 26203 13348
rect 26145 13339 26203 13345
rect 26694 13336 26700 13348
rect 26752 13336 26758 13388
rect 22373 13311 22431 13317
rect 22373 13277 22385 13311
rect 22419 13277 22431 13311
rect 22373 13271 22431 13277
rect 21192 13144 22094 13172
rect 22388 13172 22416 13271
rect 22554 13268 22560 13320
rect 22612 13268 22618 13320
rect 23290 13268 23296 13320
rect 23348 13268 23354 13320
rect 23382 13268 23388 13320
rect 23440 13317 23446 13320
rect 23440 13311 23468 13317
rect 23456 13277 23468 13311
rect 23440 13271 23468 13277
rect 24857 13311 24915 13317
rect 24857 13277 24869 13311
rect 24903 13308 24915 13311
rect 25498 13308 25504 13320
rect 24903 13280 25504 13308
rect 24903 13277 24915 13280
rect 24857 13271 24915 13277
rect 23440 13268 23446 13271
rect 25498 13268 25504 13280
rect 25556 13268 25562 13320
rect 25869 13311 25927 13317
rect 25869 13277 25881 13311
rect 25915 13308 25927 13311
rect 26510 13308 26516 13320
rect 25915 13280 26516 13308
rect 25915 13277 25927 13280
rect 25869 13271 25927 13277
rect 26510 13268 26516 13280
rect 26568 13268 26574 13320
rect 24044 13212 24808 13240
rect 23014 13172 23020 13184
rect 22388 13144 23020 13172
rect 23014 13132 23020 13144
rect 23072 13172 23078 13184
rect 24044 13172 24072 13212
rect 23072 13144 24072 13172
rect 24397 13175 24455 13181
rect 23072 13132 23078 13144
rect 24397 13141 24409 13175
rect 24443 13172 24455 13175
rect 24670 13172 24676 13184
rect 24443 13144 24676 13172
rect 24443 13141 24455 13144
rect 24397 13135 24455 13141
rect 24670 13132 24676 13144
rect 24728 13132 24734 13184
rect 24780 13181 24808 13212
rect 25038 13200 25044 13252
rect 25096 13240 25102 13252
rect 25961 13243 26019 13249
rect 25961 13240 25973 13243
rect 25096 13212 25973 13240
rect 25096 13200 25102 13212
rect 25961 13209 25973 13212
rect 26007 13240 26019 13243
rect 27356 13240 27384 13416
rect 27430 13404 27436 13416
rect 27488 13404 27494 13456
rect 29089 13447 29147 13453
rect 29089 13413 29101 13447
rect 29135 13444 29147 13447
rect 29546 13444 29552 13456
rect 29135 13416 29552 13444
rect 29135 13413 29147 13416
rect 29089 13407 29147 13413
rect 29546 13404 29552 13416
rect 29604 13404 29610 13456
rect 30282 13404 30288 13456
rect 30340 13444 30346 13456
rect 30561 13447 30619 13453
rect 30561 13444 30573 13447
rect 30340 13416 30573 13444
rect 30340 13404 30346 13416
rect 30561 13413 30573 13416
rect 30607 13413 30619 13447
rect 30561 13407 30619 13413
rect 33134 13404 33140 13456
rect 33192 13444 33198 13456
rect 33428 13444 33456 13484
rect 33192 13416 33456 13444
rect 33505 13447 33563 13453
rect 33192 13404 33198 13416
rect 33505 13413 33517 13447
rect 33551 13444 33563 13447
rect 33551 13416 34744 13444
rect 33551 13413 33563 13416
rect 33505 13407 33563 13413
rect 29822 13376 29828 13388
rect 28460 13348 29828 13376
rect 27433 13311 27491 13317
rect 27433 13277 27445 13311
rect 27479 13308 27491 13311
rect 27522 13308 27528 13320
rect 27479 13280 27528 13308
rect 27479 13277 27491 13280
rect 27433 13271 27491 13277
rect 27522 13268 27528 13280
rect 27580 13268 27586 13320
rect 28460 13308 28488 13348
rect 29822 13336 29828 13348
rect 29880 13336 29886 13388
rect 30098 13336 30104 13388
rect 30156 13336 30162 13388
rect 30650 13336 30656 13388
rect 30708 13376 30714 13388
rect 30837 13379 30895 13385
rect 30837 13376 30849 13379
rect 30708 13348 30849 13376
rect 30708 13336 30714 13348
rect 30837 13345 30849 13348
rect 30883 13345 30895 13379
rect 30837 13339 30895 13345
rect 30926 13336 30932 13388
rect 30984 13385 30990 13388
rect 30984 13379 31012 13385
rect 31000 13345 31012 13379
rect 30984 13339 31012 13345
rect 31113 13379 31171 13385
rect 31113 13345 31125 13379
rect 31159 13376 31171 13379
rect 31294 13376 31300 13388
rect 31159 13348 31300 13376
rect 31159 13345 31171 13348
rect 31113 13339 31171 13345
rect 30984 13336 30990 13339
rect 31294 13336 31300 13348
rect 31352 13336 31358 13388
rect 31662 13336 31668 13388
rect 31720 13376 31726 13388
rect 31849 13379 31907 13385
rect 31849 13376 31861 13379
rect 31720 13348 31861 13376
rect 31720 13336 31726 13348
rect 27632 13280 28488 13308
rect 29273 13311 29331 13317
rect 27632 13240 27660 13280
rect 29273 13277 29285 13311
rect 29319 13308 29331 13311
rect 29917 13311 29975 13317
rect 29319 13280 29868 13308
rect 29319 13277 29331 13280
rect 29273 13271 29331 13277
rect 27706 13249 27712 13252
rect 26007 13212 27660 13240
rect 26007 13209 26019 13212
rect 25961 13203 26019 13209
rect 27700 13203 27712 13249
rect 27706 13200 27712 13203
rect 27764 13200 27770 13252
rect 24765 13175 24823 13181
rect 24765 13141 24777 13175
rect 24811 13172 24823 13175
rect 25774 13172 25780 13184
rect 24811 13144 25780 13172
rect 24811 13141 24823 13144
rect 24765 13135 24823 13141
rect 25774 13132 25780 13144
rect 25832 13132 25838 13184
rect 26326 13132 26332 13184
rect 26384 13172 26390 13184
rect 28718 13172 28724 13184
rect 26384 13144 28724 13172
rect 26384 13132 26390 13144
rect 28718 13132 28724 13144
rect 28776 13132 28782 13184
rect 29840 13172 29868 13280
rect 29917 13277 29929 13311
rect 29963 13308 29975 13311
rect 30006 13308 30012 13320
rect 29963 13280 30012 13308
rect 29963 13277 29975 13280
rect 29917 13271 29975 13277
rect 30006 13268 30012 13280
rect 30064 13268 30070 13320
rect 31772 13240 31800 13348
rect 31849 13345 31861 13348
rect 31895 13345 31907 13379
rect 31849 13339 31907 13345
rect 33040 13348 33916 13376
rect 31938 13268 31944 13320
rect 31996 13308 32002 13320
rect 32105 13311 32163 13317
rect 32105 13308 32117 13311
rect 31996 13280 32117 13308
rect 31996 13268 32002 13280
rect 32105 13277 32117 13280
rect 32151 13277 32163 13311
rect 32105 13271 32163 13277
rect 33040 13240 33068 13348
rect 33689 13311 33747 13317
rect 33689 13277 33701 13311
rect 33735 13308 33747 13311
rect 33888 13308 33916 13348
rect 34238 13336 34244 13388
rect 34296 13336 34302 13388
rect 34330 13336 34336 13388
rect 34388 13336 34394 13388
rect 34716 13376 34744 13416
rect 34716 13348 34836 13376
rect 34701 13311 34759 13317
rect 34701 13308 34713 13311
rect 33735 13280 33824 13308
rect 33888 13280 34713 13308
rect 33735 13277 33747 13280
rect 33689 13271 33747 13277
rect 31772 13212 33068 13240
rect 33410 13172 33416 13184
rect 29840 13144 33416 13172
rect 33410 13132 33416 13144
rect 33468 13132 33474 13184
rect 33796 13181 33824 13280
rect 34701 13277 34713 13280
rect 34747 13277 34759 13311
rect 34808 13308 34836 13348
rect 34957 13311 35015 13317
rect 34957 13308 34969 13311
rect 34808 13280 34969 13308
rect 34701 13271 34759 13277
rect 34957 13277 34969 13280
rect 35003 13277 35015 13311
rect 35728 13308 35756 13484
rect 36173 13481 36185 13515
rect 36219 13512 36231 13515
rect 36262 13512 36268 13524
rect 36219 13484 36268 13512
rect 36219 13481 36231 13484
rect 36173 13475 36231 13481
rect 36262 13472 36268 13484
rect 36320 13472 36326 13524
rect 36354 13472 36360 13524
rect 36412 13512 36418 13524
rect 46106 13512 46112 13524
rect 36412 13484 46112 13512
rect 36412 13472 36418 13484
rect 46106 13472 46112 13484
rect 46164 13472 46170 13524
rect 42981 13447 43039 13453
rect 42981 13413 42993 13447
rect 43027 13444 43039 13447
rect 43714 13444 43720 13456
rect 43027 13416 43720 13444
rect 43027 13413 43039 13416
rect 42981 13407 43039 13413
rect 43714 13404 43720 13416
rect 43772 13404 43778 13456
rect 36817 13379 36875 13385
rect 36817 13345 36829 13379
rect 36863 13376 36875 13379
rect 36998 13376 37004 13388
rect 36863 13348 37004 13376
rect 36863 13345 36875 13348
rect 36817 13339 36875 13345
rect 36998 13336 37004 13348
rect 37056 13336 37062 13388
rect 36541 13311 36599 13317
rect 36541 13308 36553 13311
rect 35728 13280 36553 13308
rect 34957 13271 35015 13277
rect 36541 13277 36553 13280
rect 36587 13308 36599 13311
rect 37090 13308 37096 13320
rect 36587 13280 37096 13308
rect 36587 13277 36599 13280
rect 36541 13271 36599 13277
rect 37090 13268 37096 13280
rect 37148 13268 37154 13320
rect 37369 13311 37427 13317
rect 37369 13277 37381 13311
rect 37415 13308 37427 13311
rect 37550 13308 37556 13320
rect 37415 13280 37556 13308
rect 37415 13277 37427 13280
rect 37369 13271 37427 13277
rect 37550 13268 37556 13280
rect 37608 13308 37614 13320
rect 38378 13308 38384 13320
rect 37608 13280 38384 13308
rect 37608 13268 37614 13280
rect 38378 13268 38384 13280
rect 38436 13268 38442 13320
rect 42518 13268 42524 13320
rect 42576 13308 42582 13320
rect 43165 13311 43223 13317
rect 43165 13308 43177 13311
rect 42576 13280 43177 13308
rect 42576 13268 42582 13280
rect 43165 13277 43177 13280
rect 43211 13277 43223 13311
rect 43165 13271 43223 13277
rect 43254 13268 43260 13320
rect 43312 13268 43318 13320
rect 45462 13268 45468 13320
rect 45520 13268 45526 13320
rect 46198 13268 46204 13320
rect 46256 13308 46262 13320
rect 46477 13311 46535 13317
rect 46477 13308 46489 13311
rect 46256 13280 46489 13308
rect 46256 13268 46262 13280
rect 46477 13277 46489 13280
rect 46523 13277 46535 13311
rect 46477 13271 46535 13277
rect 33870 13200 33876 13252
rect 33928 13240 33934 13252
rect 34149 13243 34207 13249
rect 34149 13240 34161 13243
rect 33928 13212 34161 13240
rect 33928 13200 33934 13212
rect 34149 13209 34161 13212
rect 34195 13240 34207 13243
rect 38010 13240 38016 13252
rect 34195 13212 36124 13240
rect 34195 13209 34207 13212
rect 34149 13203 34207 13209
rect 33781 13175 33839 13181
rect 33781 13141 33793 13175
rect 33827 13141 33839 13175
rect 33781 13135 33839 13141
rect 33962 13132 33968 13184
rect 34020 13172 34026 13184
rect 34330 13172 34336 13184
rect 34020 13144 34336 13172
rect 34020 13132 34026 13144
rect 34330 13132 34336 13144
rect 34388 13132 34394 13184
rect 36096 13181 36124 13212
rect 36648 13212 38016 13240
rect 36648 13184 36676 13212
rect 38010 13200 38016 13212
rect 38068 13200 38074 13252
rect 42981 13243 43039 13249
rect 42981 13209 42993 13243
rect 43027 13209 43039 13243
rect 42981 13203 43039 13209
rect 36081 13175 36139 13181
rect 36081 13141 36093 13175
rect 36127 13141 36139 13175
rect 36081 13135 36139 13141
rect 36630 13132 36636 13184
rect 36688 13132 36694 13184
rect 37458 13132 37464 13184
rect 37516 13132 37522 13184
rect 42996 13172 43024 13203
rect 43070 13172 43076 13184
rect 42996 13144 43076 13172
rect 43070 13132 43076 13144
rect 43128 13172 43134 13184
rect 43254 13172 43260 13184
rect 43128 13144 43260 13172
rect 43128 13132 43134 13144
rect 43254 13132 43260 13144
rect 43312 13132 43318 13184
rect 45094 13132 45100 13184
rect 45152 13172 45158 13184
rect 45281 13175 45339 13181
rect 45281 13172 45293 13175
rect 45152 13144 45293 13172
rect 45152 13132 45158 13144
rect 45281 13141 45293 13144
rect 45327 13141 45339 13175
rect 45281 13135 45339 13141
rect 46658 13132 46664 13184
rect 46716 13132 46722 13184
rect 1104 13082 47104 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 47104 13082
rect 1104 13008 47104 13030
rect 4430 12928 4436 12980
rect 4488 12968 4494 12980
rect 5169 12971 5227 12977
rect 5169 12968 5181 12971
rect 4488 12940 5181 12968
rect 4488 12928 4494 12940
rect 5169 12937 5181 12940
rect 5215 12937 5227 12971
rect 5169 12931 5227 12937
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 9858 12968 9864 12980
rect 7708 12940 9864 12968
rect 7708 12928 7714 12940
rect 9858 12928 9864 12940
rect 9916 12968 9922 12980
rect 9916 12940 9996 12968
rect 9916 12928 9922 12940
rect 3964 12903 4022 12909
rect 3964 12869 3976 12903
rect 4010 12900 4022 12903
rect 4246 12900 4252 12912
rect 4010 12872 4252 12900
rect 4010 12869 4022 12872
rect 3964 12863 4022 12869
rect 4246 12860 4252 12872
rect 4304 12860 4310 12912
rect 6270 12900 6276 12912
rect 5920 12872 6276 12900
rect 1486 12792 1492 12844
rect 1544 12792 1550 12844
rect 5537 12835 5595 12841
rect 5537 12801 5549 12835
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 1670 12724 1676 12776
rect 1728 12724 1734 12776
rect 3694 12724 3700 12776
rect 3752 12724 3758 12776
rect 5077 12699 5135 12705
rect 5077 12665 5089 12699
rect 5123 12696 5135 12699
rect 5552 12696 5580 12795
rect 5626 12724 5632 12776
rect 5684 12724 5690 12776
rect 5813 12767 5871 12773
rect 5813 12733 5825 12767
rect 5859 12764 5871 12767
rect 5920 12764 5948 12872
rect 6270 12860 6276 12872
rect 6328 12900 6334 12912
rect 6454 12900 6460 12912
rect 6328 12872 6460 12900
rect 6328 12860 6334 12872
rect 6454 12860 6460 12872
rect 6512 12860 6518 12912
rect 9208 12903 9266 12909
rect 9208 12869 9220 12903
rect 9254 12900 9266 12903
rect 9306 12900 9312 12912
rect 9254 12872 9312 12900
rect 9254 12869 9266 12872
rect 9208 12863 9266 12869
rect 9306 12860 9312 12872
rect 9364 12860 9370 12912
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12832 6423 12835
rect 6730 12832 6736 12844
rect 6411 12804 6736 12832
rect 6411 12801 6423 12804
rect 6365 12795 6423 12801
rect 6730 12792 6736 12804
rect 6788 12792 6794 12844
rect 8938 12792 8944 12844
rect 8996 12792 9002 12844
rect 5859 12736 5948 12764
rect 5859 12733 5871 12736
rect 5813 12727 5871 12733
rect 5994 12724 6000 12776
rect 6052 12764 6058 12776
rect 6546 12764 6552 12776
rect 6052 12736 6552 12764
rect 6052 12724 6058 12736
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 6886 12736 7297 12764
rect 6886 12696 6914 12736
rect 7285 12733 7297 12736
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 7374 12724 7380 12776
rect 7432 12773 7438 12776
rect 7432 12767 7460 12773
rect 7448 12733 7460 12767
rect 7432 12727 7460 12733
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12764 7619 12767
rect 7742 12764 7748 12776
rect 7607 12736 7748 12764
rect 7607 12733 7619 12736
rect 7561 12727 7619 12733
rect 7432 12724 7438 12727
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 9968 12764 9996 12940
rect 10410 12928 10416 12980
rect 10468 12928 10474 12980
rect 10686 12928 10692 12980
rect 10744 12968 10750 12980
rect 10781 12971 10839 12977
rect 10781 12968 10793 12971
rect 10744 12940 10793 12968
rect 10744 12928 10750 12940
rect 10781 12937 10793 12940
rect 10827 12968 10839 12971
rect 10827 12940 11560 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 10873 12903 10931 12909
rect 10873 12869 10885 12903
rect 10919 12900 10931 12903
rect 10962 12900 10968 12912
rect 10919 12872 10968 12900
rect 10919 12869 10931 12872
rect 10873 12863 10931 12869
rect 10962 12860 10968 12872
rect 11020 12860 11026 12912
rect 11532 12841 11560 12940
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 13449 12971 13507 12977
rect 13449 12968 13461 12971
rect 11756 12940 13461 12968
rect 11756 12928 11762 12940
rect 13449 12937 13461 12940
rect 13495 12937 13507 12971
rect 13449 12931 13507 12937
rect 13814 12928 13820 12980
rect 13872 12928 13878 12980
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 15749 12971 15807 12977
rect 15749 12968 15761 12971
rect 15344 12940 15761 12968
rect 15344 12928 15350 12940
rect 15749 12937 15761 12940
rect 15795 12937 15807 12971
rect 15749 12931 15807 12937
rect 16114 12928 16120 12980
rect 16172 12928 16178 12980
rect 16853 12971 16911 12977
rect 16853 12937 16865 12971
rect 16899 12968 16911 12971
rect 16942 12968 16948 12980
rect 16899 12940 16948 12968
rect 16899 12937 16911 12940
rect 16853 12931 16911 12937
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 19061 12971 19119 12977
rect 19061 12968 19073 12971
rect 17052 12940 19073 12968
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12832 11575 12835
rect 11606 12832 11612 12844
rect 11563 12804 11612 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12832 11759 12835
rect 11882 12832 11888 12844
rect 11747 12804 11888 12832
rect 11747 12801 11759 12804
rect 11701 12795 11759 12801
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 12710 12792 12716 12844
rect 12768 12792 12774 12844
rect 14274 12792 14280 12844
rect 14332 12792 14338 12844
rect 14550 12841 14556 12844
rect 14544 12832 14556 12841
rect 14511 12804 14556 12832
rect 14544 12795 14556 12804
rect 14550 12792 14556 12795
rect 14608 12792 14614 12844
rect 17052 12841 17080 12940
rect 19061 12937 19073 12940
rect 19107 12937 19119 12971
rect 19061 12931 19119 12937
rect 19150 12928 19156 12980
rect 19208 12968 19214 12980
rect 19429 12971 19487 12977
rect 19429 12968 19441 12971
rect 19208 12940 19441 12968
rect 19208 12928 19214 12940
rect 19429 12937 19441 12940
rect 19475 12937 19487 12971
rect 19429 12931 19487 12937
rect 24670 12928 24676 12980
rect 24728 12928 24734 12980
rect 24854 12928 24860 12980
rect 24912 12928 24918 12980
rect 24946 12928 24952 12980
rect 25004 12968 25010 12980
rect 29914 12968 29920 12980
rect 25004 12940 29920 12968
rect 25004 12928 25010 12940
rect 29914 12928 29920 12940
rect 29972 12928 29978 12980
rect 30193 12971 30251 12977
rect 30193 12937 30205 12971
rect 30239 12968 30251 12971
rect 30742 12968 30748 12980
rect 30239 12940 30748 12968
rect 30239 12937 30251 12940
rect 30193 12931 30251 12937
rect 30742 12928 30748 12940
rect 30800 12928 30806 12980
rect 33134 12968 33140 12980
rect 30852 12940 33140 12968
rect 19889 12903 19947 12909
rect 19889 12869 19901 12903
rect 19935 12900 19947 12903
rect 20162 12900 20168 12912
rect 19935 12872 20168 12900
rect 19935 12869 19947 12872
rect 19889 12863 19947 12869
rect 20162 12860 20168 12872
rect 20220 12860 20226 12912
rect 24688 12900 24716 12928
rect 30852 12900 30880 12940
rect 33134 12928 33140 12940
rect 33192 12928 33198 12980
rect 33870 12968 33876 12980
rect 33244 12940 33876 12968
rect 24688 12872 25176 12900
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 17310 12792 17316 12844
rect 17368 12792 17374 12844
rect 18138 12792 18144 12844
rect 18196 12841 18202 12844
rect 18196 12835 18224 12841
rect 18212 12801 18224 12835
rect 18196 12795 18224 12801
rect 18196 12792 18202 12795
rect 18322 12792 18328 12844
rect 18380 12792 18386 12844
rect 19521 12835 19579 12841
rect 19521 12801 19533 12835
rect 19567 12832 19579 12835
rect 19702 12832 19708 12844
rect 19567 12804 19708 12832
rect 19567 12801 19579 12804
rect 19521 12795 19579 12801
rect 19702 12792 19708 12804
rect 19760 12792 19766 12844
rect 20898 12792 20904 12844
rect 20956 12792 20962 12844
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 12618 12773 12624 12776
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 9968 12736 10977 12764
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 10965 12727 11023 12733
rect 12268 12736 12449 12764
rect 5123 12668 6914 12696
rect 7009 12699 7067 12705
rect 5123 12665 5135 12668
rect 5077 12659 5135 12665
rect 6564 12640 6592 12668
rect 7009 12665 7021 12699
rect 7055 12665 7067 12699
rect 12161 12699 12219 12705
rect 12161 12696 12173 12699
rect 7009 12659 7067 12665
rect 7944 12668 8892 12696
rect 6546 12588 6552 12640
rect 6604 12588 6610 12640
rect 7024 12628 7052 12659
rect 7466 12628 7472 12640
rect 7024 12600 7472 12628
rect 7466 12588 7472 12600
rect 7524 12628 7530 12640
rect 7944 12628 7972 12668
rect 7524 12600 7972 12628
rect 7524 12588 7530 12600
rect 8202 12588 8208 12640
rect 8260 12588 8266 12640
rect 8864 12628 8892 12668
rect 10152 12668 12173 12696
rect 10152 12628 10180 12668
rect 12161 12665 12173 12668
rect 12207 12665 12219 12699
rect 12161 12659 12219 12665
rect 8864 12600 10180 12628
rect 10318 12588 10324 12640
rect 10376 12628 10382 12640
rect 12268 12628 12296 12736
rect 12437 12733 12449 12736
rect 12483 12733 12495 12767
rect 12437 12727 12495 12733
rect 12575 12767 12624 12773
rect 12575 12733 12587 12767
rect 12621 12733 12624 12767
rect 12575 12727 12624 12733
rect 12618 12724 12624 12727
rect 12676 12724 12682 12776
rect 13906 12724 13912 12776
rect 13964 12724 13970 12776
rect 13998 12724 14004 12776
rect 14056 12724 14062 12776
rect 16206 12724 16212 12776
rect 16264 12724 16270 12776
rect 16393 12767 16451 12773
rect 16393 12733 16405 12767
rect 16439 12764 16451 12767
rect 16482 12764 16488 12776
rect 16439 12736 16488 12764
rect 16439 12733 16451 12736
rect 16393 12727 16451 12733
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 16942 12724 16948 12776
rect 17000 12764 17006 12776
rect 17129 12767 17187 12773
rect 17129 12764 17141 12767
rect 17000 12736 17141 12764
rect 17000 12724 17006 12736
rect 17129 12733 17141 12736
rect 17175 12733 17187 12767
rect 17129 12727 17187 12733
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 17770 12764 17776 12776
rect 17552 12736 17776 12764
rect 17552 12724 17558 12736
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 17862 12724 17868 12776
rect 17920 12764 17926 12776
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 17920 12736 18061 12764
rect 17920 12724 17926 12736
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 18874 12724 18880 12776
rect 18932 12764 18938 12776
rect 19334 12764 19340 12776
rect 18932 12736 19340 12764
rect 18932 12724 18938 12736
rect 19334 12724 19340 12736
rect 19392 12764 19398 12776
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19392 12736 19625 12764
rect 19392 12724 19398 12736
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 18969 12699 19027 12705
rect 15580 12668 17264 12696
rect 12526 12628 12532 12640
rect 10376 12600 12532 12628
rect 10376 12588 10382 12600
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 13357 12631 13415 12637
rect 13357 12597 13369 12631
rect 13403 12628 13415 12631
rect 15580 12628 15608 12668
rect 13403 12600 15608 12628
rect 13403 12597 13415 12600
rect 13357 12591 13415 12597
rect 15654 12588 15660 12640
rect 15712 12588 15718 12640
rect 17236 12628 17264 12668
rect 18969 12665 18981 12699
rect 19015 12696 19027 12699
rect 20165 12699 20223 12705
rect 20165 12696 20177 12699
rect 19015 12668 20177 12696
rect 19015 12665 19027 12668
rect 18969 12659 19027 12665
rect 20165 12665 20177 12668
rect 20211 12665 20223 12699
rect 21100 12696 21128 12795
rect 21174 12792 21180 12844
rect 21232 12792 21238 12844
rect 22554 12792 22560 12844
rect 22612 12832 22618 12844
rect 25148 12841 25176 12872
rect 25792 12872 29224 12900
rect 25133 12835 25191 12841
rect 22612 12804 23244 12832
rect 22612 12792 22618 12804
rect 23014 12724 23020 12776
rect 23072 12724 23078 12776
rect 23216 12773 23244 12804
rect 25133 12801 25145 12835
rect 25179 12801 25191 12835
rect 25133 12795 25191 12801
rect 23201 12767 23259 12773
rect 23201 12733 23213 12767
rect 23247 12733 23259 12767
rect 23201 12727 23259 12733
rect 20165 12659 20223 12665
rect 20272 12668 21128 12696
rect 23216 12696 23244 12727
rect 23290 12724 23296 12776
rect 23348 12764 23354 12776
rect 23934 12764 23940 12776
rect 23348 12736 23940 12764
rect 23348 12724 23354 12736
rect 23934 12724 23940 12736
rect 23992 12724 23998 12776
rect 24026 12724 24032 12776
rect 24084 12773 24090 12776
rect 24084 12767 24112 12773
rect 24100 12733 24112 12767
rect 24084 12727 24112 12733
rect 24213 12767 24271 12773
rect 24213 12733 24225 12767
rect 24259 12764 24271 12767
rect 24578 12764 24584 12776
rect 24259 12736 24584 12764
rect 24259 12733 24271 12736
rect 24213 12727 24271 12733
rect 24084 12724 24090 12727
rect 24578 12724 24584 12736
rect 24636 12724 24642 12776
rect 25792 12764 25820 12872
rect 25958 12792 25964 12844
rect 26016 12832 26022 12844
rect 27706 12832 27712 12844
rect 26016 12804 27712 12832
rect 26016 12792 26022 12804
rect 27706 12792 27712 12804
rect 27764 12792 27770 12844
rect 27893 12835 27951 12841
rect 27893 12801 27905 12835
rect 27939 12832 27951 12835
rect 28902 12832 28908 12844
rect 27939 12804 28908 12832
rect 27939 12801 27951 12804
rect 27893 12795 27951 12801
rect 28902 12792 28908 12804
rect 28960 12792 28966 12844
rect 29086 12841 29092 12844
rect 29080 12832 29092 12841
rect 29047 12804 29092 12832
rect 29080 12795 29092 12804
rect 29086 12792 29092 12795
rect 29144 12792 29150 12844
rect 29196 12832 29224 12872
rect 30024 12872 30880 12900
rect 30024 12832 30052 12872
rect 31018 12860 31024 12912
rect 31076 12900 31082 12912
rect 32674 12900 32680 12912
rect 31076 12872 32680 12900
rect 31076 12860 31082 12872
rect 32674 12860 32680 12872
rect 32732 12860 32738 12912
rect 29196 12804 30052 12832
rect 30098 12792 30104 12844
rect 30156 12832 30162 12844
rect 30282 12832 30288 12844
rect 30156 12804 30288 12832
rect 30156 12792 30162 12804
rect 30282 12792 30288 12804
rect 30340 12792 30346 12844
rect 30374 12792 30380 12844
rect 30432 12832 30438 12844
rect 33244 12841 33272 12940
rect 33870 12928 33876 12940
rect 33928 12928 33934 12980
rect 34514 12928 34520 12980
rect 34572 12968 34578 12980
rect 35069 12971 35127 12977
rect 35069 12968 35081 12971
rect 34572 12940 35081 12968
rect 34572 12928 34578 12940
rect 35069 12937 35081 12940
rect 35115 12937 35127 12971
rect 35069 12931 35127 12937
rect 36078 12928 36084 12980
rect 36136 12928 36142 12980
rect 39669 12971 39727 12977
rect 39669 12937 39681 12971
rect 39715 12968 39727 12971
rect 39850 12968 39856 12980
rect 39715 12940 39856 12968
rect 39715 12937 39727 12940
rect 39669 12931 39727 12937
rect 39850 12928 39856 12940
rect 39908 12928 39914 12980
rect 42797 12971 42855 12977
rect 42797 12937 42809 12971
rect 42843 12968 42855 12971
rect 43162 12968 43168 12980
rect 42843 12940 43168 12968
rect 42843 12937 42855 12940
rect 42797 12931 42855 12937
rect 43162 12928 43168 12940
rect 43220 12928 43226 12980
rect 39316 12872 39804 12900
rect 33229 12835 33287 12841
rect 30432 12804 33180 12832
rect 30432 12792 30438 12804
rect 24688 12736 25820 12764
rect 23216 12668 23336 12696
rect 20272 12628 20300 12668
rect 17236 12600 20300 12628
rect 20346 12588 20352 12640
rect 20404 12588 20410 12640
rect 20717 12631 20775 12637
rect 20717 12597 20729 12631
rect 20763 12628 20775 12631
rect 23198 12628 23204 12640
rect 20763 12600 23204 12628
rect 20763 12597 20775 12600
rect 20717 12591 20775 12597
rect 23198 12588 23204 12600
rect 23256 12588 23262 12640
rect 23308 12628 23336 12668
rect 23658 12656 23664 12708
rect 23716 12656 23722 12708
rect 24688 12628 24716 12736
rect 27798 12724 27804 12776
rect 27856 12764 27862 12776
rect 28626 12764 28632 12776
rect 27856 12736 28632 12764
rect 27856 12724 27862 12736
rect 28626 12724 28632 12736
rect 28684 12764 28690 12776
rect 28813 12767 28871 12773
rect 28813 12764 28825 12767
rect 28684 12736 28825 12764
rect 28684 12724 28690 12736
rect 28813 12733 28825 12736
rect 28859 12733 28871 12767
rect 28813 12727 28871 12733
rect 29914 12724 29920 12776
rect 29972 12764 29978 12776
rect 33152 12764 33180 12804
rect 33229 12801 33241 12835
rect 33275 12801 33287 12835
rect 33229 12795 33287 12801
rect 33336 12804 33640 12832
rect 33336 12764 33364 12804
rect 29972 12736 31754 12764
rect 33152 12736 33364 12764
rect 33413 12767 33471 12773
rect 29972 12724 29978 12736
rect 24762 12656 24768 12708
rect 24820 12696 24826 12708
rect 24820 12668 25084 12696
rect 24820 12656 24826 12668
rect 23308 12600 24716 12628
rect 24946 12588 24952 12640
rect 25004 12588 25010 12640
rect 25056 12628 25084 12668
rect 27614 12656 27620 12708
rect 27672 12696 27678 12708
rect 27709 12699 27767 12705
rect 27709 12696 27721 12699
rect 27672 12668 27721 12696
rect 27672 12656 27678 12668
rect 27709 12665 27721 12668
rect 27755 12665 27767 12699
rect 27709 12659 27767 12665
rect 29822 12656 29828 12708
rect 29880 12696 29886 12708
rect 31726 12696 31754 12736
rect 33413 12733 33425 12767
rect 33459 12764 33471 12767
rect 33502 12764 33508 12776
rect 33459 12736 33508 12764
rect 33459 12733 33471 12736
rect 33413 12727 33471 12733
rect 33502 12724 33508 12736
rect 33560 12724 33566 12776
rect 33612 12764 33640 12804
rect 34146 12792 34152 12844
rect 34204 12792 34210 12844
rect 34330 12841 34336 12844
rect 34287 12835 34336 12841
rect 34287 12801 34299 12835
rect 34333 12801 34336 12835
rect 34287 12795 34336 12801
rect 34330 12792 34336 12795
rect 34388 12792 34394 12844
rect 36265 12835 36323 12841
rect 36265 12801 36277 12835
rect 36311 12832 36323 12835
rect 37274 12832 37280 12844
rect 36311 12804 37280 12832
rect 36311 12801 36323 12804
rect 36265 12795 36323 12801
rect 37274 12792 37280 12804
rect 37332 12792 37338 12844
rect 39206 12792 39212 12844
rect 39264 12792 39270 12844
rect 33778 12764 33784 12776
rect 33612 12736 33784 12764
rect 33778 12724 33784 12736
rect 33836 12724 33842 12776
rect 33962 12724 33968 12776
rect 34020 12764 34026 12776
rect 34425 12767 34483 12773
rect 34425 12764 34437 12767
rect 34020 12736 34437 12764
rect 34020 12724 34026 12736
rect 34425 12733 34437 12736
rect 34471 12733 34483 12767
rect 39316 12764 39344 12872
rect 39393 12835 39451 12841
rect 39393 12801 39405 12835
rect 39439 12801 39451 12835
rect 39393 12795 39451 12801
rect 39485 12835 39543 12841
rect 39485 12801 39497 12835
rect 39531 12801 39543 12835
rect 39485 12795 39543 12801
rect 34425 12727 34483 12733
rect 39224 12736 39344 12764
rect 33226 12696 33232 12708
rect 29880 12668 31616 12696
rect 31726 12668 33232 12696
rect 29880 12656 29886 12668
rect 31478 12628 31484 12640
rect 25056 12600 31484 12628
rect 31478 12588 31484 12600
rect 31536 12588 31542 12640
rect 31588 12628 31616 12668
rect 33226 12656 33232 12668
rect 33284 12696 33290 12708
rect 39224 12705 39252 12736
rect 33873 12699 33931 12705
rect 33873 12696 33885 12699
rect 33284 12668 33885 12696
rect 33284 12656 33290 12668
rect 33873 12665 33885 12668
rect 33919 12665 33931 12699
rect 33873 12659 33931 12665
rect 39209 12699 39267 12705
rect 39209 12665 39221 12699
rect 39255 12665 39267 12699
rect 39408 12696 39436 12795
rect 39500 12764 39528 12795
rect 39574 12792 39580 12844
rect 39632 12792 39638 12844
rect 39776 12841 39804 12872
rect 39761 12835 39819 12841
rect 39761 12801 39773 12835
rect 39807 12801 39819 12835
rect 39761 12795 39819 12801
rect 39942 12792 39948 12844
rect 40000 12832 40006 12844
rect 40405 12835 40463 12841
rect 40405 12832 40417 12835
rect 40000 12804 40417 12832
rect 40000 12792 40006 12804
rect 40405 12801 40417 12804
rect 40451 12801 40463 12835
rect 40405 12795 40463 12801
rect 45094 12792 45100 12844
rect 45152 12792 45158 12844
rect 40497 12767 40555 12773
rect 40497 12764 40509 12767
rect 39500 12736 40509 12764
rect 40497 12733 40509 12736
rect 40543 12733 40555 12767
rect 40497 12727 40555 12733
rect 40773 12767 40831 12773
rect 40773 12733 40785 12767
rect 40819 12764 40831 12767
rect 40954 12764 40960 12776
rect 40819 12736 40960 12764
rect 40819 12733 40831 12736
rect 40773 12727 40831 12733
rect 39942 12696 39948 12708
rect 39408 12668 39948 12696
rect 39209 12659 39267 12665
rect 39942 12656 39948 12668
rect 40000 12656 40006 12708
rect 40512 12696 40540 12727
rect 40954 12724 40960 12736
rect 41012 12724 41018 12776
rect 41046 12724 41052 12776
rect 41104 12764 41110 12776
rect 42794 12764 42800 12776
rect 41104 12736 42800 12764
rect 41104 12724 41110 12736
rect 42794 12724 42800 12736
rect 42852 12764 42858 12776
rect 42981 12767 43039 12773
rect 42981 12764 42993 12767
rect 42852 12736 42993 12764
rect 42852 12724 42858 12736
rect 42981 12733 42993 12736
rect 43027 12733 43039 12767
rect 42981 12727 43039 12733
rect 43070 12724 43076 12776
rect 43128 12724 43134 12776
rect 43162 12724 43168 12776
rect 43220 12724 43226 12776
rect 44910 12724 44916 12776
rect 44968 12724 44974 12776
rect 41598 12696 41604 12708
rect 40512 12668 41604 12696
rect 41598 12656 41604 12668
rect 41656 12656 41662 12708
rect 36630 12628 36636 12640
rect 31588 12600 36636 12628
rect 36630 12588 36636 12600
rect 36688 12588 36694 12640
rect 40034 12588 40040 12640
rect 40092 12628 40098 12640
rect 43530 12628 43536 12640
rect 40092 12600 43536 12628
rect 40092 12588 40098 12600
rect 43530 12588 43536 12600
rect 43588 12628 43594 12640
rect 44082 12628 44088 12640
rect 43588 12600 44088 12628
rect 43588 12588 43594 12600
rect 44082 12588 44088 12600
rect 44140 12588 44146 12640
rect 44542 12588 44548 12640
rect 44600 12628 44606 12640
rect 45281 12631 45339 12637
rect 45281 12628 45293 12631
rect 44600 12600 45293 12628
rect 44600 12588 44606 12600
rect 45281 12597 45293 12600
rect 45327 12597 45339 12631
rect 45281 12591 45339 12597
rect 1104 12538 47104 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 47104 12538
rect 1104 12464 47104 12486
rect 5169 12427 5227 12433
rect 5169 12393 5181 12427
rect 5215 12424 5227 12427
rect 5258 12424 5264 12436
rect 5215 12396 5264 12424
rect 5215 12393 5227 12396
rect 5169 12387 5227 12393
rect 5258 12384 5264 12396
rect 5316 12424 5322 12436
rect 6914 12424 6920 12436
rect 5316 12396 6920 12424
rect 5316 12384 5322 12396
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 7745 12427 7803 12433
rect 7745 12424 7757 12427
rect 7156 12396 7757 12424
rect 7156 12384 7162 12396
rect 7745 12393 7757 12396
rect 7791 12393 7803 12427
rect 7745 12387 7803 12393
rect 9674 12384 9680 12436
rect 9732 12384 9738 12436
rect 14553 12427 14611 12433
rect 14553 12393 14565 12427
rect 14599 12424 14611 12427
rect 14642 12424 14648 12436
rect 14599 12396 14648 12424
rect 14599 12393 14611 12396
rect 14553 12387 14611 12393
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 15654 12384 15660 12436
rect 15712 12424 15718 12436
rect 17862 12424 17868 12436
rect 15712 12396 17868 12424
rect 15712 12384 15718 12396
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 19705 12427 19763 12433
rect 19705 12393 19717 12427
rect 19751 12424 19763 12427
rect 20346 12424 20352 12436
rect 19751 12396 20352 12424
rect 19751 12393 19763 12396
rect 19705 12387 19763 12393
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 20548 12396 25360 12424
rect 7653 12359 7711 12365
rect 7653 12325 7665 12359
rect 7699 12356 7711 12359
rect 11054 12356 11060 12368
rect 7699 12328 11060 12356
rect 7699 12325 7711 12328
rect 7653 12319 7711 12325
rect 11054 12316 11060 12328
rect 11112 12316 11118 12368
rect 12250 12316 12256 12368
rect 12308 12316 12314 12368
rect 17402 12356 17408 12368
rect 16960 12328 17408 12356
rect 16960 12300 16988 12328
rect 17402 12316 17408 12328
rect 17460 12316 17466 12368
rect 3694 12248 3700 12300
rect 3752 12288 3758 12300
rect 3789 12291 3847 12297
rect 3789 12288 3801 12291
rect 3752 12260 3801 12288
rect 3752 12248 3758 12260
rect 3789 12257 3801 12260
rect 3835 12257 3847 12291
rect 3789 12251 3847 12257
rect 5994 12248 6000 12300
rect 6052 12248 6058 12300
rect 6454 12248 6460 12300
rect 6512 12248 6518 12300
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 6914 12297 6920 12300
rect 6733 12291 6791 12297
rect 6733 12288 6745 12291
rect 6604 12260 6745 12288
rect 6604 12248 6610 12260
rect 6733 12257 6745 12260
rect 6779 12257 6791 12291
rect 6733 12251 6791 12257
rect 6871 12291 6920 12297
rect 6871 12257 6883 12291
rect 6917 12257 6920 12291
rect 6871 12251 6920 12257
rect 6914 12248 6920 12251
rect 6972 12288 6978 12300
rect 7374 12288 7380 12300
rect 6972 12260 7380 12288
rect 6972 12248 6978 12260
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 8018 12248 8024 12300
rect 8076 12288 8082 12300
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 8076 12260 8401 12288
rect 8076 12248 8082 12260
rect 8389 12257 8401 12260
rect 8435 12288 8447 12291
rect 8478 12288 8484 12300
rect 8435 12260 8484 12288
rect 8435 12257 8447 12260
rect 8389 12251 8447 12257
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12288 10287 12291
rect 10410 12288 10416 12300
rect 10275 12260 10416 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 11606 12248 11612 12300
rect 11664 12248 11670 12300
rect 11793 12291 11851 12297
rect 11793 12257 11805 12291
rect 11839 12288 11851 12291
rect 11882 12288 11888 12300
rect 11839 12260 11888 12288
rect 11839 12257 11851 12260
rect 11793 12251 11851 12257
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 12526 12248 12532 12300
rect 12584 12248 12590 12300
rect 12618 12248 12624 12300
rect 12676 12297 12682 12300
rect 12676 12291 12704 12297
rect 12692 12257 12704 12291
rect 12676 12251 12704 12257
rect 12676 12248 12682 12251
rect 15102 12248 15108 12300
rect 15160 12248 15166 12300
rect 16942 12248 16948 12300
rect 17000 12248 17006 12300
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12288 17187 12291
rect 17310 12288 17316 12300
rect 17175 12260 17316 12288
rect 17175 12257 17187 12260
rect 17129 12251 17187 12257
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12288 17647 12291
rect 17678 12288 17684 12300
rect 17635 12260 17684 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 17862 12248 17868 12300
rect 17920 12248 17926 12300
rect 18046 12297 18052 12300
rect 18003 12291 18052 12297
rect 18003 12257 18015 12291
rect 18049 12257 18052 12291
rect 18003 12251 18052 12257
rect 18046 12248 18052 12251
rect 18104 12248 18110 12300
rect 18141 12291 18199 12297
rect 18141 12257 18153 12291
rect 18187 12288 18199 12291
rect 19058 12288 19064 12300
rect 18187 12260 19064 12288
rect 18187 12257 18199 12260
rect 18141 12251 18199 12257
rect 19058 12248 19064 12260
rect 19116 12248 19122 12300
rect 19242 12248 19248 12300
rect 19300 12288 19306 12300
rect 19300 12260 19840 12288
rect 19300 12248 19306 12260
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 4056 12155 4114 12161
rect 4056 12121 4068 12155
rect 4102 12152 4114 12155
rect 4154 12152 4160 12164
rect 4102 12124 4160 12152
rect 4102 12121 4114 12124
rect 4056 12115 4114 12121
rect 4154 12112 4160 12124
rect 4212 12112 4218 12164
rect 5828 12084 5856 12183
rect 7006 12180 7012 12232
rect 7064 12180 7070 12232
rect 7834 12180 7840 12232
rect 7892 12220 7898 12232
rect 8113 12223 8171 12229
rect 8113 12220 8125 12223
rect 7892 12192 8125 12220
rect 7892 12180 7898 12192
rect 8113 12189 8125 12192
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12220 10103 12223
rect 10318 12220 10324 12232
rect 10091 12192 10324 12220
rect 10091 12189 10103 12192
rect 10045 12183 10103 12189
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 12802 12180 12808 12232
rect 12860 12180 12866 12232
rect 14921 12223 14979 12229
rect 14921 12189 14933 12223
rect 14967 12220 14979 12223
rect 15654 12220 15660 12232
rect 14967 12192 15660 12220
rect 14967 12189 14979 12192
rect 14921 12183 14979 12189
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 19426 12180 19432 12232
rect 19484 12180 19490 12232
rect 19518 12180 19524 12232
rect 19576 12180 19582 12232
rect 19812 12229 19840 12260
rect 19797 12223 19855 12229
rect 19797 12189 19809 12223
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 19886 12180 19892 12232
rect 19944 12180 19950 12232
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12189 20223 12223
rect 20165 12183 20223 12189
rect 15013 12155 15071 12161
rect 15013 12152 15025 12155
rect 8220 12124 11836 12152
rect 8220 12096 8248 12124
rect 6730 12084 6736 12096
rect 5828 12056 6736 12084
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 8202 12044 8208 12096
rect 8260 12044 8266 12096
rect 10137 12087 10195 12093
rect 10137 12053 10149 12087
rect 10183 12084 10195 12087
rect 10962 12084 10968 12096
rect 10183 12056 10968 12084
rect 10183 12053 10195 12056
rect 10137 12047 10195 12053
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 11808 12084 11836 12124
rect 13372 12124 15025 12152
rect 13372 12084 13400 12124
rect 15013 12121 15025 12124
rect 15059 12121 15071 12155
rect 15013 12115 15071 12121
rect 16669 12155 16727 12161
rect 16669 12121 16681 12155
rect 16715 12152 16727 12155
rect 19245 12155 19303 12161
rect 16715 12124 17172 12152
rect 16715 12121 16727 12124
rect 16669 12115 16727 12121
rect 11808 12056 13400 12084
rect 13449 12087 13507 12093
rect 13449 12053 13461 12087
rect 13495 12084 13507 12087
rect 14458 12084 14464 12096
rect 13495 12056 14464 12084
rect 13495 12053 13507 12056
rect 13449 12047 13507 12053
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 15028 12084 15056 12115
rect 16206 12084 16212 12096
rect 15028 12056 16212 12084
rect 16206 12044 16212 12056
rect 16264 12084 16270 12096
rect 16761 12087 16819 12093
rect 16761 12084 16773 12087
rect 16264 12056 16773 12084
rect 16264 12044 16270 12056
rect 16761 12053 16773 12056
rect 16807 12053 16819 12087
rect 17144 12084 17172 12124
rect 19245 12121 19257 12155
rect 19291 12152 19303 12155
rect 20180 12152 20208 12183
rect 19291 12124 20208 12152
rect 19291 12121 19303 12124
rect 19245 12115 19303 12121
rect 18690 12084 18696 12096
rect 17144 12056 18696 12084
rect 16761 12047 16819 12053
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 18785 12087 18843 12093
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 20548 12084 20576 12396
rect 23017 12359 23075 12365
rect 23017 12325 23029 12359
rect 23063 12356 23075 12359
rect 23382 12356 23388 12368
rect 23063 12328 23388 12356
rect 23063 12325 23075 12328
rect 23017 12319 23075 12325
rect 23382 12316 23388 12328
rect 23440 12356 23446 12368
rect 24026 12356 24032 12368
rect 23440 12328 24032 12356
rect 23440 12316 23446 12328
rect 24026 12316 24032 12328
rect 24084 12316 24090 12368
rect 25332 12356 25360 12396
rect 25774 12384 25780 12436
rect 25832 12384 25838 12436
rect 25958 12384 25964 12436
rect 26016 12424 26022 12436
rect 33686 12424 33692 12436
rect 26016 12396 33692 12424
rect 26016 12384 26022 12396
rect 33686 12384 33692 12396
rect 33744 12384 33750 12436
rect 38746 12424 38752 12436
rect 37936 12396 38752 12424
rect 26145 12359 26203 12365
rect 26145 12356 26157 12359
rect 25332 12328 26157 12356
rect 26145 12325 26157 12328
rect 26191 12325 26203 12359
rect 30009 12359 30067 12365
rect 30009 12356 30021 12359
rect 26145 12319 26203 12325
rect 28966 12328 30021 12356
rect 22922 12248 22928 12300
rect 22980 12288 22986 12300
rect 23753 12291 23811 12297
rect 23753 12288 23765 12291
rect 22980 12260 23765 12288
rect 22980 12248 22986 12260
rect 23753 12257 23765 12260
rect 23799 12257 23811 12291
rect 27709 12291 27767 12297
rect 23753 12251 23811 12257
rect 25424 12260 27660 12288
rect 21637 12223 21695 12229
rect 21637 12189 21649 12223
rect 21683 12220 21695 12223
rect 22462 12220 22468 12232
rect 21683 12192 22468 12220
rect 21683 12189 21695 12192
rect 21637 12183 21695 12189
rect 22462 12180 22468 12192
rect 22520 12180 22526 12232
rect 22738 12180 22744 12232
rect 22796 12220 22802 12232
rect 23290 12220 23296 12232
rect 22796 12192 23296 12220
rect 22796 12180 22802 12192
rect 23290 12180 23296 12192
rect 23348 12220 23354 12232
rect 23348 12192 23612 12220
rect 23348 12180 23354 12192
rect 21904 12155 21962 12161
rect 21904 12121 21916 12155
rect 21950 12152 21962 12155
rect 22002 12152 22008 12164
rect 21950 12124 22008 12152
rect 21950 12121 21962 12124
rect 21904 12115 21962 12121
rect 22002 12112 22008 12124
rect 22060 12112 22066 12164
rect 23584 12161 23612 12192
rect 23569 12155 23627 12161
rect 23569 12121 23581 12155
rect 23615 12152 23627 12155
rect 23768 12152 23796 12251
rect 24397 12223 24455 12229
rect 24397 12189 24409 12223
rect 24443 12220 24455 12223
rect 24486 12220 24492 12232
rect 24443 12192 24492 12220
rect 24443 12189 24455 12192
rect 24397 12183 24455 12189
rect 24486 12180 24492 12192
rect 24544 12180 24550 12232
rect 24670 12229 24676 12232
rect 24664 12183 24676 12229
rect 24670 12180 24676 12183
rect 24728 12180 24734 12232
rect 25424 12220 25452 12260
rect 24780 12192 25452 12220
rect 24780 12152 24808 12192
rect 25498 12180 25504 12232
rect 25556 12220 25562 12232
rect 25556 12192 27200 12220
rect 25556 12180 25562 12192
rect 23615 12124 23704 12152
rect 23768 12124 24808 12152
rect 23615 12121 23627 12124
rect 23569 12115 23627 12121
rect 18831 12056 20576 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 20714 12044 20720 12096
rect 20772 12084 20778 12096
rect 20901 12087 20959 12093
rect 20901 12084 20913 12087
rect 20772 12056 20913 12084
rect 20772 12044 20778 12056
rect 20901 12053 20913 12056
rect 20947 12053 20959 12087
rect 20901 12047 20959 12053
rect 23106 12044 23112 12096
rect 23164 12044 23170 12096
rect 23474 12044 23480 12096
rect 23532 12044 23538 12096
rect 23676 12084 23704 12124
rect 25038 12112 25044 12164
rect 25096 12152 25102 12164
rect 25866 12152 25872 12164
rect 25096 12124 25872 12152
rect 25096 12112 25102 12124
rect 25866 12112 25872 12124
rect 25924 12112 25930 12164
rect 25498 12084 25504 12096
rect 23676 12056 25504 12084
rect 25498 12044 25504 12056
rect 25556 12044 25562 12096
rect 26329 12087 26387 12093
rect 26329 12053 26341 12087
rect 26375 12084 26387 12087
rect 26694 12084 26700 12096
rect 26375 12056 26700 12084
rect 26375 12053 26387 12056
rect 26329 12047 26387 12053
rect 26694 12044 26700 12056
rect 26752 12044 26758 12096
rect 26786 12044 26792 12096
rect 26844 12084 26850 12096
rect 27065 12087 27123 12093
rect 27065 12084 27077 12087
rect 26844 12056 27077 12084
rect 26844 12044 26850 12056
rect 27065 12053 27077 12056
rect 27111 12053 27123 12087
rect 27172 12084 27200 12192
rect 27246 12112 27252 12164
rect 27304 12152 27310 12164
rect 27433 12155 27491 12161
rect 27433 12152 27445 12155
rect 27304 12124 27445 12152
rect 27304 12112 27310 12124
rect 27433 12121 27445 12124
rect 27479 12121 27491 12155
rect 27632 12152 27660 12260
rect 27709 12257 27721 12291
rect 27755 12288 27767 12291
rect 28966 12288 28994 12328
rect 30009 12325 30021 12328
rect 30055 12356 30067 12359
rect 30466 12356 30472 12368
rect 30055 12328 30472 12356
rect 30055 12325 30067 12328
rect 30009 12319 30067 12325
rect 30466 12316 30472 12328
rect 30524 12316 30530 12368
rect 36446 12316 36452 12368
rect 36504 12316 36510 12368
rect 27755 12260 28994 12288
rect 27755 12257 27767 12260
rect 27709 12251 27767 12257
rect 30282 12248 30288 12300
rect 30340 12288 30346 12300
rect 30340 12260 36216 12288
rect 30340 12248 30346 12260
rect 29825 12223 29883 12229
rect 29825 12189 29837 12223
rect 29871 12220 29883 12223
rect 29914 12220 29920 12232
rect 29871 12192 29920 12220
rect 29871 12189 29883 12192
rect 29825 12183 29883 12189
rect 29914 12180 29920 12192
rect 29972 12180 29978 12232
rect 32493 12223 32551 12229
rect 32493 12189 32505 12223
rect 32539 12220 32551 12223
rect 32766 12220 32772 12232
rect 32539 12192 32772 12220
rect 32539 12189 32551 12192
rect 32493 12183 32551 12189
rect 32766 12180 32772 12192
rect 32824 12180 32830 12232
rect 36188 12229 36216 12260
rect 35897 12223 35955 12229
rect 35897 12189 35909 12223
rect 35943 12189 35955 12223
rect 35897 12183 35955 12189
rect 36173 12223 36231 12229
rect 36173 12189 36185 12223
rect 36219 12189 36231 12223
rect 36173 12183 36231 12189
rect 36317 12223 36375 12229
rect 36317 12189 36329 12223
rect 36363 12220 36375 12223
rect 36538 12220 36544 12232
rect 36363 12192 36544 12220
rect 36363 12189 36375 12192
rect 36317 12183 36375 12189
rect 33594 12152 33600 12164
rect 27632 12124 33600 12152
rect 27433 12115 27491 12121
rect 33594 12112 33600 12124
rect 33652 12112 33658 12164
rect 27525 12087 27583 12093
rect 27525 12084 27537 12087
rect 27172 12056 27537 12084
rect 27065 12047 27123 12053
rect 27525 12053 27537 12056
rect 27571 12084 27583 12087
rect 29270 12084 29276 12096
rect 27571 12056 29276 12084
rect 27571 12053 27583 12056
rect 27525 12047 27583 12053
rect 29270 12044 29276 12056
rect 29328 12044 29334 12096
rect 32677 12087 32735 12093
rect 32677 12053 32689 12087
rect 32723 12084 32735 12087
rect 33686 12084 33692 12096
rect 32723 12056 33692 12084
rect 32723 12053 32735 12056
rect 32677 12047 32735 12053
rect 33686 12044 33692 12056
rect 33744 12044 33750 12096
rect 35912 12084 35940 12183
rect 36538 12180 36544 12192
rect 36596 12220 36602 12232
rect 36722 12220 36728 12232
rect 36596 12192 36728 12220
rect 36596 12180 36602 12192
rect 36722 12180 36728 12192
rect 36780 12180 36786 12232
rect 36081 12155 36139 12161
rect 36081 12121 36093 12155
rect 36127 12152 36139 12155
rect 37936 12152 37964 12396
rect 38746 12384 38752 12396
rect 38804 12384 38810 12436
rect 38838 12384 38844 12436
rect 38896 12424 38902 12436
rect 39117 12427 39175 12433
rect 39117 12424 39129 12427
rect 38896 12396 39129 12424
rect 38896 12384 38902 12396
rect 39117 12393 39129 12396
rect 39163 12393 39175 12427
rect 39117 12387 39175 12393
rect 39206 12384 39212 12436
rect 39264 12424 39270 12436
rect 39577 12427 39635 12433
rect 39577 12424 39589 12427
rect 39264 12396 39589 12424
rect 39264 12384 39270 12396
rect 39577 12393 39589 12396
rect 39623 12393 39635 12427
rect 39577 12387 39635 12393
rect 40034 12384 40040 12436
rect 40092 12384 40098 12436
rect 41598 12384 41604 12436
rect 41656 12384 41662 12436
rect 41690 12384 41696 12436
rect 41748 12424 41754 12436
rect 41748 12396 42564 12424
rect 41748 12384 41754 12396
rect 38657 12359 38715 12365
rect 38657 12325 38669 12359
rect 38703 12356 38715 12359
rect 39482 12356 39488 12368
rect 38703 12328 39488 12356
rect 38703 12325 38715 12328
rect 38657 12319 38715 12325
rect 39482 12316 39488 12328
rect 39540 12316 39546 12368
rect 40862 12316 40868 12368
rect 40920 12356 40926 12368
rect 41233 12359 41291 12365
rect 41233 12356 41245 12359
rect 40920 12328 41245 12356
rect 40920 12316 40926 12328
rect 41233 12325 41245 12328
rect 41279 12356 41291 12359
rect 42536 12356 42564 12396
rect 43070 12384 43076 12436
rect 43128 12424 43134 12436
rect 43441 12427 43499 12433
rect 43441 12424 43453 12427
rect 43128 12396 43453 12424
rect 43128 12384 43134 12396
rect 43441 12393 43453 12396
rect 43487 12393 43499 12427
rect 43441 12387 43499 12393
rect 41279 12328 42472 12356
rect 42536 12328 43116 12356
rect 41279 12325 41291 12328
rect 41233 12319 41291 12325
rect 38010 12248 38016 12300
rect 38068 12288 38074 12300
rect 38933 12291 38991 12297
rect 38933 12288 38945 12291
rect 38068 12260 38945 12288
rect 38068 12248 38074 12260
rect 38933 12257 38945 12260
rect 38979 12257 38991 12291
rect 38933 12251 38991 12257
rect 41417 12291 41475 12297
rect 41417 12257 41429 12291
rect 41463 12288 41475 12291
rect 42444 12288 42472 12328
rect 43088 12297 43116 12328
rect 44082 12316 44088 12368
rect 44140 12316 44146 12368
rect 43073 12291 43131 12297
rect 41463 12260 42380 12288
rect 42444 12260 42840 12288
rect 41463 12257 41475 12260
rect 41417 12251 41475 12257
rect 38381 12223 38439 12229
rect 38381 12189 38393 12223
rect 38427 12189 38439 12223
rect 38381 12183 38439 12189
rect 38565 12223 38623 12229
rect 38565 12189 38577 12223
rect 38611 12220 38623 12223
rect 38838 12220 38844 12232
rect 38611 12192 38844 12220
rect 38611 12189 38623 12192
rect 38565 12183 38623 12189
rect 36127 12124 37964 12152
rect 36127 12121 36139 12124
rect 36081 12115 36139 12121
rect 37458 12084 37464 12096
rect 35912 12056 37464 12084
rect 37458 12044 37464 12056
rect 37516 12044 37522 12096
rect 38396 12084 38424 12183
rect 38838 12180 38844 12192
rect 38896 12180 38902 12232
rect 38948 12220 38976 12251
rect 39025 12223 39083 12229
rect 39025 12220 39037 12223
rect 38948 12192 39037 12220
rect 39025 12189 39037 12192
rect 39071 12189 39083 12223
rect 39025 12183 39083 12189
rect 39301 12223 39359 12229
rect 39301 12189 39313 12223
rect 39347 12189 39359 12223
rect 39301 12183 39359 12189
rect 39114 12152 39120 12164
rect 38764 12124 39120 12152
rect 38764 12084 38792 12124
rect 39114 12112 39120 12124
rect 39172 12152 39178 12164
rect 39316 12152 39344 12183
rect 39758 12180 39764 12232
rect 39816 12220 39822 12232
rect 39853 12223 39911 12229
rect 39853 12220 39865 12223
rect 39816 12192 39865 12220
rect 39816 12180 39822 12192
rect 39853 12189 39865 12192
rect 39899 12189 39911 12223
rect 39853 12183 39911 12189
rect 40037 12223 40095 12229
rect 40037 12189 40049 12223
rect 40083 12220 40095 12223
rect 40402 12220 40408 12232
rect 40083 12192 40408 12220
rect 40083 12189 40095 12192
rect 40037 12183 40095 12189
rect 40402 12180 40408 12192
rect 40460 12180 40466 12232
rect 41141 12223 41199 12229
rect 41141 12189 41153 12223
rect 41187 12220 41199 12223
rect 41690 12220 41696 12232
rect 41187 12192 41696 12220
rect 41187 12189 41199 12192
rect 41141 12183 41199 12189
rect 41690 12180 41696 12192
rect 41748 12180 41754 12232
rect 41800 12229 41828 12260
rect 41785 12223 41843 12229
rect 41785 12189 41797 12223
rect 41831 12189 41843 12223
rect 41785 12183 41843 12189
rect 42242 12180 42248 12232
rect 42300 12180 42306 12232
rect 41046 12152 41052 12164
rect 39172 12124 39344 12152
rect 40144 12124 41052 12152
rect 39172 12112 39178 12124
rect 38396 12056 38792 12084
rect 38838 12044 38844 12096
rect 38896 12044 38902 12096
rect 38930 12044 38936 12096
rect 38988 12084 38994 12096
rect 40144 12084 40172 12124
rect 41046 12112 41052 12124
rect 41104 12112 41110 12164
rect 42352 12152 42380 12260
rect 42429 12223 42487 12229
rect 42429 12189 42441 12223
rect 42475 12220 42487 12223
rect 42702 12220 42708 12232
rect 42475 12192 42708 12220
rect 42475 12189 42487 12192
rect 42429 12183 42487 12189
rect 42702 12180 42708 12192
rect 42760 12180 42766 12232
rect 42812 12229 42840 12260
rect 43073 12257 43085 12291
rect 43119 12257 43131 12291
rect 43073 12251 43131 12257
rect 43346 12248 43352 12300
rect 43404 12288 43410 12300
rect 44100 12288 44128 12316
rect 43404 12260 43944 12288
rect 44100 12260 44496 12288
rect 43404 12248 43410 12260
rect 42797 12223 42855 12229
rect 42797 12189 42809 12223
rect 42843 12189 42855 12223
rect 42797 12183 42855 12189
rect 43622 12180 43628 12232
rect 43680 12220 43686 12232
rect 43717 12223 43775 12229
rect 43717 12220 43729 12223
rect 43680 12192 43729 12220
rect 43680 12180 43686 12192
rect 43717 12189 43729 12192
rect 43763 12189 43775 12223
rect 43717 12183 43775 12189
rect 43806 12180 43812 12232
rect 43864 12180 43870 12232
rect 43916 12229 43944 12260
rect 43901 12223 43959 12229
rect 43901 12189 43913 12223
rect 43947 12189 43959 12223
rect 43901 12183 43959 12189
rect 43990 12180 43996 12232
rect 44048 12220 44054 12232
rect 44085 12223 44143 12229
rect 44085 12220 44097 12223
rect 44048 12192 44097 12220
rect 44048 12180 44054 12192
rect 44085 12189 44097 12192
rect 44131 12189 44143 12223
rect 44085 12183 44143 12189
rect 44174 12180 44180 12232
rect 44232 12180 44238 12232
rect 44468 12229 44496 12260
rect 44453 12223 44511 12229
rect 44453 12189 44465 12223
rect 44499 12189 44511 12223
rect 44453 12183 44511 12189
rect 44542 12180 44548 12232
rect 44600 12180 44606 12232
rect 43162 12152 43168 12164
rect 42352 12124 43168 12152
rect 43162 12112 43168 12124
rect 43220 12112 43226 12164
rect 43254 12112 43260 12164
rect 43312 12152 43318 12164
rect 44361 12155 44419 12161
rect 44361 12152 44373 12155
rect 43312 12124 44373 12152
rect 43312 12112 43318 12124
rect 44361 12121 44373 12124
rect 44407 12121 44419 12155
rect 44361 12115 44419 12121
rect 38988 12056 40172 12084
rect 38988 12044 38994 12056
rect 40218 12044 40224 12096
rect 40276 12044 40282 12096
rect 41414 12044 41420 12096
rect 41472 12044 41478 12096
rect 43530 12044 43536 12096
rect 43588 12084 43594 12096
rect 44729 12087 44787 12093
rect 44729 12084 44741 12087
rect 43588 12056 44741 12084
rect 43588 12044 43594 12056
rect 44729 12053 44741 12056
rect 44775 12053 44787 12087
rect 44729 12047 44787 12053
rect 1104 11994 47104 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 47104 11994
rect 1104 11920 47104 11942
rect 4154 11840 4160 11892
rect 4212 11840 4218 11892
rect 4801 11883 4859 11889
rect 4801 11849 4813 11883
rect 4847 11849 4859 11883
rect 4801 11843 4859 11849
rect 5169 11883 5227 11889
rect 5169 11849 5181 11883
rect 5215 11880 5227 11883
rect 5258 11880 5264 11892
rect 5215 11852 5264 11880
rect 5215 11849 5227 11852
rect 5169 11843 5227 11849
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11744 4399 11747
rect 4816 11744 4844 11843
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 8202 11880 8208 11892
rect 6840 11852 8208 11880
rect 6840 11821 6868 11852
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 10413 11883 10471 11889
rect 10413 11849 10425 11883
rect 10459 11880 10471 11883
rect 10873 11883 10931 11889
rect 10873 11880 10885 11883
rect 10459 11852 10885 11880
rect 10459 11849 10471 11852
rect 10413 11843 10471 11849
rect 10873 11849 10885 11852
rect 10919 11880 10931 11883
rect 12618 11880 12624 11892
rect 10919 11852 12624 11880
rect 10919 11849 10931 11852
rect 10873 11843 10931 11849
rect 12618 11840 12624 11852
rect 12676 11840 12682 11892
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 21266 11880 21272 11892
rect 19576 11852 21272 11880
rect 19576 11840 19582 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 22002 11840 22008 11892
rect 22060 11840 22066 11892
rect 23385 11883 23443 11889
rect 23385 11849 23397 11883
rect 23431 11880 23443 11883
rect 23934 11880 23940 11892
rect 23431 11852 23940 11880
rect 23431 11849 23443 11852
rect 23385 11843 23443 11849
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 26605 11883 26663 11889
rect 26605 11849 26617 11883
rect 26651 11849 26663 11883
rect 26605 11843 26663 11849
rect 6825 11815 6883 11821
rect 6825 11812 6837 11815
rect 5644 11784 6837 11812
rect 5644 11756 5672 11784
rect 6825 11781 6837 11784
rect 6871 11781 6883 11815
rect 6825 11775 6883 11781
rect 7006 11772 7012 11824
rect 7064 11812 7070 11824
rect 8846 11812 8852 11824
rect 7064 11784 8852 11812
rect 7064 11772 7070 11784
rect 8846 11772 8852 11784
rect 8904 11772 8910 11824
rect 23290 11772 23296 11824
rect 23348 11812 23354 11824
rect 23477 11815 23535 11821
rect 23477 11812 23489 11815
rect 23348 11784 23489 11812
rect 23348 11772 23354 11784
rect 23477 11781 23489 11784
rect 23523 11781 23535 11815
rect 23477 11775 23535 11781
rect 23842 11772 23848 11824
rect 23900 11812 23906 11824
rect 25958 11812 25964 11824
rect 23900 11784 25964 11812
rect 23900 11772 23906 11784
rect 25958 11772 25964 11784
rect 26016 11772 26022 11824
rect 26620 11812 26648 11843
rect 26694 11840 26700 11892
rect 26752 11880 26758 11892
rect 30377 11883 30435 11889
rect 26752 11852 29776 11880
rect 26752 11840 26758 11852
rect 27218 11815 27276 11821
rect 27218 11812 27230 11815
rect 26620 11784 27230 11812
rect 27218 11781 27230 11784
rect 27264 11781 27276 11815
rect 27218 11775 27276 11781
rect 4387 11716 4844 11744
rect 5261 11747 5319 11753
rect 4387 11713 4399 11716
rect 4341 11707 4399 11713
rect 5261 11713 5273 11747
rect 5307 11744 5319 11747
rect 5626 11744 5632 11756
rect 5307 11716 5632 11744
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 5997 11747 6055 11753
rect 5997 11713 6009 11747
rect 6043 11744 6055 11747
rect 6043 11716 6408 11744
rect 6043 11713 6055 11716
rect 5997 11707 6055 11713
rect 5445 11679 5503 11685
rect 5445 11645 5457 11679
rect 5491 11676 5503 11679
rect 5491 11648 6132 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 5626 11500 5632 11552
rect 5684 11540 5690 11552
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 5684 11512 5825 11540
rect 5684 11500 5690 11512
rect 5813 11509 5825 11512
rect 5859 11509 5871 11543
rect 6104 11540 6132 11648
rect 6380 11617 6408 11716
rect 6730 11704 6736 11756
rect 6788 11704 6794 11756
rect 8938 11704 8944 11756
rect 8996 11744 9002 11756
rect 9306 11753 9312 11756
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8996 11716 9045 11744
rect 8996 11704 9002 11716
rect 9033 11713 9045 11716
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 9300 11707 9312 11753
rect 9306 11704 9312 11707
rect 9364 11704 9370 11756
rect 10962 11704 10968 11756
rect 11020 11744 11026 11756
rect 14182 11744 14188 11756
rect 11020 11716 14188 11744
rect 11020 11704 11026 11716
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11744 22247 11747
rect 23106 11744 23112 11756
rect 22235 11716 23112 11744
rect 22235 11713 22247 11716
rect 22189 11707 22247 11713
rect 23106 11704 23112 11716
rect 23164 11704 23170 11756
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11676 7067 11679
rect 7650 11676 7656 11688
rect 7055 11648 7656 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 7650 11636 7656 11648
rect 7708 11636 7714 11688
rect 11057 11679 11115 11685
rect 11057 11676 11069 11679
rect 10980 11648 11069 11676
rect 10980 11620 11008 11648
rect 11057 11645 11069 11648
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 23661 11679 23719 11685
rect 23661 11645 23673 11679
rect 23707 11676 23719 11679
rect 23860 11676 23888 11772
rect 26786 11704 26792 11756
rect 26844 11704 26850 11756
rect 26973 11747 27031 11753
rect 26973 11713 26985 11747
rect 27019 11744 27031 11747
rect 27522 11744 27528 11756
rect 27019 11716 27528 11744
rect 27019 11713 27031 11716
rect 26973 11707 27031 11713
rect 23707 11648 23888 11676
rect 23707 11645 23719 11648
rect 23661 11639 23719 11645
rect 24486 11636 24492 11688
rect 24544 11676 24550 11688
rect 26988 11676 27016 11707
rect 27522 11704 27528 11716
rect 27580 11704 27586 11756
rect 29270 11704 29276 11756
rect 29328 11744 29334 11756
rect 29748 11753 29776 11852
rect 30377 11849 30389 11883
rect 30423 11880 30435 11883
rect 31846 11880 31852 11892
rect 30423 11852 31852 11880
rect 30423 11849 30435 11852
rect 30377 11843 30435 11849
rect 31846 11840 31852 11852
rect 31904 11840 31910 11892
rect 33413 11883 33471 11889
rect 33413 11880 33425 11883
rect 33244 11852 33425 11880
rect 30006 11772 30012 11824
rect 30064 11812 30070 11824
rect 31570 11812 31576 11824
rect 30064 11784 31576 11812
rect 30064 11772 30070 11784
rect 31570 11772 31576 11784
rect 31628 11772 31634 11824
rect 31665 11815 31723 11821
rect 31665 11781 31677 11815
rect 31711 11812 31723 11815
rect 33244 11812 33272 11852
rect 33413 11849 33425 11852
rect 33459 11880 33471 11883
rect 34238 11880 34244 11892
rect 33459 11852 34244 11880
rect 33459 11849 33471 11852
rect 33413 11843 33471 11849
rect 34238 11840 34244 11852
rect 34296 11840 34302 11892
rect 38010 11840 38016 11892
rect 38068 11840 38074 11892
rect 41414 11880 41420 11892
rect 38580 11852 41420 11880
rect 31711 11784 33272 11812
rect 33321 11815 33379 11821
rect 31711 11781 31723 11784
rect 31665 11775 31723 11781
rect 33321 11781 33333 11815
rect 33367 11812 33379 11815
rect 34330 11812 34336 11824
rect 33367 11784 34336 11812
rect 33367 11781 33379 11784
rect 33321 11775 33379 11781
rect 34330 11772 34336 11784
rect 34388 11772 34394 11824
rect 37826 11812 37832 11824
rect 37568 11784 37832 11812
rect 29365 11747 29423 11753
rect 29365 11744 29377 11747
rect 29328 11716 29377 11744
rect 29328 11704 29334 11716
rect 29365 11713 29377 11716
rect 29411 11713 29423 11747
rect 29365 11707 29423 11713
rect 29457 11747 29515 11753
rect 29457 11713 29469 11747
rect 29503 11713 29515 11747
rect 29457 11707 29515 11713
rect 29733 11747 29791 11753
rect 29733 11713 29745 11747
rect 29779 11713 29791 11747
rect 29733 11707 29791 11713
rect 24544 11648 27016 11676
rect 29472 11676 29500 11707
rect 29822 11704 29828 11756
rect 29880 11744 29886 11756
rect 30190 11744 30196 11756
rect 29880 11716 30196 11744
rect 29880 11704 29886 11716
rect 30190 11704 30196 11716
rect 30248 11704 30254 11756
rect 30374 11704 30380 11756
rect 30432 11744 30438 11756
rect 30469 11747 30527 11753
rect 30469 11744 30481 11747
rect 30432 11716 30481 11744
rect 30432 11704 30438 11716
rect 30469 11713 30481 11716
rect 30515 11744 30527 11747
rect 31386 11744 31392 11756
rect 30515 11716 31392 11744
rect 30515 11713 30527 11716
rect 30469 11707 30527 11713
rect 31386 11704 31392 11716
rect 31444 11704 31450 11756
rect 32217 11747 32275 11753
rect 32217 11713 32229 11747
rect 32263 11744 32275 11747
rect 32490 11744 32496 11756
rect 32263 11716 32496 11744
rect 32263 11713 32275 11716
rect 32217 11707 32275 11713
rect 32490 11704 32496 11716
rect 32548 11704 32554 11756
rect 32585 11747 32643 11753
rect 32585 11713 32597 11747
rect 32631 11744 32643 11747
rect 32631 11716 33640 11744
rect 32631 11713 32643 11716
rect 32585 11707 32643 11713
rect 33612 11688 33640 11716
rect 34146 11704 34152 11756
rect 34204 11704 34210 11756
rect 37568 11753 37596 11784
rect 37826 11772 37832 11784
rect 37884 11812 37890 11824
rect 37884 11784 38332 11812
rect 37884 11772 37890 11784
rect 38304 11753 38332 11784
rect 37553 11747 37611 11753
rect 37553 11713 37565 11747
rect 37599 11713 37611 11747
rect 37553 11707 37611 11713
rect 38105 11747 38163 11753
rect 38105 11713 38117 11747
rect 38151 11713 38163 11747
rect 38105 11707 38163 11713
rect 38289 11747 38347 11753
rect 38289 11713 38301 11747
rect 38335 11744 38347 11747
rect 38470 11744 38476 11756
rect 38335 11716 38476 11744
rect 38335 11713 38347 11716
rect 38289 11707 38347 11713
rect 30009 11679 30067 11685
rect 30009 11676 30021 11679
rect 29472 11648 30021 11676
rect 24544 11636 24550 11648
rect 30009 11645 30021 11648
rect 30055 11645 30067 11679
rect 30009 11639 30067 11645
rect 30558 11636 30564 11688
rect 30616 11676 30622 11688
rect 31757 11679 31815 11685
rect 31757 11676 31769 11679
rect 30616 11648 31769 11676
rect 30616 11636 30622 11648
rect 31757 11645 31769 11648
rect 31803 11645 31815 11679
rect 31757 11639 31815 11645
rect 33594 11636 33600 11688
rect 33652 11636 33658 11688
rect 33686 11636 33692 11688
rect 33744 11676 33750 11688
rect 34333 11679 34391 11685
rect 34333 11676 34345 11679
rect 33744 11648 34345 11676
rect 33744 11636 33750 11648
rect 34333 11645 34345 11648
rect 34379 11645 34391 11679
rect 34333 11639 34391 11645
rect 38120 11620 38148 11707
rect 38470 11704 38476 11716
rect 38528 11704 38534 11756
rect 38580 11744 38608 11852
rect 41414 11840 41420 11852
rect 41472 11840 41478 11892
rect 41601 11883 41659 11889
rect 41601 11849 41613 11883
rect 41647 11880 41659 11883
rect 41690 11880 41696 11892
rect 41647 11852 41696 11880
rect 41647 11849 41659 11852
rect 41601 11843 41659 11849
rect 41690 11840 41696 11852
rect 41748 11840 41754 11892
rect 42245 11883 42303 11889
rect 42245 11849 42257 11883
rect 42291 11849 42303 11883
rect 42245 11843 42303 11849
rect 42613 11883 42671 11889
rect 42613 11849 42625 11883
rect 42659 11880 42671 11883
rect 43162 11880 43168 11892
rect 42659 11852 43168 11880
rect 42659 11849 42671 11852
rect 42613 11843 42671 11849
rect 38727 11815 38785 11821
rect 38727 11781 38739 11815
rect 38773 11812 38785 11815
rect 38838 11812 38844 11824
rect 38773 11784 38844 11812
rect 38773 11781 38785 11784
rect 38727 11775 38785 11781
rect 38838 11772 38844 11784
rect 38896 11772 38902 11824
rect 39117 11815 39175 11821
rect 39117 11781 39129 11815
rect 39163 11812 39175 11815
rect 42260 11812 42288 11843
rect 43162 11840 43168 11852
rect 43220 11840 43226 11892
rect 43990 11812 43996 11824
rect 39163 11784 39528 11812
rect 42260 11784 43996 11812
rect 39163 11781 39175 11784
rect 39117 11775 39175 11781
rect 39025 11747 39083 11753
rect 38580 11716 38792 11744
rect 38197 11679 38255 11685
rect 38197 11645 38209 11679
rect 38243 11645 38255 11679
rect 38197 11639 38255 11645
rect 38657 11679 38715 11685
rect 38657 11645 38669 11679
rect 38703 11676 38715 11679
rect 38764 11676 38792 11716
rect 39025 11713 39037 11747
rect 39071 11744 39083 11747
rect 39301 11747 39359 11753
rect 39301 11744 39313 11747
rect 39071 11716 39313 11744
rect 39071 11713 39083 11716
rect 39025 11707 39083 11713
rect 39301 11713 39313 11716
rect 39347 11744 39359 11747
rect 39390 11744 39396 11756
rect 39347 11716 39396 11744
rect 39347 11713 39359 11716
rect 39301 11707 39359 11713
rect 39390 11704 39396 11716
rect 39448 11704 39454 11756
rect 38703 11648 38792 11676
rect 38703 11645 38715 11648
rect 38657 11639 38715 11645
rect 6365 11611 6423 11617
rect 6365 11577 6377 11611
rect 6411 11577 6423 11611
rect 6365 11571 6423 11577
rect 6454 11568 6460 11620
rect 6512 11608 6518 11620
rect 8294 11608 8300 11620
rect 6512 11580 8300 11608
rect 6512 11568 6518 11580
rect 8294 11568 8300 11580
rect 8352 11568 8358 11620
rect 10962 11568 10968 11620
rect 11020 11568 11026 11620
rect 29181 11611 29239 11617
rect 22066 11580 27016 11608
rect 7558 11540 7564 11552
rect 6104 11512 7564 11540
rect 5813 11503 5871 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 10502 11500 10508 11552
rect 10560 11500 10566 11552
rect 18690 11500 18696 11552
rect 18748 11540 18754 11552
rect 19702 11540 19708 11552
rect 18748 11512 19708 11540
rect 18748 11500 18754 11512
rect 19702 11500 19708 11512
rect 19760 11540 19766 11552
rect 22066 11540 22094 11580
rect 19760 11512 22094 11540
rect 19760 11500 19766 11512
rect 23014 11500 23020 11552
rect 23072 11500 23078 11552
rect 23198 11500 23204 11552
rect 23256 11540 23262 11552
rect 25866 11540 25872 11552
rect 23256 11512 25872 11540
rect 23256 11500 23262 11512
rect 25866 11500 25872 11512
rect 25924 11500 25930 11552
rect 26988 11540 27016 11580
rect 29181 11577 29193 11611
rect 29227 11608 29239 11611
rect 35894 11608 35900 11620
rect 29227 11580 35900 11608
rect 29227 11577 29239 11580
rect 29181 11571 29239 11577
rect 35894 11568 35900 11580
rect 35952 11568 35958 11620
rect 38102 11608 38108 11620
rect 37844 11580 38108 11608
rect 27246 11540 27252 11552
rect 26988 11512 27252 11540
rect 27246 11500 27252 11512
rect 27304 11500 27310 11552
rect 27338 11500 27344 11552
rect 27396 11540 27402 11552
rect 28353 11543 28411 11549
rect 28353 11540 28365 11543
rect 27396 11512 28365 11540
rect 27396 11500 27402 11512
rect 28353 11509 28365 11512
rect 28399 11509 28411 11543
rect 28353 11503 28411 11509
rect 28718 11500 28724 11552
rect 28776 11540 28782 11552
rect 29641 11543 29699 11549
rect 29641 11540 29653 11543
rect 28776 11512 29653 11540
rect 28776 11500 28782 11512
rect 29641 11509 29653 11512
rect 29687 11509 29699 11543
rect 29641 11503 29699 11509
rect 31205 11543 31263 11549
rect 31205 11509 31217 11543
rect 31251 11540 31263 11543
rect 31386 11540 31392 11552
rect 31251 11512 31392 11540
rect 31251 11509 31263 11512
rect 31205 11503 31263 11509
rect 31386 11500 31392 11512
rect 31444 11500 31450 11552
rect 32674 11500 32680 11552
rect 32732 11540 32738 11552
rect 32953 11543 33011 11549
rect 32953 11540 32965 11543
rect 32732 11512 32965 11540
rect 32732 11500 32738 11512
rect 32953 11509 32965 11512
rect 32999 11509 33011 11543
rect 32953 11503 33011 11509
rect 33781 11543 33839 11549
rect 33781 11509 33793 11543
rect 33827 11540 33839 11543
rect 34422 11540 34428 11552
rect 33827 11512 34428 11540
rect 33827 11509 33839 11512
rect 33781 11503 33839 11509
rect 34422 11500 34428 11512
rect 34480 11500 34486 11552
rect 37844 11549 37872 11580
rect 38102 11568 38108 11580
rect 38160 11568 38166 11620
rect 38212 11608 38240 11639
rect 38838 11636 38844 11688
rect 38896 11636 38902 11688
rect 39500 11676 39528 11784
rect 43990 11772 43996 11784
rect 44048 11772 44054 11824
rect 40402 11704 40408 11756
rect 40460 11744 40466 11756
rect 41509 11747 41567 11753
rect 41509 11744 41521 11747
rect 40460 11716 41521 11744
rect 40460 11704 40466 11716
rect 41509 11713 41521 11716
rect 41555 11713 41567 11747
rect 41509 11707 41567 11713
rect 41785 11747 41843 11753
rect 41785 11713 41797 11747
rect 41831 11744 41843 11747
rect 42058 11744 42064 11756
rect 41831 11716 42064 11744
rect 41831 11713 41843 11716
rect 41785 11707 41843 11713
rect 42058 11704 42064 11716
rect 42116 11704 42122 11756
rect 43162 11704 43168 11756
rect 43220 11744 43226 11756
rect 43349 11747 43407 11753
rect 43349 11744 43361 11747
rect 43220 11716 43361 11744
rect 43220 11704 43226 11716
rect 43349 11713 43361 11716
rect 43395 11713 43407 11747
rect 43349 11707 43407 11713
rect 43530 11704 43536 11756
rect 43588 11704 43594 11756
rect 43622 11704 43628 11756
rect 43680 11744 43686 11756
rect 44085 11747 44143 11753
rect 44085 11744 44097 11747
rect 43680 11716 44097 11744
rect 43680 11704 43686 11716
rect 44085 11713 44097 11716
rect 44131 11713 44143 11747
rect 44085 11707 44143 11713
rect 39040 11648 39528 11676
rect 38933 11611 38991 11617
rect 38933 11608 38945 11611
rect 38212 11580 38945 11608
rect 38933 11577 38945 11580
rect 38979 11608 38991 11611
rect 39040 11608 39068 11648
rect 42426 11636 42432 11688
rect 42484 11636 42490 11688
rect 42797 11679 42855 11685
rect 42797 11645 42809 11679
rect 42843 11676 42855 11679
rect 42978 11676 42984 11688
rect 42843 11648 42984 11676
rect 42843 11645 42855 11648
rect 42797 11639 42855 11645
rect 42812 11608 42840 11639
rect 42978 11636 42984 11648
rect 43036 11636 43042 11688
rect 43254 11636 43260 11688
rect 43312 11636 43318 11688
rect 43438 11636 43444 11688
rect 43496 11636 43502 11688
rect 43990 11636 43996 11688
rect 44048 11636 44054 11688
rect 44453 11679 44511 11685
rect 44453 11645 44465 11679
rect 44499 11676 44511 11679
rect 44910 11676 44916 11688
rect 44499 11648 44916 11676
rect 44499 11645 44511 11648
rect 44453 11639 44511 11645
rect 44910 11636 44916 11648
rect 44968 11636 44974 11688
rect 43346 11608 43352 11620
rect 38979 11580 39068 11608
rect 39408 11580 42840 11608
rect 42996 11580 43352 11608
rect 38979 11577 38991 11580
rect 38933 11571 38991 11577
rect 37829 11543 37887 11549
rect 37829 11509 37841 11543
rect 37875 11509 37887 11543
rect 37829 11503 37887 11509
rect 38562 11500 38568 11552
rect 38620 11540 38626 11552
rect 39408 11540 39436 11580
rect 38620 11512 39436 11540
rect 39485 11543 39543 11549
rect 38620 11500 38626 11512
rect 39485 11509 39497 11543
rect 39531 11540 39543 11543
rect 40034 11540 40040 11552
rect 39531 11512 40040 11540
rect 39531 11509 39543 11512
rect 39485 11503 39543 11509
rect 40034 11500 40040 11512
rect 40092 11500 40098 11552
rect 41892 11549 41920 11580
rect 41877 11543 41935 11549
rect 41877 11509 41889 11543
rect 41923 11509 41935 11543
rect 41877 11503 41935 11509
rect 42702 11500 42708 11552
rect 42760 11540 42766 11552
rect 42996 11549 43024 11580
rect 43346 11568 43352 11580
rect 43404 11568 43410 11620
rect 42981 11543 43039 11549
rect 42981 11540 42993 11543
rect 42760 11512 42993 11540
rect 42760 11500 42766 11512
rect 42981 11509 42993 11512
rect 43027 11509 43039 11543
rect 42981 11503 43039 11509
rect 43070 11500 43076 11552
rect 43128 11500 43134 11552
rect 1104 11450 47104 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 47104 11450
rect 1104 11376 47104 11398
rect 6730 11296 6736 11348
rect 6788 11296 6794 11348
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 9364 11308 9413 11336
rect 9364 11296 9370 11308
rect 9401 11305 9413 11308
rect 9447 11305 9459 11339
rect 9401 11299 9459 11305
rect 13541 11339 13599 11345
rect 13541 11305 13553 11339
rect 13587 11336 13599 11339
rect 23198 11336 23204 11348
rect 13587 11308 23204 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 23198 11296 23204 11308
rect 23256 11296 23262 11348
rect 23845 11339 23903 11345
rect 23845 11305 23857 11339
rect 23891 11336 23903 11339
rect 23934 11336 23940 11348
rect 23891 11308 23940 11336
rect 23891 11305 23903 11308
rect 23845 11299 23903 11305
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 26513 11339 26571 11345
rect 26513 11336 26525 11339
rect 25700 11308 26525 11336
rect 15473 11271 15531 11277
rect 15473 11237 15485 11271
rect 15519 11237 15531 11271
rect 15473 11231 15531 11237
rect 3694 11160 3700 11212
rect 3752 11200 3758 11212
rect 5353 11203 5411 11209
rect 5353 11200 5365 11203
rect 3752 11172 5365 11200
rect 3752 11160 3758 11172
rect 5353 11169 5365 11172
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 5368 11064 5396 11163
rect 7558 11160 7564 11212
rect 7616 11200 7622 11212
rect 10962 11200 10968 11212
rect 7616 11172 10968 11200
rect 7616 11160 7622 11172
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 12897 11203 12955 11209
rect 12897 11200 12909 11203
rect 12492 11172 12909 11200
rect 12492 11160 12498 11172
rect 12897 11169 12909 11172
rect 12943 11169 12955 11203
rect 12897 11163 12955 11169
rect 14458 11160 14464 11212
rect 14516 11160 14522 11212
rect 14553 11203 14611 11209
rect 14553 11169 14565 11203
rect 14599 11200 14611 11203
rect 14734 11200 14740 11212
rect 14599 11172 14740 11200
rect 14599 11169 14611 11172
rect 14553 11163 14611 11169
rect 5626 11141 5632 11144
rect 5620 11132 5632 11141
rect 5587 11104 5632 11132
rect 5620 11095 5632 11104
rect 5626 11092 5632 11095
rect 5684 11092 5690 11144
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11132 9643 11135
rect 10502 11132 10508 11144
rect 9631 11104 10508 11132
rect 9631 11101 9643 11104
rect 9585 11095 9643 11101
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 13265 11135 13323 11141
rect 13265 11132 13277 11135
rect 12860 11104 13277 11132
rect 12860 11092 12866 11104
rect 13265 11101 13277 11104
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 13538 11132 13544 11144
rect 13403 11104 13544 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 13538 11092 13544 11104
rect 13596 11132 13602 11144
rect 14568 11132 14596 11163
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 13596 11104 14596 11132
rect 15381 11135 15439 11141
rect 13596 11092 13602 11104
rect 15381 11101 15393 11135
rect 15427 11132 15439 11135
rect 15488 11132 15516 11231
rect 19702 11228 19708 11280
rect 19760 11268 19766 11280
rect 20073 11271 20131 11277
rect 20073 11268 20085 11271
rect 19760 11240 20085 11268
rect 19760 11228 19766 11240
rect 20073 11237 20085 11240
rect 20119 11237 20131 11271
rect 20073 11231 20131 11237
rect 25130 11228 25136 11280
rect 25188 11228 25194 11280
rect 16117 11203 16175 11209
rect 16117 11169 16129 11203
rect 16163 11200 16175 11203
rect 16482 11200 16488 11212
rect 16163 11172 16488 11200
rect 16163 11169 16175 11172
rect 16117 11163 16175 11169
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 18141 11203 18199 11209
rect 18141 11169 18153 11203
rect 18187 11200 18199 11203
rect 19334 11200 19340 11212
rect 18187 11172 19340 11200
rect 18187 11169 18199 11172
rect 18141 11163 18199 11169
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 19794 11160 19800 11212
rect 19852 11200 19858 11212
rect 20162 11200 20168 11212
rect 19852 11172 20168 11200
rect 19852 11160 19858 11172
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 24857 11203 24915 11209
rect 24857 11169 24869 11203
rect 24903 11200 24915 11203
rect 25038 11200 25044 11212
rect 24903 11172 25044 11200
rect 24903 11169 24915 11172
rect 24857 11163 24915 11169
rect 25038 11160 25044 11172
rect 25096 11160 25102 11212
rect 25700 11200 25728 11308
rect 26513 11305 26525 11308
rect 26559 11305 26571 11339
rect 26513 11299 26571 11305
rect 29270 11296 29276 11348
rect 29328 11336 29334 11348
rect 30009 11339 30067 11345
rect 30009 11336 30021 11339
rect 29328 11308 30021 11336
rect 29328 11296 29334 11308
rect 30009 11305 30021 11308
rect 30055 11305 30067 11339
rect 30009 11299 30067 11305
rect 31570 11296 31576 11348
rect 31628 11336 31634 11348
rect 32217 11339 32275 11345
rect 32217 11336 32229 11339
rect 31628 11308 32229 11336
rect 31628 11296 31634 11308
rect 32217 11305 32229 11308
rect 32263 11305 32275 11339
rect 32217 11299 32275 11305
rect 34149 11339 34207 11345
rect 34149 11305 34161 11339
rect 34195 11336 34207 11339
rect 34330 11336 34336 11348
rect 34195 11308 34336 11336
rect 34195 11305 34207 11308
rect 34149 11299 34207 11305
rect 34330 11296 34336 11308
rect 34388 11296 34394 11348
rect 36906 11336 36912 11348
rect 35636 11308 36912 11336
rect 25866 11228 25872 11280
rect 25924 11228 25930 11280
rect 26326 11228 26332 11280
rect 26384 11228 26390 11280
rect 29822 11268 29828 11280
rect 26804 11240 29828 11268
rect 25608 11172 25728 11200
rect 15427 11104 15516 11132
rect 15427 11101 15439 11104
rect 15381 11095 15439 11101
rect 15930 11092 15936 11144
rect 15988 11092 15994 11144
rect 17310 11092 17316 11144
rect 17368 11132 17374 11144
rect 17957 11135 18015 11141
rect 17957 11132 17969 11135
rect 17368 11104 17969 11132
rect 17368 11092 17374 11104
rect 17957 11101 17969 11104
rect 18003 11101 18015 11135
rect 17957 11095 18015 11101
rect 22462 11092 22468 11144
rect 22520 11132 22526 11144
rect 24486 11132 24492 11144
rect 22520 11104 24492 11132
rect 22520 11092 22526 11104
rect 24486 11092 24492 11104
rect 24544 11092 24550 11144
rect 25608 11141 25636 11172
rect 26050 11160 26056 11212
rect 26108 11200 26114 11212
rect 26108 11172 26740 11200
rect 26108 11160 26114 11172
rect 25593 11135 25651 11141
rect 25593 11101 25605 11135
rect 25639 11101 25651 11135
rect 25593 11095 25651 11101
rect 25685 11135 25743 11141
rect 25685 11101 25697 11135
rect 25731 11101 25743 11135
rect 25685 11095 25743 11101
rect 6178 11064 6184 11076
rect 5368 11036 6184 11064
rect 6178 11024 6184 11036
rect 6236 11024 6242 11076
rect 8846 11024 8852 11076
rect 8904 11064 8910 11076
rect 10042 11064 10048 11076
rect 8904 11036 10048 11064
rect 8904 11024 8910 11036
rect 10042 11024 10048 11036
rect 10100 11024 10106 11076
rect 10873 11067 10931 11073
rect 10873 11033 10885 11067
rect 10919 11064 10931 11067
rect 10962 11064 10968 11076
rect 10919 11036 10968 11064
rect 10919 11033 10931 11036
rect 10873 11027 10931 11033
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 13630 11064 13636 11076
rect 13504 11036 13636 11064
rect 13504 11024 13510 11036
rect 13630 11024 13636 11036
rect 13688 11064 13694 11076
rect 14093 11067 14151 11073
rect 14093 11064 14105 11067
rect 13688 11036 14105 11064
rect 13688 11024 13694 11036
rect 14093 11033 14105 11036
rect 14139 11033 14151 11067
rect 14093 11027 14151 11033
rect 14737 11067 14795 11073
rect 14737 11033 14749 11067
rect 14783 11064 14795 11067
rect 16298 11064 16304 11076
rect 14783 11036 16304 11064
rect 14783 11033 14795 11036
rect 14737 11027 14795 11033
rect 16298 11024 16304 11036
rect 16356 11024 16362 11076
rect 17865 11067 17923 11073
rect 17865 11033 17877 11067
rect 17911 11064 17923 11067
rect 18046 11064 18052 11076
rect 17911 11036 18052 11064
rect 17911 11033 17923 11036
rect 17865 11027 17923 11033
rect 18046 11024 18052 11036
rect 18104 11024 18110 11076
rect 22732 11067 22790 11073
rect 22732 11033 22744 11067
rect 22778 11064 22790 11067
rect 22830 11064 22836 11076
rect 22778 11036 22836 11064
rect 22778 11033 22790 11036
rect 22732 11027 22790 11033
rect 22830 11024 22836 11036
rect 22888 11024 22894 11076
rect 25406 11024 25412 11076
rect 25464 11024 25470 11076
rect 25700 11064 25728 11095
rect 25866 11092 25872 11144
rect 25924 11132 25930 11144
rect 25961 11135 26019 11141
rect 25961 11132 25973 11135
rect 25924 11104 25973 11132
rect 25924 11092 25930 11104
rect 25961 11101 25973 11104
rect 26007 11101 26019 11135
rect 25961 11095 26019 11101
rect 26605 11067 26663 11073
rect 26605 11064 26617 11067
rect 25700 11036 26004 11064
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 10413 10999 10471 11005
rect 10413 10996 10425 10999
rect 9732 10968 10425 10996
rect 9732 10956 9738 10968
rect 10413 10965 10425 10968
rect 10459 10965 10471 10999
rect 10413 10959 10471 10965
rect 10778 10956 10784 11008
rect 10836 10956 10842 11008
rect 15194 10956 15200 11008
rect 15252 10956 15258 11008
rect 15838 10956 15844 11008
rect 15896 10956 15902 11008
rect 17497 10999 17555 11005
rect 17497 10965 17509 10999
rect 17543 10996 17555 10999
rect 17770 10996 17776 11008
rect 17543 10968 17776 10996
rect 17543 10965 17555 10968
rect 17497 10959 17555 10965
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 20254 10956 20260 11008
rect 20312 10956 20318 11008
rect 25317 10999 25375 11005
rect 25317 10965 25329 10999
rect 25363 10996 25375 10999
rect 25866 10996 25872 11008
rect 25363 10968 25872 10996
rect 25363 10965 25375 10968
rect 25317 10959 25375 10965
rect 25866 10956 25872 10968
rect 25924 10956 25930 11008
rect 25976 10996 26004 11036
rect 26160 11036 26617 11064
rect 26160 10996 26188 11036
rect 26605 11033 26617 11036
rect 26651 11033 26663 11067
rect 26712 11064 26740 11172
rect 26804 11141 26832 11240
rect 29822 11228 29828 11240
rect 29880 11228 29886 11280
rect 29917 11271 29975 11277
rect 29917 11237 29929 11271
rect 29963 11268 29975 11271
rect 30466 11268 30472 11280
rect 29963 11240 30472 11268
rect 29963 11237 29975 11240
rect 29917 11231 29975 11237
rect 30466 11228 30472 11240
rect 30524 11228 30530 11280
rect 32493 11271 32551 11277
rect 32493 11237 32505 11271
rect 32539 11237 32551 11271
rect 32493 11231 32551 11237
rect 29549 11203 29607 11209
rect 29549 11200 29561 11203
rect 26896 11172 29561 11200
rect 26789 11135 26847 11141
rect 26789 11101 26801 11135
rect 26835 11101 26847 11135
rect 26789 11095 26847 11101
rect 26896 11064 26924 11172
rect 29549 11169 29561 11172
rect 29595 11169 29607 11203
rect 32508 11200 32536 11231
rect 32508 11172 32904 11200
rect 29549 11163 29607 11169
rect 27065 11135 27123 11141
rect 27065 11101 27077 11135
rect 27111 11132 27123 11135
rect 30374 11132 30380 11144
rect 27111 11104 30380 11132
rect 27111 11101 27123 11104
rect 27065 11095 27123 11101
rect 30374 11092 30380 11104
rect 30432 11092 30438 11144
rect 30837 11135 30895 11141
rect 30837 11101 30849 11135
rect 30883 11132 30895 11135
rect 31662 11132 31668 11144
rect 30883 11104 31668 11132
rect 30883 11101 30895 11104
rect 30837 11095 30895 11101
rect 31662 11092 31668 11104
rect 31720 11132 31726 11144
rect 31720 11104 32628 11132
rect 31720 11092 31726 11104
rect 26712 11036 26924 11064
rect 26973 11067 27031 11073
rect 26605 11027 26663 11033
rect 26973 11033 26985 11067
rect 27019 11064 27031 11067
rect 27430 11064 27436 11076
rect 27019 11036 27436 11064
rect 27019 11033 27031 11036
rect 26973 11027 27031 11033
rect 27430 11024 27436 11036
rect 27488 11024 27494 11076
rect 31104 11067 31162 11073
rect 31104 11033 31116 11067
rect 31150 11064 31162 11067
rect 31202 11064 31208 11076
rect 31150 11036 31208 11064
rect 31150 11033 31162 11036
rect 31104 11027 31162 11033
rect 31202 11024 31208 11036
rect 31260 11024 31266 11076
rect 32600 11064 32628 11104
rect 32674 11092 32680 11144
rect 32732 11092 32738 11144
rect 32769 11135 32827 11141
rect 32769 11101 32781 11135
rect 32815 11101 32827 11135
rect 32876 11132 32904 11172
rect 35342 11160 35348 11212
rect 35400 11200 35406 11212
rect 35636 11209 35664 11308
rect 36906 11296 36912 11308
rect 36964 11296 36970 11348
rect 38197 11339 38255 11345
rect 38197 11305 38209 11339
rect 38243 11336 38255 11339
rect 38746 11336 38752 11348
rect 38243 11308 38752 11336
rect 38243 11305 38255 11308
rect 38197 11299 38255 11305
rect 38746 11296 38752 11308
rect 38804 11336 38810 11348
rect 39022 11336 39028 11348
rect 38804 11308 39028 11336
rect 38804 11296 38810 11308
rect 39022 11296 39028 11308
rect 39080 11296 39086 11348
rect 42518 11296 42524 11348
rect 42576 11336 42582 11348
rect 42797 11339 42855 11345
rect 42797 11336 42809 11339
rect 42576 11308 42809 11336
rect 42576 11296 42582 11308
rect 42797 11305 42809 11308
rect 42843 11305 42855 11339
rect 42797 11299 42855 11305
rect 43349 11339 43407 11345
rect 43349 11305 43361 11339
rect 43395 11336 43407 11339
rect 43438 11336 43444 11348
rect 43395 11308 43444 11336
rect 43395 11305 43407 11308
rect 43349 11299 43407 11305
rect 43438 11296 43444 11308
rect 43496 11296 43502 11348
rect 36633 11271 36691 11277
rect 36633 11237 36645 11271
rect 36679 11268 36691 11271
rect 38562 11268 38568 11280
rect 36679 11240 38568 11268
rect 36679 11237 36691 11240
rect 36633 11231 36691 11237
rect 38562 11228 38568 11240
rect 38620 11228 38626 11280
rect 39482 11268 39488 11280
rect 38672 11240 39488 11268
rect 35621 11203 35679 11209
rect 35621 11200 35633 11203
rect 35400 11172 35633 11200
rect 35400 11160 35406 11172
rect 35621 11169 35633 11172
rect 35667 11169 35679 11203
rect 35621 11163 35679 11169
rect 33025 11135 33083 11141
rect 33025 11132 33037 11135
rect 32876 11104 33037 11132
rect 32769 11095 32827 11101
rect 33025 11101 33037 11104
rect 33071 11101 33083 11135
rect 33025 11095 33083 11101
rect 32784 11064 32812 11095
rect 34422 11092 34428 11144
rect 34480 11092 34486 11144
rect 35894 11092 35900 11144
rect 35952 11092 35958 11144
rect 37734 11092 37740 11144
rect 37792 11092 37798 11144
rect 37918 11092 37924 11144
rect 37976 11132 37982 11144
rect 38197 11135 38255 11141
rect 38197 11132 38209 11135
rect 37976 11104 38209 11132
rect 37976 11092 37982 11104
rect 38197 11101 38209 11104
rect 38243 11101 38255 11135
rect 38197 11095 38255 11101
rect 38378 11092 38384 11144
rect 38436 11092 38442 11144
rect 38672 11132 38700 11240
rect 39482 11228 39488 11240
rect 39540 11228 39546 11280
rect 43990 11268 43996 11280
rect 42996 11240 43996 11268
rect 42996 11200 43024 11240
rect 43990 11228 43996 11240
rect 44048 11268 44054 11280
rect 44269 11271 44327 11277
rect 44269 11268 44281 11271
rect 44048 11240 44281 11268
rect 44048 11228 44054 11240
rect 44269 11237 44281 11240
rect 44315 11237 44327 11271
rect 44269 11231 44327 11237
rect 42536 11172 43024 11200
rect 38749 11135 38807 11141
rect 38749 11132 38761 11135
rect 38672 11104 38761 11132
rect 38749 11101 38761 11104
rect 38795 11101 38807 11135
rect 38749 11095 38807 11101
rect 38838 11092 38844 11144
rect 38896 11092 38902 11144
rect 39114 11092 39120 11144
rect 39172 11092 39178 11144
rect 39209 11135 39267 11141
rect 39209 11101 39221 11135
rect 39255 11101 39267 11135
rect 39209 11095 39267 11101
rect 33226 11064 33232 11076
rect 32600 11036 33232 11064
rect 33226 11024 33232 11036
rect 33284 11024 33290 11076
rect 38105 11067 38163 11073
rect 34072 11036 34376 11064
rect 25976 10968 26188 10996
rect 26234 10956 26240 11008
rect 26292 10996 26298 11008
rect 34072 10996 34100 11036
rect 26292 10968 34100 10996
rect 26292 10956 26298 10968
rect 34238 10956 34244 11008
rect 34296 10956 34302 11008
rect 34348 10996 34376 11036
rect 38105 11033 38117 11067
rect 38151 11064 38163 11067
rect 38856 11064 38884 11092
rect 39224 11064 39252 11095
rect 39298 11092 39304 11144
rect 39356 11141 39362 11144
rect 39356 11135 39405 11141
rect 39356 11101 39359 11135
rect 39393 11101 39405 11135
rect 39356 11095 39405 11101
rect 39669 11135 39727 11141
rect 39669 11101 39681 11135
rect 39715 11132 39727 11135
rect 40770 11132 40776 11144
rect 39715 11104 40776 11132
rect 39715 11101 39727 11104
rect 39669 11095 39727 11101
rect 39356 11092 39362 11095
rect 40770 11092 40776 11104
rect 40828 11092 40834 11144
rect 42536 11141 42564 11172
rect 43622 11160 43628 11212
rect 43680 11200 43686 11212
rect 43901 11203 43959 11209
rect 43901 11200 43913 11203
rect 43680 11172 43913 11200
rect 43680 11160 43686 11172
rect 43901 11169 43913 11172
rect 43947 11169 43959 11203
rect 43901 11163 43959 11169
rect 42521 11135 42579 11141
rect 42521 11101 42533 11135
rect 42567 11101 42579 11135
rect 42521 11095 42579 11101
rect 42610 11092 42616 11144
rect 42668 11132 42674 11144
rect 42705 11135 42763 11141
rect 42705 11132 42717 11135
rect 42668 11104 42717 11132
rect 42668 11092 42674 11104
rect 42705 11101 42717 11104
rect 42751 11101 42763 11135
rect 42705 11095 42763 11101
rect 42794 11092 42800 11144
rect 42852 11132 42858 11144
rect 42981 11135 43039 11141
rect 42981 11132 42993 11135
rect 42852 11104 42993 11132
rect 42852 11092 42858 11104
rect 42981 11101 42993 11104
rect 43027 11101 43039 11135
rect 42981 11095 43039 11101
rect 43162 11092 43168 11144
rect 43220 11092 43226 11144
rect 43257 11135 43315 11141
rect 43257 11101 43269 11135
rect 43303 11134 43315 11135
rect 43303 11106 43392 11134
rect 43303 11101 43315 11106
rect 43257 11095 43315 11101
rect 43180 11064 43208 11092
rect 43364 11076 43392 11106
rect 43530 11092 43536 11144
rect 43588 11092 43594 11144
rect 43809 11135 43867 11141
rect 43809 11101 43821 11135
rect 43855 11132 43867 11135
rect 44085 11135 44143 11141
rect 44085 11132 44097 11135
rect 43855 11104 44097 11132
rect 43855 11101 43867 11104
rect 43809 11095 43867 11101
rect 44085 11101 44097 11104
rect 44131 11101 44143 11135
rect 44085 11095 44143 11101
rect 38151 11036 38792 11064
rect 38856 11036 39252 11064
rect 38151 11033 38163 11036
rect 38105 11027 38163 11033
rect 35434 10996 35440 11008
rect 34348 10968 35440 10996
rect 35434 10956 35440 10968
rect 35492 10956 35498 11008
rect 38378 10956 38384 11008
rect 38436 10996 38442 11008
rect 38565 10999 38623 11005
rect 38565 10996 38577 10999
rect 38436 10968 38577 10996
rect 38436 10956 38442 10968
rect 38565 10965 38577 10968
rect 38611 10965 38623 10999
rect 38764 10996 38792 11036
rect 39114 10996 39120 11008
rect 38764 10968 39120 10996
rect 38565 10959 38623 10965
rect 39114 10956 39120 10968
rect 39172 10956 39178 11008
rect 39224 10996 39252 11036
rect 43088 11036 43208 11064
rect 39390 10996 39396 11008
rect 39224 10968 39396 10996
rect 39390 10956 39396 10968
rect 39448 10956 39454 11008
rect 39574 10956 39580 11008
rect 39632 10956 39638 11008
rect 42705 10999 42763 11005
rect 42705 10965 42717 10999
rect 42751 10996 42763 10999
rect 43088 10996 43116 11036
rect 43346 11024 43352 11076
rect 43404 11064 43410 11076
rect 43824 11064 43852 11095
rect 43404 11036 43852 11064
rect 43404 11024 43410 11036
rect 42751 10968 43116 10996
rect 42751 10965 42763 10968
rect 42705 10959 42763 10965
rect 43162 10956 43168 11008
rect 43220 10996 43226 11008
rect 43622 10996 43628 11008
rect 43220 10968 43628 10996
rect 43220 10956 43226 10968
rect 43622 10956 43628 10968
rect 43680 10996 43686 11008
rect 43717 10999 43775 11005
rect 43717 10996 43729 10999
rect 43680 10968 43729 10996
rect 43680 10956 43686 10968
rect 43717 10965 43729 10968
rect 43763 10965 43775 10999
rect 43717 10959 43775 10965
rect 1104 10906 47104 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 47104 10906
rect 1104 10832 47104 10854
rect 6733 10795 6791 10801
rect 6733 10761 6745 10795
rect 6779 10761 6791 10795
rect 6733 10755 6791 10761
rect 7101 10795 7159 10801
rect 7101 10761 7113 10795
rect 7147 10792 7159 10795
rect 7742 10792 7748 10804
rect 7147 10764 7748 10792
rect 7147 10761 7159 10764
rect 7101 10755 7159 10761
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 6748 10656 6776 10755
rect 7742 10752 7748 10764
rect 7800 10792 7806 10804
rect 8662 10792 8668 10804
rect 7800 10764 8668 10792
rect 7800 10752 7806 10764
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 10778 10752 10784 10804
rect 10836 10792 10842 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 10836 10764 10977 10792
rect 10836 10752 10842 10764
rect 10965 10761 10977 10764
rect 11011 10792 11023 10795
rect 12618 10792 12624 10804
rect 11011 10764 12624 10792
rect 11011 10761 11023 10764
rect 10965 10755 11023 10761
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 14093 10795 14151 10801
rect 14093 10761 14105 10795
rect 14139 10761 14151 10795
rect 14093 10755 14151 10761
rect 6595 10628 6776 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 8662 10616 8668 10668
rect 8720 10665 8726 10668
rect 8720 10659 8748 10665
rect 8736 10625 8748 10659
rect 8720 10619 8748 10625
rect 8720 10616 8726 10619
rect 8846 10616 8852 10668
rect 8904 10616 8910 10668
rect 9490 10616 9496 10668
rect 9548 10656 9554 10668
rect 9841 10659 9899 10665
rect 9841 10656 9853 10659
rect 9548 10628 9853 10656
rect 9548 10616 9554 10628
rect 9841 10625 9853 10628
rect 9887 10625 9899 10659
rect 9841 10619 9899 10625
rect 12710 10616 12716 10668
rect 12768 10616 12774 10668
rect 14001 10659 14059 10665
rect 14001 10625 14013 10659
rect 14047 10656 14059 10659
rect 14108 10656 14136 10755
rect 14182 10752 14188 10804
rect 14240 10792 14246 10804
rect 14553 10795 14611 10801
rect 14553 10792 14565 10795
rect 14240 10764 14565 10792
rect 14240 10752 14246 10764
rect 14553 10761 14565 10764
rect 14599 10792 14611 10795
rect 14599 10764 15332 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 14274 10684 14280 10736
rect 14332 10724 14338 10736
rect 15194 10733 15200 10736
rect 15188 10724 15200 10733
rect 14332 10696 14964 10724
rect 15155 10696 15200 10724
rect 14332 10684 14338 10696
rect 14936 10665 14964 10696
rect 15188 10687 15200 10696
rect 15194 10684 15200 10687
rect 15252 10684 15258 10736
rect 15304 10724 15332 10764
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 15896 10764 16313 10792
rect 15896 10752 15902 10764
rect 16301 10761 16313 10764
rect 16347 10792 16359 10795
rect 18874 10792 18880 10804
rect 16347 10764 18880 10792
rect 16347 10761 16359 10764
rect 16301 10755 16359 10761
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 20806 10752 20812 10804
rect 20864 10792 20870 10804
rect 21177 10795 21235 10801
rect 21177 10792 21189 10795
rect 20864 10764 21189 10792
rect 20864 10752 20870 10764
rect 21177 10761 21189 10764
rect 21223 10761 21235 10795
rect 21177 10755 21235 10761
rect 22830 10752 22836 10804
rect 22888 10752 22894 10804
rect 30466 10752 30472 10804
rect 30524 10752 30530 10804
rect 31202 10752 31208 10804
rect 31260 10752 31266 10804
rect 34146 10752 34152 10804
rect 34204 10792 34210 10804
rect 34609 10795 34667 10801
rect 34609 10792 34621 10795
rect 34204 10764 34621 10792
rect 34204 10752 34210 10764
rect 34609 10761 34621 10764
rect 34655 10761 34667 10795
rect 34609 10755 34667 10761
rect 36725 10795 36783 10801
rect 36725 10761 36737 10795
rect 36771 10792 36783 10795
rect 37918 10792 37924 10804
rect 36771 10764 37924 10792
rect 36771 10761 36783 10764
rect 36725 10755 36783 10761
rect 37918 10752 37924 10764
rect 37976 10752 37982 10804
rect 38289 10795 38347 10801
rect 38289 10761 38301 10795
rect 38335 10792 38347 10795
rect 38838 10792 38844 10804
rect 38335 10764 38844 10792
rect 38335 10761 38347 10764
rect 38289 10755 38347 10761
rect 38838 10752 38844 10764
rect 38896 10752 38902 10804
rect 39117 10795 39175 10801
rect 39117 10761 39129 10795
rect 39163 10792 39175 10795
rect 39298 10792 39304 10804
rect 39163 10764 39304 10792
rect 39163 10761 39175 10764
rect 39117 10755 39175 10761
rect 39298 10752 39304 10764
rect 39356 10752 39362 10804
rect 40402 10752 40408 10804
rect 40460 10792 40466 10804
rect 40589 10795 40647 10801
rect 40589 10792 40601 10795
rect 40460 10764 40601 10792
rect 40460 10752 40466 10764
rect 40589 10761 40601 10764
rect 40635 10792 40647 10795
rect 41046 10792 41052 10804
rect 40635 10764 41052 10792
rect 40635 10761 40647 10764
rect 40589 10755 40647 10761
rect 41046 10752 41052 10764
rect 41104 10792 41110 10804
rect 41233 10795 41291 10801
rect 41233 10792 41245 10795
rect 41104 10764 41245 10792
rect 41104 10752 41110 10764
rect 41233 10761 41245 10764
rect 41279 10761 41291 10795
rect 41233 10755 41291 10761
rect 42426 10752 42432 10804
rect 42484 10792 42490 10804
rect 42484 10764 43208 10792
rect 42484 10752 42490 10764
rect 15930 10724 15936 10736
rect 15304 10696 15936 10724
rect 15930 10684 15936 10696
rect 15988 10684 15994 10736
rect 19705 10727 19763 10733
rect 19705 10693 19717 10727
rect 19751 10724 19763 10727
rect 25130 10724 25136 10736
rect 19751 10696 25136 10724
rect 19751 10693 19763 10696
rect 19705 10687 19763 10693
rect 25130 10684 25136 10696
rect 25188 10684 25194 10736
rect 33496 10727 33554 10733
rect 33496 10693 33508 10727
rect 33542 10724 33554 10727
rect 34238 10724 34244 10736
rect 33542 10696 34244 10724
rect 33542 10693 33554 10696
rect 33496 10687 33554 10693
rect 34238 10684 34244 10696
rect 34296 10684 34302 10736
rect 39574 10724 39580 10736
rect 38488 10696 39580 10724
rect 14047 10628 14136 10656
rect 14461 10659 14519 10665
rect 14047 10625 14059 10628
rect 14001 10619 14059 10625
rect 14461 10625 14473 10659
rect 14507 10625 14519 10659
rect 14461 10619 14519 10625
rect 14921 10659 14979 10665
rect 14921 10625 14933 10659
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 7190 10548 7196 10600
rect 7248 10548 7254 10600
rect 7377 10591 7435 10597
rect 7377 10557 7389 10591
rect 7423 10588 7435 10591
rect 7558 10588 7564 10600
rect 7423 10560 7564 10588
rect 7423 10557 7435 10560
rect 7377 10551 7435 10557
rect 7558 10548 7564 10560
rect 7616 10548 7622 10600
rect 7650 10548 7656 10600
rect 7708 10548 7714 10600
rect 7834 10548 7840 10600
rect 7892 10548 7898 10600
rect 8294 10548 8300 10600
rect 8352 10548 8358 10600
rect 8570 10548 8576 10600
rect 8628 10548 8634 10600
rect 9030 10548 9036 10600
rect 9088 10588 9094 10600
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 9088 10560 9597 10588
rect 9088 10548 9094 10560
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 11296 10560 11529 10588
rect 11296 10548 11302 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 11606 10548 11612 10600
rect 11664 10588 11670 10600
rect 11701 10591 11759 10597
rect 11701 10588 11713 10591
rect 11664 10560 11713 10588
rect 11664 10548 11670 10560
rect 11701 10557 11713 10560
rect 11747 10557 11759 10591
rect 11701 10551 11759 10557
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 12250 10588 12256 10600
rect 12207 10560 12256 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 12250 10548 12256 10560
rect 12308 10548 12314 10600
rect 12434 10548 12440 10600
rect 12492 10548 12498 10600
rect 12618 10597 12624 10600
rect 12575 10591 12624 10597
rect 12575 10557 12587 10591
rect 12621 10557 12624 10591
rect 12575 10551 12624 10557
rect 12618 10548 12624 10551
rect 12676 10548 12682 10600
rect 6362 10412 6368 10464
rect 6420 10412 6426 10464
rect 9493 10455 9551 10461
rect 9493 10421 9505 10455
rect 9539 10452 9551 10455
rect 12802 10452 12808 10464
rect 9539 10424 12808 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13357 10455 13415 10461
rect 13357 10421 13369 10455
rect 13403 10452 13415 10455
rect 13630 10452 13636 10464
rect 13403 10424 13636 10452
rect 13403 10421 13415 10424
rect 13357 10415 13415 10421
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 13817 10455 13875 10461
rect 13817 10421 13829 10455
rect 13863 10452 13875 10455
rect 14182 10452 14188 10464
rect 13863 10424 14188 10452
rect 13863 10421 13875 10424
rect 13817 10415 13875 10421
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 14476 10452 14504 10619
rect 15010 10616 15016 10668
rect 15068 10616 15074 10668
rect 17310 10616 17316 10668
rect 17368 10616 17374 10668
rect 17770 10616 17776 10668
rect 17828 10616 17834 10668
rect 18046 10616 18052 10668
rect 18104 10616 18110 10668
rect 18874 10616 18880 10668
rect 18932 10665 18938 10668
rect 18932 10659 18960 10665
rect 18948 10625 18960 10659
rect 18932 10619 18960 10625
rect 18932 10616 18938 10619
rect 19058 10616 19064 10668
rect 19116 10616 19122 10668
rect 20070 10616 20076 10668
rect 20128 10656 20134 10668
rect 20441 10659 20499 10665
rect 20441 10656 20453 10659
rect 20128 10628 20453 10656
rect 20128 10616 20134 10628
rect 20441 10625 20453 10628
rect 20487 10625 20499 10659
rect 20441 10619 20499 10625
rect 23014 10616 23020 10668
rect 23072 10616 23078 10668
rect 28629 10659 28687 10665
rect 28629 10625 28641 10659
rect 28675 10656 28687 10659
rect 28994 10656 29000 10668
rect 28675 10628 29000 10656
rect 28675 10625 28687 10628
rect 28629 10619 28687 10625
rect 28994 10616 29000 10628
rect 29052 10616 29058 10668
rect 29638 10616 29644 10668
rect 29696 10665 29702 10668
rect 29696 10659 29724 10665
rect 29712 10625 29724 10659
rect 29696 10619 29724 10625
rect 29696 10616 29702 10619
rect 29822 10616 29828 10668
rect 29880 10616 29886 10668
rect 31386 10616 31392 10668
rect 31444 10616 31450 10668
rect 33226 10616 33232 10668
rect 33284 10656 33290 10668
rect 34606 10656 34612 10668
rect 33284 10628 34612 10656
rect 33284 10616 33290 10628
rect 34606 10616 34612 10628
rect 34664 10616 34670 10668
rect 35342 10616 35348 10668
rect 35400 10656 35406 10668
rect 35713 10659 35771 10665
rect 35713 10656 35725 10659
rect 35400 10628 35725 10656
rect 35400 10616 35406 10628
rect 35713 10625 35725 10628
rect 35759 10625 35771 10659
rect 35713 10619 35771 10625
rect 35986 10616 35992 10668
rect 36044 10616 36050 10668
rect 37826 10616 37832 10668
rect 37884 10656 37890 10668
rect 37921 10659 37979 10665
rect 37921 10656 37933 10659
rect 37884 10628 37933 10656
rect 37884 10616 37890 10628
rect 37921 10625 37933 10628
rect 37967 10625 37979 10659
rect 37921 10619 37979 10625
rect 38102 10616 38108 10668
rect 38160 10616 38166 10668
rect 38378 10616 38384 10668
rect 38436 10616 38442 10668
rect 38488 10665 38516 10696
rect 39574 10684 39580 10696
rect 39632 10684 39638 10736
rect 40221 10727 40279 10733
rect 40221 10693 40233 10727
rect 40267 10724 40279 10727
rect 40494 10724 40500 10736
rect 40267 10696 40500 10724
rect 40267 10693 40279 10696
rect 40221 10687 40279 10693
rect 40494 10684 40500 10696
rect 40552 10724 40558 10736
rect 42797 10727 42855 10733
rect 42797 10724 42809 10727
rect 40552 10696 42809 10724
rect 40552 10684 40558 10696
rect 42797 10693 42809 10696
rect 42843 10693 42855 10727
rect 42797 10687 42855 10693
rect 42981 10727 43039 10733
rect 42981 10693 42993 10727
rect 43027 10724 43039 10727
rect 43070 10724 43076 10736
rect 43027 10696 43076 10724
rect 43027 10693 43039 10696
rect 42981 10687 43039 10693
rect 43070 10684 43076 10696
rect 43128 10684 43134 10736
rect 38473 10659 38531 10665
rect 38473 10625 38485 10659
rect 38519 10625 38531 10659
rect 38473 10619 38531 10625
rect 38746 10616 38752 10668
rect 38804 10616 38810 10668
rect 38933 10659 38991 10665
rect 38933 10625 38945 10659
rect 38979 10656 38991 10659
rect 39114 10656 39120 10668
rect 38979 10628 39120 10656
rect 38979 10625 38991 10628
rect 38933 10619 38991 10625
rect 39114 10616 39120 10628
rect 39172 10616 39178 10668
rect 40034 10616 40040 10668
rect 40092 10616 40098 10668
rect 40313 10659 40371 10665
rect 40313 10625 40325 10659
rect 40359 10625 40371 10659
rect 40313 10619 40371 10625
rect 14737 10591 14795 10597
rect 14737 10557 14749 10591
rect 14783 10588 14795 10591
rect 15028 10588 15056 10616
rect 14783 10560 15056 10588
rect 14783 10557 14795 10560
rect 14737 10551 14795 10557
rect 15930 10548 15936 10600
rect 15988 10588 15994 10600
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 15988 10560 17509 10588
rect 15988 10548 15994 10560
rect 17497 10557 17509 10560
rect 17543 10557 17555 10591
rect 17497 10551 17555 10557
rect 17862 10548 17868 10600
rect 17920 10548 17926 10600
rect 18782 10588 18788 10600
rect 18616 10560 18788 10588
rect 17586 10480 17592 10532
rect 17644 10480 17650 10532
rect 17678 10480 17684 10532
rect 17736 10520 17742 10532
rect 18509 10523 18567 10529
rect 18509 10520 18521 10523
rect 17736 10492 18521 10520
rect 17736 10480 17742 10492
rect 18509 10489 18521 10492
rect 18555 10489 18567 10523
rect 18509 10483 18567 10489
rect 15286 10452 15292 10464
rect 14476 10424 15292 10452
rect 15286 10412 15292 10424
rect 15344 10452 15350 10464
rect 18616 10452 18644 10560
rect 18782 10548 18788 10560
rect 18840 10548 18846 10600
rect 19886 10548 19892 10600
rect 19944 10588 19950 10600
rect 20165 10591 20223 10597
rect 20165 10588 20177 10591
rect 19944 10560 20177 10588
rect 19944 10548 19950 10560
rect 20165 10557 20177 10560
rect 20211 10557 20223 10591
rect 20165 10551 20223 10557
rect 28813 10591 28871 10597
rect 28813 10557 28825 10591
rect 28859 10588 28871 10591
rect 29178 10588 29184 10600
rect 28859 10560 29184 10588
rect 28859 10557 28871 10560
rect 28813 10551 28871 10557
rect 29178 10548 29184 10560
rect 29236 10548 29242 10600
rect 29273 10591 29331 10597
rect 29273 10557 29285 10591
rect 29319 10588 29331 10591
rect 29362 10588 29368 10600
rect 29319 10560 29368 10588
rect 29319 10557 29331 10560
rect 29273 10551 29331 10557
rect 29362 10548 29368 10560
rect 29420 10548 29426 10600
rect 29546 10548 29552 10600
rect 29604 10548 29610 10600
rect 38654 10548 38660 10600
rect 38712 10548 38718 10600
rect 40328 10532 40356 10619
rect 40402 10616 40408 10668
rect 40460 10616 40466 10668
rect 40681 10659 40739 10665
rect 40681 10625 40693 10659
rect 40727 10656 40739 10659
rect 40770 10656 40776 10668
rect 40727 10628 40776 10656
rect 40727 10625 40739 10628
rect 40681 10619 40739 10625
rect 40770 10616 40776 10628
rect 40828 10616 40834 10668
rect 41049 10659 41107 10665
rect 41049 10656 41061 10659
rect 40880 10628 41061 10656
rect 22002 10520 22008 10532
rect 21192 10492 22008 10520
rect 15344 10424 18644 10452
rect 15344 10412 15350 10424
rect 20530 10412 20536 10464
rect 20588 10452 20594 10464
rect 21192 10452 21220 10492
rect 22002 10480 22008 10492
rect 22060 10480 22066 10532
rect 38378 10480 38384 10532
rect 38436 10520 38442 10532
rect 38565 10523 38623 10529
rect 38565 10520 38577 10523
rect 38436 10492 38577 10520
rect 38436 10480 38442 10492
rect 38565 10489 38577 10492
rect 38611 10489 38623 10523
rect 38565 10483 38623 10489
rect 39482 10480 39488 10532
rect 39540 10520 39546 10532
rect 40037 10523 40095 10529
rect 40037 10520 40049 10523
rect 39540 10492 40049 10520
rect 39540 10480 39546 10492
rect 40037 10489 40049 10492
rect 40083 10489 40095 10523
rect 40037 10483 40095 10489
rect 40310 10480 40316 10532
rect 40368 10520 40374 10532
rect 40405 10523 40463 10529
rect 40405 10520 40417 10523
rect 40368 10492 40417 10520
rect 40368 10480 40374 10492
rect 40405 10489 40417 10492
rect 40451 10489 40463 10523
rect 40405 10483 40463 10489
rect 20588 10424 21220 10452
rect 20588 10412 20594 10424
rect 21266 10412 21272 10464
rect 21324 10452 21330 10464
rect 31478 10452 31484 10464
rect 21324 10424 31484 10452
rect 21324 10412 21330 10424
rect 31478 10412 31484 10424
rect 31536 10412 31542 10464
rect 38286 10412 38292 10464
rect 38344 10452 38350 10464
rect 40880 10452 40908 10628
rect 41049 10625 41061 10628
rect 41095 10625 41107 10659
rect 41049 10619 41107 10625
rect 42705 10659 42763 10665
rect 42705 10625 42717 10659
rect 42751 10625 42763 10659
rect 42705 10619 42763 10625
rect 42720 10520 42748 10619
rect 42886 10616 42892 10668
rect 42944 10616 42950 10668
rect 43180 10665 43208 10764
rect 43346 10752 43352 10804
rect 43404 10752 43410 10804
rect 43622 10752 43628 10804
rect 43680 10801 43686 10804
rect 43680 10795 43699 10801
rect 43687 10761 43699 10795
rect 43680 10755 43699 10761
rect 43680 10752 43686 10755
rect 43438 10684 43444 10736
rect 43496 10684 43502 10736
rect 43165 10659 43223 10665
rect 43165 10625 43177 10659
rect 43211 10656 43223 10659
rect 44174 10656 44180 10668
rect 43211 10628 44180 10656
rect 43211 10625 43223 10628
rect 43165 10619 43223 10625
rect 44174 10616 44180 10628
rect 44232 10616 44238 10668
rect 46474 10616 46480 10668
rect 46532 10616 46538 10668
rect 43809 10523 43867 10529
rect 43809 10520 43821 10523
rect 42720 10492 43821 10520
rect 43809 10489 43821 10492
rect 43855 10489 43867 10523
rect 43809 10483 43867 10489
rect 38344 10424 40908 10452
rect 38344 10412 38350 10424
rect 43346 10412 43352 10464
rect 43404 10452 43410 10464
rect 43625 10455 43683 10461
rect 43625 10452 43637 10455
rect 43404 10424 43637 10452
rect 43404 10412 43410 10424
rect 43625 10421 43637 10424
rect 43671 10421 43683 10455
rect 43625 10415 43683 10421
rect 46658 10412 46664 10464
rect 46716 10412 46722 10464
rect 1104 10362 47104 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 47104 10362
rect 1104 10288 47104 10310
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 6104 10220 7665 10248
rect 6104 10053 6132 10220
rect 7653 10217 7665 10220
rect 7699 10217 7711 10251
rect 8478 10248 8484 10260
rect 7653 10211 7711 10217
rect 8128 10220 8484 10248
rect 6178 10072 6184 10124
rect 6236 10072 6242 10124
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 8128 10121 8156 10220
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 9217 10251 9275 10257
rect 9217 10217 9229 10251
rect 9263 10248 9275 10251
rect 9490 10248 9496 10260
rect 9263 10220 9496 10248
rect 9263 10217 9275 10220
rect 9217 10211 9275 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 10410 10248 10416 10260
rect 9600 10220 10416 10248
rect 9600 10180 9628 10220
rect 10410 10208 10416 10220
rect 10468 10208 10474 10260
rect 13909 10251 13967 10257
rect 13909 10217 13921 10251
rect 13955 10248 13967 10251
rect 13955 10220 18000 10248
rect 13955 10217 13967 10220
rect 13909 10211 13967 10217
rect 8220 10152 9628 10180
rect 8220 10121 8248 10152
rect 9674 10140 9680 10192
rect 9732 10140 9738 10192
rect 11885 10183 11943 10189
rect 11885 10180 11897 10183
rect 10796 10152 11897 10180
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 7248 10084 8125 10112
rect 7248 10072 7254 10084
rect 8113 10081 8125 10084
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10081 8263 10115
rect 9692 10112 9720 10140
rect 8205 10075 8263 10081
rect 9416 10084 9720 10112
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10013 6147 10047
rect 6089 10007 6147 10013
rect 6270 10004 6276 10056
rect 6328 10044 6334 10056
rect 8220 10044 8248 10075
rect 9416 10053 9444 10084
rect 6328 10016 8248 10044
rect 9401 10047 9459 10053
rect 6328 10004 6334 10016
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 9674 10004 9680 10056
rect 9732 10004 9738 10056
rect 9769 10047 9827 10053
rect 9769 10013 9781 10047
rect 9815 10044 9827 10047
rect 9815 10016 10180 10044
rect 9815 10013 9827 10016
rect 9769 10007 9827 10013
rect 10152 9988 10180 10016
rect 1489 9979 1547 9985
rect 1489 9945 1501 9979
rect 1535 9976 1547 9979
rect 2222 9976 2228 9988
rect 1535 9948 2228 9976
rect 1535 9945 1547 9948
rect 1489 9939 1547 9945
rect 2222 9936 2228 9948
rect 2280 9936 2286 9988
rect 6426 9979 6484 9985
rect 6426 9976 6438 9979
rect 5920 9948 6438 9976
rect 1578 9868 1584 9920
rect 1636 9868 1642 9920
rect 5920 9917 5948 9948
rect 6426 9945 6438 9948
rect 6472 9945 6484 9979
rect 6426 9939 6484 9945
rect 8021 9979 8079 9985
rect 8021 9945 8033 9979
rect 8067 9976 8079 9979
rect 8570 9976 8576 9988
rect 8067 9948 8576 9976
rect 8067 9945 8079 9948
rect 8021 9939 8079 9945
rect 5905 9911 5963 9917
rect 5905 9877 5917 9911
rect 5951 9877 5963 9911
rect 5905 9871 5963 9877
rect 7561 9911 7619 9917
rect 7561 9877 7573 9911
rect 7607 9908 7619 9911
rect 8036 9908 8064 9939
rect 8570 9936 8576 9948
rect 8628 9976 8634 9988
rect 8846 9976 8852 9988
rect 8628 9948 8852 9976
rect 8628 9936 8634 9948
rect 8846 9936 8852 9948
rect 8904 9936 8910 9988
rect 10014 9979 10072 9985
rect 10014 9976 10026 9979
rect 9508 9948 10026 9976
rect 9508 9917 9536 9948
rect 10014 9945 10026 9948
rect 10060 9945 10072 9979
rect 10014 9939 10072 9945
rect 10134 9936 10140 9988
rect 10192 9936 10198 9988
rect 7607 9880 8064 9908
rect 9493 9911 9551 9917
rect 7607 9877 7619 9880
rect 7561 9871 7619 9877
rect 9493 9877 9505 9911
rect 9539 9877 9551 9911
rect 9493 9871 9551 9877
rect 9582 9868 9588 9920
rect 9640 9908 9646 9920
rect 10796 9908 10824 10152
rect 11885 10149 11897 10152
rect 11931 10149 11943 10183
rect 11885 10143 11943 10149
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 15473 10183 15531 10189
rect 15473 10180 15485 10183
rect 15344 10152 15485 10180
rect 15344 10140 15350 10152
rect 15473 10149 15485 10152
rect 15519 10149 15531 10183
rect 17972 10180 18000 10220
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 18325 10251 18383 10257
rect 18325 10248 18337 10251
rect 18104 10220 18337 10248
rect 18104 10208 18110 10220
rect 18325 10217 18337 10220
rect 18371 10217 18383 10251
rect 18325 10211 18383 10217
rect 20070 10208 20076 10260
rect 20128 10208 20134 10260
rect 20254 10208 20260 10260
rect 20312 10248 20318 10260
rect 20533 10251 20591 10257
rect 20533 10248 20545 10251
rect 20312 10220 20545 10248
rect 20312 10208 20318 10220
rect 20533 10217 20545 10220
rect 20579 10217 20591 10251
rect 20533 10211 20591 10217
rect 20717 10251 20775 10257
rect 20717 10217 20729 10251
rect 20763 10248 20775 10251
rect 37366 10248 37372 10260
rect 20763 10220 34192 10248
rect 20763 10217 20775 10220
rect 20717 10211 20775 10217
rect 22649 10183 22707 10189
rect 17972 10152 21312 10180
rect 15473 10143 15531 10149
rect 11238 10072 11244 10124
rect 11296 10072 11302 10124
rect 11425 10115 11483 10121
rect 11425 10081 11437 10115
rect 11471 10112 11483 10115
rect 11606 10112 11612 10124
rect 11471 10084 11612 10112
rect 11471 10081 11483 10084
rect 11425 10075 11483 10081
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 12299 10115 12357 10121
rect 12299 10081 12311 10115
rect 12345 10112 12357 10115
rect 12618 10112 12624 10124
rect 12345 10084 12624 10112
rect 12345 10081 12357 10084
rect 12299 10075 12357 10081
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10112 13323 10115
rect 13446 10112 13452 10124
rect 13311 10084 13452 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 13630 10072 13636 10124
rect 13688 10072 13694 10124
rect 14090 10072 14096 10124
rect 14148 10072 14154 10124
rect 20530 10112 20536 10124
rect 20272 10084 20536 10112
rect 12158 10004 12164 10056
rect 12216 10004 12222 10056
rect 12434 10004 12440 10056
rect 12492 10004 12498 10056
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 13725 10047 13783 10053
rect 13725 10044 13737 10047
rect 13596 10016 13737 10044
rect 13596 10004 13602 10016
rect 13725 10013 13737 10016
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 14349 10047 14407 10053
rect 14349 10044 14361 10047
rect 14240 10016 14361 10044
rect 14240 10004 14246 10016
rect 14349 10013 14361 10016
rect 14395 10013 14407 10047
rect 14349 10007 14407 10013
rect 16666 10004 16672 10056
rect 16724 10044 16730 10056
rect 16945 10047 17003 10053
rect 16945 10044 16957 10047
rect 16724 10016 16957 10044
rect 16724 10004 16730 10016
rect 16945 10013 16957 10016
rect 16991 10044 17003 10047
rect 17034 10044 17040 10056
rect 16991 10016 17040 10044
rect 16991 10013 17003 10016
rect 16945 10007 17003 10013
rect 17034 10004 17040 10016
rect 17092 10004 17098 10056
rect 17212 10047 17270 10053
rect 17212 10013 17224 10047
rect 17258 10044 17270 10047
rect 17586 10044 17592 10056
rect 17258 10016 17592 10044
rect 17258 10013 17270 10016
rect 17212 10007 17270 10013
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 19426 10004 19432 10056
rect 19484 10044 19490 10056
rect 20272 10053 20300 10084
rect 20530 10072 20536 10084
rect 20588 10112 20594 10124
rect 20588 10084 20760 10112
rect 20588 10072 20594 10084
rect 20257 10047 20315 10053
rect 20257 10044 20269 10047
rect 19484 10016 20269 10044
rect 19484 10004 19490 10016
rect 20257 10013 20269 10016
rect 20303 10013 20315 10047
rect 20257 10007 20315 10013
rect 20346 10004 20352 10056
rect 20404 10004 20410 10056
rect 20438 10004 20444 10056
rect 20496 10040 20502 10056
rect 20625 10047 20683 10053
rect 20625 10044 20637 10047
rect 20548 10040 20637 10044
rect 20496 10016 20637 10040
rect 20496 10012 20576 10016
rect 20625 10013 20637 10016
rect 20671 10013 20683 10047
rect 20732 10044 20760 10084
rect 21082 10072 21088 10124
rect 21140 10112 21146 10124
rect 21177 10115 21235 10121
rect 21177 10112 21189 10115
rect 21140 10084 21189 10112
rect 21140 10072 21146 10084
rect 21177 10081 21189 10084
rect 21223 10081 21235 10115
rect 21177 10075 21235 10081
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 20732 10016 20913 10044
rect 20496 10004 20502 10012
rect 20625 10007 20683 10013
rect 20901 10013 20913 10016
rect 20947 10013 20959 10047
rect 20901 10007 20959 10013
rect 20990 10004 20996 10056
rect 21048 10004 21054 10056
rect 21284 10053 21312 10152
rect 21836 10152 22416 10180
rect 21269 10047 21327 10053
rect 21269 10013 21281 10047
rect 21315 10013 21327 10047
rect 21269 10007 21327 10013
rect 21634 10004 21640 10056
rect 21692 10004 21698 10056
rect 21836 10040 21864 10152
rect 22388 10124 22416 10152
rect 22649 10149 22661 10183
rect 22695 10180 22707 10183
rect 26234 10180 26240 10192
rect 22695 10152 26240 10180
rect 22695 10149 22707 10152
rect 22649 10143 22707 10149
rect 26234 10140 26240 10152
rect 26292 10140 26298 10192
rect 27525 10183 27583 10189
rect 27525 10149 27537 10183
rect 27571 10149 27583 10183
rect 29914 10180 29920 10192
rect 27525 10143 27583 10149
rect 29564 10152 29920 10180
rect 22005 10115 22063 10121
rect 22005 10081 22017 10115
rect 22051 10112 22063 10115
rect 22278 10112 22284 10124
rect 22051 10084 22284 10112
rect 22051 10081 22063 10084
rect 22005 10075 22063 10081
rect 22278 10072 22284 10084
rect 22336 10072 22342 10124
rect 22370 10072 22376 10124
rect 22428 10072 22434 10124
rect 23106 10072 23112 10124
rect 23164 10072 23170 10124
rect 21897 10041 21955 10047
rect 21897 10040 21909 10041
rect 21836 10012 21909 10040
rect 21897 10007 21909 10012
rect 21943 10007 21955 10041
rect 21897 10001 21955 10007
rect 22186 10004 22192 10056
rect 22244 10004 22250 10056
rect 22388 10044 22416 10072
rect 22465 10047 22523 10053
rect 22465 10044 22477 10047
rect 22388 10016 22477 10044
rect 22465 10013 22477 10016
rect 22511 10013 22523 10047
rect 22465 10007 22523 10013
rect 22833 10047 22891 10053
rect 22833 10013 22845 10047
rect 22879 10013 22891 10047
rect 22833 10007 22891 10013
rect 22925 10047 22983 10053
rect 22925 10013 22937 10047
rect 22971 10013 22983 10047
rect 22925 10007 22983 10013
rect 13081 9979 13139 9985
rect 13081 9945 13093 9979
rect 13127 9976 13139 9979
rect 20070 9976 20076 9988
rect 13127 9948 20076 9976
rect 13127 9945 13139 9948
rect 13081 9939 13139 9945
rect 20070 9936 20076 9948
rect 20128 9936 20134 9988
rect 22848 9976 22876 10007
rect 22296 9948 22876 9976
rect 9640 9880 10824 9908
rect 9640 9868 9646 9880
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 11149 9911 11207 9917
rect 11149 9908 11161 9911
rect 11112 9880 11161 9908
rect 11112 9868 11118 9880
rect 11149 9877 11161 9880
rect 11195 9908 11207 9911
rect 12158 9908 12164 9920
rect 11195 9880 12164 9908
rect 11195 9877 11207 9880
rect 11149 9871 11207 9877
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 16298 9868 16304 9920
rect 16356 9908 16362 9920
rect 20162 9908 20168 9920
rect 16356 9880 20168 9908
rect 16356 9868 16362 9880
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 21450 9868 21456 9920
rect 21508 9868 21514 9920
rect 21542 9868 21548 9920
rect 21600 9908 21606 9920
rect 21821 9911 21879 9917
rect 21821 9908 21833 9911
rect 21600 9880 21833 9908
rect 21600 9868 21606 9880
rect 21821 9877 21833 9880
rect 21867 9877 21879 9911
rect 21821 9871 21879 9877
rect 22002 9868 22008 9920
rect 22060 9908 22066 9920
rect 22296 9908 22324 9948
rect 22060 9880 22324 9908
rect 22060 9868 22066 9880
rect 22370 9868 22376 9920
rect 22428 9868 22434 9920
rect 22940 9908 22968 10007
rect 23198 10004 23204 10056
rect 23256 10004 23262 10056
rect 27540 10044 27568 10143
rect 27798 10072 27804 10124
rect 27856 10072 27862 10124
rect 28994 10072 29000 10124
rect 29052 10112 29058 10124
rect 29564 10121 29592 10152
rect 29914 10140 29920 10152
rect 29972 10140 29978 10192
rect 30098 10140 30104 10192
rect 30156 10180 30162 10192
rect 30193 10183 30251 10189
rect 30193 10180 30205 10183
rect 30156 10152 30205 10180
rect 30156 10140 30162 10152
rect 30193 10149 30205 10152
rect 30239 10149 30251 10183
rect 30193 10143 30251 10149
rect 31478 10140 31484 10192
rect 31536 10140 31542 10192
rect 29549 10115 29607 10121
rect 29549 10112 29561 10115
rect 29052 10084 29561 10112
rect 29052 10072 29058 10084
rect 29549 10081 29561 10084
rect 29595 10081 29607 10115
rect 29549 10075 29607 10081
rect 29638 10072 29644 10124
rect 29696 10112 29702 10124
rect 30469 10115 30527 10121
rect 30469 10112 30481 10115
rect 29696 10084 30481 10112
rect 29696 10072 29702 10084
rect 30469 10081 30481 10084
rect 30515 10081 30527 10115
rect 30469 10075 30527 10081
rect 30742 10072 30748 10124
rect 30800 10112 30806 10124
rect 31110 10112 31116 10124
rect 30800 10084 31116 10112
rect 30800 10072 30806 10084
rect 31110 10072 31116 10084
rect 31168 10072 31174 10124
rect 32030 10072 32036 10124
rect 32088 10072 32094 10124
rect 27540 10016 27660 10044
rect 27632 9976 27660 10016
rect 27706 10004 27712 10056
rect 27764 10004 27770 10056
rect 29178 10004 29184 10056
rect 29236 10044 29242 10056
rect 29362 10044 29368 10056
rect 29236 10016 29368 10044
rect 29236 10004 29242 10016
rect 29362 10004 29368 10016
rect 29420 10044 29426 10056
rect 29733 10047 29791 10053
rect 29733 10044 29745 10047
rect 29420 10016 29745 10044
rect 29420 10004 29426 10016
rect 29733 10013 29745 10016
rect 29779 10013 29791 10047
rect 29733 10007 29791 10013
rect 30558 10004 30564 10056
rect 30616 10053 30622 10056
rect 30616 10047 30644 10053
rect 30632 10013 30644 10047
rect 30616 10007 30644 10013
rect 30616 10004 30622 10007
rect 28046 9979 28104 9985
rect 28046 9976 28058 9979
rect 27632 9948 28058 9976
rect 28046 9945 28058 9948
rect 28092 9945 28104 9979
rect 28046 9939 28104 9945
rect 29454 9936 29460 9988
rect 29512 9976 29518 9988
rect 31389 9979 31447 9985
rect 29512 9948 29776 9976
rect 29512 9936 29518 9948
rect 29086 9908 29092 9920
rect 22940 9880 29092 9908
rect 29086 9868 29092 9880
rect 29144 9868 29150 9920
rect 29178 9868 29184 9920
rect 29236 9908 29242 9920
rect 29546 9908 29552 9920
rect 29236 9880 29552 9908
rect 29236 9868 29242 9880
rect 29546 9868 29552 9880
rect 29604 9868 29610 9920
rect 29748 9908 29776 9948
rect 31389 9945 31401 9979
rect 31435 9976 31447 9979
rect 31849 9979 31907 9985
rect 31849 9976 31861 9979
rect 31435 9948 31861 9976
rect 31435 9945 31447 9948
rect 31389 9939 31447 9945
rect 31849 9945 31861 9948
rect 31895 9945 31907 9979
rect 34164 9976 34192 10220
rect 35176 10220 37372 10248
rect 35176 10121 35204 10220
rect 36280 10121 36308 10220
rect 37366 10208 37372 10220
rect 37424 10208 37430 10260
rect 40402 10208 40408 10260
rect 40460 10248 40466 10260
rect 40773 10251 40831 10257
rect 40773 10248 40785 10251
rect 40460 10220 40785 10248
rect 40460 10208 40466 10220
rect 40773 10217 40785 10220
rect 40819 10217 40831 10251
rect 40773 10211 40831 10217
rect 37277 10183 37335 10189
rect 37277 10149 37289 10183
rect 37323 10180 37335 10183
rect 37826 10180 37832 10192
rect 37323 10152 37832 10180
rect 37323 10149 37335 10152
rect 37277 10143 37335 10149
rect 37826 10140 37832 10152
rect 37884 10140 37890 10192
rect 42705 10183 42763 10189
rect 42705 10149 42717 10183
rect 42751 10180 42763 10183
rect 43070 10180 43076 10192
rect 42751 10152 43076 10180
rect 42751 10149 42763 10152
rect 42705 10143 42763 10149
rect 43070 10140 43076 10152
rect 43128 10140 43134 10192
rect 35161 10115 35219 10121
rect 35161 10081 35173 10115
rect 35207 10081 35219 10115
rect 35161 10075 35219 10081
rect 36265 10115 36323 10121
rect 36265 10081 36277 10115
rect 36311 10081 36323 10115
rect 36265 10075 36323 10081
rect 39206 10072 39212 10124
rect 39264 10112 39270 10124
rect 39669 10115 39727 10121
rect 39264 10084 39620 10112
rect 39264 10072 39270 10084
rect 35434 10004 35440 10056
rect 35492 10004 35498 10056
rect 36541 10047 36599 10053
rect 36541 10013 36553 10047
rect 36587 10013 36599 10047
rect 36541 10007 36599 10013
rect 36556 9976 36584 10007
rect 39390 10004 39396 10056
rect 39448 10004 39454 10056
rect 39482 10004 39488 10056
rect 39540 10004 39546 10056
rect 39592 10044 39620 10084
rect 39669 10081 39681 10115
rect 39715 10112 39727 10115
rect 40586 10112 40592 10124
rect 39715 10084 40592 10112
rect 39715 10081 39727 10084
rect 39669 10075 39727 10081
rect 40586 10072 40592 10084
rect 40644 10072 40650 10124
rect 40862 10072 40868 10124
rect 40920 10112 40926 10124
rect 42889 10115 42947 10121
rect 40920 10084 41184 10112
rect 40920 10072 40926 10084
rect 39853 10047 39911 10053
rect 39853 10044 39865 10047
rect 39592 10016 39865 10044
rect 39853 10013 39865 10016
rect 39899 10013 39911 10047
rect 39853 10007 39911 10013
rect 40129 10047 40187 10053
rect 40129 10013 40141 10047
rect 40175 10013 40187 10047
rect 40129 10007 40187 10013
rect 38286 9976 38292 9988
rect 34164 9948 36584 9976
rect 37292 9948 38292 9976
rect 31849 9939 31907 9945
rect 30558 9908 30564 9920
rect 29748 9880 30564 9908
rect 30558 9868 30564 9880
rect 30616 9868 30622 9920
rect 31941 9911 31999 9917
rect 31941 9877 31953 9911
rect 31987 9908 31999 9911
rect 33318 9908 33324 9920
rect 31987 9880 33324 9908
rect 31987 9877 31999 9880
rect 31941 9871 31999 9877
rect 33318 9868 33324 9880
rect 33376 9868 33382 9920
rect 36173 9911 36231 9917
rect 36173 9877 36185 9911
rect 36219 9908 36231 9911
rect 37292 9908 37320 9948
rect 38286 9936 38292 9948
rect 38344 9936 38350 9988
rect 40144 9976 40172 10007
rect 41046 10004 41052 10056
rect 41104 10004 41110 10056
rect 41156 10053 41184 10084
rect 41248 10084 42748 10112
rect 41248 10053 41276 10084
rect 41141 10047 41199 10053
rect 41141 10013 41153 10047
rect 41187 10013 41199 10047
rect 41141 10007 41199 10013
rect 41233 10047 41291 10053
rect 41233 10013 41245 10047
rect 41279 10013 41291 10047
rect 41233 10007 41291 10013
rect 41417 10047 41475 10053
rect 41417 10013 41429 10047
rect 41463 10044 41475 10047
rect 42426 10044 42432 10056
rect 41463 10016 42432 10044
rect 41463 10013 41475 10016
rect 41417 10007 41475 10013
rect 41432 9976 41460 10007
rect 42426 10004 42432 10016
rect 42484 10004 42490 10056
rect 42613 10047 42671 10053
rect 42613 10013 42625 10047
rect 42659 10013 42671 10047
rect 42720 10044 42748 10084
rect 42889 10081 42901 10115
rect 42935 10112 42947 10115
rect 43714 10112 43720 10124
rect 42935 10084 43720 10112
rect 42935 10081 42947 10084
rect 42889 10075 42947 10081
rect 43714 10072 43720 10084
rect 43772 10072 43778 10124
rect 42978 10044 42984 10056
rect 42720 10016 42984 10044
rect 42613 10007 42671 10013
rect 40144 9948 41460 9976
rect 42628 9976 42656 10007
rect 42978 10004 42984 10016
rect 43036 10004 43042 10056
rect 43165 10047 43223 10053
rect 43165 10013 43177 10047
rect 43211 10044 43223 10047
rect 44174 10044 44180 10056
rect 43211 10016 44180 10044
rect 43211 10013 43223 10016
rect 43165 10007 43223 10013
rect 44174 10004 44180 10016
rect 44232 10004 44238 10056
rect 42794 9976 42800 9988
rect 42628 9948 42800 9976
rect 42794 9936 42800 9948
rect 42852 9936 42858 9988
rect 36219 9880 37320 9908
rect 36219 9877 36231 9880
rect 36173 9871 36231 9877
rect 37366 9868 37372 9920
rect 37424 9908 37430 9920
rect 39669 9911 39727 9917
rect 39669 9908 39681 9911
rect 37424 9880 39681 9908
rect 37424 9868 37430 9880
rect 39669 9877 39681 9880
rect 39715 9877 39727 9911
rect 39669 9871 39727 9877
rect 39758 9868 39764 9920
rect 39816 9908 39822 9920
rect 42889 9911 42947 9917
rect 42889 9908 42901 9911
rect 39816 9880 42901 9908
rect 39816 9868 39822 9880
rect 42889 9877 42901 9880
rect 42935 9877 42947 9911
rect 42889 9871 42947 9877
rect 43162 9868 43168 9920
rect 43220 9868 43226 9920
rect 1104 9818 47104 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 47104 9818
rect 1104 9744 47104 9766
rect 7742 9664 7748 9716
rect 7800 9664 7806 9716
rect 12434 9704 12440 9716
rect 10980 9676 12440 9704
rect 6362 9596 6368 9648
rect 6420 9636 6426 9648
rect 6610 9639 6668 9645
rect 6610 9636 6622 9639
rect 6420 9608 6622 9636
rect 6420 9596 6426 9608
rect 6610 9605 6622 9608
rect 6656 9605 6668 9639
rect 6610 9599 6668 9605
rect 10042 9596 10048 9648
rect 10100 9596 10106 9648
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 7892 9540 8125 9568
rect 7892 9528 7898 9540
rect 8113 9537 8125 9540
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 8846 9528 8852 9580
rect 8904 9528 8910 9580
rect 6178 9460 6184 9512
rect 6236 9500 6242 9512
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 6236 9472 6377 9500
rect 6236 9460 6242 9472
rect 6365 9469 6377 9472
rect 6411 9469 6423 9503
rect 6365 9463 6423 9469
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 7929 9503 7987 9509
rect 7929 9500 7941 9503
rect 7708 9472 7941 9500
rect 7708 9460 7714 9472
rect 7929 9469 7941 9472
rect 7975 9469 7987 9503
rect 7929 9463 7987 9469
rect 8662 9460 8668 9512
rect 8720 9500 8726 9512
rect 8966 9503 9024 9509
rect 8966 9500 8978 9503
rect 8720 9472 8978 9500
rect 8720 9460 8726 9472
rect 8966 9469 8978 9472
rect 9012 9469 9024 9503
rect 8966 9463 9024 9469
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9500 9183 9503
rect 10594 9500 10600 9512
rect 9171 9472 10600 9500
rect 9171 9469 9183 9472
rect 9125 9463 9183 9469
rect 10594 9460 10600 9472
rect 10652 9500 10658 9512
rect 10980 9500 11008 9676
rect 12434 9664 12440 9676
rect 12492 9664 12498 9716
rect 17034 9664 17040 9716
rect 17092 9704 17098 9716
rect 20254 9704 20260 9716
rect 17092 9676 20260 9704
rect 17092 9664 17098 9676
rect 20254 9664 20260 9676
rect 20312 9664 20318 9716
rect 20346 9664 20352 9716
rect 20404 9704 20410 9716
rect 25130 9704 25136 9716
rect 20404 9676 25136 9704
rect 20404 9664 20410 9676
rect 25130 9664 25136 9676
rect 25188 9664 25194 9716
rect 27706 9664 27712 9716
rect 27764 9704 27770 9716
rect 28445 9707 28503 9713
rect 28445 9704 28457 9707
rect 27764 9676 28457 9704
rect 27764 9664 27770 9676
rect 28445 9673 28457 9676
rect 28491 9673 28503 9707
rect 28905 9707 28963 9713
rect 28905 9704 28917 9707
rect 28445 9667 28503 9673
rect 28736 9676 28917 9704
rect 19702 9596 19708 9648
rect 19760 9596 19766 9648
rect 19794 9596 19800 9648
rect 19852 9636 19858 9648
rect 20809 9639 20867 9645
rect 20809 9636 20821 9639
rect 19852 9608 20821 9636
rect 19852 9596 19858 9608
rect 20809 9605 20821 9608
rect 20855 9605 20867 9639
rect 20809 9599 20867 9605
rect 25869 9639 25927 9645
rect 25869 9605 25881 9639
rect 25915 9636 25927 9639
rect 26326 9636 26332 9648
rect 25915 9608 26332 9636
rect 25915 9605 25927 9608
rect 25869 9599 25927 9605
rect 26326 9596 26332 9608
rect 26384 9596 26390 9648
rect 26436 9608 27384 9636
rect 17862 9528 17868 9580
rect 17920 9528 17926 9580
rect 18046 9528 18052 9580
rect 18104 9528 18110 9580
rect 18782 9528 18788 9580
rect 18840 9528 18846 9580
rect 18874 9528 18880 9580
rect 18932 9577 18938 9580
rect 18932 9571 18960 9577
rect 18948 9537 18960 9571
rect 18932 9531 18960 9537
rect 18932 9528 18938 9531
rect 19058 9528 19064 9580
rect 19116 9528 19122 9580
rect 21082 9568 21088 9580
rect 20272 9540 21088 9568
rect 10652 9472 11008 9500
rect 17880 9500 17908 9528
rect 19794 9500 19800 9512
rect 17880 9472 19800 9500
rect 10652 9460 10658 9472
rect 19794 9460 19800 9472
rect 19852 9460 19858 9512
rect 20272 9509 20300 9540
rect 21082 9528 21088 9540
rect 21140 9528 21146 9580
rect 21450 9528 21456 9580
rect 21508 9568 21514 9580
rect 22278 9568 22284 9580
rect 21508 9540 22284 9568
rect 21508 9528 21514 9540
rect 22278 9528 22284 9540
rect 22336 9528 22342 9580
rect 24029 9571 24087 9577
rect 24029 9537 24041 9571
rect 24075 9568 24087 9571
rect 24394 9568 24400 9580
rect 24075 9540 24400 9568
rect 24075 9537 24087 9540
rect 24029 9531 24087 9537
rect 24394 9528 24400 9540
rect 24452 9528 24458 9580
rect 25222 9528 25228 9580
rect 25280 9528 25286 9580
rect 20257 9503 20315 9509
rect 20257 9469 20269 9503
rect 20303 9469 20315 9503
rect 20257 9463 20315 9469
rect 21269 9503 21327 9509
rect 21269 9469 21281 9503
rect 21315 9500 21327 9503
rect 23106 9500 23112 9512
rect 21315 9472 23112 9500
rect 21315 9469 21327 9472
rect 21269 9463 21327 9469
rect 23106 9460 23112 9472
rect 23164 9460 23170 9512
rect 24213 9503 24271 9509
rect 24213 9469 24225 9503
rect 24259 9500 24271 9503
rect 24578 9500 24584 9512
rect 24259 9472 24584 9500
rect 24259 9469 24271 9472
rect 24213 9463 24271 9469
rect 24578 9460 24584 9472
rect 24636 9460 24642 9512
rect 24946 9460 24952 9512
rect 25004 9460 25010 9512
rect 25087 9503 25145 9509
rect 25087 9469 25099 9503
rect 25133 9500 25145 9503
rect 25406 9500 25412 9512
rect 25133 9472 25412 9500
rect 25133 9469 25145 9472
rect 25087 9463 25145 9469
rect 25406 9460 25412 9472
rect 25464 9460 25470 9512
rect 8573 9435 8631 9441
rect 8573 9401 8585 9435
rect 8619 9401 8631 9435
rect 8573 9395 8631 9401
rect 8588 9364 8616 9395
rect 17494 9392 17500 9444
rect 17552 9432 17558 9444
rect 18509 9435 18567 9441
rect 18509 9432 18521 9435
rect 17552 9404 18521 9432
rect 17552 9392 17558 9404
rect 18509 9401 18521 9404
rect 18555 9401 18567 9435
rect 18509 9395 18567 9401
rect 9582 9364 9588 9376
rect 8588 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 9766 9324 9772 9376
rect 9824 9324 9830 9376
rect 10134 9324 10140 9376
rect 10192 9324 10198 9376
rect 16574 9324 16580 9376
rect 16632 9364 16638 9376
rect 17034 9364 17040 9376
rect 16632 9336 17040 9364
rect 16632 9324 16638 9336
rect 17034 9324 17040 9336
rect 17092 9324 17098 9376
rect 18524 9364 18552 9395
rect 20070 9392 20076 9444
rect 20128 9392 20134 9444
rect 21082 9392 21088 9444
rect 21140 9392 21146 9444
rect 24118 9392 24124 9444
rect 24176 9432 24182 9444
rect 24673 9435 24731 9441
rect 24673 9432 24685 9435
rect 24176 9404 24685 9432
rect 24176 9392 24182 9404
rect 24673 9401 24685 9404
rect 24719 9401 24731 9435
rect 24673 9395 24731 9401
rect 19886 9364 19892 9376
rect 18524 9336 19892 9364
rect 19886 9324 19892 9336
rect 19944 9324 19950 9376
rect 22554 9324 22560 9376
rect 22612 9364 22618 9376
rect 26436 9364 26464 9608
rect 26786 9528 26792 9580
rect 26844 9528 26850 9580
rect 27229 9571 27287 9577
rect 27229 9568 27241 9571
rect 26896 9540 27241 9568
rect 26605 9435 26663 9441
rect 26605 9401 26617 9435
rect 26651 9432 26663 9435
rect 26896 9432 26924 9540
rect 27229 9537 27241 9540
rect 27275 9537 27287 9571
rect 27356 9568 27384 9608
rect 27522 9596 27528 9648
rect 27580 9636 27586 9648
rect 28736 9636 28764 9676
rect 28905 9673 28917 9676
rect 28951 9673 28963 9707
rect 28905 9667 28963 9673
rect 29086 9664 29092 9716
rect 29144 9704 29150 9716
rect 30745 9707 30803 9713
rect 30745 9704 30757 9707
rect 29144 9676 30757 9704
rect 29144 9664 29150 9676
rect 30745 9673 30757 9676
rect 30791 9673 30803 9707
rect 30745 9667 30803 9673
rect 35250 9664 35256 9716
rect 35308 9704 35314 9716
rect 36170 9704 36176 9716
rect 35308 9676 36176 9704
rect 35308 9664 35314 9676
rect 36170 9664 36176 9676
rect 36228 9664 36234 9716
rect 39850 9664 39856 9716
rect 39908 9704 39914 9716
rect 46474 9704 46480 9716
rect 39908 9676 46480 9704
rect 39908 9664 39914 9676
rect 46474 9664 46480 9676
rect 46532 9664 46538 9716
rect 27580 9608 28764 9636
rect 28813 9639 28871 9645
rect 27580 9596 27586 9608
rect 28813 9605 28825 9639
rect 28859 9636 28871 9639
rect 29178 9636 29184 9648
rect 28859 9608 29184 9636
rect 28859 9605 28871 9608
rect 28813 9599 28871 9605
rect 29178 9596 29184 9608
rect 29236 9596 29242 9648
rect 29546 9596 29552 9648
rect 29604 9636 29610 9648
rect 29604 9608 31754 9636
rect 29604 9596 29610 9608
rect 31113 9571 31171 9577
rect 27356 9540 29592 9568
rect 27229 9531 27287 9537
rect 26973 9503 27031 9509
rect 26973 9469 26985 9503
rect 27019 9469 27031 9503
rect 26973 9463 27031 9469
rect 28997 9503 29055 9509
rect 28997 9469 29009 9503
rect 29043 9469 29055 9503
rect 28997 9463 29055 9469
rect 26651 9404 26924 9432
rect 26651 9401 26663 9404
rect 26605 9395 26663 9401
rect 22612 9336 26464 9364
rect 26988 9364 27016 9463
rect 28258 9392 28264 9444
rect 28316 9432 28322 9444
rect 29012 9432 29040 9463
rect 29270 9432 29276 9444
rect 28316 9404 29276 9432
rect 28316 9392 28322 9404
rect 29270 9392 29276 9404
rect 29328 9392 29334 9444
rect 27706 9364 27712 9376
rect 26988 9336 27712 9364
rect 22612 9324 22618 9336
rect 27706 9324 27712 9336
rect 27764 9324 27770 9376
rect 28350 9324 28356 9376
rect 28408 9364 28414 9376
rect 29454 9364 29460 9376
rect 28408 9336 29460 9364
rect 28408 9324 28414 9336
rect 29454 9324 29460 9336
rect 29512 9324 29518 9376
rect 29564 9364 29592 9540
rect 31113 9537 31125 9571
rect 31159 9568 31171 9571
rect 31294 9568 31300 9580
rect 31159 9540 31300 9568
rect 31159 9537 31171 9540
rect 31113 9531 31171 9537
rect 31294 9528 31300 9540
rect 31352 9528 31358 9580
rect 31726 9568 31754 9608
rect 31938 9596 31944 9648
rect 31996 9636 32002 9648
rect 35986 9636 35992 9648
rect 31996 9608 35992 9636
rect 31996 9596 32002 9608
rect 35986 9596 35992 9608
rect 36044 9636 36050 9648
rect 36446 9636 36452 9648
rect 36044 9608 36452 9636
rect 36044 9596 36050 9608
rect 36446 9596 36452 9608
rect 36504 9596 36510 9648
rect 40494 9596 40500 9648
rect 40552 9596 40558 9648
rect 41046 9596 41052 9648
rect 41104 9636 41110 9648
rect 42245 9639 42303 9645
rect 41104 9608 41276 9636
rect 41104 9596 41110 9608
rect 36173 9571 36231 9577
rect 36173 9568 36185 9571
rect 31726 9540 36185 9568
rect 36173 9537 36185 9540
rect 36219 9537 36231 9571
rect 36173 9531 36231 9537
rect 38378 9528 38384 9580
rect 38436 9528 38442 9580
rect 38565 9571 38623 9577
rect 38565 9537 38577 9571
rect 38611 9568 38623 9571
rect 38654 9568 38660 9580
rect 38611 9540 38660 9568
rect 38611 9537 38623 9540
rect 38565 9531 38623 9537
rect 38654 9528 38660 9540
rect 38712 9528 38718 9580
rect 40034 9528 40040 9580
rect 40092 9568 40098 9580
rect 40092 9540 40264 9568
rect 40092 9528 40098 9540
rect 31205 9503 31263 9509
rect 31205 9469 31217 9503
rect 31251 9469 31263 9503
rect 31205 9463 31263 9469
rect 31389 9503 31447 9509
rect 31389 9469 31401 9503
rect 31435 9500 31447 9503
rect 32030 9500 32036 9512
rect 31435 9472 32036 9500
rect 31435 9469 31447 9472
rect 31389 9463 31447 9469
rect 31220 9432 31248 9463
rect 32030 9460 32036 9472
rect 32088 9460 32094 9512
rect 32122 9460 32128 9512
rect 32180 9500 32186 9512
rect 32217 9503 32275 9509
rect 32217 9500 32229 9503
rect 32180 9472 32229 9500
rect 32180 9460 32186 9472
rect 32217 9469 32229 9472
rect 32263 9469 32275 9503
rect 32217 9463 32275 9469
rect 32306 9460 32312 9512
rect 32364 9500 32370 9512
rect 32493 9503 32551 9509
rect 32493 9500 32505 9503
rect 32364 9472 32505 9500
rect 32364 9460 32370 9472
rect 32493 9469 32505 9472
rect 32539 9469 32551 9503
rect 32493 9463 32551 9469
rect 35342 9460 35348 9512
rect 35400 9500 35406 9512
rect 35802 9500 35808 9512
rect 35400 9472 35808 9500
rect 35400 9460 35406 9472
rect 35802 9460 35808 9472
rect 35860 9500 35866 9512
rect 35897 9503 35955 9509
rect 35897 9500 35909 9503
rect 35860 9472 35909 9500
rect 35860 9460 35866 9472
rect 35897 9469 35909 9472
rect 35943 9469 35955 9503
rect 35897 9463 35955 9469
rect 39482 9460 39488 9512
rect 39540 9500 39546 9512
rect 40129 9503 40187 9509
rect 40129 9500 40141 9503
rect 39540 9472 40141 9500
rect 39540 9460 39546 9472
rect 40129 9469 40141 9472
rect 40175 9469 40187 9503
rect 40236 9500 40264 9540
rect 40310 9528 40316 9580
rect 40368 9528 40374 9580
rect 40405 9571 40463 9577
rect 40405 9537 40417 9571
rect 40451 9568 40463 9571
rect 40512 9568 40540 9596
rect 40451 9540 40540 9568
rect 40589 9571 40647 9577
rect 40451 9537 40463 9540
rect 40405 9531 40463 9537
rect 40589 9537 40601 9571
rect 40635 9568 40647 9571
rect 40678 9568 40684 9580
rect 40635 9540 40684 9568
rect 40635 9537 40647 9540
rect 40589 9531 40647 9537
rect 40678 9528 40684 9540
rect 40736 9568 40742 9580
rect 41138 9568 41144 9580
rect 40736 9540 41144 9568
rect 40736 9528 40742 9540
rect 41138 9528 41144 9540
rect 41196 9528 41202 9580
rect 41248 9577 41276 9608
rect 42245 9605 42257 9639
rect 42291 9636 42303 9639
rect 43346 9636 43352 9648
rect 42291 9608 43352 9636
rect 42291 9605 42303 9608
rect 42245 9599 42303 9605
rect 43346 9596 43352 9608
rect 43404 9596 43410 9648
rect 41233 9571 41291 9577
rect 41233 9537 41245 9571
rect 41279 9537 41291 9571
rect 42613 9571 42671 9577
rect 41233 9531 41291 9537
rect 40497 9503 40555 9509
rect 40497 9500 40509 9503
rect 40236 9472 40509 9500
rect 40129 9463 40187 9469
rect 40497 9469 40509 9472
rect 40543 9469 40555 9503
rect 40497 9463 40555 9469
rect 40770 9460 40776 9512
rect 40828 9500 40834 9512
rect 41340 9500 41368 9554
rect 42613 9537 42625 9571
rect 42659 9537 42671 9571
rect 42613 9531 42671 9537
rect 42521 9503 42579 9509
rect 42521 9500 42533 9503
rect 40828 9472 42533 9500
rect 40828 9460 40834 9472
rect 42521 9469 42533 9472
rect 42567 9469 42579 9503
rect 42521 9463 42579 9469
rect 34790 9432 34796 9444
rect 31220 9404 34796 9432
rect 34790 9392 34796 9404
rect 34848 9392 34854 9444
rect 37734 9432 37740 9444
rect 36556 9404 37740 9432
rect 36556 9364 36584 9404
rect 37734 9392 37740 9404
rect 37792 9392 37798 9444
rect 41046 9392 41052 9444
rect 41104 9432 41110 9444
rect 42628 9432 42656 9531
rect 42886 9528 42892 9580
rect 42944 9568 42950 9580
rect 43162 9568 43168 9580
rect 42944 9540 43168 9568
rect 42944 9528 42950 9540
rect 43162 9528 43168 9540
rect 43220 9568 43226 9580
rect 43441 9571 43499 9577
rect 43441 9568 43453 9571
rect 43220 9540 43453 9568
rect 43220 9528 43226 9540
rect 43441 9537 43453 9540
rect 43487 9537 43499 9571
rect 43441 9531 43499 9537
rect 43070 9460 43076 9512
rect 43128 9460 43134 9512
rect 43254 9460 43260 9512
rect 43312 9460 43318 9512
rect 43349 9503 43407 9509
rect 43349 9469 43361 9503
rect 43395 9469 43407 9503
rect 43349 9463 43407 9469
rect 43533 9503 43591 9509
rect 43533 9469 43545 9503
rect 43579 9469 43591 9503
rect 43533 9463 43591 9469
rect 41104 9404 42656 9432
rect 41104 9392 41110 9404
rect 42702 9392 42708 9444
rect 42760 9432 42766 9444
rect 42981 9435 43039 9441
rect 42981 9432 42993 9435
rect 42760 9404 42993 9432
rect 42760 9392 42766 9404
rect 42981 9401 42993 9404
rect 43027 9432 43039 9435
rect 43364 9432 43392 9463
rect 43027 9404 43392 9432
rect 43027 9401 43039 9404
rect 42981 9395 43039 9401
rect 29564 9336 36584 9364
rect 36909 9367 36967 9373
rect 36909 9333 36921 9367
rect 36955 9364 36967 9367
rect 38102 9364 38108 9376
rect 36955 9336 38108 9364
rect 36955 9333 36967 9336
rect 36909 9327 36967 9333
rect 38102 9324 38108 9336
rect 38160 9324 38166 9376
rect 38378 9324 38384 9376
rect 38436 9324 38442 9376
rect 41414 9324 41420 9376
rect 41472 9364 41478 9376
rect 43548 9364 43576 9463
rect 41472 9336 43576 9364
rect 41472 9324 41478 9336
rect 1104 9274 47104 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 47104 9274
rect 1104 9200 47104 9222
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 6236 9132 6914 9160
rect 6236 9120 6242 9132
rect 6886 9024 6914 9132
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 22370 9160 22376 9172
rect 9824 9132 22376 9160
rect 9824 9120 9830 9132
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 26329 9163 26387 9169
rect 26329 9160 26341 9163
rect 24228 9132 26341 9160
rect 9674 9052 9680 9104
rect 9732 9092 9738 9104
rect 10597 9095 10655 9101
rect 10597 9092 10609 9095
rect 9732 9064 10609 9092
rect 9732 9052 9738 9064
rect 10597 9061 10609 9064
rect 10643 9061 10655 9095
rect 10597 9055 10655 9061
rect 13173 9095 13231 9101
rect 13173 9061 13185 9095
rect 13219 9092 13231 9095
rect 14550 9092 14556 9104
rect 13219 9064 14556 9092
rect 13219 9061 13231 9064
rect 13173 9055 13231 9061
rect 14550 9052 14556 9064
rect 14608 9052 14614 9104
rect 20898 9052 20904 9104
rect 20956 9092 20962 9104
rect 21453 9095 21511 9101
rect 21453 9092 21465 9095
rect 20956 9064 21465 9092
rect 20956 9052 20962 9064
rect 21453 9061 21465 9064
rect 21499 9061 21511 9095
rect 21453 9055 21511 9061
rect 21637 9095 21695 9101
rect 21637 9061 21649 9095
rect 21683 9092 21695 9095
rect 22833 9095 22891 9101
rect 22833 9092 22845 9095
rect 21683 9064 22845 9092
rect 21683 9061 21695 9064
rect 21637 9055 21695 9061
rect 22833 9061 22845 9064
rect 22879 9061 22891 9095
rect 22833 9055 22891 9061
rect 10134 9024 10140 9036
rect 6886 8996 10140 9024
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 10468 8996 11161 9024
rect 10468 8984 10474 8996
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 13725 9027 13783 9033
rect 13725 8993 13737 9027
rect 13771 9024 13783 9027
rect 14182 9024 14188 9036
rect 13771 8996 14188 9024
rect 13771 8993 13783 8996
rect 13725 8987 13783 8993
rect 14182 8984 14188 8996
rect 14240 9024 14246 9036
rect 15010 9024 15016 9036
rect 14240 8996 15016 9024
rect 14240 8984 14246 8996
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 15841 9027 15899 9033
rect 15841 8993 15853 9027
rect 15887 9024 15899 9027
rect 16482 9024 16488 9036
rect 15887 8996 16488 9024
rect 15887 8993 15899 8996
rect 15841 8987 15899 8993
rect 16482 8984 16488 8996
rect 16540 9024 16546 9036
rect 16577 9027 16635 9033
rect 16577 9024 16589 9027
rect 16540 8996 16589 9024
rect 16540 8984 16546 8996
rect 16577 8993 16589 8996
rect 16623 8993 16635 9027
rect 16577 8987 16635 8993
rect 21177 9027 21235 9033
rect 21177 8993 21189 9027
rect 21223 9024 21235 9027
rect 21818 9024 21824 9036
rect 21223 8996 21824 9024
rect 21223 8993 21235 8996
rect 21177 8987 21235 8993
rect 21818 8984 21824 8996
rect 21876 8984 21882 9036
rect 22186 8984 22192 9036
rect 22244 8984 22250 9036
rect 22462 8984 22468 9036
rect 22520 9024 22526 9036
rect 22520 8996 22968 9024
rect 22520 8984 22526 8996
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8956 11023 8959
rect 11054 8956 11060 8968
rect 11011 8928 11060 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 19610 8916 19616 8968
rect 19668 8956 19674 8968
rect 20346 8956 20352 8968
rect 19668 8928 20352 8956
rect 19668 8916 19674 8928
rect 20346 8916 20352 8928
rect 20404 8916 20410 8968
rect 21913 8959 21971 8965
rect 21913 8925 21925 8959
rect 21959 8925 21971 8959
rect 21913 8919 21971 8925
rect 12618 8848 12624 8900
rect 12676 8888 12682 8900
rect 13633 8891 13691 8897
rect 13633 8888 13645 8891
rect 12676 8860 13645 8888
rect 12676 8848 12682 8860
rect 13633 8857 13645 8860
rect 13679 8857 13691 8891
rect 13633 8851 13691 8857
rect 13998 8848 14004 8900
rect 14056 8888 14062 8900
rect 16393 8891 16451 8897
rect 14056 8860 16252 8888
rect 14056 8848 14062 8860
rect 10962 8780 10968 8832
rect 11020 8820 11026 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 11020 8792 11069 8820
rect 11020 8780 11026 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11057 8783 11115 8789
rect 13541 8823 13599 8829
rect 13541 8789 13553 8823
rect 13587 8820 13599 8823
rect 13814 8820 13820 8832
rect 13587 8792 13820 8820
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 14826 8780 14832 8832
rect 14884 8820 14890 8832
rect 15197 8823 15255 8829
rect 15197 8820 15209 8823
rect 14884 8792 15209 8820
rect 14884 8780 14890 8792
rect 15197 8789 15209 8792
rect 15243 8789 15255 8823
rect 15197 8783 15255 8789
rect 15562 8780 15568 8832
rect 15620 8780 15626 8832
rect 15654 8780 15660 8832
rect 15712 8780 15718 8832
rect 16025 8823 16083 8829
rect 16025 8789 16037 8823
rect 16071 8820 16083 8823
rect 16114 8820 16120 8832
rect 16071 8792 16120 8820
rect 16071 8789 16083 8792
rect 16025 8783 16083 8789
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 16224 8820 16252 8860
rect 16393 8857 16405 8891
rect 16439 8888 16451 8891
rect 17126 8888 17132 8900
rect 16439 8860 17132 8888
rect 16439 8857 16451 8860
rect 16393 8851 16451 8857
rect 17126 8848 17132 8860
rect 17184 8848 17190 8900
rect 19334 8848 19340 8900
rect 19392 8888 19398 8900
rect 20622 8888 20628 8900
rect 19392 8860 20628 8888
rect 19392 8848 19398 8860
rect 20622 8848 20628 8860
rect 20680 8848 20686 8900
rect 21928 8888 21956 8919
rect 22002 8916 22008 8968
rect 22060 8916 22066 8968
rect 22278 8916 22284 8968
rect 22336 8916 22342 8968
rect 22940 8965 22968 8996
rect 24228 8965 24256 9132
rect 26329 9129 26341 9132
rect 26375 9129 26387 9163
rect 26329 9123 26387 9129
rect 26786 9120 26792 9172
rect 26844 9160 26850 9172
rect 27249 9163 27307 9169
rect 27249 9160 27261 9163
rect 26844 9132 27261 9160
rect 26844 9120 26850 9132
rect 27249 9129 27261 9132
rect 27295 9129 27307 9163
rect 27249 9123 27307 9129
rect 27522 9120 27528 9172
rect 27580 9160 27586 9172
rect 31938 9160 31944 9172
rect 27580 9132 31944 9160
rect 27580 9120 27586 9132
rect 31938 9120 31944 9132
rect 31996 9120 32002 9172
rect 36725 9163 36783 9169
rect 36725 9160 36737 9163
rect 32048 9132 36737 9160
rect 24854 9092 24860 9104
rect 24596 9064 24860 9092
rect 24596 9036 24624 9064
rect 24854 9052 24860 9064
rect 24912 9052 24918 9104
rect 24946 9052 24952 9104
rect 25004 9092 25010 9104
rect 28258 9092 28264 9104
rect 25004 9064 25176 9092
rect 25004 9052 25010 9064
rect 24394 8984 24400 9036
rect 24452 8984 24458 9036
rect 24578 8984 24584 9036
rect 24636 8984 24642 9036
rect 25038 8984 25044 9036
rect 25096 8984 25102 9036
rect 25148 9024 25176 9064
rect 26988 9064 28264 9092
rect 25317 9027 25375 9033
rect 25317 9024 25329 9027
rect 25148 8996 25329 9024
rect 25317 8993 25329 8996
rect 25363 9024 25375 9027
rect 25958 9024 25964 9036
rect 25363 8996 25964 9024
rect 25363 8993 25375 8996
rect 25317 8987 25375 8993
rect 25958 8984 25964 8996
rect 26016 9024 26022 9036
rect 26988 9033 27016 9064
rect 28258 9052 28264 9064
rect 28316 9052 28322 9104
rect 30377 9095 30435 9101
rect 30377 9061 30389 9095
rect 30423 9061 30435 9095
rect 30377 9055 30435 9061
rect 26973 9027 27031 9033
rect 26016 8996 26740 9024
rect 26016 8984 26022 8996
rect 22557 8959 22615 8965
rect 22557 8925 22569 8959
rect 22603 8925 22615 8959
rect 22557 8919 22615 8925
rect 22649 8959 22707 8965
rect 22649 8925 22661 8959
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8925 22983 8959
rect 22925 8919 22983 8925
rect 24213 8959 24271 8965
rect 24213 8925 24225 8959
rect 24259 8925 24271 8959
rect 24213 8919 24271 8925
rect 22572 8888 22600 8919
rect 21928 8860 22600 8888
rect 22664 8888 22692 8919
rect 25406 8916 25412 8968
rect 25464 8965 25470 8968
rect 25464 8959 25492 8965
rect 25480 8925 25492 8959
rect 25464 8919 25492 8925
rect 25464 8916 25470 8919
rect 25590 8916 25596 8968
rect 25648 8916 25654 8968
rect 26712 8965 26740 8996
rect 26973 8993 26985 9027
rect 27019 8993 27031 9027
rect 26973 8987 27031 8993
rect 27246 8984 27252 9036
rect 27304 9024 27310 9036
rect 27522 9024 27528 9036
rect 27304 8996 27528 9024
rect 27304 8984 27310 8996
rect 27522 8984 27528 8996
rect 27580 9024 27586 9036
rect 27709 9027 27767 9033
rect 27709 9024 27721 9027
rect 27580 8996 27721 9024
rect 27580 8984 27586 8996
rect 27709 8993 27721 8996
rect 27755 8993 27767 9027
rect 27709 8987 27767 8993
rect 27798 8984 27804 9036
rect 27856 8984 27862 9036
rect 26697 8959 26755 8965
rect 26697 8925 26709 8959
rect 26743 8925 26755 8959
rect 26697 8919 26755 8925
rect 27617 8959 27675 8965
rect 27617 8925 27629 8959
rect 27663 8956 27675 8959
rect 28350 8956 28356 8968
rect 27663 8928 28356 8956
rect 27663 8925 27675 8928
rect 27617 8919 27675 8925
rect 28350 8916 28356 8928
rect 28408 8916 28414 8968
rect 30392 8956 30420 9055
rect 30834 8984 30840 9036
rect 30892 9024 30898 9036
rect 30929 9027 30987 9033
rect 30929 9024 30941 9027
rect 30892 8996 30941 9024
rect 30892 8984 30898 8996
rect 30929 8993 30941 8996
rect 30975 8993 30987 9027
rect 30929 8987 30987 8993
rect 28460 8928 30420 8956
rect 28460 8888 28488 8928
rect 31018 8916 31024 8968
rect 31076 8956 31082 8968
rect 32048 8956 32076 9132
rect 36725 9129 36737 9132
rect 36771 9129 36783 9163
rect 38378 9160 38384 9172
rect 36725 9123 36783 9129
rect 36832 9132 38384 9160
rect 36832 9092 36860 9132
rect 38378 9120 38384 9132
rect 38436 9120 38442 9172
rect 38473 9163 38531 9169
rect 38473 9129 38485 9163
rect 38519 9160 38531 9163
rect 40770 9160 40776 9172
rect 38519 9132 40776 9160
rect 38519 9129 38531 9132
rect 38473 9123 38531 9129
rect 40770 9120 40776 9132
rect 40828 9120 40834 9172
rect 42705 9163 42763 9169
rect 42705 9129 42717 9163
rect 42751 9160 42763 9163
rect 42794 9160 42800 9172
rect 42751 9132 42800 9160
rect 42751 9129 42763 9132
rect 42705 9123 42763 9129
rect 42794 9120 42800 9132
rect 42852 9120 42858 9172
rect 33152 9064 36860 9092
rect 31076 8928 32076 8956
rect 32125 8959 32183 8965
rect 31076 8916 31082 8928
rect 32125 8925 32137 8959
rect 32171 8956 32183 8959
rect 32214 8956 32220 8968
rect 32171 8928 32220 8956
rect 32171 8925 32183 8928
rect 32125 8919 32183 8925
rect 32214 8916 32220 8928
rect 32272 8916 32278 8968
rect 33152 8956 33180 9064
rect 37366 9024 37372 9036
rect 36372 8996 37372 9024
rect 36372 8965 36400 8996
rect 37366 8984 37372 8996
rect 37424 8984 37430 9036
rect 32324 8928 33180 8956
rect 36173 8959 36231 8965
rect 32324 8888 32352 8928
rect 36173 8925 36185 8959
rect 36219 8925 36231 8959
rect 36173 8919 36231 8925
rect 36357 8959 36415 8965
rect 36357 8925 36369 8959
rect 36403 8925 36415 8959
rect 36357 8919 36415 8925
rect 32398 8897 32404 8900
rect 22664 8860 24164 8888
rect 16485 8823 16543 8829
rect 16485 8820 16497 8823
rect 16224 8792 16497 8820
rect 16485 8789 16497 8792
rect 16531 8820 16543 8823
rect 16574 8820 16580 8832
rect 16531 8792 16580 8820
rect 16531 8789 16543 8792
rect 16485 8783 16543 8789
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 16942 8780 16948 8832
rect 17000 8820 17006 8832
rect 18874 8820 18880 8832
rect 17000 8792 18880 8820
rect 17000 8780 17006 8792
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 19058 8780 19064 8832
rect 19116 8820 19122 8832
rect 20438 8820 20444 8832
rect 19116 8792 20444 8820
rect 19116 8780 19122 8792
rect 20438 8780 20444 8792
rect 20496 8780 20502 8832
rect 21726 8780 21732 8832
rect 21784 8780 21790 8832
rect 22373 8823 22431 8829
rect 22373 8789 22385 8823
rect 22419 8820 22431 8823
rect 22462 8820 22468 8832
rect 22419 8792 22468 8820
rect 22419 8789 22431 8792
rect 22373 8783 22431 8789
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 22572 8820 22600 8860
rect 23566 8820 23572 8832
rect 22572 8792 23572 8820
rect 23566 8780 23572 8792
rect 23624 8780 23630 8832
rect 24026 8780 24032 8832
rect 24084 8780 24090 8832
rect 24136 8820 24164 8860
rect 26068 8860 28488 8888
rect 28644 8860 32352 8888
rect 26068 8820 26096 8860
rect 24136 8792 26096 8820
rect 26234 8780 26240 8832
rect 26292 8780 26298 8832
rect 26789 8823 26847 8829
rect 26789 8789 26801 8823
rect 26835 8820 26847 8823
rect 27522 8820 27528 8832
rect 26835 8792 27528 8820
rect 26835 8789 26847 8792
rect 26789 8783 26847 8789
rect 27522 8780 27528 8792
rect 27580 8820 27586 8832
rect 28644 8820 28672 8860
rect 32392 8851 32404 8897
rect 32398 8848 32404 8851
rect 32456 8848 32462 8900
rect 36188 8888 36216 8919
rect 36446 8916 36452 8968
rect 36504 8916 36510 8968
rect 36538 8916 36544 8968
rect 36596 8965 36602 8968
rect 36596 8919 36604 8965
rect 37461 8959 37519 8965
rect 37461 8925 37473 8959
rect 37507 8925 37519 8959
rect 37461 8919 37519 8925
rect 36596 8916 36602 8919
rect 37366 8888 37372 8900
rect 36188 8860 37372 8888
rect 37366 8848 37372 8860
rect 37424 8848 37430 8900
rect 27580 8792 28672 8820
rect 27580 8780 27586 8792
rect 30742 8780 30748 8832
rect 30800 8780 30806 8832
rect 30837 8823 30895 8829
rect 30837 8789 30849 8823
rect 30883 8820 30895 8823
rect 33042 8820 33048 8832
rect 30883 8792 33048 8820
rect 30883 8789 30895 8792
rect 30837 8783 30895 8789
rect 33042 8780 33048 8792
rect 33100 8780 33106 8832
rect 33505 8823 33563 8829
rect 33505 8789 33517 8823
rect 33551 8820 33563 8823
rect 33594 8820 33600 8832
rect 33551 8792 33600 8820
rect 33551 8789 33563 8792
rect 33505 8783 33563 8789
rect 33594 8780 33600 8792
rect 33652 8780 33658 8832
rect 35802 8780 35808 8832
rect 35860 8820 35866 8832
rect 37476 8820 37504 8919
rect 37734 8916 37740 8968
rect 37792 8916 37798 8968
rect 39666 8916 39672 8968
rect 39724 8916 39730 8968
rect 42702 8916 42708 8968
rect 42760 8916 42766 8968
rect 42886 8916 42892 8968
rect 42944 8916 42950 8968
rect 42981 8959 43039 8965
rect 42981 8925 42993 8959
rect 43027 8956 43039 8959
rect 43254 8956 43260 8968
rect 43027 8928 43260 8956
rect 43027 8925 43039 8928
rect 42981 8919 43039 8925
rect 43254 8916 43260 8928
rect 43312 8916 43318 8968
rect 37918 8848 37924 8900
rect 37976 8888 37982 8900
rect 38657 8891 38715 8897
rect 38657 8888 38669 8891
rect 37976 8860 38669 8888
rect 37976 8848 37982 8860
rect 38657 8857 38669 8860
rect 38703 8857 38715 8891
rect 38657 8851 38715 8857
rect 35860 8792 37504 8820
rect 35860 8780 35866 8792
rect 38470 8780 38476 8832
rect 38528 8820 38534 8832
rect 38749 8823 38807 8829
rect 38749 8820 38761 8823
rect 38528 8792 38761 8820
rect 38528 8780 38534 8792
rect 38749 8789 38761 8792
rect 38795 8789 38807 8823
rect 38749 8783 38807 8789
rect 1104 8730 47104 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 47104 8730
rect 1104 8656 47104 8678
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 7892 8588 8401 8616
rect 7892 8576 7898 8588
rect 8389 8585 8401 8588
rect 8435 8616 8447 8619
rect 8754 8616 8760 8628
rect 8435 8588 8760 8616
rect 8435 8585 8447 8588
rect 8389 8579 8447 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9398 8576 9404 8628
rect 9456 8616 9462 8628
rect 13998 8616 14004 8628
rect 9456 8588 14004 8616
rect 9456 8576 9462 8588
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 14645 8619 14703 8625
rect 14108 8588 14596 8616
rect 8018 8508 8024 8560
rect 8076 8548 8082 8560
rect 8076 8520 8616 8548
rect 8076 8508 8082 8520
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8480 7987 8483
rect 8294 8480 8300 8492
rect 7975 8452 8300 8480
rect 7975 8449 7987 8452
rect 7929 8443 7987 8449
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 8478 8440 8484 8492
rect 8536 8440 8542 8492
rect 8588 8421 8616 8520
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8480 10747 8483
rect 11698 8480 11704 8492
rect 10735 8452 11704 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 12434 8440 12440 8492
rect 12492 8480 12498 8492
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12492 8452 12909 8480
rect 12492 8440 12498 8452
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 13906 8440 13912 8492
rect 13964 8440 13970 8492
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 12250 8412 12256 8424
rect 8619 8384 12256 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 12621 8415 12679 8421
rect 12621 8381 12633 8415
rect 12667 8412 12679 8415
rect 14108 8412 14136 8588
rect 12667 8384 14136 8412
rect 12667 8381 12679 8384
rect 12621 8375 12679 8381
rect 14182 8372 14188 8424
rect 14240 8372 14246 8424
rect 14568 8412 14596 8588
rect 14645 8585 14657 8619
rect 14691 8616 14703 8619
rect 14691 8588 14964 8616
rect 14691 8585 14703 8588
rect 14645 8579 14703 8585
rect 14936 8548 14964 8588
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 16301 8619 16359 8625
rect 16301 8616 16313 8619
rect 15620 8588 16313 8616
rect 15620 8576 15626 8588
rect 16301 8585 16313 8588
rect 16347 8616 16359 8619
rect 18138 8616 18144 8628
rect 16347 8588 18144 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 18138 8576 18144 8588
rect 18196 8576 18202 8628
rect 18969 8619 19027 8625
rect 18969 8585 18981 8619
rect 19015 8616 19027 8619
rect 20070 8616 20076 8628
rect 19015 8588 20076 8616
rect 19015 8585 19027 8588
rect 18969 8579 19027 8585
rect 20070 8576 20076 8588
rect 20128 8576 20134 8628
rect 20898 8576 20904 8628
rect 20956 8576 20962 8628
rect 22186 8576 22192 8628
rect 22244 8616 22250 8628
rect 22281 8619 22339 8625
rect 22281 8616 22293 8619
rect 22244 8588 22293 8616
rect 22244 8576 22250 8588
rect 22281 8585 22293 8588
rect 22327 8585 22339 8619
rect 22281 8579 22339 8585
rect 24394 8576 24400 8628
rect 24452 8616 24458 8628
rect 25590 8616 25596 8628
rect 24452 8588 25596 8616
rect 24452 8576 24458 8588
rect 25590 8576 25596 8588
rect 25648 8576 25654 8628
rect 25958 8576 25964 8628
rect 26016 8616 26022 8628
rect 26053 8619 26111 8625
rect 26053 8616 26065 8619
rect 26016 8588 26065 8616
rect 26016 8576 26022 8588
rect 26053 8585 26065 8588
rect 26099 8585 26111 8619
rect 26053 8579 26111 8585
rect 31294 8576 31300 8628
rect 31352 8576 31358 8628
rect 32309 8619 32367 8625
rect 32309 8585 32321 8619
rect 32355 8616 32367 8619
rect 32398 8616 32404 8628
rect 32355 8588 32404 8616
rect 32355 8585 32367 8588
rect 32309 8579 32367 8585
rect 32398 8576 32404 8588
rect 32456 8576 32462 8628
rect 34790 8576 34796 8628
rect 34848 8576 34854 8628
rect 37918 8616 37924 8628
rect 36096 8588 37924 8616
rect 36096 8560 36124 8588
rect 37918 8576 37924 8588
rect 37976 8576 37982 8628
rect 38013 8619 38071 8625
rect 38013 8585 38025 8619
rect 38059 8616 38071 8619
rect 39758 8616 39764 8628
rect 38059 8588 39764 8616
rect 38059 8585 38071 8588
rect 38013 8579 38071 8585
rect 39758 8576 39764 8588
rect 39816 8576 39822 8628
rect 39850 8576 39856 8628
rect 39908 8576 39914 8628
rect 15166 8551 15224 8557
rect 15166 8548 15178 8551
rect 14936 8520 15178 8548
rect 15166 8517 15178 8520
rect 15212 8517 15224 8551
rect 15166 8511 15224 8517
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 21784 8520 23980 8548
rect 21784 8508 21790 8520
rect 14826 8440 14832 8492
rect 14884 8440 14890 8492
rect 16942 8480 16948 8492
rect 14936 8452 16948 8480
rect 14936 8421 14964 8452
rect 16942 8440 16948 8452
rect 17000 8440 17006 8492
rect 18138 8440 18144 8492
rect 18196 8489 18202 8492
rect 18196 8483 18224 8489
rect 18212 8449 18224 8483
rect 18196 8443 18224 8449
rect 18196 8440 18202 8443
rect 21818 8440 21824 8492
rect 21876 8440 21882 8492
rect 23106 8440 23112 8492
rect 23164 8440 23170 8492
rect 23952 8480 23980 8520
rect 24026 8508 24032 8560
rect 24084 8548 24090 8560
rect 24918 8551 24976 8557
rect 24918 8548 24930 8551
rect 24084 8520 24930 8548
rect 24084 8508 24090 8520
rect 24918 8517 24930 8520
rect 24964 8517 24976 8551
rect 24918 8511 24976 8517
rect 35989 8551 36047 8557
rect 35989 8517 36001 8551
rect 36035 8548 36047 8551
rect 36078 8548 36084 8560
rect 36035 8520 36084 8548
rect 36035 8517 36047 8520
rect 35989 8511 36047 8517
rect 36078 8508 36084 8520
rect 36136 8508 36142 8560
rect 37550 8508 37556 8560
rect 37608 8548 37614 8560
rect 38740 8551 38798 8557
rect 37608 8520 38240 8548
rect 37608 8508 37614 8520
rect 29546 8480 29552 8492
rect 23952 8452 29552 8480
rect 29546 8440 29552 8452
rect 29604 8440 29610 8492
rect 30650 8440 30656 8492
rect 30708 8440 30714 8492
rect 32490 8440 32496 8492
rect 32548 8440 32554 8492
rect 34146 8440 34152 8492
rect 34204 8440 34210 8492
rect 37642 8440 37648 8492
rect 37700 8440 37706 8492
rect 37901 8483 37959 8489
rect 37901 8449 37913 8483
rect 37947 8480 37959 8483
rect 38010 8480 38016 8492
rect 37947 8452 38016 8480
rect 37947 8449 37959 8452
rect 37901 8443 37959 8449
rect 38010 8440 38016 8452
rect 38068 8440 38074 8492
rect 38212 8489 38240 8520
rect 38740 8517 38752 8551
rect 38786 8548 38798 8551
rect 39666 8548 39672 8560
rect 38786 8520 39672 8548
rect 38786 8517 38798 8520
rect 38740 8511 38798 8517
rect 39666 8508 39672 8520
rect 39724 8508 39730 8560
rect 38197 8483 38255 8489
rect 38197 8449 38209 8483
rect 38243 8449 38255 8483
rect 40218 8480 40224 8492
rect 38197 8443 38255 8449
rect 38396 8452 40224 8480
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14568 8384 14933 8412
rect 14921 8381 14933 8384
rect 14967 8381 14979 8415
rect 14921 8375 14979 8381
rect 17129 8415 17187 8421
rect 17129 8381 17141 8415
rect 17175 8412 17187 8415
rect 17218 8412 17224 8424
rect 17175 8384 17224 8412
rect 17175 8381 17187 8384
rect 17129 8375 17187 8381
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8412 17371 8415
rect 17678 8412 17684 8424
rect 17359 8384 17684 8412
rect 17359 8381 17371 8384
rect 17313 8375 17371 8381
rect 17678 8372 17684 8384
rect 17736 8372 17742 8424
rect 18046 8412 18052 8424
rect 17880 8384 18052 8412
rect 7282 8304 7288 8356
rect 7340 8344 7346 8356
rect 8021 8347 8079 8353
rect 8021 8344 8033 8347
rect 7340 8316 8033 8344
rect 7340 8304 7346 8316
rect 8021 8313 8033 8316
rect 8067 8313 8079 8347
rect 8021 8307 8079 8313
rect 13541 8347 13599 8353
rect 13541 8313 13553 8347
rect 13587 8344 13599 8347
rect 14274 8344 14280 8356
rect 13587 8316 14280 8344
rect 13587 8313 13599 8316
rect 13541 8307 13599 8313
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 17494 8304 17500 8356
rect 17552 8344 17558 8356
rect 17773 8347 17831 8353
rect 17773 8344 17785 8347
rect 17552 8316 17785 8344
rect 17552 8304 17558 8316
rect 17773 8313 17785 8316
rect 17819 8313 17831 8347
rect 17773 8307 17831 8313
rect 7742 8236 7748 8288
rect 7800 8236 7806 8288
rect 10502 8236 10508 8288
rect 10560 8236 10566 8288
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 17880 8276 17908 8384
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 18325 8415 18383 8421
rect 18325 8381 18337 8415
rect 18371 8412 18383 8415
rect 18966 8412 18972 8424
rect 18371 8384 18972 8412
rect 18371 8381 18383 8384
rect 18325 8375 18383 8381
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 19058 8372 19064 8424
rect 19116 8372 19122 8424
rect 19245 8415 19303 8421
rect 19245 8381 19257 8415
rect 19291 8412 19303 8415
rect 19291 8384 19564 8412
rect 19291 8381 19303 8384
rect 19245 8375 19303 8381
rect 19536 8356 19564 8384
rect 19610 8372 19616 8424
rect 19668 8412 19674 8424
rect 19981 8415 20039 8421
rect 19981 8412 19993 8415
rect 19668 8384 19993 8412
rect 19668 8372 19674 8384
rect 19518 8304 19524 8356
rect 19576 8304 19582 8356
rect 19702 8304 19708 8356
rect 19760 8304 19766 8356
rect 13872 8248 17908 8276
rect 19812 8276 19840 8384
rect 19981 8381 19993 8384
rect 20027 8381 20039 8415
rect 19981 8375 20039 8381
rect 20070 8372 20076 8424
rect 20128 8421 20134 8424
rect 20128 8415 20156 8421
rect 20144 8381 20156 8415
rect 20128 8375 20156 8381
rect 20257 8415 20315 8421
rect 20257 8381 20269 8415
rect 20303 8412 20315 8415
rect 20622 8412 20628 8424
rect 20303 8384 20628 8412
rect 20303 8381 20315 8384
rect 20257 8375 20315 8381
rect 20128 8372 20134 8375
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 24486 8372 24492 8424
rect 24544 8412 24550 8424
rect 24673 8415 24731 8421
rect 24673 8412 24685 8415
rect 24544 8384 24685 8412
rect 24544 8372 24550 8384
rect 24673 8381 24685 8384
rect 24719 8381 24731 8415
rect 24673 8375 24731 8381
rect 29454 8372 29460 8424
rect 29512 8372 29518 8424
rect 29638 8372 29644 8424
rect 29696 8372 29702 8424
rect 30098 8372 30104 8424
rect 30156 8372 30162 8424
rect 30374 8372 30380 8424
rect 30432 8372 30438 8424
rect 30558 8421 30564 8424
rect 30515 8415 30564 8421
rect 30515 8381 30527 8415
rect 30561 8381 30564 8415
rect 30515 8375 30564 8381
rect 30558 8372 30564 8375
rect 30616 8372 30622 8424
rect 32674 8372 32680 8424
rect 32732 8412 32738 8424
rect 32953 8415 33011 8421
rect 32953 8412 32965 8415
rect 32732 8384 32965 8412
rect 32732 8372 32738 8384
rect 32953 8381 32965 8384
rect 32999 8381 33011 8415
rect 32953 8375 33011 8381
rect 33137 8415 33195 8421
rect 33137 8381 33149 8415
rect 33183 8381 33195 8415
rect 33137 8375 33195 8381
rect 22094 8304 22100 8356
rect 22152 8304 22158 8356
rect 23014 8304 23020 8356
rect 23072 8344 23078 8356
rect 23658 8344 23664 8356
rect 23072 8316 23664 8344
rect 23072 8304 23078 8316
rect 23658 8304 23664 8316
rect 23716 8304 23722 8356
rect 20162 8276 20168 8288
rect 19812 8248 20168 8276
rect 13872 8236 13878 8248
rect 20162 8236 20168 8248
rect 20220 8236 20226 8288
rect 22830 8236 22836 8288
rect 22888 8276 22894 8288
rect 22925 8279 22983 8285
rect 22925 8276 22937 8279
rect 22888 8248 22937 8276
rect 22888 8236 22894 8248
rect 22925 8245 22937 8248
rect 22971 8245 22983 8279
rect 22925 8239 22983 8245
rect 23474 8236 23480 8288
rect 23532 8276 23538 8288
rect 30834 8276 30840 8288
rect 23532 8248 30840 8276
rect 23532 8236 23538 8248
rect 30834 8236 30840 8248
rect 30892 8236 30898 8288
rect 32950 8236 32956 8288
rect 33008 8276 33014 8288
rect 33152 8276 33180 8375
rect 33686 8372 33692 8424
rect 33744 8412 33750 8424
rect 33873 8415 33931 8421
rect 33873 8412 33885 8415
rect 33744 8384 33885 8412
rect 33744 8372 33750 8384
rect 33873 8381 33885 8384
rect 33919 8381 33931 8415
rect 33873 8375 33931 8381
rect 33962 8372 33968 8424
rect 34020 8421 34026 8424
rect 34020 8415 34048 8421
rect 34036 8381 34048 8415
rect 38105 8415 38163 8421
rect 34020 8375 34048 8381
rect 34624 8384 36308 8412
rect 34020 8372 34026 8375
rect 34624 8356 34652 8384
rect 33410 8304 33416 8356
rect 33468 8344 33474 8356
rect 33597 8347 33655 8353
rect 33597 8344 33609 8347
rect 33468 8316 33609 8344
rect 33468 8304 33474 8316
rect 33597 8313 33609 8316
rect 33643 8313 33655 8347
rect 33597 8307 33655 8313
rect 34606 8304 34612 8356
rect 34664 8304 34670 8356
rect 35342 8304 35348 8356
rect 35400 8344 35406 8356
rect 36173 8347 36231 8353
rect 36173 8344 36185 8347
rect 35400 8316 36185 8344
rect 35400 8304 35406 8316
rect 36173 8313 36185 8316
rect 36219 8313 36231 8347
rect 36280 8344 36308 8384
rect 38105 8381 38117 8415
rect 38151 8412 38163 8415
rect 38396 8412 38424 8452
rect 40218 8440 40224 8452
rect 40276 8440 40282 8492
rect 46106 8440 46112 8492
rect 46164 8480 46170 8492
rect 46201 8483 46259 8489
rect 46201 8480 46213 8483
rect 46164 8452 46213 8480
rect 46164 8440 46170 8452
rect 46201 8449 46213 8452
rect 46247 8449 46259 8483
rect 46201 8443 46259 8449
rect 38151 8384 38424 8412
rect 38151 8381 38163 8384
rect 38105 8375 38163 8381
rect 38470 8372 38476 8424
rect 38528 8372 38534 8424
rect 45922 8372 45928 8424
rect 45980 8372 45986 8424
rect 38488 8344 38516 8372
rect 36280 8316 38516 8344
rect 36173 8307 36231 8313
rect 34330 8276 34336 8288
rect 33008 8248 34336 8276
rect 33008 8236 33014 8248
rect 34330 8236 34336 8248
rect 34388 8236 34394 8288
rect 37458 8236 37464 8288
rect 37516 8236 37522 8288
rect 1104 8186 47104 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 47104 8186
rect 1104 8112 47104 8134
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8352 8044 8953 8072
rect 8352 8032 8358 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 11606 8032 11612 8084
rect 11664 8032 11670 8084
rect 11698 8032 11704 8084
rect 11756 8032 11762 8084
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 13964 8044 17080 8072
rect 13964 8032 13970 8044
rect 8754 7964 8760 8016
rect 8812 7964 8818 8016
rect 8478 7896 8484 7948
rect 8536 7936 8542 7948
rect 9398 7936 9404 7948
rect 8536 7908 9404 7936
rect 8536 7896 8542 7908
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 9585 7939 9643 7945
rect 9585 7905 9597 7939
rect 9631 7936 9643 7939
rect 9858 7936 9864 7948
rect 9631 7908 9864 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 9858 7896 9864 7908
rect 9916 7896 9922 7948
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10226 7936 10232 7948
rect 10008 7908 10232 7936
rect 10008 7896 10014 7908
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 12250 7896 12256 7948
rect 12308 7896 12314 7948
rect 15013 7939 15071 7945
rect 15013 7936 15025 7939
rect 14200 7908 15025 7936
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 7374 7828 7380 7880
rect 7432 7828 7438 7880
rect 10502 7877 10508 7880
rect 10496 7868 10508 7877
rect 10463 7840 10508 7868
rect 10496 7831 10508 7840
rect 10502 7828 10508 7831
rect 10560 7828 10566 7880
rect 11606 7828 11612 7880
rect 11664 7868 11670 7880
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 11664 7840 12081 7868
rect 11664 7828 11670 7840
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12492 7840 12541 7868
rect 12492 7828 12498 7840
rect 12529 7837 12541 7840
rect 12575 7837 12587 7871
rect 14200 7868 14228 7908
rect 15013 7905 15025 7908
rect 15059 7936 15071 7939
rect 15654 7936 15660 7948
rect 15059 7908 15660 7936
rect 15059 7905 15071 7908
rect 15013 7899 15071 7905
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 12529 7831 12587 7837
rect 12636 7840 14228 7868
rect 12636 7812 12664 7840
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 14550 7828 14556 7880
rect 14608 7828 14614 7880
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7868 15807 7871
rect 16758 7868 16764 7880
rect 15795 7840 16764 7868
rect 15795 7837 15807 7840
rect 15749 7831 15807 7837
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 7622 7803 7680 7809
rect 7622 7800 7634 7803
rect 7116 7772 7634 7800
rect 7116 7741 7144 7772
rect 7622 7769 7634 7772
rect 7668 7769 7680 7803
rect 7622 7763 7680 7769
rect 10962 7760 10968 7812
rect 11020 7800 11026 7812
rect 11974 7800 11980 7812
rect 11020 7772 11980 7800
rect 11020 7760 11026 7772
rect 11974 7760 11980 7772
rect 12032 7800 12038 7812
rect 12161 7803 12219 7809
rect 12161 7800 12173 7803
rect 12032 7772 12173 7800
rect 12032 7760 12038 7772
rect 12161 7769 12173 7772
rect 12207 7800 12219 7803
rect 12618 7800 12624 7812
rect 12207 7772 12624 7800
rect 12207 7769 12219 7772
rect 12161 7763 12219 7769
rect 12618 7760 12624 7772
rect 12676 7760 12682 7812
rect 12796 7803 12854 7809
rect 12796 7769 12808 7803
rect 12842 7800 12854 7803
rect 12842 7772 14136 7800
rect 12842 7769 12854 7772
rect 12796 7763 12854 7769
rect 7101 7735 7159 7741
rect 7101 7701 7113 7735
rect 7147 7701 7159 7735
rect 7101 7695 7159 7701
rect 9306 7692 9312 7744
rect 9364 7692 9370 7744
rect 14108 7741 14136 7772
rect 14182 7760 14188 7812
rect 14240 7800 14246 7812
rect 16022 7809 16028 7812
rect 14829 7803 14887 7809
rect 14829 7800 14841 7803
rect 14240 7772 14841 7800
rect 14240 7760 14246 7772
rect 14829 7769 14841 7772
rect 14875 7769 14887 7803
rect 14829 7763 14887 7769
rect 16016 7763 16028 7809
rect 16022 7760 16028 7763
rect 16080 7760 16086 7812
rect 14093 7735 14151 7741
rect 14093 7701 14105 7735
rect 14139 7701 14151 7735
rect 14093 7695 14151 7701
rect 14366 7692 14372 7744
rect 14424 7692 14430 7744
rect 17052 7732 17080 8044
rect 17126 8032 17132 8084
rect 17184 8072 17190 8084
rect 19061 8075 19119 8081
rect 17184 8044 19012 8072
rect 17184 8032 17190 8044
rect 17862 7964 17868 8016
rect 17920 7964 17926 8016
rect 18984 8004 19012 8044
rect 19061 8041 19073 8075
rect 19107 8072 19119 8075
rect 19107 8044 20852 8072
rect 19107 8041 19119 8044
rect 19061 8035 19119 8041
rect 19978 8004 19984 8016
rect 18984 7976 19984 8004
rect 19978 7964 19984 7976
rect 20036 7964 20042 8016
rect 20824 8004 20852 8044
rect 21082 8032 21088 8084
rect 21140 8032 21146 8084
rect 21174 8032 21180 8084
rect 21232 8072 21238 8084
rect 21232 8044 25544 8072
rect 21232 8032 21238 8044
rect 22094 8004 22100 8016
rect 20824 7976 22100 8004
rect 22094 7964 22100 7976
rect 22152 7964 22158 8016
rect 24949 8007 25007 8013
rect 24949 7973 24961 8007
rect 24995 8004 25007 8007
rect 25130 8004 25136 8016
rect 24995 7976 25136 8004
rect 24995 7973 25007 7976
rect 24949 7967 25007 7973
rect 25130 7964 25136 7976
rect 25188 7964 25194 8016
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 17770 7936 17776 7948
rect 17276 7908 17776 7936
rect 17276 7896 17282 7908
rect 17770 7896 17776 7908
rect 17828 7896 17834 7948
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 18012 7908 18153 7936
rect 18012 7896 18018 7908
rect 18141 7905 18153 7908
rect 18187 7905 18199 7939
rect 18141 7899 18199 7905
rect 18230 7896 18236 7948
rect 18288 7945 18294 7948
rect 18288 7939 18316 7945
rect 18304 7905 18316 7939
rect 18288 7899 18316 7905
rect 18417 7939 18475 7945
rect 18417 7905 18429 7939
rect 18463 7936 18475 7939
rect 18463 7908 19012 7936
rect 18463 7905 18475 7908
rect 18417 7899 18475 7905
rect 18288 7896 18294 7899
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7868 17463 7871
rect 17586 7868 17592 7880
rect 17451 7840 17592 7868
rect 17451 7837 17463 7840
rect 17405 7831 17463 7837
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 18984 7868 19012 7908
rect 19058 7896 19064 7948
rect 19116 7936 19122 7948
rect 19245 7939 19303 7945
rect 19245 7936 19257 7939
rect 19116 7908 19257 7936
rect 19116 7896 19122 7908
rect 19245 7905 19257 7908
rect 19291 7936 19303 7939
rect 19334 7936 19340 7948
rect 19291 7908 19340 7936
rect 19291 7905 19303 7908
rect 19245 7899 19303 7905
rect 19334 7896 19340 7908
rect 19392 7896 19398 7948
rect 19429 7939 19487 7945
rect 19429 7905 19441 7939
rect 19475 7936 19487 7939
rect 19518 7936 19524 7948
rect 19475 7908 19524 7936
rect 19475 7905 19487 7908
rect 19429 7899 19487 7905
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 19886 7896 19892 7948
rect 19944 7896 19950 7948
rect 19996 7936 20024 7964
rect 20282 7939 20340 7945
rect 20282 7936 20294 7939
rect 19996 7908 20294 7936
rect 20282 7905 20294 7908
rect 20328 7905 20340 7939
rect 20282 7899 20340 7905
rect 20438 7896 20444 7948
rect 20496 7896 20502 7948
rect 25516 7945 25544 8044
rect 30742 8032 30748 8084
rect 30800 8072 30806 8084
rect 31389 8075 31447 8081
rect 31389 8072 31401 8075
rect 30800 8044 31401 8072
rect 30800 8032 30806 8044
rect 31389 8041 31401 8044
rect 31435 8041 31447 8075
rect 31389 8035 31447 8041
rect 31849 8075 31907 8081
rect 31849 8041 31861 8075
rect 31895 8072 31907 8075
rect 32490 8072 32496 8084
rect 31895 8044 32496 8072
rect 31895 8041 31907 8044
rect 31849 8035 31907 8041
rect 32490 8032 32496 8044
rect 32548 8032 32554 8084
rect 33042 8032 33048 8084
rect 33100 8072 33106 8084
rect 34517 8075 34575 8081
rect 34517 8072 34529 8075
rect 33100 8044 34529 8072
rect 33100 8032 33106 8044
rect 34517 8041 34529 8044
rect 34563 8041 34575 8075
rect 36262 8072 36268 8084
rect 34517 8035 34575 8041
rect 34716 8044 36268 8072
rect 29380 7976 30328 8004
rect 25501 7939 25559 7945
rect 22066 7908 22692 7936
rect 19150 7868 19156 7880
rect 18984 7840 19156 7868
rect 19150 7828 19156 7840
rect 19208 7828 19214 7880
rect 19610 7868 19616 7880
rect 19444 7840 19616 7868
rect 19444 7732 19472 7840
rect 19610 7828 19616 7840
rect 19668 7828 19674 7880
rect 20162 7828 20168 7880
rect 20220 7828 20226 7880
rect 17052 7704 19472 7732
rect 19610 7692 19616 7744
rect 19668 7732 19674 7744
rect 22066 7732 22094 7908
rect 22557 7871 22615 7877
rect 22557 7837 22569 7871
rect 22603 7837 22615 7871
rect 22557 7831 22615 7837
rect 19668 7704 22094 7732
rect 22572 7732 22600 7831
rect 22664 7800 22692 7908
rect 25501 7905 25513 7939
rect 25547 7905 25559 7939
rect 25501 7899 25559 7905
rect 26510 7896 26516 7948
rect 26568 7936 26574 7948
rect 27798 7936 27804 7948
rect 26568 7908 27804 7936
rect 26568 7896 26574 7908
rect 27798 7896 27804 7908
rect 27856 7936 27862 7948
rect 28077 7939 28135 7945
rect 28077 7936 28089 7939
rect 27856 7908 28089 7936
rect 27856 7896 27862 7908
rect 28077 7905 28089 7908
rect 28123 7905 28135 7939
rect 28077 7899 28135 7905
rect 22830 7877 22836 7880
rect 22824 7868 22836 7877
rect 22791 7840 22836 7868
rect 22824 7831 22836 7840
rect 22830 7828 22836 7831
rect 22888 7828 22894 7880
rect 25317 7871 25375 7877
rect 25317 7837 25329 7871
rect 25363 7868 25375 7871
rect 26234 7868 26240 7880
rect 25363 7840 26240 7868
rect 25363 7837 25375 7840
rect 25317 7831 25375 7837
rect 26234 7828 26240 7840
rect 26292 7828 26298 7880
rect 27893 7871 27951 7877
rect 27893 7837 27905 7871
rect 27939 7868 27951 7871
rect 28534 7868 28540 7880
rect 27939 7840 28540 7868
rect 27939 7837 27951 7840
rect 27893 7831 27951 7837
rect 28534 7828 28540 7840
rect 28592 7868 28598 7880
rect 29380 7868 29408 7976
rect 29454 7896 29460 7948
rect 29512 7936 29518 7948
rect 29549 7939 29607 7945
rect 29549 7936 29561 7939
rect 29512 7908 29561 7936
rect 29512 7896 29518 7908
rect 29549 7905 29561 7908
rect 29595 7936 29607 7939
rect 30098 7936 30104 7948
rect 29595 7908 30104 7936
rect 29595 7905 29607 7908
rect 29549 7899 29607 7905
rect 30098 7896 30104 7908
rect 30156 7896 30162 7948
rect 30190 7896 30196 7948
rect 30248 7896 30254 7948
rect 30300 7936 30328 7976
rect 32232 7976 33456 8004
rect 30558 7936 30564 7948
rect 30616 7945 30622 7948
rect 30616 7939 30644 7945
rect 30300 7908 30564 7936
rect 30558 7896 30564 7908
rect 30632 7905 30644 7939
rect 30616 7899 30644 7905
rect 30616 7896 30622 7899
rect 28592 7840 29408 7868
rect 28592 7828 28598 7840
rect 29638 7828 29644 7880
rect 29696 7868 29702 7880
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 29696 7840 29745 7868
rect 29696 7828 29702 7840
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 30466 7828 30472 7880
rect 30524 7828 30530 7880
rect 30742 7828 30748 7880
rect 30800 7828 30806 7880
rect 32232 7877 32260 7976
rect 32493 7939 32551 7945
rect 32493 7905 32505 7939
rect 32539 7936 32551 7939
rect 32766 7936 32772 7948
rect 32539 7908 32772 7936
rect 32539 7905 32551 7908
rect 32493 7899 32551 7905
rect 32766 7896 32772 7908
rect 32824 7896 32830 7948
rect 32861 7939 32919 7945
rect 32861 7905 32873 7939
rect 32907 7936 32919 7939
rect 32950 7936 32956 7948
rect 32907 7908 32956 7936
rect 32907 7905 32919 7908
rect 32861 7899 32919 7905
rect 32950 7896 32956 7908
rect 33008 7896 33014 7948
rect 33321 7939 33379 7945
rect 33321 7936 33333 7939
rect 33060 7908 33333 7936
rect 33060 7880 33088 7908
rect 33321 7905 33333 7908
rect 33367 7905 33379 7939
rect 33428 7936 33456 7976
rect 34330 7964 34336 8016
rect 34388 8004 34394 8016
rect 34716 8004 34744 8044
rect 36262 8032 36268 8044
rect 36320 8072 36326 8084
rect 36633 8075 36691 8081
rect 36633 8072 36645 8075
rect 36320 8044 36645 8072
rect 36320 8032 36326 8044
rect 36633 8041 36645 8044
rect 36679 8041 36691 8075
rect 36633 8035 36691 8041
rect 38654 8032 38660 8084
rect 38712 8032 38718 8084
rect 34388 7976 34744 8004
rect 34388 7964 34394 7976
rect 33594 7936 33600 7948
rect 33428 7908 33600 7936
rect 33321 7899 33379 7905
rect 33594 7896 33600 7908
rect 33652 7896 33658 7948
rect 34514 7936 34520 7948
rect 33868 7908 34520 7936
rect 33868 7880 33896 7908
rect 34514 7896 34520 7908
rect 34572 7896 34578 7948
rect 34606 7896 34612 7948
rect 34664 7936 34670 7948
rect 35250 7936 35256 7948
rect 34664 7908 35256 7936
rect 34664 7896 34670 7908
rect 35250 7896 35256 7908
rect 35308 7896 35314 7948
rect 32217 7871 32275 7877
rect 32217 7837 32229 7871
rect 32263 7837 32275 7871
rect 32217 7831 32275 7837
rect 32674 7828 32680 7880
rect 32732 7828 32738 7880
rect 33042 7828 33048 7880
rect 33100 7828 33106 7880
rect 33686 7828 33692 7880
rect 33744 7877 33750 7880
rect 33744 7871 33772 7877
rect 33760 7837 33772 7871
rect 33744 7831 33772 7837
rect 33744 7828 33750 7831
rect 33850 7828 33856 7880
rect 33908 7877 33914 7880
rect 33908 7871 33931 7877
rect 33919 7837 33931 7871
rect 33908 7831 33931 7837
rect 33908 7828 33914 7831
rect 35158 7828 35164 7880
rect 35216 7828 35222 7880
rect 38010 7828 38016 7880
rect 38068 7868 38074 7880
rect 38565 7871 38623 7877
rect 38565 7868 38577 7871
rect 38068 7840 38577 7868
rect 38068 7828 38074 7840
rect 38565 7837 38577 7840
rect 38611 7837 38623 7871
rect 38565 7831 38623 7837
rect 38746 7828 38752 7880
rect 38804 7828 38810 7880
rect 27985 7803 28043 7809
rect 27985 7800 27997 7803
rect 22664 7772 27997 7800
rect 27985 7769 27997 7772
rect 28031 7800 28043 7803
rect 29178 7800 29184 7812
rect 28031 7772 29184 7800
rect 28031 7769 28043 7772
rect 27985 7763 28043 7769
rect 29178 7760 29184 7772
rect 29236 7760 29242 7812
rect 35498 7803 35556 7809
rect 35498 7800 35510 7803
rect 34992 7772 35510 7800
rect 23842 7732 23848 7744
rect 22572 7704 23848 7732
rect 19668 7692 19674 7704
rect 23842 7692 23848 7704
rect 23900 7692 23906 7744
rect 23934 7692 23940 7744
rect 23992 7692 23998 7744
rect 25409 7735 25467 7741
rect 25409 7701 25421 7735
rect 25455 7732 25467 7735
rect 26786 7732 26792 7744
rect 25455 7704 26792 7732
rect 25455 7701 25467 7704
rect 25409 7695 25467 7701
rect 26786 7692 26792 7704
rect 26844 7692 26850 7744
rect 27154 7692 27160 7744
rect 27212 7732 27218 7744
rect 27525 7735 27583 7741
rect 27525 7732 27537 7735
rect 27212 7704 27537 7732
rect 27212 7692 27218 7704
rect 27525 7701 27537 7704
rect 27571 7701 27583 7735
rect 29196 7732 29224 7760
rect 31202 7732 31208 7744
rect 29196 7704 31208 7732
rect 27525 7695 27583 7701
rect 31202 7692 31208 7704
rect 31260 7692 31266 7744
rect 32309 7735 32367 7741
rect 32309 7701 32321 7735
rect 32355 7732 32367 7735
rect 33134 7732 33140 7744
rect 32355 7704 33140 7732
rect 32355 7701 32367 7704
rect 32309 7695 32367 7701
rect 33134 7692 33140 7704
rect 33192 7692 33198 7744
rect 34992 7741 35020 7772
rect 35498 7769 35510 7772
rect 35544 7769 35556 7803
rect 35498 7763 35556 7769
rect 34977 7735 35035 7741
rect 34977 7701 34989 7735
rect 35023 7701 35035 7735
rect 34977 7695 35035 7701
rect 1104 7642 47104 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 47104 7642
rect 1104 7568 47104 7590
rect 7650 7488 7656 7540
rect 7708 7528 7714 7540
rect 8849 7531 8907 7537
rect 8849 7528 8861 7531
rect 7708 7500 8861 7528
rect 7708 7488 7714 7500
rect 8849 7497 8861 7500
rect 8895 7528 8907 7531
rect 9306 7528 9312 7540
rect 8895 7500 9312 7528
rect 8895 7497 8907 7500
rect 8849 7491 8907 7497
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 9858 7488 9864 7540
rect 9916 7528 9922 7540
rect 10962 7528 10968 7540
rect 9916 7500 10968 7528
rect 9916 7488 9922 7500
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11333 7531 11391 7537
rect 11333 7528 11345 7531
rect 11296 7500 11345 7528
rect 11296 7488 11302 7500
rect 11333 7497 11345 7500
rect 11379 7528 11391 7531
rect 11885 7531 11943 7537
rect 11885 7528 11897 7531
rect 11379 7500 11897 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 11885 7497 11897 7500
rect 11931 7497 11943 7531
rect 11885 7491 11943 7497
rect 11974 7488 11980 7540
rect 12032 7488 12038 7540
rect 13814 7488 13820 7540
rect 13872 7488 13878 7540
rect 15933 7531 15991 7537
rect 15933 7497 15945 7531
rect 15979 7528 15991 7531
rect 16022 7528 16028 7540
rect 15979 7500 16028 7528
rect 15979 7497 15991 7500
rect 15933 7491 15991 7497
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 16632 7500 18061 7528
rect 16632 7488 16638 7500
rect 18049 7497 18061 7500
rect 18095 7497 18107 7531
rect 18049 7491 18107 7497
rect 18524 7500 18736 7528
rect 7742 7469 7748 7472
rect 7736 7460 7748 7469
rect 7703 7432 7748 7460
rect 7736 7423 7748 7432
rect 7742 7420 7748 7423
rect 7800 7420 7806 7472
rect 12704 7463 12762 7469
rect 9646 7432 10364 7460
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7392 1547 7395
rect 9646 7392 9674 7432
rect 10226 7401 10232 7404
rect 1535 7364 9674 7392
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 10220 7355 10232 7401
rect 10226 7352 10232 7355
rect 10284 7352 10290 7404
rect 10336 7392 10364 7432
rect 12704 7429 12716 7463
rect 12750 7460 12762 7463
rect 14366 7460 14372 7472
rect 12750 7432 14372 7460
rect 12750 7429 12762 7432
rect 12704 7423 12762 7429
rect 14366 7420 14372 7432
rect 14424 7420 14430 7472
rect 17957 7463 18015 7469
rect 14476 7432 16252 7460
rect 14476 7392 14504 7432
rect 10336 7364 14504 7392
rect 16114 7352 16120 7404
rect 16172 7352 16178 7404
rect 16224 7392 16252 7432
rect 17957 7429 17969 7463
rect 18003 7460 18015 7463
rect 18524 7460 18552 7500
rect 18003 7432 18552 7460
rect 18708 7460 18736 7500
rect 18782 7488 18788 7540
rect 18840 7528 18846 7540
rect 20714 7528 20720 7540
rect 18840 7500 20720 7528
rect 18840 7488 18846 7500
rect 20714 7488 20720 7500
rect 20772 7488 20778 7540
rect 20901 7531 20959 7537
rect 20901 7497 20913 7531
rect 20947 7528 20959 7531
rect 20990 7528 20996 7540
rect 20947 7500 20996 7528
rect 20947 7497 20959 7500
rect 20901 7491 20959 7497
rect 20990 7488 20996 7500
rect 21048 7488 21054 7540
rect 22002 7488 22008 7540
rect 22060 7488 22066 7540
rect 23106 7488 23112 7540
rect 23164 7488 23170 7540
rect 23477 7531 23535 7537
rect 23477 7497 23489 7531
rect 23523 7528 23535 7531
rect 23934 7528 23940 7540
rect 23523 7500 23940 7528
rect 23523 7497 23535 7500
rect 23477 7491 23535 7497
rect 23934 7488 23940 7500
rect 23992 7528 23998 7540
rect 25406 7528 25412 7540
rect 23992 7500 25412 7528
rect 23992 7488 23998 7500
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 28721 7531 28779 7537
rect 28721 7528 28733 7531
rect 26804 7500 28733 7528
rect 19610 7460 19616 7472
rect 18708 7432 19616 7460
rect 18003 7429 18015 7432
rect 17957 7423 18015 7429
rect 19610 7420 19616 7432
rect 19668 7420 19674 7472
rect 19702 7420 19708 7472
rect 19760 7460 19766 7472
rect 22373 7463 22431 7469
rect 22373 7460 22385 7463
rect 19760 7432 22385 7460
rect 19760 7420 19766 7432
rect 22373 7429 22385 7432
rect 22419 7429 22431 7463
rect 22373 7423 22431 7429
rect 22465 7463 22523 7469
rect 22465 7429 22477 7463
rect 22511 7460 22523 7463
rect 23658 7460 23664 7472
rect 22511 7432 23664 7460
rect 22511 7429 22523 7432
rect 22465 7423 22523 7429
rect 23658 7420 23664 7432
rect 23716 7420 23722 7472
rect 26510 7460 26516 7472
rect 23768 7432 26516 7460
rect 18782 7392 18788 7404
rect 16224 7364 18788 7392
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 18874 7352 18880 7404
rect 18932 7392 18938 7404
rect 19061 7395 19119 7401
rect 19061 7392 19073 7395
rect 18932 7364 19073 7392
rect 18932 7352 18938 7364
rect 19061 7361 19073 7364
rect 19107 7392 19119 7395
rect 19107 7364 19380 7392
rect 19107 7361 19119 7364
rect 19061 7355 19119 7361
rect 7374 7284 7380 7336
rect 7432 7324 7438 7336
rect 7469 7327 7527 7333
rect 7469 7324 7481 7327
rect 7432 7296 7481 7324
rect 7432 7284 7438 7296
rect 7469 7293 7481 7296
rect 7515 7293 7527 7327
rect 7469 7287 7527 7293
rect 1578 7148 1584 7200
rect 1636 7148 1642 7200
rect 7484 7188 7512 7287
rect 9950 7284 9956 7336
rect 10008 7284 10014 7336
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 12069 7327 12127 7333
rect 12069 7324 12081 7327
rect 11020 7296 12081 7324
rect 11020 7284 11026 7296
rect 12069 7293 12081 7296
rect 12115 7293 12127 7327
rect 12069 7287 12127 7293
rect 12434 7284 12440 7336
rect 12492 7284 12498 7336
rect 17310 7284 17316 7336
rect 17368 7324 17374 7336
rect 17368 7296 19288 7324
rect 17368 7284 17374 7296
rect 16758 7216 16764 7268
rect 16816 7256 16822 7268
rect 18877 7259 18935 7265
rect 18877 7256 18889 7259
rect 16816 7228 18889 7256
rect 16816 7216 16822 7228
rect 18877 7225 18889 7228
rect 18923 7256 18935 7259
rect 18966 7256 18972 7268
rect 18923 7228 18972 7256
rect 18923 7225 18935 7228
rect 18877 7219 18935 7225
rect 18966 7216 18972 7228
rect 19024 7216 19030 7268
rect 9950 7188 9956 7200
rect 7484 7160 9956 7188
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 11514 7148 11520 7200
rect 11572 7148 11578 7200
rect 19058 7148 19064 7200
rect 19116 7188 19122 7200
rect 19153 7191 19211 7197
rect 19153 7188 19165 7191
rect 19116 7160 19165 7188
rect 19116 7148 19122 7160
rect 19153 7157 19165 7160
rect 19199 7157 19211 7191
rect 19260 7188 19288 7296
rect 19352 7256 19380 7364
rect 19518 7352 19524 7404
rect 19576 7352 19582 7404
rect 19886 7352 19892 7404
rect 19944 7392 19950 7404
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 19944 7364 21281 7392
rect 19944 7352 19950 7364
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 23382 7392 23388 7404
rect 21407 7364 23388 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 23382 7352 23388 7364
rect 23440 7352 23446 7404
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 19797 7327 19855 7333
rect 19797 7324 19809 7327
rect 19484 7296 19809 7324
rect 19484 7284 19490 7296
rect 19797 7293 19809 7296
rect 19843 7293 19855 7327
rect 19797 7287 19855 7293
rect 19981 7327 20039 7333
rect 19981 7293 19993 7327
rect 20027 7324 20039 7327
rect 20162 7324 20168 7336
rect 20027 7296 20168 7324
rect 20027 7293 20039 7296
rect 19981 7287 20039 7293
rect 20162 7284 20168 7296
rect 20220 7284 20226 7336
rect 20257 7327 20315 7333
rect 20257 7293 20269 7327
rect 20303 7293 20315 7327
rect 20257 7287 20315 7293
rect 20272 7256 20300 7287
rect 21174 7284 21180 7336
rect 21232 7324 21238 7336
rect 21453 7327 21511 7333
rect 21453 7324 21465 7327
rect 21232 7296 21465 7324
rect 21232 7284 21238 7296
rect 21453 7293 21465 7296
rect 21499 7293 21511 7327
rect 21453 7287 21511 7293
rect 22649 7327 22707 7333
rect 22649 7293 22661 7327
rect 22695 7324 22707 7327
rect 23474 7324 23480 7336
rect 22695 7296 23480 7324
rect 22695 7293 22707 7296
rect 22649 7287 22707 7293
rect 23474 7284 23480 7296
rect 23532 7284 23538 7336
rect 23768 7333 23796 7432
rect 26510 7420 26516 7432
rect 26568 7420 26574 7472
rect 23842 7352 23848 7404
rect 23900 7392 23906 7404
rect 24305 7395 24363 7401
rect 24305 7392 24317 7395
rect 23900 7364 24317 7392
rect 23900 7352 23906 7364
rect 24305 7361 24317 7364
rect 24351 7392 24363 7395
rect 24670 7392 24676 7404
rect 24351 7364 24676 7392
rect 24351 7361 24363 7364
rect 24305 7355 24363 7361
rect 24670 7352 24676 7364
rect 24728 7352 24734 7404
rect 26804 7401 26832 7500
rect 28721 7497 28733 7500
rect 28767 7497 28779 7531
rect 28721 7491 28779 7497
rect 29178 7488 29184 7540
rect 29236 7488 29242 7540
rect 31757 7531 31815 7537
rect 31757 7497 31769 7531
rect 31803 7497 31815 7531
rect 31757 7491 31815 7497
rect 27494 7463 27552 7469
rect 27494 7460 27506 7463
rect 26988 7432 27506 7460
rect 26789 7395 26847 7401
rect 26789 7361 26801 7395
rect 26835 7361 26847 7395
rect 26789 7355 26847 7361
rect 23569 7327 23627 7333
rect 23569 7293 23581 7327
rect 23615 7293 23627 7327
rect 23569 7287 23627 7293
rect 23753 7327 23811 7333
rect 23753 7293 23765 7327
rect 23799 7293 23811 7327
rect 23753 7287 23811 7293
rect 19352 7228 20300 7256
rect 23584 7256 23612 7287
rect 24210 7284 24216 7336
rect 24268 7324 24274 7336
rect 24581 7327 24639 7333
rect 24581 7324 24593 7327
rect 24268 7296 24593 7324
rect 24268 7284 24274 7296
rect 24581 7293 24593 7296
rect 24627 7293 24639 7327
rect 26988 7324 27016 7432
rect 27494 7429 27506 7432
rect 27540 7429 27552 7463
rect 27494 7423 27552 7429
rect 30101 7463 30159 7469
rect 30101 7429 30113 7463
rect 30147 7460 30159 7463
rect 30190 7460 30196 7472
rect 30147 7432 30196 7460
rect 30147 7429 30159 7432
rect 30101 7423 30159 7429
rect 30190 7420 30196 7432
rect 30248 7420 30254 7472
rect 31772 7460 31800 7491
rect 35158 7488 35164 7540
rect 35216 7528 35222 7540
rect 35897 7531 35955 7537
rect 35897 7528 35909 7531
rect 35216 7500 35909 7528
rect 35216 7488 35222 7500
rect 35897 7497 35909 7500
rect 35943 7497 35955 7531
rect 35897 7491 35955 7497
rect 36357 7531 36415 7537
rect 36357 7497 36369 7531
rect 36403 7528 36415 7531
rect 37458 7528 37464 7540
rect 36403 7500 37464 7528
rect 36403 7497 36415 7500
rect 36357 7491 36415 7497
rect 37458 7488 37464 7500
rect 37516 7488 37522 7540
rect 32370 7463 32428 7469
rect 32370 7460 32382 7463
rect 31772 7432 32382 7460
rect 32370 7429 32382 7432
rect 32416 7429 32428 7463
rect 32370 7423 32428 7429
rect 36262 7420 36268 7472
rect 36320 7420 36326 7472
rect 27154 7352 27160 7404
rect 27212 7352 27218 7404
rect 29089 7395 29147 7401
rect 29089 7361 29101 7395
rect 29135 7361 29147 7395
rect 29089 7355 29147 7361
rect 24581 7287 24639 7293
rect 26620 7296 27016 7324
rect 26234 7256 26240 7268
rect 23584 7228 26240 7256
rect 23584 7188 23612 7228
rect 26234 7216 26240 7228
rect 26292 7216 26298 7268
rect 26620 7265 26648 7296
rect 27062 7284 27068 7336
rect 27120 7324 27126 7336
rect 27249 7327 27307 7333
rect 27249 7324 27261 7327
rect 27120 7296 27261 7324
rect 27120 7284 27126 7296
rect 27249 7293 27261 7296
rect 27295 7293 27307 7327
rect 27249 7287 27307 7293
rect 26605 7259 26663 7265
rect 26605 7225 26617 7259
rect 26651 7225 26663 7259
rect 26605 7219 26663 7225
rect 28629 7259 28687 7265
rect 28629 7225 28641 7259
rect 28675 7256 28687 7259
rect 29104 7256 29132 7355
rect 29546 7352 29552 7404
rect 29604 7392 29610 7404
rect 30006 7392 30012 7404
rect 29604 7364 30012 7392
rect 29604 7352 29610 7364
rect 30006 7352 30012 7364
rect 30064 7392 30070 7404
rect 30064 7364 30328 7392
rect 30064 7352 30070 7364
rect 29270 7284 29276 7336
rect 29328 7284 29334 7336
rect 29822 7284 29828 7336
rect 29880 7324 29886 7336
rect 30300 7333 30328 7364
rect 31938 7352 31944 7404
rect 31996 7352 32002 7404
rect 32125 7395 32183 7401
rect 32125 7361 32137 7395
rect 32171 7392 32183 7395
rect 32214 7392 32220 7404
rect 32171 7364 32220 7392
rect 32171 7361 32183 7364
rect 32125 7355 32183 7361
rect 32214 7352 32220 7364
rect 32272 7352 32278 7404
rect 32674 7352 32680 7404
rect 32732 7392 32738 7404
rect 33965 7395 34023 7401
rect 33965 7392 33977 7395
rect 32732 7364 33977 7392
rect 32732 7352 32738 7364
rect 33965 7361 33977 7364
rect 34011 7361 34023 7395
rect 33965 7355 34023 7361
rect 30193 7327 30251 7333
rect 30193 7324 30205 7327
rect 29880 7296 30205 7324
rect 29880 7284 29886 7296
rect 30193 7293 30205 7296
rect 30239 7293 30251 7327
rect 30193 7287 30251 7293
rect 30285 7327 30343 7333
rect 30285 7293 30297 7327
rect 30331 7293 30343 7327
rect 30285 7287 30343 7293
rect 30466 7256 30472 7268
rect 28675 7228 30472 7256
rect 28675 7225 28687 7228
rect 28629 7219 28687 7225
rect 30466 7216 30472 7228
rect 30524 7216 30530 7268
rect 33980 7256 34008 7355
rect 34422 7352 34428 7404
rect 34480 7352 34486 7404
rect 34514 7352 34520 7404
rect 34572 7392 34578 7404
rect 34681 7395 34739 7401
rect 34681 7392 34693 7395
rect 34572 7364 34693 7392
rect 34572 7352 34578 7364
rect 34681 7361 34693 7364
rect 34727 7361 34739 7395
rect 34681 7355 34739 7361
rect 34054 7284 34060 7336
rect 34112 7284 34118 7336
rect 34238 7284 34244 7336
rect 34296 7284 34302 7336
rect 36538 7284 36544 7336
rect 36596 7284 36602 7336
rect 33980 7228 34468 7256
rect 19260 7160 23612 7188
rect 26973 7191 27031 7197
rect 19153 7151 19211 7157
rect 26973 7157 26985 7191
rect 27019 7188 27031 7191
rect 27246 7188 27252 7200
rect 27019 7160 27252 7188
rect 27019 7157 27031 7160
rect 26973 7151 27031 7157
rect 27246 7148 27252 7160
rect 27304 7148 27310 7200
rect 29733 7191 29791 7197
rect 29733 7157 29745 7191
rect 29779 7188 29791 7191
rect 30834 7188 30840 7200
rect 29779 7160 30840 7188
rect 29779 7157 29791 7160
rect 29733 7151 29791 7157
rect 30834 7148 30840 7160
rect 30892 7148 30898 7200
rect 31202 7148 31208 7200
rect 31260 7188 31266 7200
rect 33226 7188 33232 7200
rect 31260 7160 33232 7188
rect 31260 7148 31266 7160
rect 33226 7148 33232 7160
rect 33284 7148 33290 7200
rect 33502 7148 33508 7200
rect 33560 7148 33566 7200
rect 33597 7191 33655 7197
rect 33597 7157 33609 7191
rect 33643 7188 33655 7191
rect 34330 7188 34336 7200
rect 33643 7160 34336 7188
rect 33643 7157 33655 7160
rect 33597 7151 33655 7157
rect 34330 7148 34336 7160
rect 34388 7148 34394 7200
rect 34440 7188 34468 7228
rect 35805 7191 35863 7197
rect 35805 7188 35817 7191
rect 34440 7160 35817 7188
rect 35805 7157 35817 7160
rect 35851 7157 35863 7191
rect 35805 7151 35863 7157
rect 1104 7098 47104 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 47104 7098
rect 1104 7024 47104 7046
rect 10226 6944 10232 6996
rect 10284 6984 10290 6996
rect 10413 6987 10471 6993
rect 10413 6984 10425 6987
rect 10284 6956 10425 6984
rect 10284 6944 10290 6956
rect 10413 6953 10425 6956
rect 10459 6953 10471 6987
rect 19426 6984 19432 6996
rect 10413 6947 10471 6953
rect 18892 6956 19432 6984
rect 15120 6888 15332 6916
rect 14458 6808 14464 6860
rect 14516 6848 14522 6860
rect 15120 6848 15148 6888
rect 14516 6820 15148 6848
rect 14516 6808 14522 6820
rect 15194 6808 15200 6860
rect 15252 6808 15258 6860
rect 15304 6848 15332 6888
rect 15562 6848 15568 6860
rect 15620 6857 15626 6860
rect 15620 6851 15648 6857
rect 15304 6820 15568 6848
rect 15562 6808 15568 6820
rect 15636 6817 15648 6851
rect 15620 6811 15648 6817
rect 15620 6808 15626 6811
rect 15746 6808 15752 6860
rect 15804 6808 15810 6860
rect 17865 6851 17923 6857
rect 17865 6817 17877 6851
rect 17911 6848 17923 6851
rect 18892 6848 18920 6956
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 20625 6987 20683 6993
rect 20625 6984 20637 6987
rect 19576 6956 20637 6984
rect 19576 6944 19582 6956
rect 20625 6953 20637 6956
rect 20671 6953 20683 6987
rect 20625 6947 20683 6953
rect 24596 6956 25728 6984
rect 17911 6820 18920 6848
rect 18984 6820 19380 6848
rect 17911 6817 17923 6820
rect 17865 6811 17923 6817
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6780 10655 6783
rect 11514 6780 11520 6792
rect 10643 6752 11520 6780
rect 10643 6749 10655 6752
rect 10597 6743 10655 6749
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 14550 6740 14556 6792
rect 14608 6740 14614 6792
rect 14642 6740 14648 6792
rect 14700 6780 14706 6792
rect 14737 6783 14795 6789
rect 14737 6780 14749 6783
rect 14700 6752 14749 6780
rect 14700 6740 14706 6752
rect 14737 6749 14749 6752
rect 14783 6749 14795 6783
rect 14737 6743 14795 6749
rect 15470 6740 15476 6792
rect 15528 6740 15534 6792
rect 18984 6780 19012 6820
rect 16316 6752 19012 6780
rect 15654 6604 15660 6656
rect 15712 6644 15718 6656
rect 16316 6644 16344 6752
rect 19058 6740 19064 6792
rect 19116 6740 19122 6792
rect 19150 6740 19156 6792
rect 19208 6780 19214 6792
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 19208 6752 19257 6780
rect 19208 6740 19214 6752
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 19352 6780 19380 6820
rect 24596 6780 24624 6956
rect 24670 6808 24676 6860
rect 24728 6808 24734 6860
rect 25700 6848 25728 6956
rect 27172 6956 28120 6984
rect 27172 6848 27200 6956
rect 28092 6916 28120 6956
rect 28534 6944 28540 6996
rect 28592 6944 28598 6996
rect 31938 6944 31944 6996
rect 31996 6984 32002 6996
rect 32033 6987 32091 6993
rect 32033 6984 32045 6987
rect 31996 6956 32045 6984
rect 31996 6944 32002 6956
rect 32033 6953 32045 6956
rect 32079 6953 32091 6987
rect 32033 6947 32091 6953
rect 33042 6944 33048 6996
rect 33100 6984 33106 6996
rect 34606 6984 34612 6996
rect 33100 6956 34612 6984
rect 33100 6944 33106 6956
rect 34606 6944 34612 6956
rect 34664 6944 34670 6996
rect 28092 6888 28212 6916
rect 25700 6820 27200 6848
rect 19352 6752 24624 6780
rect 24688 6780 24716 6808
rect 27062 6780 27068 6792
rect 24688 6752 27068 6780
rect 19245 6743 19303 6749
rect 27062 6740 27068 6752
rect 27120 6780 27126 6792
rect 27157 6783 27215 6789
rect 27157 6780 27169 6783
rect 27120 6752 27169 6780
rect 27120 6740 27126 6752
rect 27157 6749 27169 6752
rect 27203 6749 27215 6783
rect 27157 6743 27215 6749
rect 27246 6740 27252 6792
rect 27304 6780 27310 6792
rect 27413 6783 27471 6789
rect 27413 6780 27425 6783
rect 27304 6752 27425 6780
rect 27304 6740 27310 6752
rect 27413 6749 27425 6752
rect 27459 6749 27471 6783
rect 27413 6743 27471 6749
rect 16393 6715 16451 6721
rect 16393 6681 16405 6715
rect 16439 6712 16451 6715
rect 18966 6712 18972 6724
rect 16439 6684 18972 6712
rect 16439 6681 16451 6684
rect 16393 6675 16451 6681
rect 18966 6672 18972 6684
rect 19024 6672 19030 6724
rect 19490 6715 19548 6721
rect 19490 6712 19502 6715
rect 19076 6684 19502 6712
rect 15712 6616 16344 6644
rect 15712 6604 15718 6616
rect 17310 6604 17316 6656
rect 17368 6604 17374 6656
rect 17678 6604 17684 6656
rect 17736 6604 17742 6656
rect 17773 6647 17831 6653
rect 17773 6613 17785 6647
rect 17819 6644 17831 6647
rect 17862 6644 17868 6656
rect 17819 6616 17868 6644
rect 17819 6613 17831 6616
rect 17773 6607 17831 6613
rect 17862 6604 17868 6616
rect 17920 6604 17926 6656
rect 18877 6647 18935 6653
rect 18877 6613 18889 6647
rect 18923 6644 18935 6647
rect 19076 6644 19104 6684
rect 19490 6681 19502 6684
rect 19536 6681 19548 6715
rect 19490 6675 19548 6681
rect 24940 6715 24998 6721
rect 24940 6681 24952 6715
rect 24986 6712 24998 6715
rect 26510 6712 26516 6724
rect 24986 6684 26516 6712
rect 24986 6681 24998 6684
rect 24940 6675 24998 6681
rect 26510 6672 26516 6684
rect 26568 6672 26574 6724
rect 28184 6712 28212 6888
rect 29822 6876 29828 6928
rect 29880 6916 29886 6928
rect 33134 6916 33140 6928
rect 29880 6888 33140 6916
rect 29880 6876 29886 6888
rect 29730 6808 29736 6860
rect 29788 6808 29794 6860
rect 32508 6857 32536 6888
rect 33134 6876 33140 6888
rect 33192 6916 33198 6928
rect 33965 6919 34023 6925
rect 33965 6916 33977 6919
rect 33192 6888 33977 6916
rect 33192 6876 33198 6888
rect 33965 6885 33977 6888
rect 34011 6916 34023 6919
rect 34054 6916 34060 6928
rect 34011 6888 34060 6916
rect 34011 6885 34023 6888
rect 33965 6879 34023 6885
rect 34054 6876 34060 6888
rect 34112 6876 34118 6928
rect 37458 6916 37464 6928
rect 34256 6888 37464 6916
rect 32493 6851 32551 6857
rect 32493 6817 32505 6851
rect 32539 6817 32551 6851
rect 32493 6811 32551 6817
rect 32582 6808 32588 6860
rect 32640 6808 32646 6860
rect 33226 6808 33232 6860
rect 33284 6848 33290 6860
rect 33284 6820 33824 6848
rect 33284 6808 33290 6820
rect 28902 6740 28908 6792
rect 28960 6780 28966 6792
rect 30009 6783 30067 6789
rect 30009 6780 30021 6783
rect 28960 6752 30021 6780
rect 28960 6740 28966 6752
rect 30009 6749 30021 6752
rect 30055 6749 30067 6783
rect 30009 6743 30067 6749
rect 30834 6740 30840 6792
rect 30892 6740 30898 6792
rect 32401 6783 32459 6789
rect 32401 6749 32413 6783
rect 32447 6780 32459 6783
rect 33502 6780 33508 6792
rect 32447 6752 33508 6780
rect 32447 6749 32459 6752
rect 32401 6743 32459 6749
rect 33502 6740 33508 6752
rect 33560 6740 33566 6792
rect 33796 6789 33824 6820
rect 33781 6783 33839 6789
rect 33781 6749 33793 6783
rect 33827 6780 33839 6783
rect 34256 6780 34284 6888
rect 37458 6876 37464 6888
rect 37516 6876 37522 6928
rect 33827 6752 34284 6780
rect 33827 6749 33839 6752
rect 33781 6743 33839 6749
rect 34330 6740 34336 6792
rect 34388 6740 34394 6792
rect 30742 6712 30748 6724
rect 28184 6684 30748 6712
rect 30742 6672 30748 6684
rect 30800 6672 30806 6724
rect 18923 6616 19104 6644
rect 18923 6613 18935 6616
rect 18877 6607 18935 6613
rect 19150 6604 19156 6656
rect 19208 6644 19214 6656
rect 19886 6644 19892 6656
rect 19208 6616 19892 6644
rect 19208 6604 19214 6616
rect 19886 6604 19892 6616
rect 19944 6604 19950 6656
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 26053 6647 26111 6653
rect 26053 6644 26065 6647
rect 24912 6616 26065 6644
rect 24912 6604 24918 6616
rect 26053 6613 26065 6616
rect 26099 6644 26111 6647
rect 26142 6644 26148 6656
rect 26099 6616 26148 6644
rect 26099 6613 26111 6616
rect 26053 6607 26111 6613
rect 26142 6604 26148 6616
rect 26200 6604 26206 6656
rect 26418 6604 26424 6656
rect 26476 6644 26482 6656
rect 30282 6644 30288 6656
rect 26476 6616 30288 6644
rect 26476 6604 26482 6616
rect 30282 6604 30288 6616
rect 30340 6604 30346 6656
rect 30650 6604 30656 6656
rect 30708 6604 30714 6656
rect 34149 6647 34207 6653
rect 34149 6613 34161 6647
rect 34195 6644 34207 6647
rect 34514 6644 34520 6656
rect 34195 6616 34520 6644
rect 34195 6613 34207 6616
rect 34149 6607 34207 6613
rect 34514 6604 34520 6616
rect 34572 6604 34578 6656
rect 1104 6554 47104 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 47104 6554
rect 1104 6480 47104 6502
rect 17678 6400 17684 6452
rect 17736 6440 17742 6452
rect 18141 6443 18199 6449
rect 18141 6440 18153 6443
rect 17736 6412 18153 6440
rect 17736 6400 17742 6412
rect 18141 6409 18153 6412
rect 18187 6409 18199 6443
rect 18141 6403 18199 6409
rect 18616 6412 23612 6440
rect 18616 6372 18644 6412
rect 19214 6375 19272 6381
rect 19214 6372 19226 6375
rect 16224 6344 18644 6372
rect 18708 6344 19226 6372
rect 13170 6264 13176 6316
rect 13228 6264 13234 6316
rect 13998 6264 14004 6316
rect 14056 6304 14062 6316
rect 15562 6313 15568 6316
rect 15519 6307 15568 6313
rect 14056 6276 14780 6304
rect 14056 6264 14062 6276
rect 14093 6239 14151 6245
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 14182 6236 14188 6248
rect 14139 6208 14188 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 14182 6196 14188 6208
rect 14240 6196 14246 6248
rect 14277 6239 14335 6245
rect 14277 6205 14289 6239
rect 14323 6236 14335 6239
rect 14461 6239 14519 6245
rect 14323 6208 14412 6236
rect 14323 6205 14335 6208
rect 14277 6199 14335 6205
rect 12986 6060 12992 6112
rect 13044 6060 13050 6112
rect 13633 6103 13691 6109
rect 13633 6069 13645 6103
rect 13679 6100 13691 6103
rect 14090 6100 14096 6112
rect 13679 6072 14096 6100
rect 13679 6069 13691 6072
rect 13633 6063 13691 6069
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 14384 6100 14412 6208
rect 14461 6205 14473 6239
rect 14507 6205 14519 6239
rect 14461 6199 14519 6205
rect 14476 6168 14504 6199
rect 14642 6196 14648 6248
rect 14700 6196 14706 6248
rect 14752 6236 14780 6276
rect 15519 6273 15531 6307
rect 15565 6273 15568 6307
rect 15519 6267 15568 6273
rect 15562 6264 15568 6267
rect 15620 6264 15626 6316
rect 15654 6264 15660 6316
rect 15712 6264 15718 6316
rect 15378 6236 15384 6248
rect 14752 6208 15384 6236
rect 15378 6196 15384 6208
rect 15436 6196 15442 6248
rect 14550 6168 14556 6180
rect 14476 6140 14556 6168
rect 14550 6128 14556 6140
rect 14608 6168 14614 6180
rect 15010 6168 15016 6180
rect 14608 6140 15016 6168
rect 14608 6128 14614 6140
rect 15010 6128 15016 6140
rect 15068 6128 15074 6180
rect 15105 6171 15163 6177
rect 15105 6137 15117 6171
rect 15151 6137 15163 6171
rect 15105 6131 15163 6137
rect 14918 6100 14924 6112
rect 14384 6072 14924 6100
rect 14918 6060 14924 6072
rect 14976 6060 14982 6112
rect 15120 6100 15148 6131
rect 16224 6100 16252 6344
rect 16758 6264 16764 6316
rect 16816 6264 16822 6316
rect 17034 6313 17040 6316
rect 17028 6267 17040 6313
rect 17034 6264 17040 6267
rect 17092 6264 17098 6316
rect 18708 6177 18736 6344
rect 19214 6341 19226 6344
rect 19260 6341 19272 6375
rect 19214 6335 19272 6341
rect 20346 6332 20352 6384
rect 20404 6372 20410 6384
rect 23584 6372 23612 6412
rect 23658 6400 23664 6452
rect 23716 6400 23722 6452
rect 24228 6412 25544 6440
rect 24228 6372 24256 6412
rect 25516 6372 25544 6412
rect 25590 6400 25596 6452
rect 25648 6400 25654 6452
rect 26418 6440 26424 6452
rect 25792 6412 26424 6440
rect 25792 6372 25820 6412
rect 26418 6400 26424 6412
rect 26476 6400 26482 6452
rect 26510 6400 26516 6452
rect 26568 6400 26574 6452
rect 27062 6400 27068 6452
rect 27120 6440 27126 6452
rect 27120 6412 27476 6440
rect 27120 6400 27126 6412
rect 27338 6372 27344 6384
rect 20404 6344 21036 6372
rect 23584 6344 24256 6372
rect 24320 6344 25360 6372
rect 25516 6344 25820 6372
rect 25884 6344 27344 6372
rect 20404 6332 20410 6344
rect 18877 6307 18935 6313
rect 18877 6273 18889 6307
rect 18923 6304 18935 6307
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 18923 6276 20484 6304
rect 18923 6273 18935 6276
rect 18877 6267 18935 6273
rect 18969 6239 19027 6245
rect 18969 6205 18981 6239
rect 19015 6205 19027 6239
rect 18969 6199 19027 6205
rect 18693 6171 18751 6177
rect 18693 6137 18705 6171
rect 18739 6137 18751 6171
rect 18693 6131 18751 6137
rect 15120 6072 16252 6100
rect 16301 6103 16359 6109
rect 16301 6069 16313 6103
rect 16347 6100 16359 6103
rect 17402 6100 17408 6112
rect 16347 6072 17408 6100
rect 16347 6069 16359 6072
rect 16301 6063 16359 6069
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 18984 6100 19012 6199
rect 20456 6177 20484 6276
rect 20548 6276 20821 6304
rect 20441 6171 20499 6177
rect 20441 6137 20453 6171
rect 20487 6137 20499 6171
rect 20441 6131 20499 6137
rect 19242 6100 19248 6112
rect 18984 6072 19248 6100
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 20349 6103 20407 6109
rect 20349 6100 20361 6103
rect 19392 6072 20361 6100
rect 19392 6060 19398 6072
rect 20349 6069 20361 6072
rect 20395 6100 20407 6103
rect 20548 6100 20576 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 21008 6245 21036 6344
rect 21821 6307 21879 6313
rect 21821 6273 21833 6307
rect 21867 6304 21879 6307
rect 22186 6304 22192 6316
rect 21867 6276 22192 6304
rect 21867 6273 21879 6276
rect 21821 6267 21879 6273
rect 22186 6264 22192 6276
rect 22244 6264 22250 6316
rect 24210 6264 24216 6316
rect 24268 6264 24274 6316
rect 20901 6239 20959 6245
rect 20901 6205 20913 6239
rect 20947 6205 20959 6239
rect 20901 6199 20959 6205
rect 20993 6239 21051 6245
rect 20993 6205 21005 6239
rect 21039 6205 21051 6239
rect 20993 6199 21051 6205
rect 22005 6239 22063 6245
rect 22005 6205 22017 6239
rect 22051 6236 22063 6239
rect 22094 6236 22100 6248
rect 22051 6208 22100 6236
rect 22051 6205 22063 6208
rect 22005 6199 22063 6205
rect 20395 6072 20576 6100
rect 20916 6100 20944 6199
rect 22094 6196 22100 6208
rect 22152 6196 22158 6248
rect 22462 6196 22468 6248
rect 22520 6196 22526 6248
rect 22554 6196 22560 6248
rect 22612 6236 22618 6248
rect 22741 6239 22799 6245
rect 22741 6236 22753 6239
rect 22612 6208 22753 6236
rect 22612 6196 22618 6208
rect 22741 6205 22753 6208
rect 22787 6205 22799 6239
rect 22741 6199 22799 6205
rect 22830 6196 22836 6248
rect 22888 6245 22894 6248
rect 22888 6239 22916 6245
rect 22904 6205 22916 6239
rect 22888 6199 22916 6205
rect 23017 6239 23075 6245
rect 23017 6205 23029 6239
rect 23063 6236 23075 6239
rect 24320 6236 24348 6344
rect 24486 6313 24492 6316
rect 24480 6267 24492 6313
rect 24486 6264 24492 6267
rect 24544 6264 24550 6316
rect 25332 6304 25360 6344
rect 25884 6304 25912 6344
rect 27338 6332 27344 6344
rect 27396 6332 27402 6384
rect 25332 6276 25912 6304
rect 25958 6264 25964 6316
rect 26016 6304 26022 6316
rect 26053 6307 26111 6313
rect 26053 6304 26065 6307
rect 26016 6276 26065 6304
rect 26016 6264 26022 6276
rect 26053 6273 26065 6276
rect 26099 6273 26111 6307
rect 26053 6267 26111 6273
rect 26142 6264 26148 6316
rect 26200 6264 26206 6316
rect 26694 6264 26700 6316
rect 26752 6264 26758 6316
rect 27448 6304 27476 6412
rect 30190 6400 30196 6452
rect 30248 6440 30254 6452
rect 31205 6443 31263 6449
rect 31205 6440 31217 6443
rect 30248 6412 31217 6440
rect 30248 6400 30254 6412
rect 31205 6409 31217 6412
rect 31251 6409 31263 6443
rect 31205 6403 31263 6409
rect 30092 6375 30150 6381
rect 30092 6341 30104 6375
rect 30138 6372 30150 6375
rect 30650 6372 30656 6384
rect 30138 6344 30656 6372
rect 30138 6341 30150 6344
rect 30092 6335 30150 6341
rect 30650 6332 30656 6344
rect 30708 6332 30714 6384
rect 32122 6372 32128 6384
rect 30760 6344 32128 6372
rect 28902 6304 28908 6316
rect 27448 6276 28908 6304
rect 28902 6264 28908 6276
rect 28960 6264 28966 6316
rect 29825 6307 29883 6313
rect 29825 6273 29837 6307
rect 29871 6304 29883 6307
rect 30760 6304 30788 6344
rect 32122 6332 32128 6344
rect 32180 6372 32186 6384
rect 33042 6372 33048 6384
rect 32180 6344 33048 6372
rect 32180 6332 32186 6344
rect 33042 6332 33048 6344
rect 33100 6332 33106 6384
rect 29871 6276 30788 6304
rect 29871 6273 29883 6276
rect 29825 6267 29883 6273
rect 31478 6264 31484 6316
rect 31536 6264 31542 6316
rect 23063 6208 24348 6236
rect 26329 6239 26387 6245
rect 23063 6205 23075 6208
rect 23017 6199 23075 6205
rect 26329 6205 26341 6239
rect 26375 6236 26387 6239
rect 28994 6236 29000 6248
rect 26375 6208 29000 6236
rect 26375 6205 26387 6208
rect 26329 6199 26387 6205
rect 22888 6196 22894 6199
rect 28994 6196 29000 6208
rect 29052 6196 29058 6248
rect 29178 6196 29184 6248
rect 29236 6196 29242 6248
rect 25685 6171 25743 6177
rect 25685 6137 25697 6171
rect 25731 6168 25743 6171
rect 26694 6168 26700 6180
rect 25731 6140 26700 6168
rect 25731 6137 25743 6140
rect 25685 6131 25743 6137
rect 26694 6128 26700 6140
rect 26752 6128 26758 6180
rect 29822 6168 29828 6180
rect 27264 6140 29828 6168
rect 27264 6100 27292 6140
rect 29822 6128 29828 6140
rect 29880 6128 29886 6180
rect 33870 6168 33876 6180
rect 31220 6140 33876 6168
rect 20916 6072 27292 6100
rect 20395 6069 20407 6072
rect 20349 6063 20407 6069
rect 27338 6060 27344 6112
rect 27396 6100 27402 6112
rect 31220 6100 31248 6140
rect 33870 6128 33876 6140
rect 33928 6128 33934 6180
rect 27396 6072 31248 6100
rect 27396 6060 27402 6072
rect 31294 6060 31300 6112
rect 31352 6060 31358 6112
rect 1104 6010 47104 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 47104 6010
rect 1104 5936 47104 5958
rect 13170 5856 13176 5908
rect 13228 5896 13234 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 13228 5868 14105 5896
rect 13228 5856 13234 5868
rect 14093 5865 14105 5868
rect 14139 5865 14151 5899
rect 14093 5859 14151 5865
rect 14642 5856 14648 5908
rect 14700 5896 14706 5908
rect 15470 5896 15476 5908
rect 14700 5868 15476 5896
rect 14700 5856 14706 5868
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 17034 5856 17040 5908
rect 17092 5896 17098 5908
rect 17129 5899 17187 5905
rect 17129 5896 17141 5899
rect 17092 5868 17141 5896
rect 17092 5856 17098 5868
rect 17129 5865 17141 5868
rect 17175 5865 17187 5899
rect 17129 5859 17187 5865
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 19702 5896 19708 5908
rect 17460 5868 19708 5896
rect 17460 5856 17466 5868
rect 19702 5856 19708 5868
rect 19760 5856 19766 5908
rect 23014 5896 23020 5908
rect 22388 5868 23020 5896
rect 13909 5831 13967 5837
rect 13909 5797 13921 5831
rect 13955 5828 13967 5831
rect 13998 5828 14004 5840
rect 13955 5800 14004 5828
rect 13955 5797 13967 5800
rect 13909 5791 13967 5797
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 14182 5788 14188 5840
rect 14240 5828 14246 5840
rect 15010 5828 15016 5840
rect 14240 5800 15016 5828
rect 14240 5788 14246 5800
rect 14568 5769 14596 5800
rect 15010 5788 15016 5800
rect 15068 5828 15074 5840
rect 17862 5828 17868 5840
rect 15068 5800 17868 5828
rect 15068 5788 15074 5800
rect 17862 5788 17868 5800
rect 17920 5828 17926 5840
rect 21726 5828 21732 5840
rect 17920 5800 21732 5828
rect 17920 5788 17926 5800
rect 21726 5788 21732 5800
rect 21784 5788 21790 5840
rect 22094 5828 22100 5840
rect 22066 5788 22100 5828
rect 22152 5788 22158 5840
rect 22388 5828 22416 5868
rect 23014 5856 23020 5868
rect 23072 5856 23078 5908
rect 23382 5856 23388 5908
rect 23440 5896 23446 5908
rect 23477 5899 23535 5905
rect 23477 5896 23489 5899
rect 23440 5868 23489 5896
rect 23440 5856 23446 5868
rect 23477 5865 23489 5868
rect 23523 5865 23535 5899
rect 23477 5859 23535 5865
rect 24486 5856 24492 5908
rect 24544 5856 24550 5908
rect 24854 5856 24860 5908
rect 24912 5896 24918 5908
rect 26234 5896 26240 5908
rect 24912 5868 26240 5896
rect 24912 5856 24918 5868
rect 26234 5856 26240 5868
rect 26292 5896 26298 5908
rect 27522 5896 27528 5908
rect 26292 5868 27528 5896
rect 26292 5856 26298 5868
rect 27522 5856 27528 5868
rect 27580 5856 27586 5908
rect 29638 5856 29644 5908
rect 29696 5896 29702 5908
rect 31021 5899 31079 5905
rect 31021 5896 31033 5899
rect 29696 5868 31033 5896
rect 29696 5856 29702 5868
rect 31021 5865 31033 5868
rect 31067 5865 31079 5899
rect 31021 5859 31079 5865
rect 22296 5800 22416 5828
rect 14553 5763 14611 5769
rect 14553 5729 14565 5763
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 14734 5720 14740 5772
rect 14792 5720 14798 5772
rect 18874 5720 18880 5772
rect 18932 5760 18938 5772
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 18932 5732 19257 5760
rect 18932 5720 18938 5732
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 19521 5763 19579 5769
rect 19521 5760 19533 5763
rect 19392 5732 19533 5760
rect 19392 5720 19398 5732
rect 19521 5729 19533 5732
rect 19567 5729 19579 5763
rect 19521 5723 19579 5729
rect 21821 5763 21879 5769
rect 21821 5729 21833 5763
rect 21867 5760 21879 5763
rect 22066 5760 22094 5788
rect 22296 5769 22324 5800
rect 24946 5788 24952 5840
rect 25004 5828 25010 5840
rect 25685 5831 25743 5837
rect 25685 5828 25697 5831
rect 25004 5800 25697 5828
rect 25004 5788 25010 5800
rect 25685 5797 25697 5800
rect 25731 5797 25743 5831
rect 25685 5791 25743 5797
rect 25774 5788 25780 5840
rect 25832 5828 25838 5840
rect 25832 5800 26280 5828
rect 25832 5788 25838 5800
rect 21867 5732 22094 5760
rect 22281 5763 22339 5769
rect 21867 5729 21879 5732
rect 21821 5723 21879 5729
rect 22281 5729 22293 5763
rect 22327 5729 22339 5763
rect 22281 5723 22339 5729
rect 22646 5720 22652 5772
rect 22704 5769 22710 5772
rect 22704 5763 22732 5769
rect 22720 5729 22732 5763
rect 22704 5723 22732 5729
rect 22833 5763 22891 5769
rect 22833 5729 22845 5763
rect 22879 5760 22891 5763
rect 23474 5760 23480 5772
rect 22879 5732 23480 5760
rect 22879 5729 22891 5732
rect 22833 5723 22891 5729
rect 22704 5720 22710 5723
rect 23474 5720 23480 5732
rect 23532 5720 23538 5772
rect 26252 5769 26280 5800
rect 26237 5763 26295 5769
rect 26237 5729 26249 5763
rect 26283 5729 26295 5763
rect 26237 5723 26295 5729
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 12529 5695 12587 5701
rect 12529 5692 12541 5695
rect 12492 5664 12541 5692
rect 12492 5652 12498 5664
rect 12529 5661 12541 5664
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 17310 5652 17316 5704
rect 17368 5652 17374 5704
rect 21637 5695 21695 5701
rect 21637 5661 21649 5695
rect 21683 5661 21695 5695
rect 21637 5655 21695 5661
rect 12796 5627 12854 5633
rect 12796 5593 12808 5627
rect 12842 5624 12854 5627
rect 13906 5624 13912 5636
rect 12842 5596 13912 5624
rect 12842 5593 12854 5596
rect 12796 5587 12854 5593
rect 13906 5584 13912 5596
rect 13964 5584 13970 5636
rect 14458 5516 14464 5568
rect 14516 5516 14522 5568
rect 21652 5556 21680 5655
rect 22554 5652 22560 5704
rect 22612 5652 22618 5704
rect 24673 5695 24731 5701
rect 24673 5661 24685 5695
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 22186 5556 22192 5568
rect 21652 5528 22192 5556
rect 22186 5516 22192 5528
rect 22244 5556 22250 5568
rect 22646 5556 22652 5568
rect 22244 5528 22652 5556
rect 22244 5516 22250 5528
rect 22646 5516 22652 5528
rect 22704 5516 22710 5568
rect 24688 5556 24716 5655
rect 25130 5652 25136 5704
rect 25188 5692 25194 5704
rect 26252 5692 26280 5723
rect 28626 5720 28632 5772
rect 28684 5760 28690 5772
rect 29178 5760 29184 5772
rect 28684 5732 29184 5760
rect 28684 5720 28690 5732
rect 29178 5720 29184 5732
rect 29236 5760 29242 5772
rect 29641 5763 29699 5769
rect 29641 5760 29653 5763
rect 29236 5732 29653 5760
rect 29236 5720 29242 5732
rect 29641 5729 29653 5732
rect 29687 5729 29699 5763
rect 29641 5723 29699 5729
rect 29546 5692 29552 5704
rect 25188 5664 26188 5692
rect 26252 5664 29552 5692
rect 25188 5652 25194 5664
rect 24854 5584 24860 5636
rect 24912 5584 24918 5636
rect 25038 5584 25044 5636
rect 25096 5584 25102 5636
rect 25590 5584 25596 5636
rect 25648 5624 25654 5636
rect 26053 5627 26111 5633
rect 26053 5624 26065 5627
rect 25648 5596 26065 5624
rect 25648 5584 25654 5596
rect 26053 5593 26065 5596
rect 26099 5593 26111 5627
rect 26160 5624 26188 5664
rect 29546 5652 29552 5664
rect 29604 5692 29610 5704
rect 29730 5692 29736 5704
rect 29604 5664 29736 5692
rect 29604 5652 29610 5664
rect 29730 5652 29736 5664
rect 29788 5652 29794 5704
rect 29908 5695 29966 5701
rect 29908 5661 29920 5695
rect 29954 5692 29966 5695
rect 31294 5692 31300 5704
rect 29954 5664 31300 5692
rect 29954 5661 29966 5664
rect 29908 5655 29966 5661
rect 31294 5652 31300 5664
rect 31352 5652 31358 5704
rect 35253 5695 35311 5701
rect 35253 5661 35265 5695
rect 35299 5692 35311 5695
rect 35342 5692 35348 5704
rect 35299 5664 35348 5692
rect 35299 5661 35311 5664
rect 35253 5655 35311 5661
rect 35342 5652 35348 5664
rect 35400 5652 35406 5704
rect 44358 5652 44364 5704
rect 44416 5692 44422 5704
rect 46385 5695 46443 5701
rect 46385 5692 46397 5695
rect 44416 5664 46397 5692
rect 44416 5652 44422 5664
rect 46385 5661 46397 5664
rect 46431 5661 46443 5695
rect 46385 5655 46443 5661
rect 31018 5624 31024 5636
rect 26160 5596 31024 5624
rect 26053 5587 26111 5593
rect 31018 5584 31024 5596
rect 31076 5584 31082 5636
rect 24946 5556 24952 5568
rect 24688 5528 24952 5556
rect 24946 5516 24952 5528
rect 25004 5516 25010 5568
rect 25056 5556 25084 5584
rect 25958 5556 25964 5568
rect 25056 5528 25964 5556
rect 25958 5516 25964 5528
rect 26016 5556 26022 5568
rect 26145 5559 26203 5565
rect 26145 5556 26157 5559
rect 26016 5528 26157 5556
rect 26016 5516 26022 5528
rect 26145 5525 26157 5528
rect 26191 5525 26203 5559
rect 26145 5519 26203 5525
rect 35066 5516 35072 5568
rect 35124 5516 35130 5568
rect 46658 5516 46664 5568
rect 46716 5516 46722 5568
rect 1104 5466 47104 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 47104 5466
rect 1104 5392 47104 5414
rect 16850 5352 16856 5364
rect 1412 5324 13768 5352
rect 1412 5225 1440 5324
rect 6086 5244 6092 5296
rect 6144 5284 6150 5296
rect 11885 5287 11943 5293
rect 11885 5284 11897 5287
rect 6144 5256 11897 5284
rect 6144 5244 6150 5256
rect 11885 5253 11897 5256
rect 11931 5253 11943 5287
rect 11885 5247 11943 5253
rect 12704 5287 12762 5293
rect 12704 5253 12716 5287
rect 12750 5284 12762 5287
rect 12986 5284 12992 5296
rect 12750 5256 12992 5284
rect 12750 5253 12762 5256
rect 12704 5247 12762 5253
rect 12986 5244 12992 5256
rect 13044 5244 13050 5296
rect 13740 5284 13768 5324
rect 13924 5324 16856 5352
rect 13924 5284 13952 5324
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 17494 5312 17500 5364
rect 17552 5352 17558 5364
rect 17862 5352 17868 5364
rect 17552 5324 17868 5352
rect 17552 5312 17558 5324
rect 17862 5312 17868 5324
rect 17920 5352 17926 5364
rect 18049 5355 18107 5361
rect 18049 5352 18061 5355
rect 17920 5324 18061 5352
rect 17920 5312 17926 5324
rect 18049 5321 18061 5324
rect 18095 5321 18107 5355
rect 18049 5315 18107 5321
rect 21453 5355 21511 5361
rect 21453 5321 21465 5355
rect 21499 5321 21511 5355
rect 21453 5315 21511 5321
rect 18782 5284 18788 5296
rect 13740 5256 13952 5284
rect 14016 5256 18788 5284
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 9858 5176 9864 5228
rect 9916 5216 9922 5228
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 9916 5188 9965 5216
rect 9916 5176 9922 5188
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 10220 5219 10278 5225
rect 10220 5185 10232 5219
rect 10266 5216 10278 5219
rect 10686 5216 10692 5228
rect 10266 5188 10692 5216
rect 10266 5185 10278 5188
rect 10220 5179 10278 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 14016 5216 14044 5256
rect 18782 5244 18788 5256
rect 18840 5244 18846 5296
rect 21468 5284 21496 5315
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 22830 5352 22836 5364
rect 22152 5324 22836 5352
rect 22152 5312 22158 5324
rect 22830 5312 22836 5324
rect 22888 5352 22894 5364
rect 23385 5355 23443 5361
rect 23385 5352 23397 5355
rect 22888 5324 23397 5352
rect 22888 5312 22894 5324
rect 23385 5321 23397 5324
rect 23431 5321 23443 5355
rect 23385 5315 23443 5321
rect 23474 5312 23480 5364
rect 23532 5352 23538 5364
rect 24762 5352 24768 5364
rect 23532 5324 24768 5352
rect 23532 5312 23538 5324
rect 24762 5312 24768 5324
rect 24820 5352 24826 5364
rect 26142 5352 26148 5364
rect 24820 5324 26148 5352
rect 24820 5312 24826 5324
rect 26142 5312 26148 5324
rect 26200 5312 26206 5364
rect 26786 5312 26792 5364
rect 26844 5312 26850 5364
rect 27522 5312 27528 5364
rect 27580 5352 27586 5364
rect 27801 5355 27859 5361
rect 27801 5352 27813 5355
rect 27580 5324 27813 5352
rect 27580 5312 27586 5324
rect 27801 5321 27813 5324
rect 27847 5321 27859 5355
rect 27801 5315 27859 5321
rect 29641 5355 29699 5361
rect 29641 5321 29653 5355
rect 29687 5352 29699 5355
rect 31478 5352 31484 5364
rect 29687 5324 31484 5352
rect 29687 5321 29699 5324
rect 29641 5315 29699 5321
rect 31478 5312 31484 5324
rect 31536 5312 31542 5364
rect 33318 5312 33324 5364
rect 33376 5352 33382 5364
rect 33965 5355 34023 5361
rect 33965 5352 33977 5355
rect 33376 5324 33977 5352
rect 33376 5312 33382 5324
rect 33965 5321 33977 5324
rect 34011 5321 34023 5355
rect 33965 5315 34023 5321
rect 22250 5287 22308 5293
rect 22250 5284 22262 5287
rect 21468 5256 22262 5284
rect 22250 5253 22262 5256
rect 22296 5253 22308 5287
rect 22250 5247 22308 5253
rect 29822 5244 29828 5296
rect 29880 5284 29886 5296
rect 35066 5293 35072 5296
rect 30009 5287 30067 5293
rect 30009 5284 30021 5287
rect 29880 5256 30021 5284
rect 29880 5244 29886 5256
rect 30009 5253 30021 5256
rect 30055 5253 30067 5287
rect 35060 5284 35072 5293
rect 35027 5256 35072 5284
rect 30009 5247 30067 5253
rect 35060 5247 35072 5256
rect 35066 5244 35072 5247
rect 35124 5244 35130 5296
rect 12176 5188 14044 5216
rect 12176 5157 12204 5188
rect 14090 5176 14096 5228
rect 14148 5176 14154 5228
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 16758 5216 16764 5228
rect 16715 5188 16764 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 16936 5219 16994 5225
rect 16936 5185 16948 5219
rect 16982 5216 16994 5219
rect 17218 5216 17224 5228
rect 16982 5188 17224 5216
rect 16982 5185 16994 5188
rect 16936 5179 16994 5185
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 18690 5176 18696 5228
rect 18748 5216 18754 5228
rect 19153 5219 19211 5225
rect 19153 5216 19165 5219
rect 18748 5188 19165 5216
rect 18748 5176 18754 5188
rect 19153 5185 19165 5188
rect 19199 5185 19211 5219
rect 19153 5179 19211 5185
rect 21634 5176 21640 5228
rect 21692 5176 21698 5228
rect 26142 5176 26148 5228
rect 26200 5176 26206 5228
rect 27709 5219 27767 5225
rect 27709 5185 27721 5219
rect 27755 5216 27767 5219
rect 28902 5216 28908 5228
rect 27755 5188 28908 5216
rect 27755 5185 27767 5188
rect 27709 5179 27767 5185
rect 11977 5151 12035 5157
rect 11977 5148 11989 5151
rect 11348 5120 11989 5148
rect 11348 5024 11376 5120
rect 11977 5117 11989 5120
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 12161 5151 12219 5157
rect 12161 5117 12173 5151
rect 12207 5117 12219 5151
rect 12161 5111 12219 5117
rect 12434 5108 12440 5160
rect 12492 5108 12498 5160
rect 21818 5108 21824 5160
rect 21876 5148 21882 5160
rect 22005 5151 22063 5157
rect 22005 5148 22017 5151
rect 21876 5120 22017 5148
rect 21876 5108 21882 5120
rect 22005 5117 22017 5120
rect 22051 5117 22063 5151
rect 22005 5111 22063 5117
rect 24946 5108 24952 5160
rect 25004 5108 25010 5160
rect 25133 5151 25191 5157
rect 25133 5117 25145 5151
rect 25179 5148 25191 5151
rect 25179 5120 25728 5148
rect 25179 5117 25191 5120
rect 25133 5111 25191 5117
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1581 5015 1639 5021
rect 1581 5012 1593 5015
rect 992 4984 1593 5012
rect 992 4972 998 4984
rect 1581 4981 1593 4984
rect 1627 4981 1639 5015
rect 1581 4975 1639 4981
rect 11330 4972 11336 5024
rect 11388 4972 11394 5024
rect 11514 4972 11520 5024
rect 11572 4972 11578 5024
rect 12452 5012 12480 5108
rect 13817 5083 13875 5089
rect 13817 5049 13829 5083
rect 13863 5080 13875 5083
rect 14458 5080 14464 5092
rect 13863 5052 14464 5080
rect 13863 5049 13875 5052
rect 13817 5043 13875 5049
rect 14458 5040 14464 5052
rect 14516 5040 14522 5092
rect 23014 5040 23020 5092
rect 23072 5080 23078 5092
rect 25593 5083 25651 5089
rect 25593 5080 25605 5083
rect 23072 5052 25605 5080
rect 23072 5040 23078 5052
rect 25593 5049 25605 5052
rect 25639 5049 25651 5083
rect 25593 5043 25651 5049
rect 13630 5012 13636 5024
rect 12452 4984 13636 5012
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 13906 4972 13912 5024
rect 13964 4972 13970 5024
rect 19242 4972 19248 5024
rect 19300 4972 19306 5024
rect 25700 5012 25728 5120
rect 25866 5108 25872 5160
rect 25924 5108 25930 5160
rect 26050 5157 26056 5160
rect 26007 5151 26056 5157
rect 26007 5117 26019 5151
rect 26053 5117 26056 5151
rect 26007 5111 26056 5117
rect 26050 5108 26056 5111
rect 26108 5108 26114 5160
rect 27724 5080 27752 5179
rect 28902 5176 28908 5188
rect 28960 5176 28966 5228
rect 28994 5176 29000 5228
rect 29052 5216 29058 5228
rect 35434 5216 35440 5228
rect 29052 5188 30236 5216
rect 29052 5176 29058 5188
rect 30208 5160 30236 5188
rect 34256 5188 35440 5216
rect 27982 5108 27988 5160
rect 28040 5108 28046 5160
rect 29638 5108 29644 5160
rect 29696 5148 29702 5160
rect 30101 5151 30159 5157
rect 30101 5148 30113 5151
rect 29696 5120 30113 5148
rect 29696 5108 29702 5120
rect 30101 5117 30113 5120
rect 30147 5117 30159 5151
rect 30101 5111 30159 5117
rect 30190 5108 30196 5160
rect 30248 5108 30254 5160
rect 32122 5108 32128 5160
rect 32180 5108 32186 5160
rect 32306 5108 32312 5160
rect 32364 5108 32370 5160
rect 33042 5108 33048 5160
rect 33100 5108 33106 5160
rect 33134 5108 33140 5160
rect 33192 5157 33198 5160
rect 33192 5151 33220 5157
rect 33208 5117 33220 5151
rect 33192 5111 33220 5117
rect 33321 5151 33379 5157
rect 33321 5117 33333 5151
rect 33367 5148 33379 5151
rect 34146 5148 34152 5160
rect 33367 5120 34152 5148
rect 33367 5117 33379 5120
rect 33321 5111 33379 5117
rect 33192 5108 33198 5111
rect 34146 5108 34152 5120
rect 34204 5108 34210 5160
rect 26528 5052 27752 5080
rect 32769 5083 32827 5089
rect 25958 5012 25964 5024
rect 25700 4984 25964 5012
rect 25958 4972 25964 4984
rect 26016 5012 26022 5024
rect 26528 5012 26556 5052
rect 32769 5049 32781 5083
rect 32815 5049 32827 5083
rect 32769 5043 32827 5049
rect 26016 4984 26556 5012
rect 27341 5015 27399 5021
rect 26016 4972 26022 4984
rect 27341 4981 27353 5015
rect 27387 5012 27399 5015
rect 27522 5012 27528 5024
rect 27387 4984 27528 5012
rect 27387 4981 27399 4984
rect 27341 4975 27399 4981
rect 27522 4972 27528 4984
rect 27580 4972 27586 5024
rect 32784 5012 32812 5043
rect 33410 5012 33416 5024
rect 32784 4984 33416 5012
rect 33410 4972 33416 4984
rect 33468 4972 33474 5024
rect 33502 4972 33508 5024
rect 33560 5012 33566 5024
rect 34256 5012 34284 5188
rect 35434 5176 35440 5188
rect 35492 5176 35498 5228
rect 34606 5108 34612 5160
rect 34664 5148 34670 5160
rect 34790 5148 34796 5160
rect 34664 5120 34796 5148
rect 34664 5108 34670 5120
rect 34790 5108 34796 5120
rect 34848 5108 34854 5160
rect 33560 4984 34284 5012
rect 33560 4972 33566 4984
rect 35434 4972 35440 5024
rect 35492 5012 35498 5024
rect 36173 5015 36231 5021
rect 36173 5012 36185 5015
rect 35492 4984 36185 5012
rect 35492 4972 35498 4984
rect 36173 4981 36185 4984
rect 36219 4981 36231 5015
rect 36173 4975 36231 4981
rect 1104 4922 47104 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 47104 4922
rect 1104 4848 47104 4870
rect 10686 4768 10692 4820
rect 10744 4768 10750 4820
rect 17218 4768 17224 4820
rect 17276 4768 17282 4820
rect 21634 4768 21640 4820
rect 21692 4808 21698 4820
rect 22465 4811 22523 4817
rect 22465 4808 22477 4811
rect 21692 4780 22477 4808
rect 21692 4768 21698 4780
rect 22465 4777 22477 4780
rect 22511 4777 22523 4811
rect 25774 4808 25780 4820
rect 22465 4771 22523 4777
rect 25700 4780 25780 4808
rect 25700 4740 25728 4780
rect 25774 4768 25780 4780
rect 25832 4768 25838 4820
rect 26252 4780 31754 4808
rect 25958 4740 25964 4752
rect 15396 4712 25728 4740
rect 25792 4712 25964 4740
rect 15396 4681 15424 4712
rect 15381 4675 15439 4681
rect 15381 4641 15393 4675
rect 15427 4641 15439 4675
rect 15381 4635 15439 4641
rect 18230 4632 18236 4684
rect 18288 4672 18294 4684
rect 18325 4675 18383 4681
rect 18325 4672 18337 4675
rect 18288 4644 18337 4672
rect 18288 4632 18294 4644
rect 18325 4641 18337 4644
rect 18371 4672 18383 4675
rect 19889 4675 19947 4681
rect 19889 4672 19901 4675
rect 18371 4644 19901 4672
rect 18371 4641 18383 4644
rect 18325 4635 18383 4641
rect 19889 4641 19901 4644
rect 19935 4672 19947 4675
rect 20346 4672 20352 4684
rect 19935 4644 20352 4672
rect 19935 4641 19947 4644
rect 19889 4635 19947 4641
rect 20346 4632 20352 4644
rect 20404 4632 20410 4684
rect 23109 4675 23167 4681
rect 23109 4641 23121 4675
rect 23155 4641 23167 4675
rect 23109 4635 23167 4641
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4604 10931 4607
rect 11514 4604 11520 4616
rect 10919 4576 11520 4604
rect 10919 4573 10931 4576
rect 10873 4567 10931 4573
rect 11514 4564 11520 4576
rect 11572 4564 11578 4616
rect 15010 4564 15016 4616
rect 15068 4604 15074 4616
rect 15565 4607 15623 4613
rect 15565 4604 15577 4607
rect 15068 4576 15577 4604
rect 15068 4564 15074 4576
rect 15565 4573 15577 4576
rect 15611 4573 15623 4607
rect 15565 4567 15623 4573
rect 15838 4564 15844 4616
rect 15896 4564 15902 4616
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4604 17463 4607
rect 17451 4576 17724 4604
rect 17451 4573 17463 4576
rect 17405 4567 17463 4573
rect 15197 4539 15255 4545
rect 15197 4505 15209 4539
rect 15243 4536 15255 4539
rect 15856 4536 15884 4564
rect 15243 4508 15884 4536
rect 15243 4505 15255 4508
rect 15197 4499 15255 4505
rect 14734 4428 14740 4480
rect 14792 4428 14798 4480
rect 15102 4428 15108 4480
rect 15160 4428 15166 4480
rect 17696 4477 17724 4576
rect 17862 4564 17868 4616
rect 17920 4604 17926 4616
rect 18049 4607 18107 4613
rect 18049 4604 18061 4607
rect 17920 4576 18061 4604
rect 17920 4564 17926 4576
rect 18049 4573 18061 4576
rect 18095 4573 18107 4607
rect 18049 4567 18107 4573
rect 18141 4607 18199 4613
rect 18141 4573 18153 4607
rect 18187 4604 18199 4607
rect 19242 4604 19248 4616
rect 18187 4576 19248 4604
rect 18187 4573 18199 4576
rect 18141 4567 18199 4573
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 22830 4564 22836 4616
rect 22888 4564 22894 4616
rect 23124 4604 23152 4635
rect 24946 4632 24952 4684
rect 25004 4672 25010 4684
rect 25590 4672 25596 4684
rect 25004 4644 25596 4672
rect 25004 4632 25010 4644
rect 25590 4632 25596 4644
rect 25648 4632 25654 4684
rect 25792 4681 25820 4712
rect 25958 4700 25964 4712
rect 26016 4700 26022 4752
rect 26252 4749 26280 4780
rect 26237 4743 26295 4749
rect 26237 4709 26249 4743
rect 26283 4709 26295 4743
rect 26237 4703 26295 4709
rect 27430 4700 27436 4752
rect 27488 4700 27494 4752
rect 28902 4700 28908 4752
rect 28960 4700 28966 4752
rect 28994 4700 29000 4752
rect 29052 4700 29058 4752
rect 29549 4743 29607 4749
rect 29549 4709 29561 4743
rect 29595 4709 29607 4743
rect 31726 4740 31754 4780
rect 31846 4768 31852 4820
rect 31904 4808 31910 4820
rect 33965 4811 34023 4817
rect 33965 4808 33977 4811
rect 31904 4780 33977 4808
rect 31904 4768 31910 4780
rect 33965 4777 33977 4780
rect 34011 4777 34023 4811
rect 33965 4771 34023 4777
rect 35069 4811 35127 4817
rect 35069 4777 35081 4811
rect 35115 4808 35127 4811
rect 35342 4808 35348 4820
rect 35115 4780 35348 4808
rect 35115 4777 35127 4780
rect 35069 4771 35127 4777
rect 35342 4768 35348 4780
rect 35400 4768 35406 4820
rect 32769 4743 32827 4749
rect 32769 4740 32781 4743
rect 31726 4712 32781 4740
rect 29549 4703 29607 4709
rect 32769 4709 32781 4712
rect 32815 4740 32827 4743
rect 32858 4740 32864 4752
rect 32815 4712 32864 4740
rect 32815 4709 32827 4712
rect 32769 4703 32827 4709
rect 25777 4675 25835 4681
rect 25777 4641 25789 4675
rect 25823 4641 25835 4675
rect 25777 4635 25835 4641
rect 25866 4632 25872 4684
rect 25924 4672 25930 4684
rect 26513 4675 26571 4681
rect 26513 4672 26525 4675
rect 25924 4644 26525 4672
rect 25924 4632 25930 4644
rect 26513 4641 26525 4644
rect 26559 4641 26571 4675
rect 26513 4635 26571 4641
rect 26789 4675 26847 4681
rect 26789 4641 26801 4675
rect 26835 4672 26847 4675
rect 26835 4644 27660 4672
rect 26835 4641 26847 4644
rect 26789 4635 26847 4641
rect 25958 4604 25964 4616
rect 23124 4576 25964 4604
rect 25958 4564 25964 4576
rect 26016 4564 26022 4616
rect 26602 4564 26608 4616
rect 26660 4613 26666 4616
rect 26660 4607 26688 4613
rect 26676 4573 26688 4607
rect 26660 4567 26688 4573
rect 26660 4564 26666 4567
rect 27430 4564 27436 4616
rect 27488 4604 27494 4616
rect 27525 4607 27583 4613
rect 27525 4604 27537 4607
rect 27488 4576 27537 4604
rect 27488 4564 27494 4576
rect 27525 4573 27537 4576
rect 27571 4573 27583 4607
rect 27632 4604 27660 4644
rect 29181 4607 29239 4613
rect 27632 4576 29132 4604
rect 27525 4567 27583 4573
rect 19613 4539 19671 4545
rect 19613 4505 19625 4539
rect 19659 4536 19671 4539
rect 19794 4536 19800 4548
rect 19659 4508 19800 4536
rect 19659 4505 19671 4508
rect 19613 4499 19671 4505
rect 19794 4496 19800 4508
rect 19852 4496 19858 4548
rect 21726 4496 21732 4548
rect 21784 4536 21790 4548
rect 22925 4539 22983 4545
rect 22925 4536 22937 4539
rect 21784 4508 22937 4536
rect 21784 4496 21790 4508
rect 22925 4505 22937 4508
rect 22971 4536 22983 4539
rect 25130 4536 25136 4548
rect 22971 4508 25136 4536
rect 22971 4505 22983 4508
rect 22925 4499 22983 4505
rect 25130 4496 25136 4508
rect 25188 4496 25194 4548
rect 27614 4496 27620 4548
rect 27672 4536 27678 4548
rect 27770 4539 27828 4545
rect 27770 4536 27782 4539
rect 27672 4508 27782 4536
rect 27672 4496 27678 4508
rect 27770 4505 27782 4508
rect 27816 4505 27828 4539
rect 29104 4536 29132 4576
rect 29181 4573 29193 4607
rect 29227 4604 29239 4607
rect 29564 4604 29592 4703
rect 32858 4700 32864 4712
rect 32916 4700 32922 4752
rect 29730 4632 29736 4684
rect 29788 4672 29794 4684
rect 30101 4675 30159 4681
rect 30101 4672 30113 4675
rect 29788 4644 30113 4672
rect 29788 4632 29794 4644
rect 30101 4641 30113 4644
rect 30147 4641 30159 4675
rect 30101 4635 30159 4641
rect 32122 4632 32128 4684
rect 32180 4632 32186 4684
rect 32674 4672 32680 4684
rect 32232 4644 32680 4672
rect 29227 4576 29592 4604
rect 29227 4573 29239 4576
rect 29181 4567 29239 4573
rect 29914 4564 29920 4616
rect 29972 4564 29978 4616
rect 32030 4564 32036 4616
rect 32088 4564 32094 4616
rect 32232 4536 32260 4644
rect 32674 4632 32680 4644
rect 32732 4632 32738 4684
rect 33045 4675 33103 4681
rect 33045 4641 33057 4675
rect 33091 4672 33103 4675
rect 33502 4672 33508 4684
rect 33091 4644 33508 4672
rect 33091 4641 33103 4644
rect 33045 4635 33103 4641
rect 33502 4632 33508 4644
rect 33560 4632 33566 4684
rect 35713 4675 35771 4681
rect 35713 4641 35725 4675
rect 35759 4672 35771 4675
rect 36078 4672 36084 4684
rect 35759 4644 36084 4672
rect 35759 4641 35771 4644
rect 35713 4635 35771 4641
rect 36078 4632 36084 4644
rect 36136 4672 36142 4684
rect 36538 4672 36544 4684
rect 36136 4644 36544 4672
rect 36136 4632 36142 4644
rect 36538 4632 36544 4644
rect 36596 4632 36602 4684
rect 32306 4564 32312 4616
rect 32364 4564 32370 4616
rect 33134 4564 33140 4616
rect 33192 4613 33198 4616
rect 33192 4607 33220 4613
rect 33208 4573 33220 4607
rect 33192 4567 33220 4573
rect 33192 4564 33198 4567
rect 33318 4564 33324 4616
rect 33376 4564 33382 4616
rect 35434 4564 35440 4616
rect 35492 4564 35498 4616
rect 35529 4607 35587 4613
rect 35529 4573 35541 4607
rect 35575 4604 35587 4607
rect 35986 4604 35992 4616
rect 35575 4576 35992 4604
rect 35575 4573 35587 4576
rect 35529 4567 35587 4573
rect 35986 4564 35992 4576
rect 36044 4564 36050 4616
rect 38286 4564 38292 4616
rect 38344 4564 38350 4616
rect 29104 4508 32260 4536
rect 27770 4499 27828 4505
rect 17681 4471 17739 4477
rect 17681 4437 17693 4471
rect 17727 4437 17739 4471
rect 17681 4431 17739 4437
rect 18598 4428 18604 4480
rect 18656 4468 18662 4480
rect 19245 4471 19303 4477
rect 19245 4468 19257 4471
rect 18656 4440 19257 4468
rect 18656 4428 18662 4440
rect 19245 4437 19257 4440
rect 19291 4437 19303 4471
rect 19245 4431 19303 4437
rect 19705 4471 19763 4477
rect 19705 4437 19717 4471
rect 19751 4468 19763 4471
rect 21358 4468 21364 4480
rect 19751 4440 21364 4468
rect 19751 4437 19763 4440
rect 19705 4431 19763 4437
rect 21358 4428 21364 4440
rect 21416 4428 21422 4480
rect 24854 4428 24860 4480
rect 24912 4468 24918 4480
rect 26050 4468 26056 4480
rect 24912 4440 26056 4468
rect 24912 4428 24918 4440
rect 26050 4428 26056 4440
rect 26108 4468 26114 4480
rect 26602 4468 26608 4480
rect 26108 4440 26608 4468
rect 26108 4428 26114 4440
rect 26602 4428 26608 4440
rect 26660 4428 26666 4480
rect 27338 4428 27344 4480
rect 27396 4468 27402 4480
rect 29822 4468 29828 4480
rect 27396 4440 29828 4468
rect 27396 4428 27402 4440
rect 29822 4428 29828 4440
rect 29880 4468 29886 4480
rect 30009 4471 30067 4477
rect 30009 4468 30021 4471
rect 29880 4440 30021 4468
rect 29880 4428 29886 4440
rect 30009 4437 30021 4440
rect 30055 4437 30067 4471
rect 30009 4431 30067 4437
rect 31846 4428 31852 4480
rect 31904 4428 31910 4480
rect 32324 4468 32352 4564
rect 35452 4536 35480 4564
rect 33796 4508 35480 4536
rect 33796 4468 33824 4508
rect 32324 4440 33824 4468
rect 1104 4378 47104 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 47104 4378
rect 1104 4304 47104 4326
rect 18417 4267 18475 4273
rect 18417 4233 18429 4267
rect 18463 4233 18475 4267
rect 18417 4227 18475 4233
rect 17497 4199 17555 4205
rect 17497 4165 17509 4199
rect 17543 4196 17555 4199
rect 17770 4196 17776 4208
rect 17543 4168 17776 4196
rect 17543 4165 17555 4168
rect 17497 4159 17555 4165
rect 17770 4156 17776 4168
rect 17828 4156 17834 4208
rect 18432 4196 18460 4227
rect 19794 4224 19800 4276
rect 19852 4264 19858 4276
rect 20073 4267 20131 4273
rect 20073 4264 20085 4267
rect 19852 4236 20085 4264
rect 19852 4224 19858 4236
rect 20073 4233 20085 4236
rect 20119 4233 20131 4267
rect 20073 4227 20131 4233
rect 22186 4224 22192 4276
rect 22244 4264 22250 4276
rect 22554 4264 22560 4276
rect 22244 4236 22560 4264
rect 22244 4224 22250 4236
rect 22554 4224 22560 4236
rect 22612 4224 22618 4276
rect 24949 4267 25007 4273
rect 24949 4233 24961 4267
rect 24995 4264 25007 4267
rect 25866 4264 25872 4276
rect 24995 4236 25872 4264
rect 24995 4233 25007 4236
rect 24949 4227 25007 4233
rect 25866 4224 25872 4236
rect 25924 4224 25930 4276
rect 25958 4224 25964 4276
rect 26016 4264 26022 4276
rect 27982 4264 27988 4276
rect 26016 4236 27988 4264
rect 26016 4224 26022 4236
rect 27982 4224 27988 4236
rect 28040 4264 28046 4276
rect 36078 4264 36084 4276
rect 28040 4236 36084 4264
rect 28040 4224 28046 4236
rect 36078 4224 36084 4236
rect 36136 4224 36142 4276
rect 18432 4168 18736 4196
rect 14366 4137 14372 4140
rect 14360 4091 14372 4137
rect 14366 4088 14372 4091
rect 14424 4088 14430 4140
rect 17034 4088 17040 4140
rect 17092 4088 17098 4140
rect 18598 4088 18604 4140
rect 18656 4088 18662 4140
rect 18708 4128 18736 4168
rect 19242 4156 19248 4208
rect 19300 4196 19306 4208
rect 27338 4196 27344 4208
rect 19300 4168 27344 4196
rect 19300 4156 19306 4168
rect 27338 4156 27344 4168
rect 27396 4156 27402 4208
rect 27430 4156 27436 4208
rect 27488 4196 27494 4208
rect 27488 4168 27660 4196
rect 27488 4156 27494 4168
rect 18949 4131 19007 4137
rect 18949 4128 18961 4131
rect 18708 4100 18961 4128
rect 18949 4097 18961 4100
rect 18995 4097 19007 4131
rect 18949 4091 19007 4097
rect 21269 4131 21327 4137
rect 21269 4097 21281 4131
rect 21315 4128 21327 4131
rect 21315 4100 21864 4128
rect 21315 4097 21327 4100
rect 21269 4091 21327 4097
rect 13630 4020 13636 4072
rect 13688 4060 13694 4072
rect 14093 4063 14151 4069
rect 14093 4060 14105 4063
rect 13688 4032 14105 4060
rect 13688 4020 13694 4032
rect 14093 4029 14105 4032
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 15838 4020 15844 4072
rect 15896 4060 15902 4072
rect 17589 4063 17647 4069
rect 17589 4060 17601 4063
rect 15896 4032 17601 4060
rect 15896 4020 15902 4032
rect 17589 4029 17601 4032
rect 17635 4029 17647 4063
rect 17589 4023 17647 4029
rect 17773 4063 17831 4069
rect 17773 4029 17785 4063
rect 17819 4060 17831 4063
rect 18230 4060 18236 4072
rect 17819 4032 18236 4060
rect 17819 4029 17831 4032
rect 17773 4023 17831 4029
rect 15102 3952 15108 4004
rect 15160 3992 15166 4004
rect 15473 3995 15531 4001
rect 15473 3992 15485 3995
rect 15160 3964 15485 3992
rect 15160 3952 15166 3964
rect 15473 3961 15485 3964
rect 15519 3961 15531 3995
rect 15473 3955 15531 3961
rect 16666 3952 16672 4004
rect 16724 3992 16730 4004
rect 17129 3995 17187 4001
rect 17129 3992 17141 3995
rect 16724 3964 17141 3992
rect 16724 3952 16730 3964
rect 17129 3961 17141 3964
rect 17175 3961 17187 3995
rect 17604 3992 17632 4023
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 18693 4063 18751 4069
rect 18693 4029 18705 4063
rect 18739 4029 18751 4063
rect 18693 4023 18751 4029
rect 18322 3992 18328 4004
rect 17604 3964 18328 3992
rect 17129 3955 17187 3961
rect 18322 3952 18328 3964
rect 18380 3952 18386 4004
rect 16853 3927 16911 3933
rect 16853 3893 16865 3927
rect 16899 3924 16911 3927
rect 16942 3924 16948 3936
rect 16899 3896 16948 3924
rect 16899 3893 16911 3896
rect 16853 3887 16911 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 18708 3924 18736 4023
rect 21836 4001 21864 4100
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 23937 4131 23995 4137
rect 23937 4128 23949 4131
rect 23532 4100 23949 4128
rect 23532 4088 23538 4100
rect 23937 4097 23949 4100
rect 23983 4097 23995 4131
rect 23937 4091 23995 4097
rect 25774 4088 25780 4140
rect 25832 4128 25838 4140
rect 26145 4131 26203 4137
rect 26145 4128 26157 4131
rect 25832 4100 26157 4128
rect 25832 4088 25838 4100
rect 26145 4097 26157 4100
rect 26191 4097 26203 4131
rect 26145 4091 26203 4097
rect 27522 4088 27528 4140
rect 27580 4088 27586 4140
rect 27632 4128 27660 4168
rect 28994 4156 29000 4208
rect 29052 4156 29058 4208
rect 31846 4156 31852 4208
rect 31904 4196 31910 4208
rect 33014 4199 33072 4205
rect 33014 4196 33026 4199
rect 31904 4168 33026 4196
rect 31904 4156 31910 4168
rect 33014 4165 33026 4168
rect 33060 4165 33072 4199
rect 33014 4159 33072 4165
rect 38096 4199 38154 4205
rect 38096 4165 38108 4199
rect 38142 4196 38154 4199
rect 38286 4196 38292 4208
rect 38142 4168 38292 4196
rect 38142 4165 38154 4168
rect 38096 4159 38154 4165
rect 38286 4156 38292 4168
rect 38344 4156 38350 4208
rect 28626 4128 28632 4140
rect 27632 4100 28632 4128
rect 28626 4088 28632 4100
rect 28684 4088 28690 4140
rect 28896 4131 28954 4137
rect 28896 4097 28908 4131
rect 28942 4128 28954 4131
rect 29012 4128 29040 4156
rect 28942 4100 29040 4128
rect 28942 4097 28954 4100
rect 28896 4091 28954 4097
rect 31018 4088 31024 4140
rect 31076 4088 31082 4140
rect 31938 4088 31944 4140
rect 31996 4128 32002 4140
rect 32214 4128 32220 4140
rect 31996 4100 32220 4128
rect 31996 4088 32002 4100
rect 32214 4088 32220 4100
rect 32272 4128 32278 4140
rect 32769 4131 32827 4137
rect 32769 4128 32781 4131
rect 32272 4100 32781 4128
rect 32272 4088 32278 4100
rect 32769 4097 32781 4100
rect 32815 4097 32827 4131
rect 32769 4091 32827 4097
rect 34790 4088 34796 4140
rect 34848 4128 34854 4140
rect 37829 4131 37887 4137
rect 37829 4128 37841 4131
rect 34848 4100 37841 4128
rect 34848 4088 34854 4100
rect 37829 4097 37841 4100
rect 37875 4097 37887 4131
rect 37829 4091 37887 4097
rect 22281 4063 22339 4069
rect 22281 4029 22293 4063
rect 22327 4029 22339 4063
rect 22281 4023 22339 4029
rect 21821 3995 21879 4001
rect 21821 3961 21833 3995
rect 21867 3961 21879 3995
rect 21821 3955 21879 3961
rect 19334 3924 19340 3936
rect 17368 3896 19340 3924
rect 17368 3884 17374 3896
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 21082 3884 21088 3936
rect 21140 3884 21146 3936
rect 21174 3884 21180 3936
rect 21232 3924 21238 3936
rect 22296 3924 22324 4023
rect 22462 4020 22468 4072
rect 22520 4060 22526 4072
rect 22520 4032 23980 4060
rect 22520 4020 22526 4032
rect 23952 3992 23980 4032
rect 24026 4020 24032 4072
rect 24084 4060 24090 4072
rect 25038 4060 25044 4072
rect 24084 4032 25044 4060
rect 24084 4020 24090 4032
rect 25038 4020 25044 4032
rect 25096 4020 25102 4072
rect 25133 4063 25191 4069
rect 25133 4029 25145 4063
rect 25179 4029 25191 4063
rect 25133 4023 25191 4029
rect 25148 3992 25176 4023
rect 27341 3995 27399 4001
rect 23952 3964 26924 3992
rect 22738 3924 22744 3936
rect 21232 3896 22744 3924
rect 21232 3884 21238 3896
rect 22738 3884 22744 3896
rect 22796 3884 22802 3936
rect 23750 3884 23756 3936
rect 23808 3884 23814 3936
rect 24581 3927 24639 3933
rect 24581 3893 24593 3927
rect 24627 3924 24639 3927
rect 25130 3924 25136 3936
rect 24627 3896 25136 3924
rect 24627 3893 24639 3896
rect 24581 3887 24639 3893
rect 25130 3884 25136 3896
rect 25188 3884 25194 3936
rect 25961 3927 26019 3933
rect 25961 3893 25973 3927
rect 26007 3924 26019 3927
rect 26050 3924 26056 3936
rect 26007 3896 26056 3924
rect 26007 3893 26019 3896
rect 25961 3887 26019 3893
rect 26050 3884 26056 3896
rect 26108 3884 26114 3936
rect 26896 3924 26924 3964
rect 27341 3961 27353 3995
rect 27387 3992 27399 3995
rect 27614 3992 27620 4004
rect 27387 3964 27620 3992
rect 27387 3961 27399 3964
rect 27341 3955 27399 3961
rect 27614 3952 27620 3964
rect 27672 3952 27678 4004
rect 29914 3952 29920 4004
rect 29972 3992 29978 4004
rect 30009 3995 30067 4001
rect 30009 3992 30021 3995
rect 29972 3964 30021 3992
rect 29972 3952 29978 3964
rect 30009 3961 30021 3964
rect 30055 3961 30067 3995
rect 32766 3992 32772 4004
rect 30009 3955 30067 3961
rect 30116 3964 32772 3992
rect 30116 3924 30144 3964
rect 32766 3952 32772 3964
rect 32824 3952 32830 4004
rect 39206 3952 39212 4004
rect 39264 3992 39270 4004
rect 44542 3992 44548 4004
rect 39264 3964 44548 3992
rect 39264 3952 39270 3964
rect 44542 3952 44548 3964
rect 44600 3952 44606 4004
rect 26896 3896 30144 3924
rect 30742 3884 30748 3936
rect 30800 3924 30806 3936
rect 30837 3927 30895 3933
rect 30837 3924 30849 3927
rect 30800 3896 30849 3924
rect 30800 3884 30806 3896
rect 30837 3893 30849 3896
rect 30883 3893 30895 3927
rect 30837 3887 30895 3893
rect 32122 3884 32128 3936
rect 32180 3924 32186 3936
rect 34149 3927 34207 3933
rect 34149 3924 34161 3927
rect 32180 3896 34161 3924
rect 32180 3884 32186 3896
rect 34149 3893 34161 3896
rect 34195 3893 34207 3927
rect 34149 3887 34207 3893
rect 1104 3834 47104 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 47104 3834
rect 1104 3760 47104 3782
rect 14366 3680 14372 3732
rect 14424 3720 14430 3732
rect 14553 3723 14611 3729
rect 14553 3720 14565 3723
rect 14424 3692 14565 3720
rect 14424 3680 14430 3692
rect 14553 3689 14565 3692
rect 14599 3689 14611 3723
rect 14553 3683 14611 3689
rect 17034 3680 17040 3732
rect 17092 3720 17098 3732
rect 18233 3723 18291 3729
rect 18233 3720 18245 3723
rect 17092 3692 18245 3720
rect 17092 3680 17098 3692
rect 18233 3689 18245 3692
rect 18279 3689 18291 3723
rect 18233 3683 18291 3689
rect 18322 3680 18328 3732
rect 18380 3720 18386 3732
rect 21174 3720 21180 3732
rect 18380 3692 21180 3720
rect 18380 3680 18386 3692
rect 17770 3612 17776 3664
rect 17828 3652 17834 3664
rect 18141 3655 18199 3661
rect 18141 3652 18153 3655
rect 17828 3624 18153 3652
rect 17828 3612 17834 3624
rect 18141 3621 18153 3624
rect 18187 3621 18199 3655
rect 18141 3615 18199 3621
rect 18524 3624 20392 3652
rect 15657 3587 15715 3593
rect 15657 3553 15669 3587
rect 15703 3584 15715 3587
rect 16390 3584 16396 3596
rect 15703 3556 16396 3584
rect 15703 3553 15715 3556
rect 15657 3547 15715 3553
rect 16390 3544 16396 3556
rect 16448 3544 16454 3596
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 14476 3448 14504 3479
rect 14734 3476 14740 3528
rect 14792 3476 14798 3528
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3516 15439 3519
rect 15838 3516 15844 3528
rect 15427 3488 15844 3516
rect 15427 3485 15439 3488
rect 15381 3479 15439 3485
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 16666 3476 16672 3528
rect 16724 3476 16730 3528
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 17310 3516 17316 3528
rect 16816 3488 17316 3516
rect 16816 3476 16822 3488
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17006 3451 17064 3457
rect 17006 3448 17018 3451
rect 14476 3420 15056 3448
rect 14274 3340 14280 3392
rect 14332 3340 14338 3392
rect 15028 3389 15056 3420
rect 16500 3420 17018 3448
rect 15013 3383 15071 3389
rect 15013 3349 15025 3383
rect 15059 3349 15071 3383
rect 15013 3343 15071 3349
rect 15470 3340 15476 3392
rect 15528 3340 15534 3392
rect 16500 3389 16528 3420
rect 17006 3417 17018 3420
rect 17052 3417 17064 3451
rect 17006 3411 17064 3417
rect 16485 3383 16543 3389
rect 16485 3349 16497 3383
rect 16531 3349 16543 3383
rect 16485 3343 16543 3349
rect 16574 3340 16580 3392
rect 16632 3380 16638 3392
rect 18524 3380 18552 3624
rect 18782 3544 18788 3596
rect 18840 3584 18846 3596
rect 18840 3556 20116 3584
rect 18840 3544 18846 3556
rect 18598 3476 18604 3528
rect 18656 3476 18662 3528
rect 19889 3519 19947 3525
rect 19889 3485 19901 3519
rect 19935 3516 19947 3519
rect 19935 3488 20024 3516
rect 19935 3485 19947 3488
rect 19889 3479 19947 3485
rect 16632 3352 18552 3380
rect 16632 3340 16638 3352
rect 18690 3340 18696 3392
rect 18748 3340 18754 3392
rect 19705 3383 19763 3389
rect 19705 3349 19717 3383
rect 19751 3380 19763 3383
rect 19794 3380 19800 3392
rect 19751 3352 19800 3380
rect 19751 3349 19763 3352
rect 19705 3343 19763 3349
rect 19794 3340 19800 3352
rect 19852 3340 19858 3392
rect 19996 3389 20024 3488
rect 19981 3383 20039 3389
rect 19981 3349 19993 3383
rect 20027 3349 20039 3383
rect 20088 3380 20116 3556
rect 20364 3516 20392 3624
rect 20456 3593 20484 3692
rect 21174 3680 21180 3692
rect 21232 3680 21238 3732
rect 22186 3680 22192 3732
rect 22244 3680 22250 3732
rect 23474 3680 23480 3732
rect 23532 3680 23538 3732
rect 25777 3723 25835 3729
rect 25777 3689 25789 3723
rect 25823 3720 25835 3723
rect 25866 3720 25872 3732
rect 25823 3692 25872 3720
rect 25823 3689 25835 3692
rect 25777 3683 25835 3689
rect 25866 3680 25872 3692
rect 25924 3680 25930 3732
rect 27430 3720 27436 3732
rect 25976 3692 27436 3720
rect 22281 3655 22339 3661
rect 22281 3621 22293 3655
rect 22327 3652 22339 3655
rect 22370 3652 22376 3664
rect 22327 3624 22376 3652
rect 22327 3621 22339 3624
rect 22281 3615 22339 3621
rect 22370 3612 22376 3624
rect 22428 3612 22434 3664
rect 20441 3587 20499 3593
rect 20441 3553 20453 3587
rect 20487 3553 20499 3587
rect 20441 3547 20499 3553
rect 20622 3544 20628 3596
rect 20680 3544 20686 3596
rect 20732 3556 20944 3584
rect 20640 3516 20668 3544
rect 20364 3488 20668 3516
rect 20349 3451 20407 3457
rect 20349 3417 20361 3451
rect 20395 3448 20407 3451
rect 20732 3448 20760 3556
rect 20916 3528 20944 3556
rect 22738 3544 22744 3596
rect 22796 3544 22802 3596
rect 22830 3544 22836 3596
rect 22888 3544 22894 3596
rect 24118 3544 24124 3596
rect 24176 3584 24182 3596
rect 25976 3593 26004 3692
rect 27430 3680 27436 3692
rect 27488 3680 27494 3732
rect 31938 3720 31944 3732
rect 30484 3692 31944 3720
rect 25961 3587 26019 3593
rect 24176 3556 24523 3584
rect 24176 3544 24182 3556
rect 20809 3519 20867 3525
rect 20809 3485 20821 3519
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 20395 3420 20760 3448
rect 20824 3448 20852 3479
rect 20898 3476 20904 3528
rect 20956 3476 20962 3528
rect 21082 3525 21088 3528
rect 21076 3516 21088 3525
rect 21043 3488 21088 3516
rect 21076 3479 21088 3488
rect 21082 3476 21088 3479
rect 21140 3476 21146 3528
rect 21358 3476 21364 3528
rect 21416 3516 21422 3528
rect 21416 3512 22232 3516
rect 21416 3488 22324 3512
rect 21416 3476 21422 3488
rect 22204 3484 22324 3488
rect 21818 3448 21824 3460
rect 20824 3420 21824 3448
rect 20395 3417 20407 3420
rect 20349 3411 20407 3417
rect 21818 3408 21824 3420
rect 21876 3408 21882 3460
rect 22296 3448 22324 3484
rect 22370 3476 22376 3528
rect 22428 3516 22434 3528
rect 23293 3519 23351 3525
rect 23293 3516 23305 3519
rect 22428 3488 23305 3516
rect 22428 3476 22434 3488
rect 23293 3485 23305 3488
rect 23339 3485 23351 3519
rect 23937 3519 23995 3525
rect 23937 3516 23949 3519
rect 23293 3479 23351 3485
rect 23768 3488 23949 3516
rect 23768 3448 23796 3488
rect 23937 3485 23949 3488
rect 23983 3516 23995 3519
rect 24026 3516 24032 3528
rect 23983 3488 24032 3516
rect 23983 3485 23995 3488
rect 23937 3479 23995 3485
rect 24026 3476 24032 3488
rect 24084 3476 24090 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 24268 3488 24409 3516
rect 24268 3476 24274 3488
rect 24397 3485 24409 3488
rect 24443 3485 24455 3519
rect 24495 3516 24523 3556
rect 25961 3553 25973 3587
rect 26007 3553 26019 3587
rect 25961 3547 26019 3553
rect 29362 3544 29368 3596
rect 29420 3584 29426 3596
rect 30006 3584 30012 3596
rect 29420 3556 30012 3584
rect 29420 3544 29426 3556
rect 30006 3544 30012 3556
rect 30064 3544 30070 3596
rect 30190 3544 30196 3596
rect 30248 3544 30254 3596
rect 30484 3593 30512 3692
rect 31938 3680 31944 3692
rect 31996 3680 32002 3732
rect 32030 3680 32036 3732
rect 32088 3720 32094 3732
rect 32585 3723 32643 3729
rect 32585 3720 32597 3723
rect 32088 3692 32597 3720
rect 32088 3680 32094 3692
rect 32585 3689 32597 3692
rect 32631 3689 32643 3723
rect 32585 3683 32643 3689
rect 32766 3680 32772 3732
rect 32824 3720 32830 3732
rect 32824 3692 34376 3720
rect 32824 3680 32830 3692
rect 31846 3612 31852 3664
rect 31904 3652 31910 3664
rect 33134 3652 33140 3664
rect 31904 3624 33140 3652
rect 31904 3612 31910 3624
rect 33134 3612 33140 3624
rect 33192 3612 33198 3664
rect 34238 3652 34244 3664
rect 33244 3624 34244 3652
rect 33244 3596 33272 3624
rect 34238 3612 34244 3624
rect 34296 3612 34302 3664
rect 30469 3587 30527 3593
rect 30469 3553 30481 3587
rect 30515 3553 30527 3587
rect 30469 3547 30527 3553
rect 31754 3544 31760 3596
rect 31812 3584 31818 3596
rect 32582 3584 32588 3596
rect 31812 3556 32588 3584
rect 31812 3544 31818 3556
rect 32582 3544 32588 3556
rect 32640 3544 32646 3596
rect 33226 3544 33232 3596
rect 33284 3544 33290 3596
rect 33870 3544 33876 3596
rect 33928 3544 33934 3596
rect 34057 3587 34115 3593
rect 34057 3553 34069 3587
rect 34103 3584 34115 3587
rect 34348 3584 34376 3692
rect 34103 3556 34376 3584
rect 34103 3553 34115 3556
rect 34057 3547 34115 3553
rect 35250 3544 35256 3596
rect 35308 3544 35314 3596
rect 24495 3488 25084 3516
rect 24397 3479 24455 3485
rect 21928 3420 22232 3448
rect 22296 3420 23796 3448
rect 23845 3451 23903 3457
rect 21928 3380 21956 3420
rect 20088 3352 21956 3380
rect 22204 3380 22232 3420
rect 23845 3417 23857 3451
rect 23891 3448 23903 3451
rect 24664 3451 24722 3457
rect 23891 3420 24624 3448
rect 23891 3417 23903 3420
rect 23845 3411 23903 3417
rect 22554 3380 22560 3392
rect 22204 3352 22560 3380
rect 19981 3343 20039 3349
rect 22554 3340 22560 3352
rect 22612 3340 22618 3392
rect 22646 3340 22652 3392
rect 22704 3340 22710 3392
rect 23106 3340 23112 3392
rect 23164 3340 23170 3392
rect 24596 3380 24624 3420
rect 24664 3417 24676 3451
rect 24710 3448 24722 3451
rect 24946 3448 24952 3460
rect 24710 3420 24952 3448
rect 24710 3417 24722 3420
rect 24664 3411 24722 3417
rect 24946 3408 24952 3420
rect 25004 3408 25010 3460
rect 25056 3448 25084 3488
rect 26050 3476 26056 3528
rect 26108 3516 26114 3528
rect 26217 3519 26275 3525
rect 26217 3516 26229 3519
rect 26108 3488 26229 3516
rect 26108 3476 26114 3488
rect 26217 3485 26229 3488
rect 26263 3485 26275 3519
rect 26217 3479 26275 3485
rect 27614 3476 27620 3528
rect 27672 3476 27678 3528
rect 29822 3476 29828 3528
rect 29880 3516 29886 3528
rect 29917 3519 29975 3525
rect 29917 3516 29929 3519
rect 29880 3488 29929 3516
rect 29880 3476 29886 3488
rect 29917 3485 29929 3488
rect 29963 3516 29975 3519
rect 30558 3516 30564 3528
rect 29963 3488 30564 3516
rect 29963 3485 29975 3488
rect 29917 3479 29975 3485
rect 30558 3476 30564 3488
rect 30616 3476 30622 3528
rect 30742 3525 30748 3528
rect 30736 3516 30748 3525
rect 30703 3488 30748 3516
rect 30736 3479 30748 3488
rect 30742 3476 30748 3479
rect 30800 3476 30806 3528
rect 32125 3519 32183 3525
rect 32125 3485 32137 3519
rect 32171 3516 32183 3519
rect 32171 3488 33364 3516
rect 32171 3485 32183 3488
rect 32125 3479 32183 3485
rect 25056 3420 29684 3448
rect 24854 3380 24860 3392
rect 24596 3352 24860 3380
rect 24854 3340 24860 3352
rect 24912 3340 24918 3392
rect 25590 3340 25596 3392
rect 25648 3380 25654 3392
rect 27341 3383 27399 3389
rect 27341 3380 27353 3383
rect 25648 3352 27353 3380
rect 25648 3340 25654 3352
rect 27341 3349 27353 3352
rect 27387 3349 27399 3383
rect 27341 3343 27399 3349
rect 29362 3340 29368 3392
rect 29420 3380 29426 3392
rect 29549 3383 29607 3389
rect 29549 3380 29561 3383
rect 29420 3352 29561 3380
rect 29420 3340 29426 3352
rect 29549 3349 29561 3352
rect 29595 3349 29607 3383
rect 29656 3380 29684 3420
rect 31478 3408 31484 3460
rect 31536 3448 31542 3460
rect 33042 3448 33048 3460
rect 31536 3420 33048 3448
rect 31536 3408 31542 3420
rect 33042 3408 33048 3420
rect 33100 3408 33106 3460
rect 31754 3380 31760 3392
rect 29656 3352 31760 3380
rect 29549 3343 29607 3349
rect 31754 3340 31760 3352
rect 31812 3340 31818 3392
rect 31938 3340 31944 3392
rect 31996 3340 32002 3392
rect 32122 3340 32128 3392
rect 32180 3380 32186 3392
rect 32953 3383 33011 3389
rect 32953 3380 32965 3383
rect 32180 3352 32965 3380
rect 32180 3340 32186 3352
rect 32953 3349 32965 3352
rect 32999 3349 33011 3383
rect 33336 3380 33364 3488
rect 33502 3476 33508 3528
rect 33560 3516 33566 3528
rect 33781 3519 33839 3525
rect 33781 3516 33793 3519
rect 33560 3488 33793 3516
rect 33560 3476 33566 3488
rect 33781 3485 33793 3488
rect 33827 3485 33839 3519
rect 33781 3479 33839 3485
rect 34698 3476 34704 3528
rect 34756 3516 34762 3528
rect 35069 3519 35127 3525
rect 35069 3516 35081 3519
rect 34756 3488 35081 3516
rect 34756 3476 34762 3488
rect 35069 3485 35081 3488
rect 35115 3485 35127 3519
rect 35069 3479 35127 3485
rect 33413 3383 33471 3389
rect 33413 3380 33425 3383
rect 33336 3352 33425 3380
rect 32953 3343 33011 3349
rect 33413 3349 33425 3352
rect 33459 3349 33471 3383
rect 33413 3343 33471 3349
rect 34698 3340 34704 3392
rect 34756 3340 34762 3392
rect 35158 3340 35164 3392
rect 35216 3340 35222 3392
rect 1104 3290 47104 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 47104 3290
rect 1104 3216 47104 3238
rect 15470 3136 15476 3188
rect 15528 3176 15534 3188
rect 15657 3179 15715 3185
rect 15657 3176 15669 3179
rect 15528 3148 15669 3176
rect 15528 3136 15534 3148
rect 15657 3145 15669 3148
rect 15703 3145 15715 3179
rect 15657 3139 15715 3145
rect 18049 3179 18107 3185
rect 18049 3145 18061 3179
rect 18095 3176 18107 3179
rect 18690 3176 18696 3188
rect 18095 3148 18696 3176
rect 18095 3145 18107 3148
rect 18049 3139 18107 3145
rect 18690 3136 18696 3148
rect 18748 3136 18754 3188
rect 20898 3136 20904 3188
rect 20956 3136 20962 3188
rect 22462 3176 22468 3188
rect 22020 3148 22468 3176
rect 14274 3068 14280 3120
rect 14332 3108 14338 3120
rect 14522 3111 14580 3117
rect 14522 3108 14534 3111
rect 14332 3080 14534 3108
rect 14332 3068 14338 3080
rect 14522 3077 14534 3080
rect 14568 3077 14580 3111
rect 14522 3071 14580 3077
rect 17126 3068 17132 3120
rect 17184 3108 17190 3120
rect 22020 3108 22048 3148
rect 22462 3136 22468 3148
rect 22520 3136 22526 3188
rect 22646 3136 22652 3188
rect 22704 3176 22710 3188
rect 23201 3179 23259 3185
rect 23201 3176 23213 3179
rect 22704 3148 23213 3176
rect 22704 3136 22710 3148
rect 23201 3145 23213 3148
rect 23247 3145 23259 3179
rect 23201 3139 23259 3145
rect 24854 3136 24860 3188
rect 24912 3136 24918 3188
rect 24946 3136 24952 3188
rect 25004 3136 25010 3188
rect 25774 3136 25780 3188
rect 25832 3136 25838 3188
rect 26326 3136 26332 3188
rect 26384 3176 26390 3188
rect 26384 3148 29960 3176
rect 26384 3136 26390 3148
rect 17184 3080 22048 3108
rect 22088 3111 22146 3117
rect 17184 3068 17190 3080
rect 22088 3077 22100 3111
rect 22134 3108 22146 3111
rect 23106 3108 23112 3120
rect 22134 3080 23112 3108
rect 22134 3077 22146 3080
rect 22088 3071 22146 3077
rect 23106 3068 23112 3080
rect 23164 3068 23170 3120
rect 23750 3117 23756 3120
rect 23744 3108 23756 3117
rect 23711 3080 23756 3108
rect 23744 3071 23756 3080
rect 23750 3068 23756 3071
rect 23808 3068 23814 3120
rect 25590 3068 25596 3120
rect 25648 3108 25654 3120
rect 26145 3111 26203 3117
rect 26145 3108 26157 3111
rect 25648 3080 26157 3108
rect 25648 3068 25654 3080
rect 26145 3077 26157 3080
rect 26191 3077 26203 3111
rect 26145 3071 26203 3077
rect 27332 3111 27390 3117
rect 27332 3077 27344 3111
rect 27378 3108 27390 3111
rect 27614 3108 27620 3120
rect 27378 3080 27620 3108
rect 27378 3077 27390 3080
rect 27332 3071 27390 3077
rect 27614 3068 27620 3080
rect 27672 3068 27678 3120
rect 1489 3043 1547 3049
rect 1489 3009 1501 3043
rect 1535 3040 1547 3043
rect 16669 3043 16727 3049
rect 1535 3012 2268 3040
rect 1535 3009 1547 3012
rect 1489 3003 1547 3009
rect 2240 2916 2268 3012
rect 16669 3009 16681 3043
rect 16715 3040 16727 3043
rect 16758 3040 16764 3052
rect 16715 3012 16764 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 16758 3000 16764 3012
rect 16816 3000 16822 3052
rect 16942 3049 16948 3052
rect 16936 3040 16948 3049
rect 16903 3012 16948 3040
rect 16936 3003 16948 3012
rect 16942 3000 16948 3003
rect 17000 3000 17006 3052
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 19794 3049 19800 3052
rect 19521 3043 19579 3049
rect 19521 3040 19533 3043
rect 19392 3012 19533 3040
rect 19392 3000 19398 3012
rect 19521 3009 19533 3012
rect 19567 3009 19579 3043
rect 19788 3040 19800 3049
rect 19755 3012 19800 3040
rect 19521 3003 19579 3009
rect 19788 3003 19800 3012
rect 19794 3000 19800 3003
rect 19852 3000 19858 3052
rect 21818 3000 21824 3052
rect 21876 3040 21882 3052
rect 22388 3040 22508 3044
rect 22756 3040 22876 3044
rect 24210 3040 24216 3052
rect 21876 3016 24216 3040
rect 21876 3012 22416 3016
rect 22480 3012 22784 3016
rect 22848 3012 24216 3016
rect 21876 3000 21882 3012
rect 13630 2932 13636 2984
rect 13688 2972 13694 2984
rect 23492 2981 23520 3012
rect 24210 3000 24216 3012
rect 24268 3000 24274 3052
rect 25130 3000 25136 3052
rect 25188 3000 25194 3052
rect 27065 3043 27123 3049
rect 27065 3009 27077 3043
rect 27111 3040 27123 3043
rect 28626 3040 28632 3052
rect 27111 3012 28632 3040
rect 27111 3009 27123 3012
rect 27065 3003 27123 3009
rect 28626 3000 28632 3012
rect 28684 3040 28690 3052
rect 29178 3049 29184 3052
rect 28905 3043 28963 3049
rect 28905 3040 28917 3043
rect 28684 3012 28917 3040
rect 28684 3000 28690 3012
rect 28905 3009 28917 3012
rect 28951 3009 28963 3043
rect 28905 3003 28963 3009
rect 29172 3003 29184 3049
rect 29178 3000 29184 3003
rect 29236 3000 29242 3052
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 13688 2944 14289 2972
rect 13688 2932 13694 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 23477 2975 23535 2981
rect 23477 2941 23489 2975
rect 23523 2941 23535 2975
rect 23477 2935 23535 2941
rect 25038 2932 25044 2984
rect 25096 2972 25102 2984
rect 26237 2975 26295 2981
rect 26237 2972 26249 2975
rect 25096 2944 26249 2972
rect 25096 2932 25102 2944
rect 26237 2941 26249 2944
rect 26283 2941 26295 2975
rect 26237 2935 26295 2941
rect 26326 2932 26332 2984
rect 26384 2932 26390 2984
rect 2222 2864 2228 2916
rect 2280 2864 2286 2916
rect 29932 2904 29960 3148
rect 30006 3136 30012 3188
rect 30064 3176 30070 3188
rect 30285 3179 30343 3185
rect 30285 3176 30297 3179
rect 30064 3148 30297 3176
rect 30064 3136 30070 3148
rect 30285 3145 30297 3148
rect 30331 3145 30343 3179
rect 30285 3139 30343 3145
rect 31018 3136 31024 3188
rect 31076 3136 31082 3188
rect 31389 3179 31447 3185
rect 31389 3145 31401 3179
rect 31435 3176 31447 3179
rect 31846 3176 31852 3188
rect 31435 3148 31852 3176
rect 31435 3145 31447 3148
rect 31389 3139 31447 3145
rect 31846 3136 31852 3148
rect 31904 3136 31910 3188
rect 33318 3136 33324 3188
rect 33376 3176 33382 3188
rect 33505 3179 33563 3185
rect 33505 3176 33517 3179
rect 33376 3148 33517 3176
rect 33376 3136 33382 3148
rect 33505 3145 33517 3148
rect 33551 3145 33563 3179
rect 33505 3139 33563 3145
rect 34606 3136 34612 3188
rect 34664 3176 34670 3188
rect 34977 3179 35035 3185
rect 34977 3176 34989 3179
rect 34664 3148 34989 3176
rect 34664 3136 34670 3148
rect 34977 3145 34989 3148
rect 35023 3176 35035 3179
rect 35158 3176 35164 3188
rect 35023 3148 35164 3176
rect 35023 3145 35035 3148
rect 34977 3139 35035 3145
rect 35158 3136 35164 3148
rect 35216 3136 35222 3188
rect 45554 3136 45560 3188
rect 45612 3176 45618 3188
rect 46661 3179 46719 3185
rect 46661 3176 46673 3179
rect 45612 3148 46673 3176
rect 45612 3136 45618 3148
rect 46661 3145 46673 3148
rect 46707 3145 46719 3179
rect 46661 3139 46719 3145
rect 30558 3068 30564 3120
rect 30616 3108 30622 3120
rect 31478 3108 31484 3120
rect 30616 3080 31484 3108
rect 30616 3068 30622 3080
rect 31478 3068 31484 3080
rect 31536 3068 31542 3120
rect 31938 3068 31944 3120
rect 31996 3108 32002 3120
rect 32370 3111 32428 3117
rect 32370 3108 32382 3111
rect 31996 3080 32382 3108
rect 31996 3068 32002 3080
rect 32370 3077 32382 3080
rect 32416 3077 32428 3111
rect 32370 3071 32428 3077
rect 32030 3000 32036 3052
rect 32088 3040 32094 3052
rect 32125 3043 32183 3049
rect 32125 3040 32137 3043
rect 32088 3012 32137 3040
rect 32088 3000 32094 3012
rect 32125 3009 32137 3012
rect 32171 3040 32183 3043
rect 32171 3012 33180 3040
rect 32171 3009 32183 3012
rect 32125 3003 32183 3009
rect 31665 2975 31723 2981
rect 31665 2941 31677 2975
rect 31711 2972 31723 2975
rect 31754 2972 31760 2984
rect 31711 2944 31760 2972
rect 31711 2941 31723 2944
rect 31665 2935 31723 2941
rect 31754 2932 31760 2944
rect 31812 2932 31818 2984
rect 33152 2972 33180 3012
rect 33410 3000 33416 3052
rect 33468 3040 33474 3052
rect 33853 3043 33911 3049
rect 33853 3040 33865 3043
rect 33468 3012 33865 3040
rect 33468 3000 33474 3012
rect 33853 3009 33865 3012
rect 33899 3009 33911 3043
rect 33853 3003 33911 3009
rect 46566 3000 46572 3052
rect 46624 3000 46630 3052
rect 33597 2975 33655 2981
rect 33597 2972 33609 2975
rect 33152 2944 33609 2972
rect 33597 2941 33609 2944
rect 33643 2941 33655 2975
rect 33597 2935 33655 2941
rect 28000 2876 28856 2904
rect 29932 2876 32168 2904
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 72 2808 1593 2836
rect 72 2796 78 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 18414 2796 18420 2848
rect 18472 2836 18478 2848
rect 22462 2836 22468 2848
rect 18472 2808 22468 2836
rect 18472 2796 18478 2808
rect 22462 2796 22468 2808
rect 22520 2796 22526 2848
rect 22554 2796 22560 2848
rect 22612 2836 22618 2848
rect 28000 2836 28028 2876
rect 22612 2808 28028 2836
rect 28445 2839 28503 2845
rect 22612 2796 22618 2808
rect 28445 2805 28457 2839
rect 28491 2836 28503 2839
rect 28626 2836 28632 2848
rect 28491 2808 28632 2836
rect 28491 2805 28503 2808
rect 28445 2799 28503 2805
rect 28626 2796 28632 2808
rect 28684 2796 28690 2848
rect 28828 2836 28856 2876
rect 31662 2836 31668 2848
rect 28828 2808 31668 2836
rect 31662 2796 31668 2808
rect 31720 2796 31726 2848
rect 32140 2836 32168 2876
rect 33226 2836 33232 2848
rect 32140 2808 33232 2836
rect 33226 2796 33232 2808
rect 33284 2796 33290 2848
rect 1104 2746 47104 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 47104 2746
rect 1104 2672 47104 2694
rect 5902 2592 5908 2644
rect 5960 2632 5966 2644
rect 6549 2635 6607 2641
rect 6549 2632 6561 2635
rect 5960 2604 6561 2632
rect 5960 2592 5966 2604
rect 6549 2601 6561 2604
rect 6595 2601 6607 2635
rect 6549 2595 6607 2601
rect 14323 2635 14381 2641
rect 14323 2601 14335 2635
rect 14369 2632 14381 2635
rect 23293 2635 23351 2641
rect 14369 2604 22094 2632
rect 14369 2601 14381 2604
rect 14323 2595 14381 2601
rect 2409 2567 2467 2573
rect 2409 2533 2421 2567
rect 2455 2564 2467 2567
rect 2682 2564 2688 2576
rect 2455 2536 2688 2564
rect 2455 2533 2467 2536
rect 2409 2527 2467 2533
rect 2682 2524 2688 2536
rect 2740 2524 2746 2576
rect 10778 2564 10784 2576
rect 4632 2536 10784 2564
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1412 2360 1440 2391
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 4632 2437 4660 2536
rect 10778 2524 10784 2536
rect 10836 2524 10842 2576
rect 13262 2524 13268 2576
rect 13320 2564 13326 2576
rect 22066 2564 22094 2604
rect 23293 2601 23305 2635
rect 23339 2632 23351 2635
rect 36446 2632 36452 2644
rect 23339 2604 36452 2632
rect 23339 2601 23351 2604
rect 23293 2595 23351 2601
rect 36446 2592 36452 2604
rect 36504 2592 36510 2644
rect 38746 2592 38752 2644
rect 38804 2632 38810 2644
rect 39393 2635 39451 2641
rect 39393 2632 39405 2635
rect 38804 2604 39405 2632
rect 38804 2592 38810 2604
rect 39393 2601 39405 2604
rect 39439 2601 39451 2635
rect 39393 2595 39451 2601
rect 37642 2564 37648 2576
rect 13320 2536 21036 2564
rect 22066 2536 37648 2564
rect 13320 2524 13326 2536
rect 9398 2456 9404 2508
rect 9456 2456 9462 2508
rect 20714 2496 20720 2508
rect 14476 2468 20720 2496
rect 2225 2431 2283 2437
rect 2225 2428 2237 2431
rect 2004 2400 2237 2428
rect 2004 2388 2010 2400
rect 2225 2397 2237 2400
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6512 2400 6745 2428
rect 6512 2388 6518 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 11330 2388 11336 2440
rect 11388 2428 11394 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11388 2400 11713 2428
rect 11388 2388 11394 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13596 2400 14105 2428
rect 13596 2388 13602 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 2041 2363 2099 2369
rect 2041 2360 2053 2363
rect 1412 2332 2053 2360
rect 2041 2329 2053 2332
rect 2087 2360 2099 2363
rect 14476 2360 14504 2468
rect 20714 2456 20720 2468
rect 20772 2456 20778 2508
rect 21008 2496 21036 2536
rect 37642 2524 37648 2536
rect 37700 2524 37706 2576
rect 25501 2499 25559 2505
rect 25501 2496 25513 2499
rect 21008 2468 25513 2496
rect 25501 2465 25513 2468
rect 25547 2465 25559 2499
rect 37182 2496 37188 2508
rect 25501 2459 25559 2465
rect 32324 2468 37188 2496
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16172 2400 16681 2428
rect 16172 2388 16178 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 16960 2360 16988 2391
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 18785 2431 18843 2437
rect 18785 2428 18797 2431
rect 18748 2400 18797 2428
rect 18748 2388 18754 2400
rect 18785 2397 18797 2400
rect 18831 2397 18843 2431
rect 18785 2391 18843 2397
rect 20990 2388 20996 2440
rect 21048 2388 21054 2440
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23477 2431 23535 2437
rect 23477 2428 23489 2431
rect 23256 2400 23489 2428
rect 23256 2388 23262 2400
rect 23477 2397 23489 2400
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 25130 2388 25136 2440
rect 25188 2428 25194 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 25188 2400 25237 2428
rect 25188 2388 25194 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 27801 2431 27859 2437
rect 27801 2397 27813 2431
rect 27847 2428 27859 2431
rect 28626 2428 28632 2440
rect 27847 2400 28632 2428
rect 27847 2397 27859 2400
rect 27801 2391 27859 2397
rect 28626 2388 28632 2400
rect 28684 2388 28690 2440
rect 29362 2388 29368 2440
rect 29420 2388 29426 2440
rect 32324 2437 32352 2468
rect 37182 2456 37188 2468
rect 37240 2456 37246 2508
rect 42702 2456 42708 2508
rect 42760 2456 42766 2508
rect 45462 2456 45468 2508
rect 45520 2496 45526 2508
rect 45925 2499 45983 2505
rect 45925 2496 45937 2499
rect 45520 2468 45937 2496
rect 45520 2456 45526 2468
rect 45925 2465 45937 2468
rect 45971 2465 45983 2499
rect 45925 2459 45983 2465
rect 46198 2456 46204 2508
rect 46256 2456 46262 2508
rect 32309 2431 32367 2437
rect 32309 2397 32321 2431
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33597 2431 33655 2437
rect 33597 2397 33609 2431
rect 33643 2428 33655 2431
rect 34698 2428 34704 2440
rect 33643 2400 34704 2428
rect 33643 2397 33655 2400
rect 33597 2391 33655 2397
rect 34698 2388 34704 2400
rect 34756 2388 34762 2440
rect 34882 2388 34888 2440
rect 34940 2388 34946 2440
rect 37458 2388 37464 2440
rect 37516 2388 37522 2440
rect 39298 2388 39304 2440
rect 39356 2428 39362 2440
rect 39577 2431 39635 2437
rect 39577 2428 39589 2431
rect 39356 2400 39589 2428
rect 39356 2388 39362 2400
rect 39577 2397 39589 2400
rect 39623 2397 39635 2431
rect 39577 2391 39635 2397
rect 41874 2388 41880 2440
rect 41932 2428 41938 2440
rect 42429 2431 42487 2437
rect 42429 2428 42441 2431
rect 41932 2400 42441 2428
rect 41932 2388 41938 2400
rect 42429 2397 42441 2400
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 44542 2388 44548 2440
rect 44600 2388 44606 2440
rect 45833 2431 45891 2437
rect 45833 2397 45845 2431
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 2087 2332 14504 2360
rect 16546 2332 16988 2360
rect 2087 2329 2099 2332
rect 2041 2323 2099 2329
rect 934 2252 940 2304
rect 992 2292 998 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 992 2264 1593 2292
rect 992 2252 998 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 4580 2264 4813 2292
rect 4580 2252 4586 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11885 2295 11943 2301
rect 11885 2292 11897 2295
rect 11664 2264 11897 2292
rect 11664 2252 11670 2264
rect 11885 2261 11897 2264
rect 11931 2261 11943 2295
rect 11885 2255 11943 2261
rect 13630 2252 13636 2304
rect 13688 2292 13694 2304
rect 16546 2292 16574 2332
rect 20622 2320 20628 2372
rect 20680 2360 20686 2372
rect 20809 2363 20867 2369
rect 20809 2360 20821 2363
rect 20680 2332 20821 2360
rect 20680 2320 20686 2332
rect 20809 2329 20821 2332
rect 20855 2329 20867 2363
rect 20809 2323 20867 2329
rect 30285 2363 30343 2369
rect 30285 2329 30297 2363
rect 30331 2360 30343 2363
rect 34606 2360 34612 2372
rect 30331 2332 34612 2360
rect 30331 2329 30343 2332
rect 30285 2323 30343 2329
rect 34606 2320 34612 2332
rect 34664 2320 34670 2372
rect 45848 2360 45876 2391
rect 46382 2360 46388 2372
rect 45848 2332 46388 2360
rect 46382 2320 46388 2332
rect 46440 2320 46446 2372
rect 13688 2264 16574 2292
rect 13688 2252 13694 2264
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18969 2295 19027 2301
rect 18969 2292 18981 2295
rect 18748 2264 18981 2292
rect 18748 2252 18754 2264
rect 18969 2261 18981 2264
rect 19015 2261 19027 2295
rect 18969 2255 19027 2261
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 27985 2295 28043 2301
rect 27985 2292 27997 2295
rect 27764 2264 27997 2292
rect 27764 2252 27770 2264
rect 27985 2261 27997 2264
rect 28031 2261 28043 2295
rect 27985 2255 28043 2261
rect 29178 2252 29184 2304
rect 29236 2252 29242 2304
rect 30374 2252 30380 2304
rect 30432 2252 30438 2304
rect 32214 2252 32220 2304
rect 32272 2292 32278 2304
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 32272 2264 32505 2292
rect 32272 2252 32278 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 32493 2255 32551 2261
rect 33410 2252 33416 2304
rect 33468 2252 33474 2304
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34848 2264 35081 2292
rect 34848 2252 34854 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 37366 2252 37372 2304
rect 37424 2292 37430 2304
rect 37645 2295 37703 2301
rect 37645 2292 37657 2295
rect 37424 2264 37657 2292
rect 37424 2252 37430 2264
rect 37645 2261 37657 2264
rect 37691 2261 37703 2295
rect 37645 2255 37703 2261
rect 44450 2252 44456 2304
rect 44508 2292 44514 2304
rect 44729 2295 44787 2301
rect 44729 2292 44741 2295
rect 44508 2264 44741 2292
rect 44508 2252 44514 2264
rect 44729 2261 44741 2264
rect 44775 2261 44787 2295
rect 44729 2255 44787 2261
rect 45646 2252 45652 2304
rect 45704 2252 45710 2304
rect 1104 2202 47104 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 47104 2202
rect 1104 2128 47104 2150
<< via1 >>
rect 6092 48016 6144 48068
rect 32128 48016 32180 48068
rect 4874 47846 4926 47898
rect 4938 47846 4990 47898
rect 5002 47846 5054 47898
rect 5066 47846 5118 47898
rect 5130 47846 5182 47898
rect 35594 47846 35646 47898
rect 35658 47846 35710 47898
rect 35722 47846 35774 47898
rect 35786 47846 35838 47898
rect 35850 47846 35902 47898
rect 1768 47787 1820 47796
rect 1768 47753 1777 47787
rect 1777 47753 1811 47787
rect 1811 47753 1820 47787
rect 1768 47744 1820 47753
rect 3240 47744 3292 47796
rect 6092 47787 6144 47796
rect 6092 47753 6101 47787
rect 6101 47753 6135 47787
rect 6135 47753 6144 47787
rect 6092 47744 6144 47753
rect 10600 47787 10652 47796
rect 10600 47753 10609 47787
rect 10609 47753 10643 47787
rect 10643 47753 10652 47787
rect 10600 47744 10652 47753
rect 13176 47787 13228 47796
rect 13176 47753 13185 47787
rect 13185 47753 13219 47787
rect 13219 47753 13228 47787
rect 13176 47744 13228 47753
rect 15752 47787 15804 47796
rect 15752 47753 15761 47787
rect 15761 47753 15795 47787
rect 15795 47753 15804 47787
rect 15752 47744 15804 47753
rect 17408 47744 17460 47796
rect 6000 47719 6052 47728
rect 6000 47685 6009 47719
rect 6009 47685 6043 47719
rect 6043 47685 6052 47719
rect 6000 47676 6052 47685
rect 2320 47608 2372 47660
rect 3056 47608 3108 47660
rect 8668 47651 8720 47660
rect 8668 47617 8677 47651
rect 8677 47617 8711 47651
rect 8711 47617 8720 47651
rect 8668 47608 8720 47617
rect 10232 47608 10284 47660
rect 15200 47608 15252 47660
rect 17316 47651 17368 47660
rect 17316 47617 17325 47651
rect 17325 47617 17359 47651
rect 17359 47617 17368 47651
rect 17316 47608 17368 47617
rect 19984 47744 20036 47796
rect 22560 47744 22612 47796
rect 29000 47744 29052 47796
rect 31760 47744 31812 47796
rect 34428 47787 34480 47796
rect 34428 47753 34437 47787
rect 34437 47753 34471 47787
rect 34471 47753 34480 47787
rect 34428 47744 34480 47753
rect 36084 47744 36136 47796
rect 41420 47744 41472 47796
rect 19248 47608 19300 47660
rect 20352 47608 20404 47660
rect 23204 47608 23256 47660
rect 24584 47651 24636 47660
rect 24584 47617 24593 47651
rect 24593 47617 24627 47651
rect 24627 47617 24636 47651
rect 24584 47608 24636 47617
rect 24860 47583 24912 47592
rect 24860 47549 24869 47583
rect 24869 47549 24903 47583
rect 24903 47549 24912 47583
rect 24860 47540 24912 47549
rect 27252 47719 27304 47728
rect 27252 47685 27261 47719
rect 27261 47685 27295 47719
rect 27295 47685 27304 47719
rect 27252 47676 27304 47685
rect 28264 47676 28316 47728
rect 38384 47676 38436 47728
rect 27344 47608 27396 47660
rect 32220 47651 32272 47660
rect 32220 47617 32229 47651
rect 32229 47617 32263 47651
rect 32263 47617 32272 47651
rect 32220 47608 32272 47617
rect 34336 47608 34388 47660
rect 36912 47608 36964 47660
rect 38660 47608 38712 47660
rect 32404 47540 32456 47592
rect 36452 47540 36504 47592
rect 43260 47651 43312 47660
rect 43260 47617 43269 47651
rect 43269 47617 43303 47651
rect 43303 47617 43312 47651
rect 43260 47608 43312 47617
rect 45836 47651 45888 47660
rect 45836 47617 45845 47651
rect 45845 47617 45879 47651
rect 45879 47617 45888 47651
rect 45836 47608 45888 47617
rect 45928 47651 45980 47660
rect 45928 47617 45937 47651
rect 45937 47617 45971 47651
rect 45971 47617 45980 47651
rect 45928 47608 45980 47617
rect 42892 47540 42944 47592
rect 46204 47583 46256 47592
rect 46204 47549 46213 47583
rect 46213 47549 46247 47583
rect 46247 47549 46256 47583
rect 46204 47540 46256 47549
rect 18236 47404 18288 47456
rect 19432 47447 19484 47456
rect 19432 47413 19441 47447
rect 19441 47413 19475 47447
rect 19475 47413 19484 47447
rect 19432 47404 19484 47413
rect 27160 47472 27212 47524
rect 27436 47515 27488 47524
rect 27436 47481 27445 47515
rect 27445 47481 27479 47515
rect 27479 47481 27488 47515
rect 27436 47472 27488 47481
rect 31392 47404 31444 47456
rect 31484 47404 31536 47456
rect 33508 47404 33560 47456
rect 38844 47404 38896 47456
rect 45652 47447 45704 47456
rect 45652 47413 45661 47447
rect 45661 47413 45695 47447
rect 45695 47413 45704 47447
rect 45652 47404 45704 47413
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 3056 47243 3108 47252
rect 3056 47209 3065 47243
rect 3065 47209 3099 47243
rect 3099 47209 3108 47243
rect 3056 47200 3108 47209
rect 17316 47200 17368 47252
rect 1124 47132 1176 47184
rect 17868 47064 17920 47116
rect 20260 47064 20312 47116
rect 25688 47200 25740 47252
rect 27344 47200 27396 47252
rect 29184 47200 29236 47252
rect 30104 47200 30156 47252
rect 1952 47039 2004 47048
rect 1952 47005 1961 47039
rect 1961 47005 1995 47039
rect 1995 47005 2004 47039
rect 1952 46996 2004 47005
rect 11336 46996 11388 47048
rect 18236 47039 18288 47048
rect 18236 47005 18245 47039
rect 18245 47005 18279 47039
rect 18279 47005 18288 47039
rect 18236 46996 18288 47005
rect 18420 46996 18472 47048
rect 19248 47039 19300 47048
rect 19248 47005 19257 47039
rect 19257 47005 19291 47039
rect 19291 47005 19300 47039
rect 19248 46996 19300 47005
rect 21364 46996 21416 47048
rect 23480 46996 23532 47048
rect 4804 46860 4856 46912
rect 20352 46928 20404 46980
rect 6000 46903 6052 46912
rect 6000 46869 6009 46903
rect 6009 46869 6043 46903
rect 6043 46869 6052 46903
rect 6000 46860 6052 46869
rect 17132 46903 17184 46912
rect 17132 46869 17141 46903
rect 17141 46869 17175 46903
rect 17175 46869 17184 46903
rect 17132 46860 17184 46869
rect 17500 46903 17552 46912
rect 17500 46869 17509 46903
rect 17509 46869 17543 46903
rect 17543 46869 17552 46903
rect 17500 46860 17552 46869
rect 17592 46903 17644 46912
rect 17592 46869 17601 46903
rect 17601 46869 17635 46903
rect 17635 46869 17644 46903
rect 17592 46860 17644 46869
rect 20904 46903 20956 46912
rect 20904 46869 20913 46903
rect 20913 46869 20947 46903
rect 20947 46869 20956 46903
rect 20904 46860 20956 46869
rect 22376 46928 22428 46980
rect 24400 47039 24452 47048
rect 24400 47005 24409 47039
rect 24409 47005 24443 47039
rect 24443 47005 24452 47039
rect 24400 46996 24452 47005
rect 28264 47107 28316 47116
rect 28264 47073 28273 47107
rect 28273 47073 28307 47107
rect 28307 47073 28316 47107
rect 28264 47064 28316 47073
rect 29828 47132 29880 47184
rect 32220 47200 32272 47252
rect 31944 47132 31996 47184
rect 26700 46996 26752 47048
rect 27068 46996 27120 47048
rect 27896 46996 27948 47048
rect 31392 47064 31444 47116
rect 22928 46860 22980 46912
rect 23204 46860 23256 46912
rect 26148 46971 26200 46980
rect 26148 46937 26182 46971
rect 26182 46937 26200 46971
rect 26148 46928 26200 46937
rect 28356 46928 28408 46980
rect 27068 46860 27120 46912
rect 29276 46903 29328 46912
rect 29276 46869 29285 46903
rect 29285 46869 29319 46903
rect 29319 46869 29328 46903
rect 29276 46860 29328 46869
rect 30104 46996 30156 47048
rect 30288 47039 30340 47048
rect 30288 47005 30297 47039
rect 30297 47005 30331 47039
rect 30331 47005 30340 47039
rect 30288 46996 30340 47005
rect 31484 47039 31536 47048
rect 31484 47005 31493 47039
rect 31493 47005 31527 47039
rect 31527 47005 31536 47039
rect 31484 46996 31536 47005
rect 30012 46971 30064 46980
rect 30012 46937 30021 46971
rect 30021 46937 30055 46971
rect 30055 46937 30064 46971
rect 30012 46928 30064 46937
rect 33324 47064 33376 47116
rect 32220 47039 32272 47048
rect 32220 47005 32229 47039
rect 32229 47005 32263 47039
rect 32263 47005 32272 47039
rect 32220 46996 32272 47005
rect 33508 46928 33560 46980
rect 34980 47039 35032 47048
rect 34980 47005 34989 47039
rect 34989 47005 35023 47039
rect 35023 47005 35032 47039
rect 34980 46996 35032 47005
rect 47676 46996 47728 47048
rect 35440 46928 35492 46980
rect 34796 46903 34848 46912
rect 34796 46869 34805 46903
rect 34805 46869 34839 46903
rect 34839 46869 34848 46903
rect 34796 46860 34848 46869
rect 46572 46903 46624 46912
rect 46572 46869 46581 46903
rect 46581 46869 46615 46903
rect 46615 46869 46624 46903
rect 46572 46860 46624 46869
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 35594 46758 35646 46810
rect 35658 46758 35710 46810
rect 35722 46758 35774 46810
rect 35786 46758 35838 46810
rect 35850 46758 35902 46810
rect 1308 46656 1360 46708
rect 17500 46656 17552 46708
rect 20260 46656 20312 46708
rect 20536 46656 20588 46708
rect 22376 46699 22428 46708
rect 22376 46665 22385 46699
rect 22385 46665 22419 46699
rect 22419 46665 22428 46699
rect 22376 46656 22428 46665
rect 6000 46588 6052 46640
rect 4804 46520 4856 46572
rect 16948 46563 17000 46572
rect 16948 46529 16982 46563
rect 16982 46529 17000 46563
rect 16948 46520 17000 46529
rect 17960 46520 18012 46572
rect 20904 46588 20956 46640
rect 22744 46520 22796 46572
rect 27344 46656 27396 46708
rect 29276 46656 29328 46708
rect 30288 46656 30340 46708
rect 32220 46656 32272 46708
rect 34980 46656 35032 46708
rect 23020 46563 23072 46572
rect 23020 46529 23029 46563
rect 23029 46529 23063 46563
rect 23063 46529 23072 46563
rect 23020 46520 23072 46529
rect 23112 46563 23164 46572
rect 23112 46529 23121 46563
rect 23121 46529 23155 46563
rect 23155 46529 23164 46563
rect 23112 46520 23164 46529
rect 23480 46563 23532 46572
rect 23480 46529 23489 46563
rect 23489 46529 23523 46563
rect 23523 46529 23532 46563
rect 23480 46520 23532 46529
rect 25320 46520 25372 46572
rect 15660 46316 15712 46368
rect 17684 46452 17736 46504
rect 20168 46495 20220 46504
rect 20168 46461 20177 46495
rect 20177 46461 20211 46495
rect 20211 46461 20220 46495
rect 20168 46452 20220 46461
rect 22652 46495 22704 46504
rect 22652 46461 22661 46495
rect 22661 46461 22695 46495
rect 22695 46461 22704 46495
rect 22652 46452 22704 46461
rect 23296 46452 23348 46504
rect 25688 46563 25740 46572
rect 25688 46529 25697 46563
rect 25697 46529 25731 46563
rect 25731 46529 25740 46563
rect 25688 46520 25740 46529
rect 28540 46588 28592 46640
rect 27068 46520 27120 46572
rect 27252 46563 27304 46572
rect 27252 46529 27286 46563
rect 27286 46529 27304 46563
rect 27252 46520 27304 46529
rect 29828 46563 29880 46572
rect 29828 46529 29837 46563
rect 29837 46529 29871 46563
rect 29871 46529 29880 46563
rect 29828 46520 29880 46529
rect 30288 46520 30340 46572
rect 19432 46316 19484 46368
rect 22928 46316 22980 46368
rect 26884 46384 26936 46436
rect 25872 46316 25924 46368
rect 26332 46316 26384 46368
rect 29184 46495 29236 46504
rect 29184 46461 29193 46495
rect 29193 46461 29227 46495
rect 29227 46461 29236 46495
rect 29184 46452 29236 46461
rect 29276 46495 29328 46504
rect 29276 46461 29285 46495
rect 29285 46461 29319 46495
rect 29319 46461 29328 46495
rect 29276 46452 29328 46461
rect 29460 46495 29512 46504
rect 29460 46461 29469 46495
rect 29469 46461 29503 46495
rect 29503 46461 29512 46495
rect 29460 46452 29512 46461
rect 34796 46588 34848 46640
rect 31944 46520 31996 46572
rect 35716 46520 35768 46572
rect 35808 46563 35860 46572
rect 35808 46529 35817 46563
rect 35817 46529 35851 46563
rect 35851 46529 35860 46563
rect 35808 46520 35860 46529
rect 33324 46495 33376 46504
rect 33324 46461 33333 46495
rect 33333 46461 33367 46495
rect 33367 46461 33376 46495
rect 33324 46452 33376 46461
rect 35440 46452 35492 46504
rect 37280 46520 37332 46572
rect 29552 46384 29604 46436
rect 30012 46384 30064 46436
rect 45652 46452 45704 46504
rect 37372 46384 37424 46436
rect 27344 46316 27396 46368
rect 27620 46316 27672 46368
rect 28356 46359 28408 46368
rect 28356 46325 28365 46359
rect 28365 46325 28399 46359
rect 28399 46325 28408 46359
rect 28356 46316 28408 46325
rect 28632 46316 28684 46368
rect 29644 46359 29696 46368
rect 29644 46325 29653 46359
rect 29653 46325 29687 46359
rect 29687 46325 29696 46359
rect 29644 46316 29696 46325
rect 30840 46316 30892 46368
rect 35348 46359 35400 46368
rect 35348 46325 35357 46359
rect 35357 46325 35391 46359
rect 35391 46325 35400 46359
rect 35348 46316 35400 46325
rect 36360 46316 36412 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 16948 46155 17000 46164
rect 16948 46121 16957 46155
rect 16957 46121 16991 46155
rect 16991 46121 17000 46155
rect 16948 46112 17000 46121
rect 21180 46155 21232 46164
rect 21180 46121 21189 46155
rect 21189 46121 21223 46155
rect 21223 46121 21232 46155
rect 21180 46112 21232 46121
rect 21364 46155 21416 46164
rect 21364 46121 21373 46155
rect 21373 46121 21407 46155
rect 21407 46121 21416 46155
rect 21364 46112 21416 46121
rect 22652 46112 22704 46164
rect 25320 46155 25372 46164
rect 25320 46121 25329 46155
rect 25329 46121 25363 46155
rect 25363 46121 25372 46155
rect 25320 46112 25372 46121
rect 26148 46155 26200 46164
rect 26148 46121 26157 46155
rect 26157 46121 26191 46155
rect 26191 46121 26200 46155
rect 26148 46112 26200 46121
rect 27252 46112 27304 46164
rect 27712 46112 27764 46164
rect 28172 46112 28224 46164
rect 18052 46044 18104 46096
rect 17868 45976 17920 46028
rect 19432 45976 19484 46028
rect 17132 45951 17184 45960
rect 17132 45917 17141 45951
rect 17141 45917 17175 45951
rect 17175 45917 17184 45951
rect 17132 45908 17184 45917
rect 17500 45908 17552 45960
rect 17684 45840 17736 45892
rect 20352 45951 20404 45960
rect 20352 45917 20361 45951
rect 20361 45917 20395 45951
rect 20395 45917 20404 45951
rect 20352 45908 20404 45917
rect 20904 45908 20956 45960
rect 15936 45772 15988 45824
rect 17592 45772 17644 45824
rect 19984 45772 20036 45824
rect 20168 45772 20220 45824
rect 20536 45815 20588 45824
rect 20536 45781 20545 45815
rect 20545 45781 20579 45815
rect 20579 45781 20588 45815
rect 20536 45772 20588 45781
rect 22376 45772 22428 45824
rect 22744 46044 22796 46096
rect 23112 46044 23164 46096
rect 23296 46044 23348 46096
rect 22744 45951 22796 45960
rect 22744 45917 22753 45951
rect 22753 45917 22787 45951
rect 22787 45917 22796 45951
rect 22744 45908 22796 45917
rect 23112 45908 23164 45960
rect 23204 45951 23256 45960
rect 23204 45917 23213 45951
rect 23213 45917 23247 45951
rect 23247 45917 23256 45951
rect 23204 45908 23256 45917
rect 23296 45951 23348 45960
rect 23296 45917 23305 45951
rect 23305 45917 23339 45951
rect 23339 45917 23348 45951
rect 23296 45908 23348 45917
rect 23572 45976 23624 46028
rect 24400 45951 24452 45960
rect 24400 45917 24409 45951
rect 24409 45917 24443 45951
rect 24443 45917 24452 45951
rect 24400 45908 24452 45917
rect 25596 45951 25648 45960
rect 25596 45917 25605 45951
rect 25605 45917 25639 45951
rect 25639 45917 25648 45951
rect 25596 45908 25648 45917
rect 25780 45951 25832 45960
rect 25780 45917 25789 45951
rect 25789 45917 25823 45951
rect 25823 45917 25832 45951
rect 25780 45908 25832 45917
rect 25964 45951 26016 45960
rect 25964 45917 25973 45951
rect 25973 45917 26007 45951
rect 26007 45917 26016 45951
rect 25964 45908 26016 45917
rect 28264 45976 28316 46028
rect 29276 45976 29328 46028
rect 30288 46112 30340 46164
rect 29460 46044 29512 46096
rect 33232 45976 33284 46028
rect 35440 45976 35492 46028
rect 35716 45976 35768 46028
rect 26332 45951 26384 45960
rect 26332 45917 26341 45951
rect 26341 45917 26375 45951
rect 26375 45917 26384 45951
rect 26332 45908 26384 45917
rect 27160 45908 27212 45960
rect 27528 45951 27580 45960
rect 27528 45917 27537 45951
rect 27537 45917 27571 45951
rect 27571 45917 27580 45951
rect 27528 45908 27580 45917
rect 27620 45951 27672 45960
rect 27620 45917 27629 45951
rect 27629 45917 27663 45951
rect 27663 45917 27672 45951
rect 27620 45908 27672 45917
rect 27988 45951 28040 45960
rect 27988 45917 27997 45951
rect 27997 45917 28031 45951
rect 28031 45917 28040 45951
rect 27988 45908 28040 45917
rect 29184 45908 29236 45960
rect 30472 45908 30524 45960
rect 30564 45951 30616 45960
rect 30564 45917 30573 45951
rect 30573 45917 30607 45951
rect 30607 45917 30616 45951
rect 30564 45908 30616 45917
rect 28356 45840 28408 45892
rect 30840 45951 30892 45960
rect 30840 45917 30849 45951
rect 30849 45917 30883 45951
rect 30883 45917 30892 45951
rect 30840 45908 30892 45917
rect 22928 45772 22980 45824
rect 27620 45772 27672 45824
rect 29552 45772 29604 45824
rect 30380 45772 30432 45824
rect 30656 45772 30708 45824
rect 33140 45840 33192 45892
rect 33692 45951 33744 45960
rect 33692 45917 33701 45951
rect 33701 45917 33735 45951
rect 33735 45917 33744 45951
rect 33692 45908 33744 45917
rect 34796 45951 34848 45960
rect 34796 45917 34805 45951
rect 34805 45917 34839 45951
rect 34839 45917 34848 45951
rect 34796 45908 34848 45917
rect 35348 45908 35400 45960
rect 36360 45951 36412 45960
rect 36360 45917 36394 45951
rect 36394 45917 36412 45951
rect 36360 45908 36412 45917
rect 33416 45815 33468 45824
rect 33416 45781 33425 45815
rect 33425 45781 33459 45815
rect 33459 45781 33468 45815
rect 33416 45772 33468 45781
rect 33692 45815 33744 45824
rect 33692 45781 33701 45815
rect 33701 45781 33735 45815
rect 33735 45781 33744 45815
rect 33692 45772 33744 45781
rect 34428 45772 34480 45824
rect 35808 45772 35860 45824
rect 36728 45772 36780 45824
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 35594 45670 35646 45722
rect 35658 45670 35710 45722
rect 35722 45670 35774 45722
rect 35786 45670 35838 45722
rect 35850 45670 35902 45722
rect 20904 45568 20956 45620
rect 25964 45568 26016 45620
rect 27988 45568 28040 45620
rect 28632 45568 28684 45620
rect 28816 45568 28868 45620
rect 22376 45500 22428 45552
rect 22836 45500 22888 45552
rect 23296 45500 23348 45552
rect 16856 45432 16908 45484
rect 17868 45432 17920 45484
rect 18052 45475 18104 45484
rect 18052 45441 18061 45475
rect 18061 45441 18095 45475
rect 18095 45441 18104 45475
rect 18052 45432 18104 45441
rect 19984 45475 20036 45484
rect 19984 45441 19993 45475
rect 19993 45441 20027 45475
rect 20027 45441 20036 45475
rect 19984 45432 20036 45441
rect 20168 45475 20220 45484
rect 20168 45441 20177 45475
rect 20177 45441 20211 45475
rect 20211 45441 20220 45475
rect 20168 45432 20220 45441
rect 17132 45407 17184 45416
rect 17132 45373 17141 45407
rect 17141 45373 17175 45407
rect 17175 45373 17184 45407
rect 17132 45364 17184 45373
rect 17316 45407 17368 45416
rect 17316 45373 17325 45407
rect 17325 45373 17359 45407
rect 17359 45373 17368 45407
rect 17316 45364 17368 45373
rect 28724 45475 28776 45484
rect 28724 45441 28733 45475
rect 28733 45441 28767 45475
rect 28767 45441 28776 45475
rect 28724 45432 28776 45441
rect 28908 45432 28960 45484
rect 29644 45500 29696 45552
rect 29276 45432 29328 45484
rect 29368 45407 29420 45416
rect 29368 45373 29377 45407
rect 29377 45373 29411 45407
rect 29411 45373 29420 45407
rect 29368 45364 29420 45373
rect 29460 45407 29512 45416
rect 29460 45373 29469 45407
rect 29469 45373 29503 45407
rect 29503 45373 29512 45407
rect 29460 45364 29512 45373
rect 30564 45568 30616 45620
rect 33140 45568 33192 45620
rect 33692 45568 33744 45620
rect 38108 45568 38160 45620
rect 33416 45543 33468 45552
rect 17960 45296 18012 45348
rect 29092 45296 29144 45348
rect 30380 45407 30432 45416
rect 30380 45373 30389 45407
rect 30389 45373 30423 45407
rect 30423 45373 30432 45407
rect 30380 45364 30432 45373
rect 30564 45364 30616 45416
rect 29736 45296 29788 45348
rect 31116 45432 31168 45484
rect 32588 45432 32640 45484
rect 33416 45509 33425 45543
rect 33425 45509 33459 45543
rect 33459 45509 33468 45543
rect 33416 45500 33468 45509
rect 32956 45475 33008 45484
rect 32956 45441 32965 45475
rect 32965 45441 32999 45475
rect 32999 45441 33008 45475
rect 32956 45432 33008 45441
rect 34796 45500 34848 45552
rect 36728 45543 36780 45552
rect 36728 45509 36737 45543
rect 36737 45509 36771 45543
rect 36771 45509 36780 45543
rect 36728 45500 36780 45509
rect 37372 45500 37424 45552
rect 46756 45475 46808 45484
rect 46756 45441 46765 45475
rect 46765 45441 46799 45475
rect 46799 45441 46808 45475
rect 46756 45432 46808 45441
rect 37280 45339 37332 45348
rect 37280 45305 37289 45339
rect 37289 45305 37323 45339
rect 37323 45305 37332 45339
rect 37280 45296 37332 45305
rect 15568 45228 15620 45280
rect 21364 45228 21416 45280
rect 28264 45228 28316 45280
rect 29184 45228 29236 45280
rect 29460 45228 29512 45280
rect 30564 45228 30616 45280
rect 31024 45228 31076 45280
rect 31576 45271 31628 45280
rect 31576 45237 31585 45271
rect 31585 45237 31619 45271
rect 31619 45237 31628 45271
rect 31576 45228 31628 45237
rect 32312 45228 32364 45280
rect 33968 45271 34020 45280
rect 33968 45237 33977 45271
rect 33977 45237 34011 45271
rect 34011 45237 34020 45271
rect 33968 45228 34020 45237
rect 38108 45228 38160 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 17132 45024 17184 45076
rect 16856 44956 16908 45008
rect 20628 45024 20680 45076
rect 21180 45024 21232 45076
rect 22744 45024 22796 45076
rect 25780 45024 25832 45076
rect 27712 45024 27764 45076
rect 27988 45024 28040 45076
rect 16580 44888 16632 44940
rect 17316 44888 17368 44940
rect 20720 44956 20772 45008
rect 20904 44999 20956 45008
rect 20904 44965 20913 44999
rect 20913 44965 20947 44999
rect 20947 44965 20956 44999
rect 20904 44956 20956 44965
rect 21272 44956 21324 45008
rect 13728 44820 13780 44872
rect 15660 44820 15712 44872
rect 16856 44863 16908 44872
rect 16856 44829 16865 44863
rect 16865 44829 16899 44863
rect 16899 44829 16908 44863
rect 16856 44820 16908 44829
rect 22652 44888 22704 44940
rect 15384 44752 15436 44804
rect 16488 44727 16540 44736
rect 16488 44693 16497 44727
rect 16497 44693 16531 44727
rect 16531 44693 16540 44727
rect 16488 44684 16540 44693
rect 20628 44863 20680 44872
rect 20628 44829 20642 44863
rect 20642 44829 20676 44863
rect 20676 44829 20680 44863
rect 20628 44820 20680 44829
rect 21180 44863 21232 44872
rect 21180 44829 21189 44863
rect 21189 44829 21223 44863
rect 21223 44829 21232 44863
rect 21180 44820 21232 44829
rect 20536 44795 20588 44804
rect 20536 44761 20545 44795
rect 20545 44761 20579 44795
rect 20579 44761 20588 44795
rect 20536 44752 20588 44761
rect 21088 44752 21140 44804
rect 21364 44863 21416 44872
rect 21364 44829 21373 44863
rect 21373 44829 21407 44863
rect 21407 44829 21416 44863
rect 21364 44820 21416 44829
rect 21548 44863 21600 44872
rect 21548 44829 21557 44863
rect 21557 44829 21591 44863
rect 21591 44829 21600 44863
rect 21548 44820 21600 44829
rect 22192 44863 22244 44872
rect 22192 44829 22201 44863
rect 22201 44829 22235 44863
rect 22235 44829 22244 44863
rect 22192 44820 22244 44829
rect 22284 44863 22336 44872
rect 22284 44829 22293 44863
rect 22293 44829 22327 44863
rect 22327 44829 22336 44863
rect 22284 44820 22336 44829
rect 22560 44820 22612 44872
rect 23204 44888 23256 44940
rect 23296 44888 23348 44940
rect 28632 44999 28684 45008
rect 28632 44965 28641 44999
rect 28641 44965 28675 44999
rect 28675 44965 28684 44999
rect 28632 44956 28684 44965
rect 26700 44931 26752 44940
rect 26700 44897 26709 44931
rect 26709 44897 26743 44931
rect 26743 44897 26752 44931
rect 26700 44888 26752 44897
rect 28448 44888 28500 44940
rect 28908 45024 28960 45076
rect 29368 45024 29420 45076
rect 30472 45024 30524 45076
rect 31024 45067 31076 45076
rect 31024 45033 31033 45067
rect 31033 45033 31067 45067
rect 31067 45033 31076 45067
rect 31024 45024 31076 45033
rect 31116 45067 31168 45076
rect 31116 45033 31125 45067
rect 31125 45033 31159 45067
rect 31159 45033 31168 45067
rect 31116 45024 31168 45033
rect 29000 44956 29052 45008
rect 29828 44956 29880 45008
rect 31576 44956 31628 45008
rect 32588 45024 32640 45076
rect 34796 44956 34848 45008
rect 32680 44931 32732 44940
rect 32680 44897 32689 44931
rect 32689 44897 32723 44931
rect 32723 44897 32732 44931
rect 32680 44888 32732 44897
rect 33968 44888 34020 44940
rect 23112 44863 23164 44872
rect 23112 44829 23121 44863
rect 23121 44829 23155 44863
rect 23155 44829 23164 44863
rect 23112 44820 23164 44829
rect 25320 44795 25372 44804
rect 25320 44761 25329 44795
rect 25329 44761 25363 44795
rect 25363 44761 25372 44795
rect 25320 44752 25372 44761
rect 25596 44820 25648 44872
rect 25780 44863 25832 44872
rect 25780 44829 25789 44863
rect 25789 44829 25823 44863
rect 25823 44829 25832 44863
rect 25780 44820 25832 44829
rect 26608 44863 26660 44872
rect 26608 44829 26617 44863
rect 26617 44829 26651 44863
rect 26651 44829 26660 44863
rect 26608 44820 26660 44829
rect 26792 44863 26844 44872
rect 26792 44829 26801 44863
rect 26801 44829 26835 44863
rect 26835 44829 26844 44863
rect 26792 44820 26844 44829
rect 26424 44795 26476 44804
rect 26424 44761 26433 44795
rect 26433 44761 26467 44795
rect 26467 44761 26476 44795
rect 26424 44752 26476 44761
rect 27804 44863 27856 44872
rect 27804 44829 27813 44863
rect 27813 44829 27847 44863
rect 27847 44829 27856 44863
rect 27804 44820 27856 44829
rect 27988 44795 28040 44804
rect 27988 44761 27997 44795
rect 27997 44761 28031 44795
rect 28031 44761 28040 44795
rect 27988 44752 28040 44761
rect 28264 44752 28316 44804
rect 28632 44820 28684 44872
rect 28816 44820 28868 44872
rect 29184 44863 29236 44872
rect 29184 44829 29193 44863
rect 29193 44829 29227 44863
rect 29227 44829 29236 44863
rect 29184 44820 29236 44829
rect 29368 44863 29420 44872
rect 29368 44829 29377 44863
rect 29377 44829 29411 44863
rect 29411 44829 29420 44863
rect 29368 44820 29420 44829
rect 29460 44752 29512 44804
rect 20352 44684 20404 44736
rect 21824 44727 21876 44736
rect 21824 44693 21833 44727
rect 21833 44693 21867 44727
rect 21867 44693 21876 44727
rect 21824 44684 21876 44693
rect 25688 44684 25740 44736
rect 27712 44727 27764 44736
rect 27712 44693 27721 44727
rect 27721 44693 27755 44727
rect 27755 44693 27764 44727
rect 27712 44684 27764 44693
rect 28632 44727 28684 44736
rect 28632 44693 28641 44727
rect 28641 44693 28675 44727
rect 28675 44693 28684 44727
rect 28632 44684 28684 44693
rect 29092 44684 29144 44736
rect 29276 44727 29328 44736
rect 29276 44693 29285 44727
rect 29285 44693 29319 44727
rect 29319 44693 29328 44727
rect 29276 44684 29328 44693
rect 29920 44684 29972 44736
rect 30472 44820 30524 44872
rect 30564 44863 30616 44872
rect 30564 44829 30573 44863
rect 30573 44829 30607 44863
rect 30607 44829 30616 44863
rect 30564 44820 30616 44829
rect 31300 44863 31352 44872
rect 31300 44829 31309 44863
rect 31309 44829 31343 44863
rect 31343 44829 31352 44863
rect 31300 44820 31352 44829
rect 31668 44820 31720 44872
rect 30104 44752 30156 44804
rect 32312 44863 32364 44872
rect 32312 44829 32321 44863
rect 32321 44829 32355 44863
rect 32355 44829 32364 44863
rect 32312 44820 32364 44829
rect 32956 44820 33008 44872
rect 38844 44863 38896 44872
rect 38844 44829 38853 44863
rect 38853 44829 38887 44863
rect 38887 44829 38896 44863
rect 38844 44820 38896 44829
rect 33324 44752 33376 44804
rect 31300 44684 31352 44736
rect 38292 44684 38344 44736
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 35594 44582 35646 44634
rect 35658 44582 35710 44634
rect 35722 44582 35774 44634
rect 35786 44582 35838 44634
rect 35850 44582 35902 44634
rect 15384 44523 15436 44532
rect 15384 44489 15393 44523
rect 15393 44489 15427 44523
rect 15427 44489 15436 44523
rect 15384 44480 15436 44489
rect 2688 44412 2740 44464
rect 20352 44480 20404 44532
rect 21548 44480 21600 44532
rect 22284 44480 22336 44532
rect 29276 44480 29328 44532
rect 29460 44480 29512 44532
rect 31760 44480 31812 44532
rect 32956 44480 33008 44532
rect 33232 44480 33284 44532
rect 34244 44480 34296 44532
rect 36452 44480 36504 44532
rect 37372 44480 37424 44532
rect 38384 44523 38436 44532
rect 38384 44489 38393 44523
rect 38393 44489 38427 44523
rect 38427 44489 38436 44523
rect 38384 44480 38436 44489
rect 1400 44387 1452 44396
rect 1400 44353 1409 44387
rect 1409 44353 1443 44387
rect 1443 44353 1452 44387
rect 1400 44344 1452 44353
rect 15568 44387 15620 44396
rect 15568 44353 15577 44387
rect 15577 44353 15611 44387
rect 15611 44353 15620 44387
rect 15568 44344 15620 44353
rect 16488 44344 16540 44396
rect 19708 44387 19760 44396
rect 19708 44353 19717 44387
rect 19717 44353 19751 44387
rect 19751 44353 19760 44387
rect 19708 44344 19760 44353
rect 20168 44344 20220 44396
rect 21824 44412 21876 44464
rect 22744 44412 22796 44464
rect 23020 44455 23072 44464
rect 23020 44421 23029 44455
rect 23029 44421 23063 44455
rect 23063 44421 23072 44455
rect 23020 44412 23072 44421
rect 20720 44344 20772 44396
rect 21088 44344 21140 44396
rect 22192 44344 22244 44396
rect 22836 44344 22888 44396
rect 940 44208 992 44260
rect 17040 44140 17092 44192
rect 22100 44251 22152 44260
rect 22100 44217 22109 44251
rect 22109 44217 22143 44251
rect 22143 44217 22152 44251
rect 22100 44208 22152 44217
rect 22284 44208 22336 44260
rect 22652 44251 22704 44260
rect 22652 44217 22661 44251
rect 22661 44217 22695 44251
rect 22695 44217 22704 44251
rect 25320 44412 25372 44464
rect 25412 44387 25464 44396
rect 25412 44353 25421 44387
rect 25421 44353 25455 44387
rect 25455 44353 25464 44387
rect 25412 44344 25464 44353
rect 25688 44344 25740 44396
rect 26424 44344 26476 44396
rect 26976 44344 27028 44396
rect 29368 44412 29420 44464
rect 27804 44344 27856 44396
rect 29000 44344 29052 44396
rect 29092 44344 29144 44396
rect 30104 44412 30156 44464
rect 35348 44412 35400 44464
rect 35440 44412 35492 44464
rect 38844 44455 38896 44464
rect 38844 44421 38853 44455
rect 38853 44421 38887 44455
rect 38887 44421 38896 44455
rect 38844 44412 38896 44421
rect 26516 44276 26568 44328
rect 28908 44276 28960 44328
rect 30288 44344 30340 44396
rect 33324 44344 33376 44396
rect 34796 44344 34848 44396
rect 37280 44387 37332 44396
rect 37280 44353 37289 44387
rect 37289 44353 37323 44387
rect 37323 44353 37332 44387
rect 37280 44344 37332 44353
rect 38292 44387 38344 44396
rect 38292 44353 38301 44387
rect 38301 44353 38335 44387
rect 38335 44353 38344 44387
rect 38292 44344 38344 44353
rect 38476 44344 38528 44396
rect 22652 44208 22704 44217
rect 26424 44208 26476 44260
rect 17776 44140 17828 44192
rect 19984 44140 20036 44192
rect 20536 44140 20588 44192
rect 23296 44140 23348 44192
rect 23388 44183 23440 44192
rect 23388 44149 23397 44183
rect 23397 44149 23431 44183
rect 23431 44149 23440 44183
rect 23388 44140 23440 44149
rect 25964 44140 26016 44192
rect 28724 44208 28776 44260
rect 29736 44276 29788 44328
rect 29920 44276 29972 44328
rect 31300 44276 31352 44328
rect 34520 44276 34572 44328
rect 27988 44140 28040 44192
rect 28080 44140 28132 44192
rect 29092 44140 29144 44192
rect 29828 44183 29880 44192
rect 29828 44149 29837 44183
rect 29837 44149 29871 44183
rect 29871 44149 29880 44183
rect 29828 44140 29880 44149
rect 32404 44140 32456 44192
rect 38384 44276 38436 44328
rect 39028 44276 39080 44328
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 4620 43936 4672 43988
rect 15936 43868 15988 43920
rect 19708 43936 19760 43988
rect 21272 43936 21324 43988
rect 23020 43936 23072 43988
rect 23112 43936 23164 43988
rect 17960 43868 18012 43920
rect 19156 43868 19208 43920
rect 21364 43868 21416 43920
rect 22652 43868 22704 43920
rect 22836 43868 22888 43920
rect 3240 43664 3292 43716
rect 15476 43732 15528 43784
rect 16764 43732 16816 43784
rect 16948 43775 17000 43784
rect 16948 43741 16957 43775
rect 16957 43741 16991 43775
rect 16991 43741 17000 43775
rect 16948 43732 17000 43741
rect 19064 43775 19116 43784
rect 19064 43741 19073 43775
rect 19073 43741 19107 43775
rect 19107 43741 19116 43775
rect 25780 43936 25832 43988
rect 24308 43868 24360 43920
rect 19064 43732 19116 43741
rect 20536 43775 20588 43784
rect 4620 43664 4672 43716
rect 20536 43741 20570 43775
rect 20570 43741 20588 43775
rect 20536 43732 20588 43741
rect 22100 43732 22152 43784
rect 22192 43775 22244 43784
rect 22192 43741 22201 43775
rect 22201 43741 22235 43775
rect 22235 43741 22244 43775
rect 22192 43732 22244 43741
rect 16028 43596 16080 43648
rect 16580 43596 16632 43648
rect 21180 43664 21232 43716
rect 21732 43664 21784 43716
rect 18328 43639 18380 43648
rect 18328 43605 18337 43639
rect 18337 43605 18371 43639
rect 18371 43605 18380 43639
rect 18328 43596 18380 43605
rect 19064 43596 19116 43648
rect 20628 43596 20680 43648
rect 21824 43596 21876 43648
rect 22192 43596 22244 43648
rect 22560 43664 22612 43716
rect 22744 43732 22796 43784
rect 23480 43732 23532 43784
rect 24216 43732 24268 43784
rect 30196 43868 30248 43920
rect 26424 43775 26476 43784
rect 26424 43741 26433 43775
rect 26433 43741 26467 43775
rect 26467 43741 26476 43775
rect 26424 43732 26476 43741
rect 25504 43664 25556 43716
rect 26240 43707 26292 43716
rect 26240 43673 26249 43707
rect 26249 43673 26283 43707
rect 26283 43673 26292 43707
rect 26240 43664 26292 43673
rect 27988 43800 28040 43852
rect 28172 43843 28224 43852
rect 28172 43809 28181 43843
rect 28181 43809 28215 43843
rect 28215 43809 28224 43843
rect 28172 43800 28224 43809
rect 28264 43843 28316 43852
rect 28264 43809 28273 43843
rect 28273 43809 28307 43843
rect 28307 43809 28316 43843
rect 28264 43800 28316 43809
rect 26976 43775 27028 43784
rect 26976 43741 26985 43775
rect 26985 43741 27019 43775
rect 27019 43741 27028 43775
rect 26976 43732 27028 43741
rect 27160 43775 27212 43784
rect 27160 43741 27169 43775
rect 27169 43741 27203 43775
rect 27203 43741 27212 43775
rect 27160 43732 27212 43741
rect 28080 43769 28132 43784
rect 28080 43735 28089 43769
rect 28089 43735 28123 43769
rect 28123 43735 28132 43769
rect 28080 43732 28132 43735
rect 28356 43775 28408 43784
rect 28356 43741 28365 43775
rect 28365 43741 28399 43775
rect 28399 43741 28408 43775
rect 28356 43732 28408 43741
rect 29828 43843 29880 43852
rect 29828 43809 29837 43843
rect 29837 43809 29871 43843
rect 29871 43809 29880 43843
rect 29828 43800 29880 43809
rect 29920 43843 29972 43852
rect 29920 43809 29929 43843
rect 29929 43809 29963 43843
rect 29963 43809 29972 43843
rect 29920 43800 29972 43809
rect 30012 43843 30064 43852
rect 30012 43809 30021 43843
rect 30021 43809 30055 43843
rect 30055 43809 30064 43843
rect 30012 43800 30064 43809
rect 28632 43732 28684 43784
rect 29092 43775 29144 43784
rect 29092 43741 29101 43775
rect 29101 43741 29135 43775
rect 29135 43741 29144 43775
rect 29092 43732 29144 43741
rect 29184 43775 29236 43784
rect 29184 43741 29193 43775
rect 29193 43741 29227 43775
rect 29227 43741 29236 43775
rect 29184 43732 29236 43741
rect 30472 43732 30524 43784
rect 33324 43936 33376 43988
rect 35348 43936 35400 43988
rect 34888 43868 34940 43920
rect 36452 43936 36504 43988
rect 37280 43936 37332 43988
rect 32036 43732 32088 43784
rect 35992 43800 36044 43852
rect 35348 43775 35400 43784
rect 35348 43741 35357 43775
rect 35357 43741 35391 43775
rect 35391 43741 35400 43775
rect 35348 43732 35400 43741
rect 22652 43596 22704 43648
rect 27712 43664 27764 43716
rect 26700 43596 26752 43648
rect 26792 43639 26844 43648
rect 26792 43605 26801 43639
rect 26801 43605 26835 43639
rect 26835 43605 26844 43639
rect 26792 43596 26844 43605
rect 27620 43596 27672 43648
rect 27988 43596 28040 43648
rect 30840 43664 30892 43716
rect 33600 43664 33652 43716
rect 34704 43664 34756 43716
rect 35440 43664 35492 43716
rect 37280 43732 37332 43784
rect 38844 43936 38896 43988
rect 35992 43664 36044 43716
rect 37832 43707 37884 43716
rect 37832 43673 37841 43707
rect 37841 43673 37875 43707
rect 37875 43673 37884 43707
rect 46572 43732 46624 43784
rect 37832 43664 37884 43673
rect 38752 43664 38804 43716
rect 29000 43596 29052 43648
rect 29092 43596 29144 43648
rect 30380 43596 30432 43648
rect 30748 43596 30800 43648
rect 38108 43596 38160 43648
rect 39212 43596 39264 43648
rect 39856 43639 39908 43648
rect 39856 43605 39865 43639
rect 39865 43605 39899 43639
rect 39899 43605 39908 43639
rect 39856 43596 39908 43605
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 35594 43494 35646 43546
rect 35658 43494 35710 43546
rect 35722 43494 35774 43546
rect 35786 43494 35838 43546
rect 35850 43494 35902 43546
rect 15200 43392 15252 43444
rect 16764 43392 16816 43444
rect 21732 43392 21784 43444
rect 17040 43324 17092 43376
rect 19708 43324 19760 43376
rect 20168 43324 20220 43376
rect 22100 43392 22152 43444
rect 15108 43256 15160 43308
rect 16580 43256 16632 43308
rect 17316 43256 17368 43308
rect 13728 43231 13780 43240
rect 13728 43197 13737 43231
rect 13737 43197 13771 43231
rect 13771 43197 13780 43231
rect 13728 43188 13780 43197
rect 18328 43256 18380 43308
rect 19616 43256 19668 43308
rect 20352 43299 20404 43308
rect 20352 43265 20361 43299
rect 20361 43265 20395 43299
rect 20395 43265 20404 43299
rect 20352 43256 20404 43265
rect 21916 43324 21968 43376
rect 25504 43435 25556 43444
rect 25504 43401 25513 43435
rect 25513 43401 25547 43435
rect 25547 43401 25556 43435
rect 25504 43392 25556 43401
rect 26240 43392 26292 43444
rect 26608 43392 26660 43444
rect 21272 43256 21324 43308
rect 21364 43299 21416 43308
rect 21364 43265 21373 43299
rect 21373 43265 21407 43299
rect 21407 43265 21416 43299
rect 21364 43256 21416 43265
rect 21456 43299 21508 43308
rect 21456 43265 21465 43299
rect 21465 43265 21499 43299
rect 21499 43265 21508 43299
rect 21456 43256 21508 43265
rect 21916 43231 21968 43240
rect 21916 43197 21925 43231
rect 21925 43197 21959 43231
rect 21959 43197 21968 43231
rect 21916 43188 21968 43197
rect 22284 43256 22336 43308
rect 22560 43256 22612 43308
rect 25596 43256 25648 43308
rect 26792 43324 26844 43376
rect 26884 43324 26936 43376
rect 25964 43299 26016 43308
rect 25964 43265 25973 43299
rect 25973 43265 26007 43299
rect 26007 43265 26016 43299
rect 25964 43256 26016 43265
rect 26056 43299 26108 43308
rect 26056 43265 26065 43299
rect 26065 43265 26099 43299
rect 26099 43265 26108 43299
rect 26056 43256 26108 43265
rect 26516 43256 26568 43308
rect 26700 43256 26752 43308
rect 28172 43324 28224 43376
rect 27252 43299 27304 43308
rect 27252 43265 27261 43299
rect 27261 43265 27295 43299
rect 27295 43265 27304 43299
rect 27252 43256 27304 43265
rect 30288 43392 30340 43444
rect 30380 43435 30432 43444
rect 30380 43401 30389 43435
rect 30389 43401 30423 43435
rect 30423 43401 30432 43435
rect 30380 43392 30432 43401
rect 30656 43435 30708 43444
rect 30656 43401 30665 43435
rect 30665 43401 30699 43435
rect 30699 43401 30708 43435
rect 30656 43392 30708 43401
rect 34796 43435 34848 43444
rect 34796 43401 34805 43435
rect 34805 43401 34839 43435
rect 34839 43401 34848 43435
rect 34796 43392 34848 43401
rect 34888 43392 34940 43444
rect 29552 43324 29604 43376
rect 30840 43324 30892 43376
rect 35992 43392 36044 43444
rect 36084 43392 36136 43444
rect 37372 43392 37424 43444
rect 37648 43435 37700 43444
rect 37648 43401 37657 43435
rect 37657 43401 37691 43435
rect 37691 43401 37700 43435
rect 37648 43392 37700 43401
rect 38568 43392 38620 43444
rect 38752 43435 38804 43444
rect 38752 43401 38761 43435
rect 38761 43401 38795 43435
rect 38795 43401 38804 43435
rect 38752 43392 38804 43401
rect 40408 43435 40460 43444
rect 40408 43401 40417 43435
rect 40417 43401 40451 43435
rect 40451 43401 40460 43435
rect 40408 43392 40460 43401
rect 29736 43299 29788 43308
rect 29736 43265 29745 43299
rect 29745 43265 29779 43299
rect 29779 43265 29788 43299
rect 29736 43256 29788 43265
rect 22192 43188 22244 43240
rect 22744 43231 22796 43240
rect 22744 43197 22753 43231
rect 22753 43197 22787 43231
rect 22787 43197 22796 43231
rect 22744 43188 22796 43197
rect 21088 43163 21140 43172
rect 21088 43129 21097 43163
rect 21097 43129 21131 43163
rect 21131 43129 21140 43163
rect 21088 43120 21140 43129
rect 18052 43095 18104 43104
rect 18052 43061 18061 43095
rect 18061 43061 18095 43095
rect 18095 43061 18104 43095
rect 18052 43052 18104 43061
rect 21824 43095 21876 43104
rect 21824 43061 21833 43095
rect 21833 43061 21867 43095
rect 21867 43061 21876 43095
rect 21824 43052 21876 43061
rect 29552 43188 29604 43240
rect 29920 43256 29972 43308
rect 30104 43299 30156 43308
rect 30104 43265 30113 43299
rect 30113 43265 30147 43299
rect 30147 43265 30156 43299
rect 30104 43256 30156 43265
rect 30748 43299 30800 43308
rect 30748 43265 30757 43299
rect 30757 43265 30791 43299
rect 30791 43265 30800 43299
rect 30748 43256 30800 43265
rect 32036 43256 32088 43308
rect 33416 43299 33468 43308
rect 33416 43265 33425 43299
rect 33425 43265 33459 43299
rect 33459 43265 33468 43299
rect 33416 43256 33468 43265
rect 34704 43256 34756 43308
rect 35072 43299 35124 43308
rect 35072 43265 35081 43299
rect 35081 43265 35115 43299
rect 35115 43265 35124 43299
rect 35072 43256 35124 43265
rect 30012 43120 30064 43172
rect 27068 43095 27120 43104
rect 27068 43061 27077 43095
rect 27077 43061 27111 43095
rect 27111 43061 27120 43095
rect 27068 43052 27120 43061
rect 28540 43052 28592 43104
rect 34520 43188 34572 43240
rect 34612 43120 34664 43172
rect 35440 43299 35492 43308
rect 35440 43265 35449 43299
rect 35449 43265 35483 43299
rect 35483 43265 35492 43299
rect 35440 43256 35492 43265
rect 35992 43299 36044 43308
rect 35992 43265 36001 43299
rect 36001 43265 36035 43299
rect 36035 43265 36044 43299
rect 35992 43256 36044 43265
rect 35532 43188 35584 43240
rect 36268 43256 36320 43308
rect 37372 43256 37424 43308
rect 39856 43324 39908 43376
rect 37740 43231 37792 43240
rect 37740 43197 37749 43231
rect 37749 43197 37783 43231
rect 37783 43197 37792 43231
rect 37740 43188 37792 43197
rect 39580 43256 39632 43308
rect 45836 43256 45888 43308
rect 38844 43188 38896 43240
rect 30380 43052 30432 43104
rect 34520 43052 34572 43104
rect 35992 43052 36044 43104
rect 36544 43095 36596 43104
rect 36544 43061 36553 43095
rect 36553 43061 36587 43095
rect 36587 43061 36596 43095
rect 36544 43052 36596 43061
rect 40408 43052 40460 43104
rect 46480 43052 46532 43104
rect 46664 43095 46716 43104
rect 46664 43061 46673 43095
rect 46673 43061 46707 43095
rect 46707 43061 46716 43095
rect 46664 43052 46716 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 15476 42891 15528 42900
rect 15476 42857 15485 42891
rect 15485 42857 15519 42891
rect 15519 42857 15528 42891
rect 15476 42848 15528 42857
rect 16580 42891 16632 42900
rect 16580 42857 16589 42891
rect 16589 42857 16623 42891
rect 16623 42857 16632 42891
rect 16580 42848 16632 42857
rect 17316 42848 17368 42900
rect 22560 42891 22612 42900
rect 22560 42857 22569 42891
rect 22569 42857 22603 42891
rect 22603 42857 22612 42891
rect 22560 42848 22612 42857
rect 30012 42848 30064 42900
rect 35440 42848 35492 42900
rect 39580 42891 39632 42900
rect 39580 42857 39589 42891
rect 39589 42857 39623 42891
rect 39623 42857 39632 42891
rect 39580 42848 39632 42857
rect 13728 42712 13780 42764
rect 15200 42712 15252 42764
rect 16212 42755 16264 42764
rect 16212 42721 16221 42755
rect 16221 42721 16255 42755
rect 16255 42721 16264 42755
rect 16212 42712 16264 42721
rect 22652 42780 22704 42832
rect 29184 42780 29236 42832
rect 30196 42780 30248 42832
rect 36544 42780 36596 42832
rect 19708 42755 19760 42764
rect 19708 42721 19717 42755
rect 19717 42721 19751 42755
rect 19751 42721 19760 42755
rect 19708 42712 19760 42721
rect 19892 42755 19944 42764
rect 19892 42721 19901 42755
rect 19901 42721 19935 42755
rect 19935 42721 19944 42755
rect 19892 42712 19944 42721
rect 26976 42755 27028 42764
rect 26976 42721 26985 42755
rect 26985 42721 27019 42755
rect 27019 42721 27028 42755
rect 26976 42712 27028 42721
rect 18052 42644 18104 42696
rect 19616 42687 19668 42696
rect 19616 42653 19625 42687
rect 19625 42653 19659 42687
rect 19659 42653 19668 42687
rect 19616 42644 19668 42653
rect 23388 42644 23440 42696
rect 27620 42644 27672 42696
rect 29460 42644 29512 42696
rect 30288 42644 30340 42696
rect 30472 42712 30524 42764
rect 32128 42644 32180 42696
rect 13268 42576 13320 42628
rect 15108 42576 15160 42628
rect 17592 42576 17644 42628
rect 20444 42576 20496 42628
rect 25872 42576 25924 42628
rect 28816 42576 28868 42628
rect 15844 42508 15896 42560
rect 19064 42508 19116 42560
rect 19248 42551 19300 42560
rect 19248 42517 19257 42551
rect 19257 42517 19291 42551
rect 19291 42517 19300 42551
rect 19248 42508 19300 42517
rect 19708 42508 19760 42560
rect 30196 42619 30248 42628
rect 30196 42585 30205 42619
rect 30205 42585 30239 42619
rect 30239 42585 30248 42619
rect 30196 42576 30248 42585
rect 32956 42687 33008 42696
rect 32956 42653 32965 42687
rect 32965 42653 32999 42687
rect 32999 42653 33008 42687
rect 32956 42644 33008 42653
rect 35072 42644 35124 42696
rect 34152 42576 34204 42628
rect 37280 42644 37332 42696
rect 38292 42644 38344 42696
rect 38476 42644 38528 42696
rect 35992 42576 36044 42628
rect 29552 42508 29604 42560
rect 29920 42508 29972 42560
rect 30840 42508 30892 42560
rect 32588 42551 32640 42560
rect 32588 42517 32597 42551
rect 32597 42517 32631 42551
rect 32631 42517 32640 42551
rect 32588 42508 32640 42517
rect 38844 42551 38896 42560
rect 38844 42517 38853 42551
rect 38853 42517 38887 42551
rect 38887 42517 38896 42551
rect 38844 42508 38896 42517
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 35594 42406 35646 42458
rect 35658 42406 35710 42458
rect 35722 42406 35774 42458
rect 35786 42406 35838 42458
rect 35850 42406 35902 42458
rect 13268 42347 13320 42356
rect 13268 42313 13277 42347
rect 13277 42313 13311 42347
rect 13311 42313 13320 42347
rect 13268 42304 13320 42313
rect 15844 42347 15896 42356
rect 15844 42313 15853 42347
rect 15853 42313 15887 42347
rect 15887 42313 15896 42347
rect 15844 42304 15896 42313
rect 18052 42304 18104 42356
rect 19064 42347 19116 42356
rect 19064 42313 19073 42347
rect 19073 42313 19107 42347
rect 19107 42313 19116 42347
rect 19064 42304 19116 42313
rect 21456 42304 21508 42356
rect 1400 42236 1452 42288
rect 29460 42279 29512 42288
rect 29460 42245 29469 42279
rect 29469 42245 29503 42279
rect 29503 42245 29512 42279
rect 29460 42236 29512 42245
rect 30012 42279 30064 42288
rect 30012 42245 30021 42279
rect 30021 42245 30055 42279
rect 30055 42245 30064 42279
rect 30012 42236 30064 42245
rect 31668 42304 31720 42356
rect 32956 42304 33008 42356
rect 33600 42347 33652 42356
rect 33600 42313 33609 42347
rect 33609 42313 33643 42347
rect 33643 42313 33652 42347
rect 33600 42304 33652 42313
rect 12716 42168 12768 42220
rect 13544 42168 13596 42220
rect 13728 42143 13780 42152
rect 13728 42109 13737 42143
rect 13737 42109 13771 42143
rect 13771 42109 13780 42143
rect 13728 42100 13780 42109
rect 19248 42168 19300 42220
rect 19892 42100 19944 42152
rect 20352 42032 20404 42084
rect 20444 42032 20496 42084
rect 26884 42032 26936 42084
rect 29552 42211 29604 42220
rect 29552 42177 29561 42211
rect 29561 42177 29595 42211
rect 29595 42177 29604 42211
rect 29552 42168 29604 42177
rect 29920 42211 29972 42220
rect 29920 42177 29929 42211
rect 29929 42177 29963 42211
rect 29963 42177 29972 42211
rect 29920 42168 29972 42177
rect 30840 42211 30892 42220
rect 30840 42177 30874 42211
rect 30874 42177 30892 42211
rect 30840 42168 30892 42177
rect 32588 42236 32640 42288
rect 34244 42279 34296 42288
rect 34244 42245 34253 42279
rect 34253 42245 34287 42279
rect 34287 42245 34296 42279
rect 34244 42236 34296 42245
rect 32036 42100 32088 42152
rect 30196 42032 30248 42084
rect 19064 41964 19116 42016
rect 19524 41964 19576 42016
rect 21640 41964 21692 42016
rect 31668 41964 31720 42016
rect 34704 42168 34756 42220
rect 35348 42211 35400 42220
rect 35348 42177 35357 42211
rect 35357 42177 35391 42211
rect 35391 42177 35400 42211
rect 35348 42168 35400 42177
rect 34244 42100 34296 42152
rect 35072 42100 35124 42152
rect 35624 42100 35676 42152
rect 35440 41964 35492 42016
rect 37096 41964 37148 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 13544 41760 13596 41812
rect 19892 41760 19944 41812
rect 21272 41692 21324 41744
rect 32128 41803 32180 41812
rect 32128 41769 32137 41803
rect 32137 41769 32171 41803
rect 32171 41769 32180 41803
rect 32128 41760 32180 41769
rect 32864 41760 32916 41812
rect 33140 41735 33192 41744
rect 33140 41701 33149 41735
rect 33149 41701 33183 41735
rect 33183 41701 33192 41735
rect 33140 41692 33192 41701
rect 11336 41667 11388 41676
rect 11336 41633 11345 41667
rect 11345 41633 11379 41667
rect 11379 41633 11388 41667
rect 11336 41624 11388 41633
rect 17040 41624 17092 41676
rect 19156 41624 19208 41676
rect 1400 41599 1452 41608
rect 1400 41565 1409 41599
rect 1409 41565 1443 41599
rect 1443 41565 1452 41599
rect 1400 41556 1452 41565
rect 940 41420 992 41472
rect 12900 41556 12952 41608
rect 17316 41556 17368 41608
rect 19064 41599 19116 41608
rect 19064 41565 19073 41599
rect 19073 41565 19107 41599
rect 19107 41565 19116 41599
rect 19064 41556 19116 41565
rect 19524 41599 19576 41608
rect 19524 41565 19558 41599
rect 19558 41565 19576 41599
rect 19524 41556 19576 41565
rect 20904 41599 20956 41608
rect 20904 41565 20913 41599
rect 20913 41565 20947 41599
rect 20947 41565 20956 41599
rect 20904 41556 20956 41565
rect 21824 41556 21876 41608
rect 24308 41556 24360 41608
rect 26884 41556 26936 41608
rect 31852 41556 31904 41608
rect 23940 41488 23992 41540
rect 27344 41488 27396 41540
rect 27988 41488 28040 41540
rect 29920 41488 29972 41540
rect 31576 41488 31628 41540
rect 31668 41488 31720 41540
rect 32680 41624 32732 41676
rect 34520 41692 34572 41744
rect 34888 41803 34940 41812
rect 34888 41769 34897 41803
rect 34897 41769 34931 41803
rect 34931 41769 34940 41803
rect 34888 41760 34940 41769
rect 35164 41803 35216 41812
rect 35164 41769 35173 41803
rect 35173 41769 35207 41803
rect 35207 41769 35216 41803
rect 35164 41760 35216 41769
rect 35440 41760 35492 41812
rect 36728 41760 36780 41812
rect 37648 41760 37700 41812
rect 38844 41760 38896 41812
rect 32036 41556 32088 41608
rect 33324 41556 33376 41608
rect 34796 41624 34848 41676
rect 35348 41624 35400 41676
rect 36360 41624 36412 41676
rect 18052 41420 18104 41472
rect 18880 41463 18932 41472
rect 18880 41429 18889 41463
rect 18889 41429 18923 41463
rect 18923 41429 18932 41463
rect 18880 41420 18932 41429
rect 20720 41463 20772 41472
rect 20720 41429 20729 41463
rect 20729 41429 20763 41463
rect 20763 41429 20772 41463
rect 20720 41420 20772 41429
rect 22100 41420 22152 41472
rect 24492 41420 24544 41472
rect 30196 41420 30248 41472
rect 32404 41420 32456 41472
rect 32588 41463 32640 41472
rect 32588 41429 32597 41463
rect 32597 41429 32631 41463
rect 32631 41429 32640 41463
rect 32588 41420 32640 41429
rect 34428 41463 34480 41472
rect 34428 41429 34437 41463
rect 34437 41429 34471 41463
rect 34471 41429 34480 41463
rect 34428 41420 34480 41429
rect 34612 41488 34664 41540
rect 34796 41488 34848 41540
rect 34980 41599 35032 41608
rect 34980 41565 34989 41599
rect 34989 41565 35023 41599
rect 35023 41565 35032 41599
rect 34980 41556 35032 41565
rect 35072 41488 35124 41540
rect 35440 41556 35492 41608
rect 35716 41556 35768 41608
rect 39396 41488 39448 41540
rect 35348 41420 35400 41472
rect 35532 41420 35584 41472
rect 35624 41420 35676 41472
rect 35992 41420 36044 41472
rect 36452 41420 36504 41472
rect 38660 41420 38712 41472
rect 38936 41463 38988 41472
rect 38936 41429 38945 41463
rect 38945 41429 38979 41463
rect 38979 41429 38988 41463
rect 38936 41420 38988 41429
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 35594 41318 35646 41370
rect 35658 41318 35710 41370
rect 35722 41318 35774 41370
rect 35786 41318 35838 41370
rect 35850 41318 35902 41370
rect 10048 41216 10100 41268
rect 11336 41148 11388 41200
rect 17408 41148 17460 41200
rect 18420 41148 18472 41200
rect 12164 41080 12216 41132
rect 13636 41080 13688 41132
rect 14464 41123 14516 41132
rect 14464 41089 14498 41123
rect 14498 41089 14516 41123
rect 14464 41080 14516 41089
rect 16948 41123 17000 41132
rect 16948 41089 16957 41123
rect 16957 41089 16991 41123
rect 16991 41089 17000 41123
rect 16948 41080 17000 41089
rect 18604 41080 18656 41132
rect 18880 41148 18932 41200
rect 20720 41148 20772 41200
rect 22100 41191 22152 41200
rect 22100 41157 22134 41191
rect 22134 41157 22152 41191
rect 23940 41259 23992 41268
rect 23940 41225 23949 41259
rect 23949 41225 23983 41259
rect 23983 41225 23992 41259
rect 23940 41216 23992 41225
rect 26056 41216 26108 41268
rect 34612 41216 34664 41268
rect 34888 41216 34940 41268
rect 35072 41216 35124 41268
rect 35348 41216 35400 41268
rect 22100 41148 22152 41157
rect 24216 41148 24268 41200
rect 34152 41148 34204 41200
rect 13268 41012 13320 41064
rect 14004 41012 14056 41064
rect 17040 41055 17092 41064
rect 17040 41021 17049 41055
rect 17049 41021 17083 41055
rect 17083 41021 17092 41055
rect 17040 41012 17092 41021
rect 21732 41012 21784 41064
rect 24032 41080 24084 41132
rect 24400 41123 24452 41132
rect 24400 41089 24409 41123
rect 24409 41089 24443 41123
rect 24443 41089 24452 41123
rect 24400 41080 24452 41089
rect 33692 41080 33744 41132
rect 34428 41080 34480 41132
rect 34980 41080 35032 41132
rect 24308 41012 24360 41064
rect 27804 41012 27856 41064
rect 28448 41012 28500 41064
rect 34796 41012 34848 41064
rect 35348 41123 35400 41132
rect 35348 41089 35357 41123
rect 35357 41089 35391 41123
rect 35391 41089 35400 41123
rect 35348 41080 35400 41089
rect 35532 41080 35584 41132
rect 36084 41148 36136 41200
rect 36728 41148 36780 41200
rect 37004 41148 37056 41200
rect 37280 41123 37332 41132
rect 37280 41089 37289 41123
rect 37289 41089 37323 41123
rect 37323 41089 37332 41123
rect 37280 41080 37332 41089
rect 35808 41012 35860 41064
rect 10692 40944 10744 40996
rect 21640 40987 21692 40996
rect 21640 40953 21649 40987
rect 21649 40953 21683 40987
rect 21683 40953 21692 40987
rect 21640 40944 21692 40953
rect 24216 40987 24268 40996
rect 24216 40953 24225 40987
rect 24225 40953 24259 40987
rect 24259 40953 24268 40987
rect 24216 40944 24268 40953
rect 34428 40944 34480 40996
rect 35348 40944 35400 40996
rect 10784 40876 10836 40928
rect 11520 40876 11572 40928
rect 15384 40876 15436 40928
rect 16580 40876 16632 40928
rect 18236 40876 18288 40928
rect 20996 40876 21048 40928
rect 22008 40876 22060 40928
rect 25872 40919 25924 40928
rect 25872 40885 25881 40919
rect 25881 40885 25915 40919
rect 25915 40885 25924 40919
rect 25872 40876 25924 40885
rect 34244 40876 34296 40928
rect 34796 40876 34848 40928
rect 36268 40944 36320 40996
rect 36544 40944 36596 40996
rect 36820 41012 36872 41064
rect 37648 41123 37700 41132
rect 37648 41089 37657 41123
rect 37657 41089 37691 41123
rect 37691 41089 37700 41123
rect 37648 41080 37700 41089
rect 39396 41148 39448 41200
rect 38384 41123 38436 41132
rect 38384 41089 38393 41123
rect 38393 41089 38427 41123
rect 38427 41089 38436 41123
rect 38384 41080 38436 41089
rect 38660 41123 38712 41132
rect 38660 41089 38669 41123
rect 38669 41089 38703 41123
rect 38703 41089 38712 41123
rect 38660 41080 38712 41089
rect 38844 41123 38896 41132
rect 38844 41089 38853 41123
rect 38853 41089 38887 41123
rect 38887 41089 38896 41123
rect 38844 41080 38896 41089
rect 38936 41012 38988 41064
rect 39212 41012 39264 41064
rect 40132 41012 40184 41064
rect 38476 40987 38528 40996
rect 38476 40953 38485 40987
rect 38485 40953 38519 40987
rect 38519 40953 38528 40987
rect 38476 40944 38528 40953
rect 36360 40876 36412 40928
rect 37096 40876 37148 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 2044 40511 2096 40520
rect 2044 40477 2053 40511
rect 2053 40477 2087 40511
rect 2087 40477 2096 40511
rect 2044 40468 2096 40477
rect 3424 40468 3476 40520
rect 2596 40332 2648 40384
rect 10232 40672 10284 40724
rect 12164 40715 12216 40724
rect 12164 40681 12173 40715
rect 12173 40681 12207 40715
rect 12207 40681 12216 40715
rect 12164 40672 12216 40681
rect 12532 40672 12584 40724
rect 14004 40672 14056 40724
rect 10784 40579 10836 40588
rect 8944 40511 8996 40520
rect 8944 40477 8953 40511
rect 8953 40477 8987 40511
rect 8987 40477 8996 40511
rect 10784 40545 10793 40579
rect 10793 40545 10827 40579
rect 10827 40545 10836 40579
rect 10784 40536 10836 40545
rect 8944 40468 8996 40477
rect 10692 40511 10744 40520
rect 10692 40477 10701 40511
rect 10701 40477 10735 40511
rect 10735 40477 10744 40511
rect 10692 40468 10744 40477
rect 12532 40511 12584 40520
rect 12532 40477 12541 40511
rect 12541 40477 12575 40511
rect 12575 40477 12584 40511
rect 12532 40468 12584 40477
rect 14004 40536 14056 40588
rect 16672 40672 16724 40724
rect 20904 40672 20956 40724
rect 21824 40715 21876 40724
rect 21824 40681 21833 40715
rect 21833 40681 21867 40715
rect 21867 40681 21876 40715
rect 21824 40672 21876 40681
rect 22560 40672 22612 40724
rect 36728 40672 36780 40724
rect 38476 40672 38528 40724
rect 18236 40579 18288 40588
rect 18236 40545 18245 40579
rect 18245 40545 18279 40579
rect 18279 40545 18288 40579
rect 18236 40536 18288 40545
rect 18696 40536 18748 40588
rect 13176 40468 13228 40520
rect 15108 40468 15160 40520
rect 16580 40511 16632 40520
rect 16580 40477 16614 40511
rect 16614 40477 16632 40511
rect 8852 40400 8904 40452
rect 6920 40375 6972 40384
rect 6920 40341 6929 40375
rect 6929 40341 6963 40375
rect 6963 40341 6972 40375
rect 6920 40332 6972 40341
rect 10416 40332 10468 40384
rect 15476 40400 15528 40452
rect 16580 40468 16632 40477
rect 37832 40604 37884 40656
rect 38844 40647 38896 40656
rect 38844 40613 38853 40647
rect 38853 40613 38887 40647
rect 38887 40613 38896 40647
rect 38844 40604 38896 40613
rect 20444 40536 20496 40588
rect 21640 40468 21692 40520
rect 17040 40400 17092 40452
rect 19064 40400 19116 40452
rect 22468 40579 22520 40588
rect 22468 40545 22477 40579
rect 22477 40545 22511 40579
rect 22511 40545 22520 40579
rect 22468 40536 22520 40545
rect 24308 40536 24360 40588
rect 22008 40468 22060 40520
rect 22560 40400 22612 40452
rect 13544 40332 13596 40384
rect 15200 40375 15252 40384
rect 15200 40341 15209 40375
rect 15209 40341 15243 40375
rect 15243 40341 15252 40375
rect 15200 40332 15252 40341
rect 15384 40332 15436 40384
rect 17684 40375 17736 40384
rect 17684 40341 17693 40375
rect 17693 40341 17727 40375
rect 17727 40341 17736 40375
rect 17684 40332 17736 40341
rect 17776 40332 17828 40384
rect 18604 40375 18656 40384
rect 18604 40341 18613 40375
rect 18613 40341 18647 40375
rect 18647 40341 18656 40375
rect 18604 40332 18656 40341
rect 20628 40375 20680 40384
rect 20628 40341 20637 40375
rect 20637 40341 20671 40375
rect 20671 40341 20680 40375
rect 20628 40332 20680 40341
rect 22284 40375 22336 40384
rect 22284 40341 22293 40375
rect 22293 40341 22327 40375
rect 22327 40341 22336 40375
rect 22284 40332 22336 40341
rect 27252 40468 27304 40520
rect 27436 40511 27488 40520
rect 27436 40477 27445 40511
rect 27445 40477 27479 40511
rect 27479 40477 27488 40511
rect 27436 40468 27488 40477
rect 36360 40536 36412 40588
rect 36544 40579 36596 40588
rect 36544 40545 36553 40579
rect 36553 40545 36587 40579
rect 36587 40545 36596 40579
rect 36544 40536 36596 40545
rect 40132 40579 40184 40588
rect 40132 40545 40141 40579
rect 40141 40545 40175 40579
rect 40175 40545 40184 40579
rect 40132 40536 40184 40545
rect 23020 40400 23072 40452
rect 26240 40400 26292 40452
rect 23572 40332 23624 40384
rect 27068 40375 27120 40384
rect 27068 40341 27077 40375
rect 27077 40341 27111 40375
rect 27111 40341 27120 40375
rect 27068 40332 27120 40341
rect 29368 40468 29420 40520
rect 30932 40468 30984 40520
rect 33048 40468 33100 40520
rect 34888 40468 34940 40520
rect 35348 40511 35400 40520
rect 35348 40477 35357 40511
rect 35357 40477 35391 40511
rect 35391 40477 35400 40511
rect 35348 40468 35400 40477
rect 35808 40511 35860 40520
rect 35808 40477 35817 40511
rect 35817 40477 35851 40511
rect 35851 40477 35860 40511
rect 35808 40468 35860 40477
rect 36728 40468 36780 40520
rect 36820 40468 36872 40520
rect 37188 40468 37240 40520
rect 38016 40468 38068 40520
rect 38660 40468 38712 40520
rect 27896 40400 27948 40452
rect 30564 40400 30616 40452
rect 34060 40400 34112 40452
rect 36268 40400 36320 40452
rect 39212 40468 39264 40520
rect 45560 40468 45612 40520
rect 38936 40400 38988 40452
rect 28264 40332 28316 40384
rect 28908 40375 28960 40384
rect 28908 40341 28917 40375
rect 28917 40341 28951 40375
rect 28951 40341 28960 40375
rect 28908 40332 28960 40341
rect 31760 40332 31812 40384
rect 33600 40332 33652 40384
rect 34796 40332 34848 40384
rect 36360 40332 36412 40384
rect 36912 40332 36964 40384
rect 37096 40332 37148 40384
rect 37464 40375 37516 40384
rect 37464 40341 37473 40375
rect 37473 40341 37507 40375
rect 37507 40341 37516 40375
rect 37464 40332 37516 40341
rect 39396 40375 39448 40384
rect 39396 40341 39405 40375
rect 39405 40341 39439 40375
rect 39439 40341 39448 40375
rect 39396 40332 39448 40341
rect 39580 40375 39632 40384
rect 39580 40341 39589 40375
rect 39589 40341 39623 40375
rect 39623 40341 39632 40375
rect 39580 40332 39632 40341
rect 39856 40332 39908 40384
rect 40408 40375 40460 40384
rect 40408 40341 40417 40375
rect 40417 40341 40451 40375
rect 40451 40341 40460 40375
rect 40408 40332 40460 40341
rect 46664 40375 46716 40384
rect 46664 40341 46673 40375
rect 46673 40341 46707 40375
rect 46707 40341 46716 40375
rect 46664 40332 46716 40341
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 35594 40230 35646 40282
rect 35658 40230 35710 40282
rect 35722 40230 35774 40282
rect 35786 40230 35838 40282
rect 35850 40230 35902 40282
rect 2044 40128 2096 40180
rect 2596 40171 2648 40180
rect 2596 40137 2605 40171
rect 2605 40137 2639 40171
rect 2639 40137 2648 40171
rect 2596 40128 2648 40137
rect 8852 40171 8904 40180
rect 8852 40137 8861 40171
rect 8861 40137 8895 40171
rect 8895 40137 8904 40171
rect 8852 40128 8904 40137
rect 2044 39992 2096 40044
rect 10048 40103 10100 40112
rect 10048 40069 10057 40103
rect 10057 40069 10091 40103
rect 10091 40069 10100 40103
rect 10048 40060 10100 40069
rect 12440 40128 12492 40180
rect 13176 40171 13228 40180
rect 13176 40137 13185 40171
rect 13185 40137 13219 40171
rect 13219 40137 13228 40171
rect 13176 40128 13228 40137
rect 13544 40171 13596 40180
rect 13544 40137 13553 40171
rect 13553 40137 13587 40171
rect 13587 40137 13596 40171
rect 13544 40128 13596 40137
rect 14464 40128 14516 40180
rect 16948 40128 17000 40180
rect 17684 40171 17736 40180
rect 17684 40137 17693 40171
rect 17693 40137 17727 40171
rect 17727 40137 17736 40171
rect 17684 40128 17736 40137
rect 23020 40171 23072 40180
rect 23020 40137 23029 40171
rect 23029 40137 23063 40171
rect 23063 40137 23072 40171
rect 23020 40128 23072 40137
rect 24032 40171 24084 40180
rect 24032 40137 24041 40171
rect 24041 40137 24075 40171
rect 24075 40137 24084 40171
rect 24032 40128 24084 40137
rect 24400 40128 24452 40180
rect 24952 40128 25004 40180
rect 25872 40128 25924 40180
rect 26240 40171 26292 40180
rect 26240 40137 26249 40171
rect 26249 40137 26283 40171
rect 26283 40137 26292 40171
rect 26240 40128 26292 40137
rect 11888 40060 11940 40112
rect 10416 39992 10468 40044
rect 10600 39992 10652 40044
rect 11336 40035 11388 40044
rect 11336 40001 11345 40035
rect 11345 40001 11379 40035
rect 11379 40001 11388 40035
rect 11336 39992 11388 40001
rect 11520 40035 11572 40044
rect 11520 40001 11529 40035
rect 11529 40001 11563 40035
rect 11563 40001 11572 40035
rect 11520 39992 11572 40001
rect 15200 40060 15252 40112
rect 22284 40060 22336 40112
rect 2688 39967 2740 39976
rect 2688 39933 2697 39967
rect 2697 39933 2731 39967
rect 2731 39933 2740 39967
rect 2688 39924 2740 39933
rect 10232 39967 10284 39976
rect 10232 39933 10241 39967
rect 10241 39933 10275 39967
rect 10275 39933 10284 39967
rect 10232 39924 10284 39933
rect 3148 39856 3200 39908
rect 13636 39967 13688 39976
rect 13636 39933 13645 39967
rect 13645 39933 13679 39967
rect 13679 39933 13688 39967
rect 13636 39924 13688 39933
rect 20444 39992 20496 40044
rect 23204 40035 23256 40044
rect 23204 40001 23213 40035
rect 23213 40001 23247 40035
rect 23247 40001 23256 40035
rect 23204 39992 23256 40001
rect 17776 39967 17828 39976
rect 17776 39933 17785 39967
rect 17785 39933 17819 39967
rect 17819 39933 17828 39967
rect 17776 39924 17828 39933
rect 24492 40060 24544 40112
rect 24676 40060 24728 40112
rect 26884 40128 26936 40180
rect 27068 40128 27120 40180
rect 29368 40171 29420 40180
rect 29368 40137 29377 40171
rect 29377 40137 29411 40171
rect 29411 40137 29420 40171
rect 29368 40128 29420 40137
rect 30564 40171 30616 40180
rect 30564 40137 30573 40171
rect 30573 40137 30607 40171
rect 30607 40137 30616 40171
rect 30564 40128 30616 40137
rect 27436 40060 27488 40112
rect 28908 40060 28960 40112
rect 31760 40128 31812 40180
rect 32772 40128 32824 40180
rect 34060 40171 34112 40180
rect 34060 40137 34069 40171
rect 34069 40137 34103 40171
rect 34103 40137 34112 40171
rect 34060 40128 34112 40137
rect 37556 40128 37608 40180
rect 38660 40128 38712 40180
rect 15016 39856 15068 39908
rect 15476 39856 15528 39908
rect 24768 39924 24820 39976
rect 940 39788 992 39840
rect 2044 39831 2096 39840
rect 2044 39797 2053 39831
rect 2053 39797 2087 39831
rect 2087 39797 2096 39831
rect 2044 39788 2096 39797
rect 6920 39831 6972 39840
rect 6920 39797 6929 39831
rect 6929 39797 6963 39831
rect 6963 39797 6972 39831
rect 6920 39788 6972 39797
rect 9036 39788 9088 39840
rect 10048 39788 10100 39840
rect 10232 39788 10284 39840
rect 17776 39788 17828 39840
rect 28448 39992 28500 40044
rect 29736 40035 29788 40044
rect 29736 40001 29745 40035
rect 29745 40001 29779 40035
rect 29779 40001 29788 40035
rect 29736 39992 29788 40001
rect 33140 40060 33192 40112
rect 33692 40103 33744 40112
rect 33692 40069 33701 40103
rect 33701 40069 33735 40103
rect 33735 40069 33744 40103
rect 33692 40060 33744 40069
rect 33784 40103 33836 40112
rect 33784 40069 33793 40103
rect 33793 40069 33827 40103
rect 33827 40069 33836 40103
rect 33784 40060 33836 40069
rect 34428 40060 34480 40112
rect 34796 40060 34848 40112
rect 34888 40060 34940 40112
rect 35992 40060 36044 40112
rect 33416 40035 33468 40044
rect 33416 40001 33425 40035
rect 33425 40001 33459 40035
rect 33459 40001 33468 40035
rect 33416 39992 33468 40001
rect 33600 40035 33652 40044
rect 33600 40001 33607 40035
rect 33607 40001 33652 40035
rect 33600 39992 33652 40001
rect 26240 39924 26292 39976
rect 27436 39967 27488 39976
rect 27436 39933 27445 39967
rect 27445 39933 27479 39967
rect 27479 39933 27488 39967
rect 27436 39924 27488 39933
rect 27528 39967 27580 39976
rect 27528 39933 27537 39967
rect 27537 39933 27571 39967
rect 27571 39933 27580 39967
rect 27528 39924 27580 39933
rect 29000 39856 29052 39908
rect 30012 39967 30064 39976
rect 30012 39933 30021 39967
rect 30021 39933 30055 39967
rect 30055 39933 30064 39967
rect 30012 39924 30064 39933
rect 31392 39967 31444 39976
rect 31392 39933 31401 39967
rect 31401 39933 31435 39967
rect 31435 39933 31444 39967
rect 31392 39924 31444 39933
rect 35256 39992 35308 40044
rect 34152 39924 34204 39976
rect 34428 39924 34480 39976
rect 34796 39924 34848 39976
rect 35440 39924 35492 39976
rect 37464 40060 37516 40112
rect 36360 39992 36412 40044
rect 36728 40035 36780 40044
rect 36728 40001 36737 40035
rect 36737 40001 36771 40035
rect 36771 40001 36780 40035
rect 36728 39992 36780 40001
rect 39396 40128 39448 40180
rect 38844 40060 38896 40112
rect 40408 40060 40460 40112
rect 36912 39924 36964 39976
rect 37832 39856 37884 39908
rect 39856 39992 39908 40044
rect 38936 39924 38988 39976
rect 39580 39924 39632 39976
rect 39856 39856 39908 39908
rect 31300 39788 31352 39840
rect 37188 39788 37240 39840
rect 37280 39788 37332 39840
rect 37648 39788 37700 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 1492 39584 1544 39636
rect 13084 39584 13136 39636
rect 2044 39559 2096 39568
rect 2044 39525 2053 39559
rect 2053 39525 2087 39559
rect 2087 39525 2096 39559
rect 2044 39516 2096 39525
rect 6920 39559 6972 39568
rect 6920 39525 6929 39559
rect 6929 39525 6963 39559
rect 6963 39525 6972 39559
rect 6920 39516 6972 39525
rect 11336 39516 11388 39568
rect 23204 39627 23256 39636
rect 23204 39593 23213 39627
rect 23213 39593 23247 39627
rect 23247 39593 23256 39627
rect 23204 39584 23256 39593
rect 27896 39627 27948 39636
rect 27896 39593 27905 39627
rect 27905 39593 27939 39627
rect 27939 39593 27948 39627
rect 27896 39584 27948 39593
rect 25688 39516 25740 39568
rect 26240 39516 26292 39568
rect 30012 39584 30064 39636
rect 30840 39584 30892 39636
rect 13084 39448 13136 39500
rect 13176 39380 13228 39432
rect 14004 39380 14056 39432
rect 17316 39448 17368 39500
rect 26792 39448 26844 39500
rect 27436 39448 27488 39500
rect 29736 39516 29788 39568
rect 36452 39516 36504 39568
rect 37188 39516 37240 39568
rect 37464 39584 37516 39636
rect 39856 39584 39908 39636
rect 37648 39516 37700 39568
rect 29092 39448 29144 39500
rect 30196 39448 30248 39500
rect 30932 39491 30984 39500
rect 30932 39457 30941 39491
rect 30941 39457 30975 39491
rect 30975 39457 30984 39491
rect 30932 39448 30984 39457
rect 31944 39448 31996 39500
rect 36912 39448 36964 39500
rect 19708 39380 19760 39432
rect 23572 39423 23624 39432
rect 23572 39389 23581 39423
rect 23581 39389 23615 39423
rect 23615 39389 23624 39423
rect 23572 39380 23624 39389
rect 27620 39380 27672 39432
rect 28264 39423 28316 39432
rect 28264 39389 28273 39423
rect 28273 39389 28307 39423
rect 28307 39389 28316 39423
rect 28264 39380 28316 39389
rect 14740 39355 14792 39364
rect 14740 39321 14749 39355
rect 14749 39321 14783 39355
rect 14783 39321 14792 39355
rect 14740 39312 14792 39321
rect 17500 39312 17552 39364
rect 27988 39312 28040 39364
rect 30748 39380 30800 39432
rect 30840 39423 30892 39432
rect 30840 39389 30849 39423
rect 30849 39389 30883 39423
rect 30883 39389 30892 39423
rect 30840 39380 30892 39389
rect 36360 39423 36412 39432
rect 36360 39389 36369 39423
rect 36369 39389 36403 39423
rect 36403 39389 36412 39423
rect 36360 39380 36412 39389
rect 36544 39423 36596 39432
rect 36544 39389 36553 39423
rect 36553 39389 36587 39423
rect 36587 39389 36596 39423
rect 36544 39380 36596 39389
rect 36636 39380 36688 39432
rect 38292 39491 38344 39500
rect 38292 39457 38301 39491
rect 38301 39457 38335 39491
rect 38335 39457 38344 39491
rect 38292 39448 38344 39457
rect 37924 39380 37976 39432
rect 9036 39244 9088 39296
rect 12164 39287 12216 39296
rect 12164 39253 12173 39287
rect 12173 39253 12207 39287
rect 12207 39253 12216 39287
rect 12164 39244 12216 39253
rect 13636 39244 13688 39296
rect 15476 39244 15528 39296
rect 16764 39287 16816 39296
rect 16764 39253 16773 39287
rect 16773 39253 16807 39287
rect 16807 39253 16816 39287
rect 16764 39244 16816 39253
rect 17132 39244 17184 39296
rect 20168 39244 20220 39296
rect 23664 39287 23716 39296
rect 23664 39253 23673 39287
rect 23673 39253 23707 39287
rect 23707 39253 23716 39287
rect 23664 39244 23716 39253
rect 24768 39244 24820 39296
rect 29092 39244 29144 39296
rect 30748 39244 30800 39296
rect 35440 39312 35492 39364
rect 35992 39355 36044 39364
rect 35992 39321 36001 39355
rect 36001 39321 36035 39355
rect 36035 39321 36044 39355
rect 35992 39312 36044 39321
rect 36912 39312 36964 39364
rect 32680 39244 32732 39296
rect 32864 39287 32916 39296
rect 32864 39253 32873 39287
rect 32873 39253 32907 39287
rect 32907 39253 32916 39287
rect 32864 39244 32916 39253
rect 34336 39244 34388 39296
rect 35164 39244 35216 39296
rect 37832 39355 37884 39364
rect 37832 39321 37841 39355
rect 37841 39321 37875 39355
rect 37875 39321 37884 39355
rect 37832 39312 37884 39321
rect 36636 39244 36688 39296
rect 36728 39287 36780 39296
rect 36728 39253 36737 39287
rect 36737 39253 36771 39287
rect 36771 39253 36780 39287
rect 36728 39244 36780 39253
rect 37740 39244 37792 39296
rect 38200 39287 38252 39296
rect 38200 39253 38209 39287
rect 38209 39253 38243 39287
rect 38243 39253 38252 39287
rect 38200 39244 38252 39253
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 35594 39142 35646 39194
rect 35658 39142 35710 39194
rect 35722 39142 35774 39194
rect 35786 39142 35838 39194
rect 35850 39142 35902 39194
rect 3516 39040 3568 39092
rect 31484 39040 31536 39092
rect 34336 39040 34388 39092
rect 34520 39040 34572 39092
rect 16396 38972 16448 39024
rect 7656 38904 7708 38956
rect 10508 38904 10560 38956
rect 15108 38947 15160 38956
rect 15108 38913 15117 38947
rect 15117 38913 15151 38947
rect 15151 38913 15160 38947
rect 15108 38904 15160 38913
rect 15936 38904 15988 38956
rect 17776 38972 17828 39024
rect 27988 38972 28040 39024
rect 29736 38972 29788 39024
rect 30288 39015 30340 39024
rect 30288 38981 30297 39015
rect 30297 38981 30331 39015
rect 30331 38981 30340 39015
rect 30288 38972 30340 38981
rect 31208 39015 31260 39024
rect 31208 38981 31217 39015
rect 31217 38981 31251 39015
rect 31251 38981 31260 39015
rect 31208 38972 31260 38981
rect 31300 38972 31352 39024
rect 32864 38972 32916 39024
rect 16856 38836 16908 38888
rect 17316 38879 17368 38888
rect 17316 38845 17325 38879
rect 17325 38845 17359 38879
rect 17359 38845 17368 38879
rect 17316 38836 17368 38845
rect 19524 38947 19576 38956
rect 19524 38913 19533 38947
rect 19533 38913 19567 38947
rect 19567 38913 19576 38947
rect 19524 38904 19576 38913
rect 20628 38904 20680 38956
rect 21732 38904 21784 38956
rect 22100 38947 22152 38956
rect 22100 38913 22134 38947
rect 22134 38913 22152 38947
rect 22100 38904 22152 38913
rect 25320 38904 25372 38956
rect 25780 38904 25832 38956
rect 30932 38904 30984 38956
rect 17960 38836 18012 38888
rect 18236 38836 18288 38888
rect 20168 38879 20220 38888
rect 20168 38845 20177 38879
rect 20177 38845 20211 38879
rect 20211 38845 20220 38879
rect 20168 38836 20220 38845
rect 7380 38743 7432 38752
rect 7380 38709 7389 38743
rect 7389 38709 7423 38743
rect 7423 38709 7432 38743
rect 7380 38700 7432 38709
rect 9312 38743 9364 38752
rect 9312 38709 9321 38743
rect 9321 38709 9355 38743
rect 9355 38709 9364 38743
rect 9312 38700 9364 38709
rect 14096 38700 14148 38752
rect 14740 38700 14792 38752
rect 17500 38811 17552 38820
rect 17500 38777 17509 38811
rect 17509 38777 17543 38811
rect 17543 38777 17552 38811
rect 17500 38768 17552 38777
rect 23664 38836 23716 38888
rect 27344 38836 27396 38888
rect 31944 38904 31996 38956
rect 34152 38972 34204 39024
rect 16672 38743 16724 38752
rect 16672 38709 16681 38743
rect 16681 38709 16715 38743
rect 16715 38709 16724 38743
rect 16672 38700 16724 38709
rect 17224 38700 17276 38752
rect 19340 38743 19392 38752
rect 19340 38709 19349 38743
rect 19349 38709 19383 38743
rect 19383 38709 19392 38743
rect 19340 38700 19392 38709
rect 20904 38700 20956 38752
rect 23204 38743 23256 38752
rect 23204 38709 23213 38743
rect 23213 38709 23247 38743
rect 23247 38709 23256 38743
rect 23204 38700 23256 38709
rect 24124 38743 24176 38752
rect 24124 38709 24133 38743
rect 24133 38709 24167 38743
rect 24167 38709 24176 38743
rect 24124 38700 24176 38709
rect 29920 38700 29972 38752
rect 31208 38700 31260 38752
rect 33048 38879 33100 38888
rect 33048 38845 33057 38879
rect 33057 38845 33091 38879
rect 33091 38845 33100 38879
rect 33048 38836 33100 38845
rect 34336 38904 34388 38956
rect 34796 38947 34848 38956
rect 34796 38913 34805 38947
rect 34805 38913 34839 38947
rect 34839 38913 34848 38947
rect 34796 38904 34848 38913
rect 34888 38947 34940 38956
rect 34888 38913 34897 38947
rect 34897 38913 34931 38947
rect 34931 38913 34940 38947
rect 34888 38904 34940 38913
rect 35164 38947 35216 38956
rect 35164 38913 35173 38947
rect 35173 38913 35207 38947
rect 35207 38913 35216 38947
rect 35164 38904 35216 38913
rect 35348 38904 35400 38956
rect 36544 38972 36596 39024
rect 36176 38947 36228 38956
rect 36176 38913 36185 38947
rect 36185 38913 36219 38947
rect 36219 38913 36228 38947
rect 36176 38904 36228 38913
rect 37280 39040 37332 39092
rect 37740 39040 37792 39092
rect 38292 38972 38344 39024
rect 35532 38836 35584 38888
rect 35808 38836 35860 38888
rect 36544 38836 36596 38888
rect 36912 38904 36964 38956
rect 37464 38947 37516 38956
rect 37464 38913 37473 38947
rect 37473 38913 37507 38947
rect 37507 38913 37516 38947
rect 37464 38904 37516 38913
rect 37648 38904 37700 38956
rect 38016 38904 38068 38956
rect 38568 38904 38620 38956
rect 37004 38700 37056 38752
rect 37464 38700 37516 38752
rect 38016 38700 38068 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 5356 38496 5408 38548
rect 10968 38496 11020 38548
rect 15936 38496 15988 38548
rect 16396 38539 16448 38548
rect 16396 38505 16405 38539
rect 16405 38505 16439 38539
rect 16439 38505 16448 38539
rect 16396 38496 16448 38505
rect 20168 38496 20220 38548
rect 20628 38539 20680 38548
rect 20628 38505 20637 38539
rect 20637 38505 20671 38539
rect 20671 38505 20680 38539
rect 20628 38496 20680 38505
rect 21456 38496 21508 38548
rect 5264 38292 5316 38344
rect 5632 38335 5684 38344
rect 5632 38301 5641 38335
rect 5641 38301 5675 38335
rect 5675 38301 5684 38335
rect 5632 38292 5684 38301
rect 7380 38335 7432 38344
rect 7380 38301 7414 38335
rect 7414 38301 7432 38335
rect 6000 38224 6052 38276
rect 7380 38292 7432 38301
rect 8944 38224 8996 38276
rect 9312 38335 9364 38344
rect 9312 38301 9346 38335
rect 9346 38301 9364 38335
rect 9312 38292 9364 38301
rect 14004 38360 14056 38412
rect 16948 38403 17000 38412
rect 16948 38369 16957 38403
rect 16957 38369 16991 38403
rect 16991 38369 17000 38403
rect 16948 38360 17000 38369
rect 17040 38360 17092 38412
rect 17684 38428 17736 38480
rect 13360 38292 13412 38344
rect 13636 38335 13688 38344
rect 13636 38301 13645 38335
rect 13645 38301 13679 38335
rect 13679 38301 13688 38335
rect 13636 38292 13688 38301
rect 13912 38335 13964 38344
rect 13912 38301 13921 38335
rect 13921 38301 13955 38335
rect 13955 38301 13964 38335
rect 13912 38292 13964 38301
rect 16672 38292 16724 38344
rect 16764 38335 16816 38344
rect 16764 38301 16773 38335
rect 16773 38301 16807 38335
rect 16807 38301 16816 38335
rect 17776 38360 17828 38412
rect 17868 38403 17920 38412
rect 17868 38369 17877 38403
rect 17877 38369 17911 38403
rect 17911 38369 17920 38403
rect 17868 38360 17920 38369
rect 18236 38403 18288 38412
rect 18236 38369 18270 38403
rect 18270 38369 18288 38403
rect 18236 38360 18288 38369
rect 21180 38403 21232 38412
rect 21180 38369 21189 38403
rect 21189 38369 21223 38403
rect 21223 38369 21232 38403
rect 21180 38360 21232 38369
rect 16764 38292 16816 38301
rect 9220 38224 9272 38276
rect 10692 38224 10744 38276
rect 4160 38199 4212 38208
rect 4160 38165 4169 38199
rect 4169 38165 4203 38199
rect 4203 38165 4212 38199
rect 4160 38156 4212 38165
rect 7012 38199 7064 38208
rect 7012 38165 7021 38199
rect 7021 38165 7055 38199
rect 7055 38165 7064 38199
rect 7012 38156 7064 38165
rect 8484 38199 8536 38208
rect 8484 38165 8493 38199
rect 8493 38165 8527 38199
rect 8527 38165 8536 38199
rect 8484 38156 8536 38165
rect 8760 38156 8812 38208
rect 10876 38156 10928 38208
rect 12532 38199 12584 38208
rect 12532 38165 12541 38199
rect 12541 38165 12575 38199
rect 12575 38165 12584 38199
rect 12532 38156 12584 38165
rect 13820 38156 13872 38208
rect 15476 38199 15528 38208
rect 15476 38165 15485 38199
rect 15485 38165 15519 38199
rect 15519 38165 15528 38199
rect 15476 38156 15528 38165
rect 16856 38199 16908 38208
rect 16856 38165 16865 38199
rect 16865 38165 16899 38199
rect 16899 38165 16908 38199
rect 16856 38156 16908 38165
rect 18420 38335 18472 38344
rect 18420 38301 18429 38335
rect 18429 38301 18463 38335
rect 18463 38301 18472 38335
rect 18420 38292 18472 38301
rect 19064 38292 19116 38344
rect 18972 38224 19024 38276
rect 20904 38335 20956 38344
rect 20904 38301 20913 38335
rect 20913 38301 20947 38335
rect 20947 38301 20956 38335
rect 20904 38292 20956 38301
rect 22744 38360 22796 38412
rect 22928 38428 22980 38480
rect 25780 38539 25832 38548
rect 25780 38505 25789 38539
rect 25789 38505 25823 38539
rect 25823 38505 25832 38539
rect 25780 38496 25832 38505
rect 30932 38539 30984 38548
rect 30932 38505 30941 38539
rect 30941 38505 30975 38539
rect 30975 38505 30984 38539
rect 30932 38496 30984 38505
rect 35440 38496 35492 38548
rect 23664 38360 23716 38412
rect 23848 38360 23900 38412
rect 24308 38360 24360 38412
rect 27344 38360 27396 38412
rect 28448 38360 28500 38412
rect 31024 38360 31076 38412
rect 31668 38403 31720 38412
rect 31668 38369 31677 38403
rect 31677 38369 31711 38403
rect 31711 38369 31720 38403
rect 31668 38360 31720 38369
rect 34428 38403 34480 38412
rect 34428 38369 34437 38403
rect 34437 38369 34471 38403
rect 34471 38369 34480 38403
rect 34428 38360 34480 38369
rect 18144 38156 18196 38208
rect 19432 38156 19484 38208
rect 22192 38335 22244 38344
rect 22192 38301 22226 38335
rect 22226 38301 22244 38335
rect 22192 38292 22244 38301
rect 22376 38335 22428 38344
rect 22376 38301 22385 38335
rect 22385 38301 22419 38335
rect 22419 38301 22428 38335
rect 22376 38292 22428 38301
rect 23204 38292 23256 38344
rect 24124 38335 24176 38344
rect 24124 38301 24133 38335
rect 24133 38301 24167 38335
rect 24167 38301 24176 38335
rect 24124 38292 24176 38301
rect 26976 38292 27028 38344
rect 27804 38292 27856 38344
rect 31576 38335 31628 38344
rect 31576 38301 31585 38335
rect 31585 38301 31619 38335
rect 31619 38301 31628 38335
rect 31576 38292 31628 38301
rect 21916 38156 21968 38208
rect 26608 38267 26660 38276
rect 26608 38233 26642 38267
rect 26642 38233 26660 38267
rect 23020 38199 23072 38208
rect 23020 38165 23029 38199
rect 23029 38165 23063 38199
rect 23063 38165 23072 38199
rect 23020 38156 23072 38165
rect 23112 38199 23164 38208
rect 23112 38165 23121 38199
rect 23121 38165 23155 38199
rect 23155 38165 23164 38199
rect 23112 38156 23164 38165
rect 26608 38224 26660 38233
rect 28080 38224 28132 38276
rect 29828 38267 29880 38276
rect 29828 38233 29862 38267
rect 29862 38233 29880 38267
rect 29828 38224 29880 38233
rect 27712 38199 27764 38208
rect 27712 38165 27721 38199
rect 27721 38165 27755 38199
rect 27755 38165 27764 38199
rect 27712 38156 27764 38165
rect 27804 38199 27856 38208
rect 27804 38165 27813 38199
rect 27813 38165 27847 38199
rect 27847 38165 27856 38199
rect 27804 38156 27856 38165
rect 28172 38199 28224 38208
rect 28172 38165 28181 38199
rect 28181 38165 28215 38199
rect 28215 38165 28224 38199
rect 28172 38156 28224 38165
rect 33232 38224 33284 38276
rect 33784 38292 33836 38344
rect 34612 38292 34664 38344
rect 35808 38428 35860 38480
rect 38200 38496 38252 38548
rect 39396 38496 39448 38548
rect 34796 38360 34848 38412
rect 35348 38292 35400 38344
rect 36728 38292 36780 38344
rect 37004 38360 37056 38412
rect 37188 38403 37240 38412
rect 37188 38369 37197 38403
rect 37197 38369 37231 38403
rect 37231 38369 37240 38403
rect 37188 38360 37240 38369
rect 37280 38403 37332 38412
rect 37280 38369 37289 38403
rect 37289 38369 37323 38403
rect 37323 38369 37332 38403
rect 37280 38360 37332 38369
rect 37372 38403 37424 38412
rect 37372 38369 37381 38403
rect 37381 38369 37415 38403
rect 37415 38369 37424 38403
rect 37372 38360 37424 38369
rect 38016 38292 38068 38344
rect 32496 38156 32548 38208
rect 34336 38156 34388 38208
rect 35532 38156 35584 38208
rect 35992 38224 36044 38276
rect 36820 38224 36872 38276
rect 36912 38199 36964 38208
rect 36912 38165 36921 38199
rect 36921 38165 36955 38199
rect 36955 38165 36964 38199
rect 36912 38156 36964 38165
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 35594 38054 35646 38106
rect 35658 38054 35710 38106
rect 35722 38054 35774 38106
rect 35786 38054 35838 38106
rect 35850 38054 35902 38106
rect 6000 37995 6052 38004
rect 6000 37961 6009 37995
rect 6009 37961 6043 37995
rect 6043 37961 6052 37995
rect 6000 37952 6052 37961
rect 7012 37952 7064 38004
rect 9588 37952 9640 38004
rect 10508 37995 10560 38004
rect 10508 37961 10517 37995
rect 10517 37961 10551 37995
rect 10551 37961 10560 37995
rect 10508 37952 10560 37961
rect 10876 37995 10928 38004
rect 10876 37961 10885 37995
rect 10885 37961 10919 37995
rect 10919 37961 10928 37995
rect 10876 37952 10928 37961
rect 10968 37995 11020 38004
rect 10968 37961 10977 37995
rect 10977 37961 11011 37995
rect 11011 37961 11020 37995
rect 10968 37952 11020 37961
rect 3424 37884 3476 37936
rect 4160 37884 4212 37936
rect 3700 37859 3752 37868
rect 3700 37825 3709 37859
rect 3709 37825 3743 37859
rect 3743 37825 3752 37859
rect 3700 37816 3752 37825
rect 3792 37859 3844 37868
rect 3792 37825 3801 37859
rect 3801 37825 3835 37859
rect 3835 37825 3844 37859
rect 6460 37884 6512 37936
rect 3792 37816 3844 37825
rect 6276 37816 6328 37868
rect 8484 37816 8536 37868
rect 8760 37859 8812 37868
rect 8760 37825 8769 37859
rect 8769 37825 8803 37859
rect 8803 37825 8812 37859
rect 8760 37816 8812 37825
rect 9588 37859 9640 37868
rect 12532 37952 12584 38004
rect 13636 37952 13688 38004
rect 15476 37952 15528 38004
rect 9588 37825 9622 37859
rect 9622 37825 9640 37859
rect 9588 37816 9640 37825
rect 12440 37859 12492 37868
rect 12440 37825 12449 37859
rect 12449 37825 12483 37859
rect 12483 37825 12492 37859
rect 12440 37816 12492 37825
rect 14004 37884 14056 37936
rect 13820 37859 13872 37868
rect 13820 37825 13854 37859
rect 13854 37825 13872 37859
rect 13820 37816 13872 37825
rect 17040 37816 17092 37868
rect 18144 37952 18196 38004
rect 18420 37952 18472 38004
rect 19800 37952 19852 38004
rect 20168 37952 20220 38004
rect 19340 37927 19392 37936
rect 19340 37893 19374 37927
rect 19374 37893 19392 37927
rect 19340 37884 19392 37893
rect 21456 37884 21508 37936
rect 17868 37859 17920 37868
rect 17868 37825 17877 37859
rect 17877 37825 17911 37859
rect 17911 37825 17920 37859
rect 17868 37816 17920 37825
rect 17960 37859 18012 37868
rect 17960 37825 17994 37859
rect 17994 37825 18012 37859
rect 17960 37816 18012 37825
rect 19064 37859 19116 37868
rect 19064 37825 19073 37859
rect 19073 37825 19107 37859
rect 19107 37825 19116 37859
rect 19064 37816 19116 37825
rect 23112 37952 23164 38004
rect 26608 37952 26660 38004
rect 22008 37884 22060 37936
rect 26148 37884 26200 37936
rect 5632 37748 5684 37800
rect 9496 37791 9548 37800
rect 4068 37612 4120 37664
rect 5172 37655 5224 37664
rect 5172 37621 5181 37655
rect 5181 37621 5215 37655
rect 5215 37621 5224 37655
rect 5172 37612 5224 37621
rect 9496 37757 9505 37791
rect 9505 37757 9539 37791
rect 9539 37757 9548 37791
rect 9496 37748 9548 37757
rect 10324 37748 10376 37800
rect 10508 37748 10560 37800
rect 11244 37748 11296 37800
rect 11888 37748 11940 37800
rect 12072 37748 12124 37800
rect 7748 37723 7800 37732
rect 7748 37689 7757 37723
rect 7757 37689 7791 37723
rect 7791 37689 7800 37723
rect 7748 37680 7800 37689
rect 9220 37723 9272 37732
rect 9220 37689 9229 37723
rect 9229 37689 9263 37723
rect 9263 37689 9272 37723
rect 9220 37680 9272 37689
rect 11428 37680 11480 37732
rect 10876 37612 10928 37664
rect 11060 37612 11112 37664
rect 13084 37748 13136 37800
rect 14740 37748 14792 37800
rect 17224 37748 17276 37800
rect 17500 37748 17552 37800
rect 17684 37748 17736 37800
rect 18328 37748 18380 37800
rect 12256 37612 12308 37664
rect 14924 37655 14976 37664
rect 14924 37621 14933 37655
rect 14933 37621 14967 37655
rect 14967 37621 14976 37655
rect 14924 37612 14976 37621
rect 18604 37612 18656 37664
rect 18696 37612 18748 37664
rect 20444 37655 20496 37664
rect 20444 37621 20453 37655
rect 20453 37621 20487 37655
rect 20487 37621 20496 37655
rect 20444 37612 20496 37621
rect 21180 37748 21232 37800
rect 22744 37859 22796 37868
rect 22744 37825 22753 37859
rect 22753 37825 22787 37859
rect 22787 37825 22796 37859
rect 22744 37816 22796 37825
rect 24492 37816 24544 37868
rect 25320 37859 25372 37868
rect 25320 37825 25329 37859
rect 25329 37825 25363 37859
rect 25363 37825 25372 37859
rect 25320 37816 25372 37825
rect 26700 37859 26752 37868
rect 26700 37825 26709 37859
rect 26709 37825 26743 37859
rect 26743 37825 26752 37859
rect 26700 37816 26752 37825
rect 27804 37884 27856 37936
rect 27620 37859 27672 37868
rect 27620 37825 27629 37859
rect 27629 37825 27663 37859
rect 27663 37825 27672 37859
rect 27620 37816 27672 37825
rect 21916 37748 21968 37800
rect 22836 37791 22888 37800
rect 22836 37757 22870 37791
rect 22870 37757 22888 37791
rect 22836 37748 22888 37757
rect 23204 37748 23256 37800
rect 24584 37791 24636 37800
rect 24584 37757 24593 37791
rect 24593 37757 24627 37791
rect 24627 37757 24636 37791
rect 24584 37748 24636 37757
rect 24952 37748 25004 37800
rect 25412 37791 25464 37800
rect 22100 37680 22152 37732
rect 22468 37723 22520 37732
rect 22468 37689 22477 37723
rect 22477 37689 22511 37723
rect 22511 37689 22520 37723
rect 22468 37680 22520 37689
rect 23572 37680 23624 37732
rect 22376 37612 22428 37664
rect 23664 37655 23716 37664
rect 23664 37621 23673 37655
rect 23673 37621 23707 37655
rect 23707 37621 23716 37655
rect 23664 37612 23716 37621
rect 25044 37723 25096 37732
rect 25044 37689 25053 37723
rect 25053 37689 25087 37723
rect 25087 37689 25096 37723
rect 25044 37680 25096 37689
rect 25412 37757 25446 37791
rect 25446 37757 25464 37791
rect 25412 37748 25464 37757
rect 25964 37748 26016 37800
rect 26148 37748 26200 37800
rect 26424 37612 26476 37664
rect 27068 37655 27120 37664
rect 27068 37621 27077 37655
rect 27077 37621 27111 37655
rect 27111 37621 27120 37655
rect 27068 37612 27120 37621
rect 28172 37748 28224 37800
rect 28724 37748 28776 37800
rect 29828 37952 29880 38004
rect 30288 37952 30340 38004
rect 31576 37952 31628 38004
rect 32496 37995 32548 38004
rect 32496 37961 32505 37995
rect 32505 37961 32539 37995
rect 32539 37961 32548 37995
rect 32496 37952 32548 37961
rect 32864 37952 32916 38004
rect 33324 37995 33376 38004
rect 33324 37961 33333 37995
rect 33333 37961 33367 37995
rect 33367 37961 33376 37995
rect 33324 37952 33376 37961
rect 36176 37952 36228 38004
rect 33232 37927 33284 37936
rect 33232 37893 33241 37927
rect 33241 37893 33275 37927
rect 33275 37893 33284 37927
rect 33232 37884 33284 37893
rect 29920 37859 29972 37868
rect 29920 37825 29929 37859
rect 29929 37825 29963 37859
rect 29963 37825 29972 37859
rect 29920 37816 29972 37825
rect 30748 37816 30800 37868
rect 36544 37859 36596 37868
rect 36544 37825 36553 37859
rect 36553 37825 36587 37859
rect 36587 37825 36596 37859
rect 36544 37816 36596 37825
rect 36728 37884 36780 37936
rect 37004 37884 37056 37936
rect 36820 37859 36872 37868
rect 36820 37825 36829 37859
rect 36829 37825 36863 37859
rect 36863 37825 36872 37859
rect 36820 37816 36872 37825
rect 37464 37995 37516 38004
rect 37464 37961 37489 37995
rect 37489 37961 37516 37995
rect 37464 37952 37516 37961
rect 37280 37927 37332 37936
rect 37280 37893 37289 37927
rect 37289 37893 37323 37927
rect 37323 37893 37332 37927
rect 37280 37884 37332 37893
rect 39580 37995 39632 38004
rect 39580 37961 39589 37995
rect 39589 37961 39623 37995
rect 39623 37961 39632 37995
rect 39580 37952 39632 37961
rect 38752 37816 38804 37868
rect 44180 37816 44232 37868
rect 32588 37748 32640 37800
rect 34428 37748 34480 37800
rect 38016 37748 38068 37800
rect 27896 37612 27948 37664
rect 28908 37612 28960 37664
rect 29000 37612 29052 37664
rect 29920 37612 29972 37664
rect 36176 37655 36228 37664
rect 36176 37621 36185 37655
rect 36185 37621 36219 37655
rect 36219 37621 36228 37655
rect 36176 37612 36228 37621
rect 37924 37680 37976 37732
rect 37648 37655 37700 37664
rect 37648 37621 37657 37655
rect 37657 37621 37691 37655
rect 37691 37621 37700 37655
rect 37648 37612 37700 37621
rect 46664 37655 46716 37664
rect 46664 37621 46673 37655
rect 46673 37621 46707 37655
rect 46707 37621 46716 37655
rect 46664 37612 46716 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 5264 37451 5316 37460
rect 5264 37417 5273 37451
rect 5273 37417 5307 37451
rect 5307 37417 5316 37451
rect 5264 37408 5316 37417
rect 3792 37315 3844 37324
rect 3792 37281 3801 37315
rect 3801 37281 3835 37315
rect 3835 37281 3844 37315
rect 3792 37272 3844 37281
rect 10508 37408 10560 37460
rect 6460 37340 6512 37392
rect 940 37204 992 37256
rect 4068 37247 4120 37256
rect 4068 37213 4102 37247
rect 4102 37213 4120 37247
rect 4068 37204 4120 37213
rect 5172 37204 5224 37256
rect 6276 37204 6328 37256
rect 6644 37204 6696 37256
rect 4712 37136 4764 37188
rect 5448 37136 5500 37188
rect 7196 37315 7248 37324
rect 7196 37281 7205 37315
rect 7205 37281 7239 37315
rect 7239 37281 7248 37315
rect 7196 37272 7248 37281
rect 9220 37340 9272 37392
rect 9496 37340 9548 37392
rect 8484 37272 8536 37324
rect 9312 37272 9364 37324
rect 9588 37315 9640 37324
rect 9588 37281 9597 37315
rect 9597 37281 9631 37315
rect 9631 37281 9640 37315
rect 9588 37272 9640 37281
rect 10692 37340 10744 37392
rect 13360 37408 13412 37460
rect 13912 37408 13964 37460
rect 14832 37408 14884 37460
rect 16212 37408 16264 37460
rect 19800 37408 19852 37460
rect 23204 37408 23256 37460
rect 25044 37408 25096 37460
rect 26148 37408 26200 37460
rect 26700 37408 26752 37460
rect 30748 37408 30800 37460
rect 19248 37340 19300 37392
rect 9956 37315 10008 37324
rect 9956 37281 9990 37315
rect 9990 37281 10008 37315
rect 9956 37272 10008 37281
rect 11244 37315 11296 37324
rect 11244 37281 11253 37315
rect 11253 37281 11287 37315
rect 11287 37281 11296 37315
rect 11244 37272 11296 37281
rect 12164 37315 12216 37324
rect 12164 37281 12173 37315
rect 12173 37281 12207 37315
rect 12207 37281 12216 37315
rect 12164 37272 12216 37281
rect 12256 37315 12308 37324
rect 12256 37281 12290 37315
rect 12290 37281 12308 37315
rect 12256 37272 12308 37281
rect 13084 37315 13136 37324
rect 13084 37281 13093 37315
rect 13093 37281 13127 37315
rect 13127 37281 13136 37315
rect 13084 37272 13136 37281
rect 7012 37247 7064 37256
rect 7012 37213 7021 37247
rect 7021 37213 7055 37247
rect 7055 37213 7064 37247
rect 7012 37204 7064 37213
rect 8760 37204 8812 37256
rect 10140 37247 10192 37256
rect 10140 37213 10149 37247
rect 10149 37213 10183 37247
rect 10183 37213 10192 37247
rect 10140 37204 10192 37213
rect 7104 37179 7156 37188
rect 7104 37145 7113 37179
rect 7113 37145 7147 37179
rect 7147 37145 7156 37179
rect 7104 37136 7156 37145
rect 2412 37068 2464 37120
rect 4436 37068 4488 37120
rect 5264 37068 5316 37120
rect 7288 37068 7340 37120
rect 7656 37111 7708 37120
rect 7656 37077 7665 37111
rect 7665 37077 7699 37111
rect 7699 37077 7708 37111
rect 7656 37068 7708 37077
rect 10968 37068 11020 37120
rect 12440 37247 12492 37256
rect 12440 37213 12449 37247
rect 12449 37213 12483 37247
rect 12483 37213 12492 37247
rect 12440 37204 12492 37213
rect 15936 37272 15988 37324
rect 17224 37272 17276 37324
rect 17776 37272 17828 37324
rect 21456 37272 21508 37324
rect 22836 37272 22888 37324
rect 24492 37272 24544 37324
rect 24584 37315 24636 37324
rect 24584 37281 24593 37315
rect 24593 37281 24627 37315
rect 24627 37281 24636 37315
rect 24584 37272 24636 37281
rect 25136 37272 25188 37324
rect 25320 37315 25372 37324
rect 25320 37281 25329 37315
rect 25329 37281 25363 37315
rect 25363 37281 25372 37315
rect 25320 37272 25372 37281
rect 25412 37315 25464 37324
rect 25412 37281 25446 37315
rect 25446 37281 25464 37315
rect 25412 37272 25464 37281
rect 26240 37315 26292 37324
rect 26240 37281 26249 37315
rect 26249 37281 26283 37315
rect 26283 37281 26292 37315
rect 26240 37272 26292 37281
rect 26792 37272 26844 37324
rect 14924 37204 14976 37256
rect 15660 37204 15712 37256
rect 20444 37204 20496 37256
rect 22192 37204 22244 37256
rect 22468 37204 22520 37256
rect 24124 37204 24176 37256
rect 25596 37247 25648 37256
rect 25596 37213 25605 37247
rect 25605 37213 25639 37247
rect 25639 37213 25648 37247
rect 25596 37204 25648 37213
rect 28080 37340 28132 37392
rect 35808 37340 35860 37392
rect 15292 37136 15344 37188
rect 20168 37136 20220 37188
rect 12532 37068 12584 37120
rect 14096 37068 14148 37120
rect 14280 37068 14332 37120
rect 14740 37111 14792 37120
rect 14740 37077 14749 37111
rect 14749 37077 14783 37111
rect 14783 37077 14792 37111
rect 14740 37068 14792 37077
rect 19524 37111 19576 37120
rect 19524 37077 19533 37111
rect 19533 37077 19567 37111
rect 19567 37077 19576 37111
rect 19524 37068 19576 37077
rect 23756 37068 23808 37120
rect 27620 37272 27672 37324
rect 27896 37272 27948 37324
rect 27988 37315 28040 37324
rect 27988 37281 27997 37315
rect 27997 37281 28031 37315
rect 28031 37281 28040 37315
rect 27988 37272 28040 37281
rect 28264 37315 28316 37324
rect 28264 37281 28273 37315
rect 28273 37281 28307 37315
rect 28307 37281 28316 37315
rect 28264 37272 28316 37281
rect 28356 37315 28408 37324
rect 28356 37281 28390 37315
rect 28390 37281 28408 37315
rect 28356 37272 28408 37281
rect 28724 37272 28776 37324
rect 29184 37315 29236 37324
rect 29184 37281 29193 37315
rect 29193 37281 29227 37315
rect 29227 37281 29236 37315
rect 29184 37272 29236 37281
rect 31668 37272 31720 37324
rect 28540 37247 28592 37256
rect 28540 37213 28549 37247
rect 28549 37213 28583 37247
rect 28583 37213 28592 37247
rect 28540 37204 28592 37213
rect 29920 37247 29972 37256
rect 29920 37213 29929 37247
rect 29929 37213 29963 37247
rect 29963 37213 29972 37247
rect 29920 37204 29972 37213
rect 33140 37204 33192 37256
rect 34428 37204 34480 37256
rect 36728 37247 36780 37256
rect 36728 37213 36737 37247
rect 36737 37213 36771 37247
rect 36771 37213 36780 37247
rect 36728 37204 36780 37213
rect 37372 37204 37424 37256
rect 27712 37068 27764 37120
rect 28356 37068 28408 37120
rect 34520 37136 34572 37188
rect 37188 37136 37240 37188
rect 36084 37111 36136 37120
rect 36084 37077 36093 37111
rect 36093 37077 36127 37111
rect 36127 37077 36136 37111
rect 36084 37068 36136 37077
rect 36544 37111 36596 37120
rect 36544 37077 36559 37111
rect 36559 37077 36593 37111
rect 36593 37077 36596 37111
rect 36544 37068 36596 37077
rect 38568 37068 38620 37120
rect 38844 37111 38896 37120
rect 38844 37077 38853 37111
rect 38853 37077 38887 37111
rect 38887 37077 38896 37111
rect 38844 37068 38896 37077
rect 39212 37111 39264 37120
rect 39212 37077 39221 37111
rect 39221 37077 39255 37111
rect 39255 37077 39264 37111
rect 39212 37068 39264 37077
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 3700 36864 3752 36916
rect 4436 36907 4488 36916
rect 4436 36873 4445 36907
rect 4445 36873 4479 36907
rect 4479 36873 4488 36907
rect 4436 36864 4488 36873
rect 5264 36864 5316 36916
rect 6644 36907 6696 36916
rect 6644 36873 6653 36907
rect 6653 36873 6687 36907
rect 6687 36873 6696 36907
rect 6644 36864 6696 36873
rect 7748 36864 7800 36916
rect 10324 36864 10376 36916
rect 12440 36864 12492 36916
rect 16488 36864 16540 36916
rect 16856 36864 16908 36916
rect 7104 36839 7156 36848
rect 7104 36805 7113 36839
rect 7113 36805 7147 36839
rect 7147 36805 7156 36839
rect 7104 36796 7156 36805
rect 7288 36796 7340 36848
rect 14464 36796 14516 36848
rect 16764 36796 16816 36848
rect 6920 36728 6972 36780
rect 10140 36728 10192 36780
rect 12992 36728 13044 36780
rect 16488 36775 16540 36780
rect 16488 36741 16505 36775
rect 16505 36741 16539 36775
rect 16539 36741 16540 36775
rect 16488 36728 16540 36741
rect 5448 36660 5500 36712
rect 8208 36660 8260 36712
rect 15844 36660 15896 36712
rect 17960 36728 18012 36780
rect 19156 36660 19208 36712
rect 20352 36660 20404 36712
rect 27068 36796 27120 36848
rect 23756 36728 23808 36780
rect 26976 36771 27028 36780
rect 26976 36737 26985 36771
rect 26985 36737 27019 36771
rect 27019 36737 27028 36771
rect 26976 36728 27028 36737
rect 28264 36864 28316 36916
rect 28080 36796 28132 36848
rect 30288 36839 30340 36848
rect 30288 36805 30297 36839
rect 30297 36805 30331 36839
rect 30331 36805 30340 36839
rect 30288 36796 30340 36805
rect 32404 36864 32456 36916
rect 32864 36864 32916 36916
rect 34520 36907 34572 36916
rect 34520 36873 34529 36907
rect 34529 36873 34563 36907
rect 34563 36873 34572 36907
rect 34520 36864 34572 36873
rect 32036 36796 32088 36848
rect 33508 36796 33560 36848
rect 34244 36796 34296 36848
rect 36084 36864 36136 36916
rect 36452 36864 36504 36916
rect 38844 36864 38896 36916
rect 44180 36864 44232 36916
rect 31576 36728 31628 36780
rect 31668 36728 31720 36780
rect 34612 36728 34664 36780
rect 34796 36771 34848 36780
rect 34796 36737 34805 36771
rect 34805 36737 34839 36771
rect 34839 36737 34848 36771
rect 34796 36728 34848 36737
rect 22008 36660 22060 36712
rect 35440 36728 35492 36780
rect 36912 36796 36964 36848
rect 39212 36796 39264 36848
rect 36176 36728 36228 36780
rect 15660 36592 15712 36644
rect 16488 36592 16540 36644
rect 19432 36592 19484 36644
rect 29276 36592 29328 36644
rect 16764 36524 16816 36576
rect 19708 36567 19760 36576
rect 19708 36533 19717 36567
rect 19717 36533 19751 36567
rect 19751 36533 19760 36567
rect 19708 36524 19760 36533
rect 34060 36524 34112 36576
rect 34520 36592 34572 36644
rect 35992 36592 36044 36644
rect 37648 36728 37700 36780
rect 38016 36728 38068 36780
rect 38660 36660 38712 36712
rect 36636 36524 36688 36576
rect 46848 36524 46900 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2136 36184 2188 36236
rect 7196 36184 7248 36236
rect 7656 36184 7708 36236
rect 9680 36184 9732 36236
rect 10508 36184 10560 36236
rect 15200 36184 15252 36236
rect 15844 36184 15896 36236
rect 19432 36320 19484 36372
rect 19524 36320 19576 36372
rect 18512 36252 18564 36304
rect 18696 36295 18748 36304
rect 18696 36261 18705 36295
rect 18705 36261 18739 36295
rect 18739 36261 18748 36295
rect 18696 36252 18748 36261
rect 20444 36252 20496 36304
rect 22100 36252 22152 36304
rect 16580 36227 16632 36236
rect 16580 36193 16614 36227
rect 16614 36193 16632 36227
rect 16580 36184 16632 36193
rect 3976 36116 4028 36168
rect 5264 36116 5316 36168
rect 9956 36116 10008 36168
rect 13728 36116 13780 36168
rect 9312 36048 9364 36100
rect 3332 35980 3384 36032
rect 4160 36023 4212 36032
rect 4160 35989 4169 36023
rect 4169 35989 4203 36023
rect 4203 35989 4212 36023
rect 4160 35980 4212 35989
rect 4528 35980 4580 36032
rect 5356 35980 5408 36032
rect 9588 35980 9640 36032
rect 11060 36023 11112 36032
rect 11060 35989 11069 36023
rect 11069 35989 11103 36023
rect 11103 35989 11112 36023
rect 11060 35980 11112 35989
rect 14096 36048 14148 36100
rect 14280 36023 14332 36032
rect 14280 35989 14289 36023
rect 14289 35989 14323 36023
rect 14323 35989 14332 36023
rect 14280 35980 14332 35989
rect 15476 36116 15528 36168
rect 16488 36159 16540 36168
rect 16488 36125 16497 36159
rect 16497 36125 16531 36159
rect 16531 36125 16540 36159
rect 16488 36116 16540 36125
rect 19616 36184 19668 36236
rect 18236 36116 18288 36168
rect 19340 36116 19392 36168
rect 19524 36116 19576 36168
rect 19892 36159 19944 36168
rect 19892 36125 19901 36159
rect 19901 36125 19935 36159
rect 19935 36125 19944 36159
rect 19892 36116 19944 36125
rect 18604 36048 18656 36100
rect 18788 36023 18840 36032
rect 18788 35989 18797 36023
rect 18797 35989 18831 36023
rect 18831 35989 18840 36023
rect 18788 35980 18840 35989
rect 19248 36048 19300 36100
rect 20260 36116 20312 36168
rect 20628 36116 20680 36168
rect 22008 36116 22060 36168
rect 22560 36227 22612 36236
rect 22560 36193 22569 36227
rect 22569 36193 22603 36227
rect 22603 36193 22612 36227
rect 22560 36184 22612 36193
rect 29092 36320 29144 36372
rect 23020 36295 23072 36304
rect 23020 36261 23029 36295
rect 23029 36261 23063 36295
rect 23063 36261 23072 36295
rect 23020 36252 23072 36261
rect 23664 36295 23716 36304
rect 23664 36261 23673 36295
rect 23673 36261 23707 36295
rect 23707 36261 23716 36295
rect 23664 36252 23716 36261
rect 23204 36184 23256 36236
rect 25504 36184 25556 36236
rect 25688 36184 25740 36236
rect 32312 36320 32364 36372
rect 34060 36320 34112 36372
rect 34612 36320 34664 36372
rect 36176 36320 36228 36372
rect 37648 36320 37700 36372
rect 38660 36320 38712 36372
rect 39028 36320 39080 36372
rect 26056 36116 26108 36168
rect 29276 36159 29328 36168
rect 29276 36125 29285 36159
rect 29285 36125 29319 36159
rect 29319 36125 29328 36159
rect 29276 36116 29328 36125
rect 23388 36048 23440 36100
rect 22284 36023 22336 36032
rect 22284 35989 22293 36023
rect 22293 35989 22327 36023
rect 22327 35989 22336 36023
rect 22284 35980 22336 35989
rect 23480 35980 23532 36032
rect 26148 35980 26200 36032
rect 29460 36048 29512 36100
rect 32496 36252 32548 36304
rect 33416 36252 33468 36304
rect 32404 36227 32456 36236
rect 32404 36193 32413 36227
rect 32413 36193 32447 36227
rect 32447 36193 32456 36227
rect 32404 36184 32456 36193
rect 32680 36227 32732 36236
rect 32680 36193 32689 36227
rect 32689 36193 32723 36227
rect 32723 36193 32732 36227
rect 32680 36184 32732 36193
rect 32772 36184 32824 36236
rect 33140 36184 33192 36236
rect 33508 36184 33560 36236
rect 34612 36184 34664 36236
rect 32128 36116 32180 36168
rect 32956 36159 33008 36168
rect 32956 36125 32965 36159
rect 32965 36125 32999 36159
rect 32999 36125 33008 36159
rect 32956 36116 33008 36125
rect 36544 36252 36596 36304
rect 35992 36159 36044 36168
rect 35992 36125 36001 36159
rect 36001 36125 36035 36159
rect 36035 36125 36044 36159
rect 35992 36116 36044 36125
rect 36268 36159 36320 36168
rect 36268 36125 36277 36159
rect 36277 36125 36311 36159
rect 36311 36125 36320 36159
rect 36268 36116 36320 36125
rect 34060 36091 34112 36100
rect 34060 36057 34069 36091
rect 34069 36057 34103 36091
rect 34103 36057 34112 36091
rect 34060 36048 34112 36057
rect 36820 36159 36872 36168
rect 36820 36125 36829 36159
rect 36829 36125 36863 36159
rect 36863 36125 36872 36159
rect 36820 36116 36872 36125
rect 37372 36159 37424 36168
rect 37372 36125 37381 36159
rect 37381 36125 37415 36159
rect 37415 36125 37424 36159
rect 37372 36116 37424 36125
rect 34152 36023 34204 36032
rect 34152 35989 34161 36023
rect 34161 35989 34195 36023
rect 34195 35989 34204 36023
rect 34152 35980 34204 35989
rect 35992 35980 36044 36032
rect 36360 36023 36412 36032
rect 36360 35989 36369 36023
rect 36369 35989 36403 36023
rect 36403 35989 36412 36023
rect 36360 35980 36412 35989
rect 36544 35980 36596 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 4160 35776 4212 35828
rect 5264 35776 5316 35828
rect 3332 35640 3384 35692
rect 3792 35683 3844 35692
rect 3792 35649 3801 35683
rect 3801 35649 3835 35683
rect 3835 35649 3844 35683
rect 3792 35640 3844 35649
rect 4620 35640 4672 35692
rect 5264 35683 5316 35692
rect 5264 35649 5298 35683
rect 5298 35649 5316 35683
rect 5264 35640 5316 35649
rect 2136 35615 2188 35624
rect 2136 35581 2145 35615
rect 2145 35581 2179 35615
rect 2179 35581 2188 35615
rect 2136 35572 2188 35581
rect 4528 35572 4580 35624
rect 4988 35572 5040 35624
rect 5172 35615 5224 35624
rect 5172 35581 5181 35615
rect 5181 35581 5215 35615
rect 5215 35581 5224 35615
rect 5172 35572 5224 35581
rect 5632 35572 5684 35624
rect 10324 35776 10376 35828
rect 13084 35776 13136 35828
rect 9312 35708 9364 35760
rect 7932 35640 7984 35692
rect 8944 35640 8996 35692
rect 7656 35615 7708 35624
rect 7656 35581 7665 35615
rect 7665 35581 7699 35615
rect 7699 35581 7708 35615
rect 7656 35572 7708 35581
rect 4712 35504 4764 35556
rect 3608 35479 3660 35488
rect 3608 35445 3617 35479
rect 3617 35445 3651 35479
rect 3651 35445 3660 35479
rect 3608 35436 3660 35445
rect 4896 35436 4948 35488
rect 9128 35504 9180 35556
rect 6092 35479 6144 35488
rect 6092 35445 6101 35479
rect 6101 35445 6135 35479
rect 6135 35445 6144 35479
rect 6092 35436 6144 35445
rect 6828 35479 6880 35488
rect 6828 35445 6837 35479
rect 6837 35445 6871 35479
rect 6871 35445 6880 35479
rect 6828 35436 6880 35445
rect 8300 35436 8352 35488
rect 9588 35683 9640 35692
rect 9588 35649 9597 35683
rect 9597 35649 9631 35683
rect 9631 35649 9640 35683
rect 9588 35640 9640 35649
rect 13820 35708 13872 35760
rect 15476 35776 15528 35828
rect 15568 35776 15620 35828
rect 16488 35776 16540 35828
rect 17960 35776 18012 35828
rect 12440 35572 12492 35624
rect 15568 35683 15620 35692
rect 15568 35649 15577 35683
rect 15577 35649 15611 35683
rect 15611 35649 15620 35683
rect 15568 35640 15620 35649
rect 15660 35683 15712 35692
rect 17408 35708 17460 35760
rect 15660 35649 15694 35683
rect 15694 35649 15712 35683
rect 15660 35640 15712 35649
rect 16764 35640 16816 35692
rect 18052 35640 18104 35692
rect 19432 35683 19484 35692
rect 19432 35649 19441 35683
rect 19441 35649 19475 35683
rect 19475 35649 19484 35683
rect 19432 35640 19484 35649
rect 19708 35683 19760 35692
rect 19708 35649 19717 35683
rect 19717 35649 19751 35683
rect 19751 35649 19760 35683
rect 19708 35640 19760 35649
rect 19892 35640 19944 35692
rect 20076 35640 20128 35692
rect 20168 35683 20220 35692
rect 20168 35649 20177 35683
rect 20177 35649 20211 35683
rect 20211 35649 20220 35683
rect 20168 35640 20220 35649
rect 22008 35776 22060 35828
rect 22284 35776 22336 35828
rect 25044 35776 25096 35828
rect 25320 35776 25372 35828
rect 22100 35751 22152 35760
rect 22100 35717 22134 35751
rect 22134 35717 22152 35751
rect 22100 35708 22152 35717
rect 23756 35751 23808 35760
rect 23756 35717 23765 35751
rect 23765 35717 23799 35751
rect 23799 35717 23808 35751
rect 23756 35708 23808 35717
rect 9588 35504 9640 35556
rect 14740 35572 14792 35624
rect 15200 35572 15252 35624
rect 15844 35615 15896 35624
rect 15844 35581 15853 35615
rect 15853 35581 15887 35615
rect 15887 35581 15896 35615
rect 15844 35572 15896 35581
rect 9956 35436 10008 35488
rect 11060 35479 11112 35488
rect 11060 35445 11069 35479
rect 11069 35445 11103 35479
rect 11103 35445 11112 35479
rect 11060 35436 11112 35445
rect 13084 35479 13136 35488
rect 13084 35445 13093 35479
rect 13093 35445 13127 35479
rect 13127 35445 13136 35479
rect 13084 35436 13136 35445
rect 14372 35436 14424 35488
rect 15292 35547 15344 35556
rect 15292 35513 15301 35547
rect 15301 35513 15335 35547
rect 15335 35513 15344 35547
rect 15292 35504 15344 35513
rect 18512 35615 18564 35624
rect 18512 35581 18521 35615
rect 18521 35581 18555 35615
rect 18555 35581 18564 35615
rect 18512 35572 18564 35581
rect 19156 35615 19208 35624
rect 19156 35581 19165 35615
rect 19165 35581 19199 35615
rect 19199 35581 19208 35615
rect 19156 35572 19208 35581
rect 21916 35640 21968 35692
rect 20628 35572 20680 35624
rect 21088 35572 21140 35624
rect 21456 35615 21508 35624
rect 21456 35581 21465 35615
rect 21465 35581 21499 35615
rect 21499 35581 21508 35615
rect 21456 35572 21508 35581
rect 21732 35572 21784 35624
rect 20444 35504 20496 35556
rect 20812 35504 20864 35556
rect 23848 35615 23900 35624
rect 23848 35581 23857 35615
rect 23857 35581 23891 35615
rect 23891 35581 23900 35615
rect 23848 35572 23900 35581
rect 24216 35572 24268 35624
rect 25044 35683 25096 35692
rect 25044 35649 25053 35683
rect 25053 35649 25087 35683
rect 25087 35649 25096 35683
rect 25044 35640 25096 35649
rect 24676 35572 24728 35624
rect 25228 35572 25280 35624
rect 25504 35572 25556 35624
rect 26148 35708 26200 35760
rect 26056 35640 26108 35692
rect 26148 35615 26200 35624
rect 26148 35581 26157 35615
rect 26157 35581 26191 35615
rect 26191 35581 26200 35615
rect 26148 35572 26200 35581
rect 19524 35436 19576 35488
rect 19800 35479 19852 35488
rect 19800 35445 19809 35479
rect 19809 35445 19843 35479
rect 19843 35445 19852 35479
rect 19800 35436 19852 35445
rect 20904 35436 20956 35488
rect 22192 35436 22244 35488
rect 24032 35436 24084 35488
rect 24124 35436 24176 35488
rect 26424 35547 26476 35556
rect 26424 35513 26433 35547
rect 26433 35513 26467 35547
rect 26467 35513 26476 35547
rect 26424 35504 26476 35513
rect 27252 35683 27304 35692
rect 27252 35649 27261 35683
rect 27261 35649 27295 35683
rect 27295 35649 27304 35683
rect 27252 35640 27304 35649
rect 30932 35776 30984 35828
rect 27896 35708 27948 35760
rect 36268 35776 36320 35828
rect 36636 35776 36688 35828
rect 36820 35776 36872 35828
rect 36360 35708 36412 35760
rect 29092 35640 29144 35692
rect 29552 35640 29604 35692
rect 30288 35640 30340 35692
rect 32128 35683 32180 35692
rect 32128 35649 32137 35683
rect 32137 35649 32171 35683
rect 32171 35649 32180 35683
rect 32128 35640 32180 35649
rect 32312 35683 32364 35692
rect 32312 35649 32321 35683
rect 32321 35649 32355 35683
rect 32355 35649 32364 35683
rect 32312 35640 32364 35649
rect 33140 35683 33192 35692
rect 33140 35649 33174 35683
rect 33174 35649 33192 35683
rect 33140 35640 33192 35649
rect 40040 35683 40092 35692
rect 40040 35649 40049 35683
rect 40049 35649 40083 35683
rect 40083 35649 40092 35683
rect 40040 35640 40092 35649
rect 46848 35640 46900 35692
rect 26976 35615 27028 35624
rect 26976 35581 26985 35615
rect 26985 35581 27019 35615
rect 27019 35581 27028 35615
rect 26976 35572 27028 35581
rect 28908 35572 28960 35624
rect 31392 35572 31444 35624
rect 32680 35572 32732 35624
rect 33324 35615 33376 35624
rect 33324 35581 33333 35615
rect 33333 35581 33367 35615
rect 33367 35581 33376 35615
rect 33324 35572 33376 35581
rect 30564 35504 30616 35556
rect 26884 35436 26936 35488
rect 29000 35436 29052 35488
rect 29736 35436 29788 35488
rect 39764 35615 39816 35624
rect 39764 35581 39773 35615
rect 39773 35581 39807 35615
rect 39807 35581 39816 35615
rect 39764 35572 39816 35581
rect 35992 35436 36044 35488
rect 41236 35436 41288 35488
rect 46664 35479 46716 35488
rect 46664 35445 46673 35479
rect 46673 35445 46707 35479
rect 46707 35445 46716 35479
rect 46664 35436 46716 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4528 35232 4580 35284
rect 4988 35232 5040 35284
rect 6092 35232 6144 35284
rect 3424 35164 3476 35216
rect 4620 35096 4672 35148
rect 4896 35139 4948 35148
rect 4896 35105 4905 35139
rect 4905 35105 4939 35139
rect 4939 35105 4948 35139
rect 4896 35096 4948 35105
rect 7932 35207 7984 35216
rect 7932 35173 7941 35207
rect 7941 35173 7975 35207
rect 7975 35173 7984 35207
rect 7932 35164 7984 35173
rect 8944 35275 8996 35284
rect 8944 35241 8953 35275
rect 8953 35241 8987 35275
rect 8987 35241 8996 35275
rect 8944 35232 8996 35241
rect 10692 35207 10744 35216
rect 10692 35173 10707 35207
rect 10707 35173 10741 35207
rect 10741 35173 10744 35207
rect 10692 35164 10744 35173
rect 5172 35139 5224 35148
rect 5172 35105 5181 35139
rect 5181 35105 5215 35139
rect 5215 35105 5224 35139
rect 5172 35096 5224 35105
rect 5264 35139 5316 35148
rect 5264 35105 5298 35139
rect 5298 35105 5316 35139
rect 5264 35096 5316 35105
rect 1768 35028 1820 35080
rect 2136 35071 2188 35080
rect 2136 35037 2145 35071
rect 2145 35037 2179 35071
rect 2179 35037 2188 35071
rect 2136 35028 2188 35037
rect 3608 35028 3660 35080
rect 6092 35139 6144 35148
rect 6092 35105 6101 35139
rect 6101 35105 6135 35139
rect 6135 35105 6144 35139
rect 6092 35096 6144 35105
rect 8208 35096 8260 35148
rect 8668 35096 8720 35148
rect 9220 35096 9272 35148
rect 10324 35096 10376 35148
rect 13728 35232 13780 35284
rect 18788 35232 18840 35284
rect 19800 35232 19852 35284
rect 17316 35164 17368 35216
rect 19616 35207 19668 35216
rect 19616 35173 19625 35207
rect 19625 35173 19659 35207
rect 19659 35173 19668 35207
rect 19616 35164 19668 35173
rect 13084 35096 13136 35148
rect 6552 35071 6604 35080
rect 6552 35037 6561 35071
rect 6561 35037 6595 35071
rect 6595 35037 6604 35071
rect 6552 35028 6604 35037
rect 6828 35071 6880 35080
rect 6828 35037 6862 35071
rect 6862 35037 6880 35071
rect 6828 35028 6880 35037
rect 9404 35028 9456 35080
rect 4712 34892 4764 34944
rect 5540 34892 5592 34944
rect 6276 34935 6328 34944
rect 6276 34901 6285 34935
rect 6285 34901 6319 34935
rect 6319 34901 6328 34935
rect 6276 34892 6328 34901
rect 6920 34892 6972 34944
rect 8392 35003 8444 35012
rect 8392 34969 8401 35003
rect 8401 34969 8435 35003
rect 8435 34969 8444 35003
rect 8392 34960 8444 34969
rect 9496 34960 9548 35012
rect 9680 34960 9732 35012
rect 10968 35071 11020 35080
rect 10968 35037 10977 35071
rect 10977 35037 11011 35071
rect 11011 35037 11020 35071
rect 10968 35028 11020 35037
rect 11244 35071 11296 35080
rect 11244 35037 11253 35071
rect 11253 35037 11287 35071
rect 11287 35037 11296 35071
rect 11244 35028 11296 35037
rect 12440 35071 12492 35080
rect 12440 35037 12449 35071
rect 12449 35037 12483 35071
rect 12483 35037 12492 35071
rect 12440 35028 12492 35037
rect 9312 34892 9364 34944
rect 11796 34960 11848 35012
rect 13636 35071 13688 35080
rect 13636 35037 13645 35071
rect 13645 35037 13679 35071
rect 13679 35037 13688 35071
rect 13636 35028 13688 35037
rect 14372 35071 14424 35080
rect 14372 35037 14381 35071
rect 14381 35037 14415 35071
rect 14415 35037 14424 35071
rect 14372 35028 14424 35037
rect 14740 35096 14792 35148
rect 17684 35071 17736 35080
rect 17684 35037 17693 35071
rect 17693 35037 17727 35071
rect 17727 35037 17736 35071
rect 17684 35028 17736 35037
rect 18512 35028 18564 35080
rect 19984 35096 20036 35148
rect 20352 35207 20404 35216
rect 20352 35173 20361 35207
rect 20361 35173 20395 35207
rect 20395 35173 20404 35207
rect 20352 35164 20404 35173
rect 21916 35164 21968 35216
rect 20444 35096 20496 35148
rect 20812 35139 20864 35148
rect 20812 35105 20821 35139
rect 20821 35105 20855 35139
rect 20855 35105 20864 35139
rect 20812 35096 20864 35105
rect 23480 35275 23532 35284
rect 23480 35241 23489 35275
rect 23489 35241 23523 35275
rect 23523 35241 23532 35275
rect 23480 35232 23532 35241
rect 27252 35232 27304 35284
rect 29092 35232 29144 35284
rect 29276 35232 29328 35284
rect 29552 35275 29604 35284
rect 29552 35241 29561 35275
rect 29561 35241 29595 35275
rect 29595 35241 29604 35275
rect 29552 35232 29604 35241
rect 37372 35275 37424 35284
rect 37372 35241 37381 35275
rect 37381 35241 37415 35275
rect 37415 35241 37424 35275
rect 37372 35232 37424 35241
rect 24400 35139 24452 35148
rect 24400 35105 24409 35139
rect 24409 35105 24443 35139
rect 24443 35105 24452 35139
rect 24400 35096 24452 35105
rect 25044 35139 25096 35148
rect 14096 35003 14148 35012
rect 14096 34969 14105 35003
rect 14105 34969 14139 35003
rect 14139 34969 14148 35003
rect 14096 34960 14148 34969
rect 18328 34960 18380 35012
rect 11060 34892 11112 34944
rect 11520 34892 11572 34944
rect 13820 34892 13872 34944
rect 16028 34892 16080 34944
rect 19984 34960 20036 35012
rect 20904 35028 20956 35080
rect 22744 35028 22796 35080
rect 23296 35071 23348 35080
rect 23296 35037 23305 35071
rect 23305 35037 23339 35071
rect 23339 35037 23348 35071
rect 23296 35028 23348 35037
rect 24032 35071 24084 35080
rect 24032 35037 24041 35071
rect 24041 35037 24075 35071
rect 24075 35037 24084 35071
rect 24032 35028 24084 35037
rect 24216 35028 24268 35080
rect 25044 35105 25053 35139
rect 25053 35105 25087 35139
rect 25087 35105 25096 35139
rect 25044 35096 25096 35105
rect 26884 35164 26936 35216
rect 24768 35028 24820 35080
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 25412 35071 25464 35080
rect 25412 35037 25446 35071
rect 25446 35037 25464 35071
rect 25412 35028 25464 35037
rect 25596 35071 25648 35080
rect 25596 35037 25605 35071
rect 25605 35037 25639 35071
rect 25639 35037 25648 35071
rect 25596 35028 25648 35037
rect 26792 35028 26844 35080
rect 27712 35071 27764 35080
rect 27712 35037 27721 35071
rect 27721 35037 27755 35071
rect 27755 35037 27764 35071
rect 27712 35028 27764 35037
rect 27896 35071 27948 35080
rect 27896 35037 27905 35071
rect 27905 35037 27939 35071
rect 27939 35037 27948 35071
rect 27896 35028 27948 35037
rect 28080 35028 28132 35080
rect 28724 35028 28776 35080
rect 28908 35028 28960 35080
rect 29000 35071 29052 35080
rect 29000 35037 29009 35071
rect 29009 35037 29043 35071
rect 29043 35037 29052 35071
rect 29000 35028 29052 35037
rect 29092 35071 29144 35080
rect 29092 35037 29101 35071
rect 29101 35037 29135 35071
rect 29135 35037 29144 35071
rect 29092 35028 29144 35037
rect 30656 35164 30708 35216
rect 30564 35139 30616 35148
rect 30564 35105 30573 35139
rect 30573 35105 30607 35139
rect 30607 35105 30616 35139
rect 30564 35096 30616 35105
rect 30840 35139 30892 35148
rect 30840 35105 30849 35139
rect 30849 35105 30883 35139
rect 30883 35105 30892 35139
rect 30840 35096 30892 35105
rect 30932 35139 30984 35148
rect 30932 35105 30966 35139
rect 30966 35105 30984 35139
rect 30932 35096 30984 35105
rect 33324 35096 33376 35148
rect 29736 35071 29788 35080
rect 29736 35037 29745 35071
rect 29745 35037 29779 35071
rect 29779 35037 29788 35071
rect 29736 35028 29788 35037
rect 29920 35071 29972 35080
rect 29920 35037 29929 35071
rect 29929 35037 29963 35071
rect 29963 35037 29972 35071
rect 29920 35028 29972 35037
rect 30288 35028 30340 35080
rect 31116 35071 31168 35080
rect 31116 35037 31125 35071
rect 31125 35037 31159 35071
rect 31159 35037 31168 35071
rect 31116 35028 31168 35037
rect 33600 35028 33652 35080
rect 34244 35071 34296 35080
rect 34244 35037 34253 35071
rect 34253 35037 34287 35071
rect 34287 35037 34296 35071
rect 34244 35028 34296 35037
rect 19064 34935 19116 34944
rect 19064 34901 19073 34935
rect 19073 34901 19107 34935
rect 19107 34901 19116 34935
rect 19064 34892 19116 34901
rect 20536 34892 20588 34944
rect 23020 34935 23072 34944
rect 23020 34901 23029 34935
rect 23029 34901 23063 34935
rect 23063 34901 23072 34935
rect 23020 34892 23072 34901
rect 23940 34892 23992 34944
rect 25872 34892 25924 34944
rect 27804 34960 27856 35012
rect 34980 35071 35032 35080
rect 34980 35037 34989 35071
rect 34989 35037 35023 35071
rect 35023 35037 35032 35071
rect 34980 35028 35032 35037
rect 35992 35071 36044 35080
rect 35992 35037 36001 35071
rect 36001 35037 36035 35071
rect 36035 35037 36044 35071
rect 35992 35028 36044 35037
rect 36544 35028 36596 35080
rect 39028 35028 39080 35080
rect 39764 35028 39816 35080
rect 40132 35071 40184 35080
rect 40132 35037 40141 35071
rect 40141 35037 40175 35071
rect 40175 35037 40184 35071
rect 40132 35028 40184 35037
rect 36636 34960 36688 35012
rect 27712 34892 27764 34944
rect 29552 34892 29604 34944
rect 29736 34892 29788 34944
rect 34428 34935 34480 34944
rect 34428 34901 34437 34935
rect 34437 34901 34471 34935
rect 34471 34901 34480 34935
rect 34428 34892 34480 34901
rect 37832 34892 37884 34944
rect 38384 34935 38436 34944
rect 38384 34901 38393 34935
rect 38393 34901 38427 34935
rect 38427 34901 38436 34935
rect 38384 34892 38436 34901
rect 41420 34892 41472 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 3792 34688 3844 34740
rect 8392 34688 8444 34740
rect 9404 34731 9456 34740
rect 9404 34697 9413 34731
rect 9413 34697 9447 34731
rect 9447 34697 9456 34731
rect 9404 34688 9456 34697
rect 9496 34688 9548 34740
rect 10416 34688 10468 34740
rect 10968 34688 11020 34740
rect 11796 34688 11848 34740
rect 14188 34688 14240 34740
rect 1492 34663 1544 34672
rect 1492 34629 1501 34663
rect 1501 34629 1535 34663
rect 1535 34629 1544 34663
rect 1492 34620 1544 34629
rect 3424 34663 3476 34672
rect 3424 34629 3433 34663
rect 3433 34629 3467 34663
rect 3467 34629 3476 34663
rect 3424 34620 3476 34629
rect 5356 34620 5408 34672
rect 6276 34620 6328 34672
rect 8024 34620 8076 34672
rect 6552 34595 6604 34604
rect 6552 34561 6561 34595
rect 6561 34561 6595 34595
rect 6595 34561 6604 34595
rect 6552 34552 6604 34561
rect 8300 34595 8352 34604
rect 8300 34561 8334 34595
rect 8334 34561 8352 34595
rect 8300 34552 8352 34561
rect 16028 34620 16080 34672
rect 17316 34688 17368 34740
rect 18512 34620 18564 34672
rect 19064 34620 19116 34672
rect 23296 34688 23348 34740
rect 26240 34688 26292 34740
rect 29092 34688 29144 34740
rect 29736 34731 29788 34740
rect 29736 34697 29745 34731
rect 29745 34697 29779 34731
rect 29779 34697 29788 34731
rect 29736 34688 29788 34697
rect 9680 34595 9732 34604
rect 9680 34561 9689 34595
rect 9689 34561 9723 34595
rect 9723 34561 9732 34595
rect 9680 34552 9732 34561
rect 10416 34595 10468 34604
rect 10416 34561 10425 34595
rect 10425 34561 10459 34595
rect 10459 34561 10468 34595
rect 10416 34552 10468 34561
rect 3700 34416 3752 34468
rect 1584 34391 1636 34400
rect 1584 34357 1593 34391
rect 1593 34357 1627 34391
rect 1627 34357 1636 34391
rect 1584 34348 1636 34357
rect 3976 34348 4028 34400
rect 10140 34527 10192 34536
rect 10140 34493 10149 34527
rect 10149 34493 10183 34527
rect 10183 34493 10192 34527
rect 10140 34484 10192 34493
rect 10232 34484 10284 34536
rect 10692 34527 10744 34536
rect 10692 34493 10701 34527
rect 10701 34493 10735 34527
rect 10735 34493 10744 34527
rect 10692 34484 10744 34493
rect 10876 34484 10928 34536
rect 13360 34595 13412 34604
rect 13360 34561 13394 34595
rect 13394 34561 13412 34595
rect 13360 34552 13412 34561
rect 15016 34595 15068 34604
rect 15016 34561 15025 34595
rect 15025 34561 15059 34595
rect 15059 34561 15068 34595
rect 15016 34552 15068 34561
rect 16304 34595 16356 34604
rect 16304 34561 16313 34595
rect 16313 34561 16347 34595
rect 16347 34561 16356 34595
rect 16304 34552 16356 34561
rect 11520 34484 11572 34536
rect 12440 34484 12492 34536
rect 12624 34484 12676 34536
rect 14096 34484 14148 34536
rect 15108 34527 15160 34536
rect 15108 34493 15117 34527
rect 15117 34493 15151 34527
rect 15151 34493 15160 34527
rect 15108 34484 15160 34493
rect 17684 34552 17736 34604
rect 20352 34552 20404 34604
rect 23296 34552 23348 34604
rect 23940 34595 23992 34604
rect 23940 34561 23974 34595
rect 23974 34561 23992 34595
rect 23940 34552 23992 34561
rect 25688 34595 25740 34604
rect 25688 34561 25697 34595
rect 25697 34561 25731 34595
rect 25731 34561 25740 34595
rect 25688 34552 25740 34561
rect 18696 34484 18748 34536
rect 23664 34527 23716 34536
rect 23664 34493 23673 34527
rect 23673 34493 23707 34527
rect 23707 34493 23716 34527
rect 23664 34484 23716 34493
rect 24768 34484 24820 34536
rect 23572 34416 23624 34468
rect 25780 34527 25832 34536
rect 25780 34493 25789 34527
rect 25789 34493 25823 34527
rect 25823 34493 25832 34527
rect 25780 34484 25832 34493
rect 37096 34688 37148 34740
rect 37556 34688 37608 34740
rect 37832 34688 37884 34740
rect 38016 34688 38068 34740
rect 39580 34688 39632 34740
rect 44180 34688 44232 34740
rect 9404 34348 9456 34400
rect 14556 34391 14608 34400
rect 14556 34357 14565 34391
rect 14565 34357 14599 34391
rect 14599 34357 14608 34391
rect 14556 34348 14608 34357
rect 16672 34348 16724 34400
rect 18512 34348 18564 34400
rect 22652 34348 22704 34400
rect 26148 34348 26200 34400
rect 27804 34552 27856 34604
rect 28356 34552 28408 34604
rect 28540 34552 28592 34604
rect 29092 34595 29144 34604
rect 29092 34561 29101 34595
rect 29101 34561 29135 34595
rect 29135 34561 29144 34595
rect 29092 34552 29144 34561
rect 29552 34595 29604 34604
rect 29552 34561 29561 34595
rect 29561 34561 29595 34595
rect 29595 34561 29604 34595
rect 29552 34552 29604 34561
rect 29736 34552 29788 34604
rect 27620 34416 27672 34468
rect 28724 34484 28776 34536
rect 29920 34595 29972 34604
rect 29920 34561 29929 34595
rect 29929 34561 29963 34595
rect 29963 34561 29972 34595
rect 29920 34552 29972 34561
rect 30840 34595 30892 34604
rect 30840 34561 30849 34595
rect 30849 34561 30883 34595
rect 30883 34561 30892 34595
rect 30840 34552 30892 34561
rect 30932 34595 30984 34604
rect 30932 34561 30966 34595
rect 30966 34561 30984 34595
rect 30932 34552 30984 34561
rect 33048 34552 33100 34604
rect 36084 34552 36136 34604
rect 37464 34552 37516 34604
rect 37832 34595 37884 34604
rect 37832 34561 37841 34595
rect 37841 34561 37875 34595
rect 37875 34561 37884 34595
rect 37832 34552 37884 34561
rect 37924 34552 37976 34604
rect 39764 34552 39816 34604
rect 39856 34595 39908 34604
rect 39856 34561 39865 34595
rect 39865 34561 39899 34595
rect 39899 34561 39908 34595
rect 39856 34552 39908 34561
rect 41236 34595 41288 34604
rect 41236 34561 41245 34595
rect 41245 34561 41279 34595
rect 41279 34561 41288 34595
rect 41788 34595 41840 34604
rect 41236 34552 41288 34561
rect 41788 34561 41797 34595
rect 41797 34561 41831 34595
rect 41831 34561 41840 34595
rect 41788 34552 41840 34561
rect 42156 34552 42208 34604
rect 30472 34484 30524 34536
rect 29184 34416 29236 34468
rect 33324 34484 33376 34536
rect 34244 34484 34296 34536
rect 35808 34527 35860 34536
rect 35808 34493 35817 34527
rect 35817 34493 35851 34527
rect 35851 34493 35860 34527
rect 35808 34484 35860 34493
rect 31760 34348 31812 34400
rect 31852 34348 31904 34400
rect 32312 34348 32364 34400
rect 42156 34459 42208 34468
rect 42156 34425 42165 34459
rect 42165 34425 42199 34459
rect 42199 34425 42208 34459
rect 42156 34416 42208 34425
rect 42708 34416 42760 34468
rect 38384 34348 38436 34400
rect 41696 34348 41748 34400
rect 41972 34348 42024 34400
rect 43812 34391 43864 34400
rect 43812 34357 43821 34391
rect 43821 34357 43855 34391
rect 43855 34357 43864 34391
rect 43812 34348 43864 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 9956 34144 10008 34196
rect 10324 34144 10376 34196
rect 10508 34144 10560 34196
rect 10876 34144 10928 34196
rect 13360 34187 13412 34196
rect 13360 34153 13369 34187
rect 13369 34153 13403 34187
rect 13403 34153 13412 34187
rect 13360 34144 13412 34153
rect 16304 34187 16356 34196
rect 16304 34153 16313 34187
rect 16313 34153 16347 34187
rect 16347 34153 16356 34187
rect 16304 34144 16356 34153
rect 18328 34187 18380 34196
rect 18328 34153 18337 34187
rect 18337 34153 18371 34187
rect 18371 34153 18380 34187
rect 18328 34144 18380 34153
rect 24124 34144 24176 34196
rect 34520 34144 34572 34196
rect 34612 34144 34664 34196
rect 11244 34076 11296 34128
rect 30932 34076 30984 34128
rect 5448 34008 5500 34060
rect 11428 34008 11480 34060
rect 15292 34008 15344 34060
rect 16764 34008 16816 34060
rect 19708 34008 19760 34060
rect 20076 34008 20128 34060
rect 21180 34008 21232 34060
rect 23572 34008 23624 34060
rect 30196 34008 30248 34060
rect 31024 34008 31076 34060
rect 3056 33940 3108 33992
rect 3608 33940 3660 33992
rect 14556 33940 14608 33992
rect 16672 33983 16724 33992
rect 16672 33949 16681 33983
rect 16681 33949 16715 33983
rect 16715 33949 16724 33983
rect 16672 33940 16724 33949
rect 18512 33983 18564 33992
rect 18512 33949 18521 33983
rect 18521 33949 18555 33983
rect 18555 33949 18564 33983
rect 18512 33940 18564 33949
rect 21272 33983 21324 33992
rect 21272 33949 21281 33983
rect 21281 33949 21315 33983
rect 21315 33949 21324 33983
rect 21272 33940 21324 33949
rect 21916 33983 21968 33992
rect 21916 33949 21925 33983
rect 21925 33949 21959 33983
rect 21959 33949 21968 33983
rect 21916 33940 21968 33949
rect 31668 33983 31720 33992
rect 31668 33949 31677 33983
rect 31677 33949 31711 33983
rect 31711 33949 31720 33983
rect 31668 33940 31720 33949
rect 31852 33940 31904 33992
rect 34612 34008 34664 34060
rect 36084 34187 36136 34196
rect 36084 34153 36093 34187
rect 36093 34153 36127 34187
rect 36127 34153 36136 34187
rect 36084 34144 36136 34153
rect 41788 34076 41840 34128
rect 42248 34119 42300 34128
rect 42248 34085 42257 34119
rect 42257 34085 42291 34119
rect 42291 34085 42300 34119
rect 42248 34076 42300 34085
rect 34520 33983 34572 33992
rect 34520 33949 34529 33983
rect 34529 33949 34563 33983
rect 34563 33949 34572 33983
rect 34520 33940 34572 33949
rect 35992 33940 36044 33992
rect 37464 33940 37516 33992
rect 42064 34008 42116 34060
rect 38660 33940 38712 33992
rect 4620 33872 4672 33924
rect 5356 33872 5408 33924
rect 15108 33872 15160 33924
rect 18328 33872 18380 33924
rect 20352 33872 20404 33924
rect 20996 33872 21048 33924
rect 21548 33915 21600 33924
rect 21548 33881 21557 33915
rect 21557 33881 21591 33915
rect 21591 33881 21600 33915
rect 21548 33872 21600 33881
rect 3884 33804 3936 33856
rect 15016 33804 15068 33856
rect 16948 33804 17000 33856
rect 22744 33804 22796 33856
rect 37740 33872 37792 33924
rect 41052 33983 41104 33992
rect 41052 33949 41061 33983
rect 41061 33949 41095 33983
rect 41095 33949 41104 33983
rect 41052 33940 41104 33949
rect 43812 34008 43864 34060
rect 44180 34008 44232 34060
rect 45192 34008 45244 34060
rect 45744 34008 45796 34060
rect 41144 33872 41196 33924
rect 41604 33872 41656 33924
rect 41972 33915 42024 33924
rect 41972 33881 41981 33915
rect 41981 33881 42015 33915
rect 42015 33881 42024 33915
rect 41972 33872 42024 33881
rect 44456 33940 44508 33992
rect 45376 33940 45428 33992
rect 32496 33804 32548 33856
rect 35808 33804 35860 33856
rect 37188 33847 37240 33856
rect 37188 33813 37197 33847
rect 37197 33813 37231 33847
rect 37231 33813 37240 33847
rect 37188 33804 37240 33813
rect 40316 33804 40368 33856
rect 41696 33804 41748 33856
rect 45008 33915 45060 33924
rect 45008 33881 45017 33915
rect 45017 33881 45051 33915
rect 45051 33881 45060 33915
rect 45008 33872 45060 33881
rect 46020 33872 46072 33924
rect 42432 33847 42484 33856
rect 42432 33813 42441 33847
rect 42441 33813 42475 33847
rect 42475 33813 42484 33847
rect 42432 33804 42484 33813
rect 42524 33804 42576 33856
rect 45376 33804 45428 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 3056 33643 3108 33652
rect 3056 33609 3065 33643
rect 3065 33609 3099 33643
rect 3099 33609 3108 33643
rect 3056 33600 3108 33609
rect 5356 33643 5408 33652
rect 5356 33609 5365 33643
rect 5365 33609 5399 33643
rect 5399 33609 5408 33643
rect 5356 33600 5408 33609
rect 13820 33600 13872 33652
rect 21916 33600 21968 33652
rect 23664 33600 23716 33652
rect 13176 33532 13228 33584
rect 15016 33532 15068 33584
rect 18604 33532 18656 33584
rect 20996 33532 21048 33584
rect 23480 33532 23532 33584
rect 2964 33507 3016 33516
rect 2964 33473 2973 33507
rect 2973 33473 3007 33507
rect 3007 33473 3016 33507
rect 2964 33464 3016 33473
rect 3884 33507 3936 33516
rect 3884 33473 3893 33507
rect 3893 33473 3927 33507
rect 3927 33473 3936 33507
rect 3884 33464 3936 33473
rect 3976 33507 4028 33516
rect 3976 33473 3985 33507
rect 3985 33473 4019 33507
rect 4019 33473 4028 33507
rect 3976 33464 4028 33473
rect 9404 33507 9456 33516
rect 9404 33473 9413 33507
rect 9413 33473 9447 33507
rect 9447 33473 9456 33507
rect 9404 33464 9456 33473
rect 3148 33439 3200 33448
rect 3148 33405 3157 33439
rect 3157 33405 3191 33439
rect 3191 33405 3200 33439
rect 3148 33396 3200 33405
rect 9680 33439 9732 33448
rect 9680 33405 9689 33439
rect 9689 33405 9723 33439
rect 9723 33405 9732 33439
rect 9680 33396 9732 33405
rect 10232 33328 10284 33380
rect 12992 33507 13044 33516
rect 12992 33473 13001 33507
rect 13001 33473 13035 33507
rect 13035 33473 13044 33507
rect 12992 33464 13044 33473
rect 13084 33396 13136 33448
rect 16580 33396 16632 33448
rect 22192 33464 22244 33516
rect 23112 33464 23164 33516
rect 27712 33600 27764 33652
rect 31668 33600 31720 33652
rect 32496 33643 32548 33652
rect 29276 33532 29328 33584
rect 30472 33532 30524 33584
rect 32496 33609 32505 33643
rect 32505 33609 32539 33643
rect 32539 33609 32548 33643
rect 32496 33600 32548 33609
rect 41052 33600 41104 33652
rect 41972 33600 42024 33652
rect 26056 33464 26108 33516
rect 27620 33464 27672 33516
rect 37188 33532 37240 33584
rect 35992 33464 36044 33516
rect 39304 33507 39356 33516
rect 39304 33473 39313 33507
rect 39313 33473 39347 33507
rect 39347 33473 39356 33507
rect 39304 33464 39356 33473
rect 2044 33260 2096 33312
rect 12164 33260 12216 33312
rect 24584 33396 24636 33448
rect 32036 33396 32088 33448
rect 31852 33328 31904 33380
rect 33508 33396 33560 33448
rect 34428 33439 34480 33448
rect 34428 33405 34437 33439
rect 34437 33405 34471 33439
rect 34471 33405 34480 33439
rect 34428 33396 34480 33405
rect 36176 33396 36228 33448
rect 37188 33396 37240 33448
rect 40316 33507 40368 33516
rect 40316 33473 40325 33507
rect 40325 33473 40359 33507
rect 40359 33473 40368 33507
rect 40316 33464 40368 33473
rect 42432 33532 42484 33584
rect 41328 33507 41380 33516
rect 41328 33473 41337 33507
rect 41337 33473 41371 33507
rect 41371 33473 41380 33507
rect 41328 33464 41380 33473
rect 41696 33507 41748 33516
rect 41696 33473 41705 33507
rect 41705 33473 41739 33507
rect 41739 33473 41748 33507
rect 41696 33464 41748 33473
rect 42064 33507 42116 33516
rect 42064 33473 42073 33507
rect 42073 33473 42107 33507
rect 42107 33473 42116 33507
rect 42064 33464 42116 33473
rect 42524 33464 42576 33516
rect 42708 33507 42760 33516
rect 42708 33473 42717 33507
rect 42717 33473 42751 33507
rect 42751 33473 42760 33507
rect 42708 33464 42760 33473
rect 43812 33532 43864 33584
rect 41880 33439 41932 33448
rect 41880 33405 41889 33439
rect 41889 33405 41923 33439
rect 41923 33405 41932 33439
rect 43904 33507 43956 33516
rect 43904 33473 43913 33507
rect 43913 33473 43947 33507
rect 43947 33473 43956 33507
rect 43904 33464 43956 33473
rect 44456 33507 44508 33516
rect 44456 33473 44465 33507
rect 44465 33473 44499 33507
rect 44499 33473 44508 33507
rect 44456 33464 44508 33473
rect 44548 33507 44600 33516
rect 44548 33473 44557 33507
rect 44557 33473 44591 33507
rect 44591 33473 44600 33507
rect 44548 33464 44600 33473
rect 44916 33507 44968 33516
rect 44916 33473 44925 33507
rect 44925 33473 44959 33507
rect 44959 33473 44968 33507
rect 44916 33464 44968 33473
rect 45008 33507 45060 33516
rect 45008 33473 45017 33507
rect 45017 33473 45051 33507
rect 45051 33473 45060 33507
rect 45008 33464 45060 33473
rect 45376 33575 45428 33584
rect 45376 33541 45385 33575
rect 45385 33541 45419 33575
rect 45419 33541 45428 33575
rect 45376 33532 45428 33541
rect 45468 33507 45520 33516
rect 45468 33473 45482 33507
rect 45482 33473 45516 33507
rect 45516 33473 45520 33507
rect 45468 33464 45520 33473
rect 45744 33507 45796 33516
rect 45744 33473 45753 33507
rect 45753 33473 45787 33507
rect 45787 33473 45796 33507
rect 45744 33464 45796 33473
rect 41880 33396 41932 33405
rect 14832 33260 14884 33312
rect 16304 33260 16356 33312
rect 18604 33303 18656 33312
rect 18604 33269 18613 33303
rect 18613 33269 18647 33303
rect 18647 33269 18656 33303
rect 18604 33260 18656 33269
rect 18972 33260 19024 33312
rect 24400 33260 24452 33312
rect 26516 33260 26568 33312
rect 37004 33260 37056 33312
rect 39212 33260 39264 33312
rect 40040 33303 40092 33312
rect 40040 33269 40049 33303
rect 40049 33269 40083 33303
rect 40083 33269 40092 33303
rect 40040 33260 40092 33269
rect 41144 33303 41196 33312
rect 41144 33269 41153 33303
rect 41153 33269 41187 33303
rect 41187 33269 41196 33303
rect 41144 33260 41196 33269
rect 41236 33303 41288 33312
rect 41236 33269 41245 33303
rect 41245 33269 41279 33303
rect 41279 33269 41288 33303
rect 41236 33260 41288 33269
rect 41696 33260 41748 33312
rect 42340 33260 42392 33312
rect 43444 33260 43496 33312
rect 44732 33260 44784 33312
rect 46112 33260 46164 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2964 33056 3016 33108
rect 4068 33056 4120 33108
rect 4712 33031 4764 33040
rect 4712 32997 4721 33031
rect 4721 32997 4755 33031
rect 4755 32997 4764 33031
rect 4712 32988 4764 32997
rect 4160 32920 4212 32972
rect 4620 32920 4672 32972
rect 6552 33056 6604 33108
rect 9312 33056 9364 33108
rect 9680 33056 9732 33108
rect 10416 33056 10468 33108
rect 5632 32920 5684 32972
rect 1676 32895 1728 32904
rect 1676 32861 1685 32895
rect 1685 32861 1719 32895
rect 1719 32861 1728 32895
rect 1676 32852 1728 32861
rect 1768 32895 1820 32904
rect 1768 32861 1777 32895
rect 1777 32861 1811 32895
rect 1811 32861 1820 32895
rect 1768 32852 1820 32861
rect 2044 32895 2096 32904
rect 2044 32861 2078 32895
rect 2078 32861 2096 32895
rect 2044 32852 2096 32861
rect 4252 32895 4304 32904
rect 4252 32861 4261 32895
rect 4261 32861 4295 32895
rect 4295 32861 4304 32895
rect 4252 32852 4304 32861
rect 4988 32895 5040 32904
rect 4988 32861 4997 32895
rect 4997 32861 5031 32895
rect 5031 32861 5040 32895
rect 4988 32852 5040 32861
rect 7104 32920 7156 32972
rect 7656 32963 7708 32972
rect 7656 32929 7665 32963
rect 7665 32929 7699 32963
rect 7699 32929 7708 32963
rect 7656 32920 7708 32929
rect 7564 32852 7616 32904
rect 8208 32920 8260 32972
rect 12992 33056 13044 33108
rect 14280 33056 14332 33108
rect 14648 32988 14700 33040
rect 9312 32895 9364 32904
rect 9312 32861 9321 32895
rect 9321 32861 9355 32895
rect 9355 32861 9364 32895
rect 9312 32852 9364 32861
rect 13912 32920 13964 32972
rect 14188 32963 14240 32972
rect 14188 32929 14197 32963
rect 14197 32929 14231 32963
rect 14231 32929 14240 32963
rect 14188 32920 14240 32929
rect 14832 32963 14884 32972
rect 14832 32929 14841 32963
rect 14841 32929 14875 32963
rect 14875 32929 14884 32963
rect 14832 32920 14884 32929
rect 16948 32963 17000 32972
rect 16948 32929 16957 32963
rect 16957 32929 16991 32963
rect 16991 32929 17000 32963
rect 16948 32920 17000 32929
rect 17040 32920 17092 32972
rect 17868 32920 17920 32972
rect 12164 32895 12216 32904
rect 12164 32861 12198 32895
rect 12198 32861 12216 32895
rect 1492 32759 1544 32768
rect 1492 32725 1501 32759
rect 1501 32725 1535 32759
rect 1535 32725 1544 32759
rect 1492 32716 1544 32725
rect 4528 32716 4580 32768
rect 5356 32716 5408 32768
rect 6736 32759 6788 32768
rect 6736 32725 6745 32759
rect 6745 32725 6779 32759
rect 6779 32725 6788 32759
rect 6736 32716 6788 32725
rect 6920 32716 6972 32768
rect 7748 32716 7800 32768
rect 7840 32759 7892 32768
rect 7840 32725 7849 32759
rect 7849 32725 7883 32759
rect 7883 32725 7892 32759
rect 7840 32716 7892 32725
rect 8208 32759 8260 32768
rect 8208 32725 8217 32759
rect 8217 32725 8251 32759
rect 8251 32725 8260 32759
rect 8208 32716 8260 32725
rect 8484 32716 8536 32768
rect 9680 32784 9732 32836
rect 9128 32716 9180 32768
rect 9864 32716 9916 32768
rect 11796 32784 11848 32836
rect 12164 32852 12216 32861
rect 14096 32852 14148 32904
rect 15200 32895 15252 32904
rect 15200 32861 15234 32895
rect 15234 32861 15252 32895
rect 15200 32852 15252 32861
rect 15384 32895 15436 32904
rect 15384 32861 15393 32895
rect 15393 32861 15427 32895
rect 15427 32861 15436 32895
rect 15384 32852 15436 32861
rect 12624 32784 12676 32836
rect 14280 32784 14332 32836
rect 15936 32784 15988 32836
rect 13912 32716 13964 32768
rect 15108 32716 15160 32768
rect 17224 32759 17276 32768
rect 17224 32725 17233 32759
rect 17233 32725 17267 32759
rect 17267 32725 17276 32759
rect 17224 32716 17276 32725
rect 18052 32784 18104 32836
rect 17960 32716 18012 32768
rect 18880 32963 18932 32972
rect 18880 32929 18889 32963
rect 18889 32929 18923 32963
rect 18923 32929 18932 32963
rect 18880 32920 18932 32929
rect 18604 32852 18656 32904
rect 20260 32920 20312 32972
rect 20996 32920 21048 32972
rect 23112 33056 23164 33108
rect 25780 33056 25832 33108
rect 26056 33099 26108 33108
rect 26056 33065 26065 33099
rect 26065 33065 26099 33099
rect 26099 33065 26108 33099
rect 26056 33056 26108 33065
rect 19800 32852 19852 32904
rect 22376 32920 22428 32972
rect 22560 32920 22612 32972
rect 23112 32920 23164 32972
rect 21640 32784 21692 32836
rect 18512 32716 18564 32768
rect 19156 32716 19208 32768
rect 20720 32759 20772 32768
rect 20720 32725 20729 32759
rect 20729 32725 20763 32759
rect 20763 32725 20772 32759
rect 20720 32716 20772 32725
rect 20812 32716 20864 32768
rect 22468 32784 22520 32836
rect 22928 32784 22980 32836
rect 24584 32852 24636 32904
rect 30012 33056 30064 33108
rect 29000 32988 29052 33040
rect 26792 32963 26844 32972
rect 26792 32929 26801 32963
rect 26801 32929 26835 32963
rect 26835 32929 26844 32963
rect 26792 32920 26844 32929
rect 26884 32920 26936 32972
rect 27160 32920 27212 32972
rect 29644 32920 29696 32972
rect 32404 33056 32456 33108
rect 33508 33056 33560 33108
rect 38660 33099 38712 33108
rect 38660 33065 38669 33099
rect 38669 33065 38703 33099
rect 38703 33065 38712 33099
rect 38660 33056 38712 33065
rect 39304 33056 39356 33108
rect 41880 33056 41932 33108
rect 42340 33056 42392 33108
rect 37372 32988 37424 33040
rect 41604 33031 41656 33040
rect 41604 32997 41613 33031
rect 41613 32997 41647 33031
rect 41647 32997 41656 33031
rect 41604 32988 41656 32997
rect 36820 32963 36872 32972
rect 36820 32929 36829 32963
rect 36829 32929 36863 32963
rect 36863 32929 36872 32963
rect 36820 32920 36872 32929
rect 41972 32963 42024 32972
rect 41972 32929 41981 32963
rect 41981 32929 42015 32963
rect 42015 32929 42024 32963
rect 41972 32920 42024 32929
rect 26516 32852 26568 32904
rect 27528 32852 27580 32904
rect 30380 32852 30432 32904
rect 32128 32895 32180 32904
rect 32128 32861 32137 32895
rect 32137 32861 32171 32895
rect 32171 32861 32180 32895
rect 32128 32852 32180 32861
rect 32312 32852 32364 32904
rect 33416 32852 33468 32904
rect 34428 32852 34480 32904
rect 24768 32827 24820 32836
rect 24768 32793 24802 32827
rect 24802 32793 24820 32827
rect 24768 32784 24820 32793
rect 24400 32716 24452 32768
rect 24584 32716 24636 32768
rect 24676 32716 24728 32768
rect 25412 32716 25464 32768
rect 26608 32784 26660 32836
rect 30748 32784 30800 32836
rect 28356 32716 28408 32768
rect 29276 32716 29328 32768
rect 29368 32716 29420 32768
rect 30656 32716 30708 32768
rect 35992 32895 36044 32904
rect 35992 32861 36001 32895
rect 36001 32861 36035 32895
rect 36035 32861 36044 32895
rect 35992 32852 36044 32861
rect 37096 32852 37148 32904
rect 36084 32784 36136 32836
rect 37832 32852 37884 32904
rect 38200 32852 38252 32904
rect 32680 32716 32732 32768
rect 39028 32784 39080 32836
rect 40500 32827 40552 32836
rect 40500 32793 40509 32827
rect 40509 32793 40543 32827
rect 40543 32793 40552 32827
rect 40500 32784 40552 32793
rect 40776 32784 40828 32836
rect 41788 32895 41840 32904
rect 41788 32861 41797 32895
rect 41797 32861 41831 32895
rect 41831 32861 41840 32895
rect 41788 32852 41840 32861
rect 42064 32895 42116 32904
rect 42064 32861 42073 32895
rect 42073 32861 42107 32895
rect 42107 32861 42116 32895
rect 42064 32852 42116 32861
rect 42248 32895 42300 32904
rect 42248 32861 42257 32895
rect 42257 32861 42291 32895
rect 42291 32861 42300 32895
rect 42248 32852 42300 32861
rect 43812 33056 43864 33108
rect 42524 33031 42576 33040
rect 42524 32997 42533 33031
rect 42533 32997 42567 33031
rect 42567 32997 42576 33031
rect 42524 32988 42576 32997
rect 44364 33099 44416 33108
rect 44364 33065 44373 33099
rect 44373 33065 44407 33099
rect 44407 33065 44416 33099
rect 44364 33056 44416 33065
rect 44548 33056 44600 33108
rect 44640 33056 44692 33108
rect 45468 33099 45520 33108
rect 45468 33065 45477 33099
rect 45477 33065 45511 33099
rect 45511 33065 45520 33099
rect 45468 33056 45520 33065
rect 46020 33099 46072 33108
rect 46020 33065 46029 33099
rect 46029 33065 46063 33099
rect 46063 33065 46072 33099
rect 46020 33056 46072 33065
rect 45836 33031 45888 33040
rect 45836 32997 45845 33031
rect 45845 32997 45879 33031
rect 45879 32997 45888 33031
rect 45836 32988 45888 32997
rect 42616 32852 42668 32904
rect 42892 32852 42944 32904
rect 42524 32827 42576 32836
rect 42524 32793 42533 32827
rect 42533 32793 42567 32827
rect 42567 32793 42576 32827
rect 42524 32784 42576 32793
rect 44640 32827 44692 32836
rect 44640 32793 44649 32827
rect 44649 32793 44683 32827
rect 44683 32793 44692 32827
rect 44640 32784 44692 32793
rect 45008 32895 45060 32904
rect 45008 32861 45017 32895
rect 45017 32861 45051 32895
rect 45051 32861 45060 32895
rect 45008 32852 45060 32861
rect 45100 32784 45152 32836
rect 37280 32759 37332 32768
rect 37280 32725 37289 32759
rect 37289 32725 37323 32759
rect 37323 32725 37332 32759
rect 37280 32716 37332 32725
rect 37648 32716 37700 32768
rect 41696 32716 41748 32768
rect 42432 32759 42484 32768
rect 42432 32725 42441 32759
rect 42441 32725 42475 32759
rect 42475 32725 42484 32759
rect 42432 32716 42484 32725
rect 42800 32716 42852 32768
rect 44916 32716 44968 32768
rect 46664 32759 46716 32768
rect 46664 32725 46673 32759
rect 46673 32725 46707 32759
rect 46707 32725 46716 32759
rect 46664 32716 46716 32725
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 1676 32512 1728 32564
rect 1492 32444 1544 32496
rect 1768 32376 1820 32428
rect 4988 32512 5040 32564
rect 3608 32487 3660 32496
rect 3608 32453 3617 32487
rect 3617 32453 3651 32487
rect 3651 32453 3660 32487
rect 3608 32444 3660 32453
rect 3976 32444 4028 32496
rect 6736 32444 6788 32496
rect 7748 32555 7800 32564
rect 7748 32521 7757 32555
rect 7757 32521 7791 32555
rect 7791 32521 7800 32555
rect 7748 32512 7800 32521
rect 10508 32512 10560 32564
rect 12072 32512 12124 32564
rect 12624 32512 12676 32564
rect 13360 32512 13412 32564
rect 14924 32512 14976 32564
rect 15200 32512 15252 32564
rect 17960 32512 18012 32564
rect 18052 32555 18104 32564
rect 18052 32521 18061 32555
rect 18061 32521 18095 32555
rect 18095 32521 18104 32555
rect 18052 32512 18104 32521
rect 18144 32512 18196 32564
rect 18788 32512 18840 32564
rect 9128 32444 9180 32496
rect 14004 32444 14056 32496
rect 4160 32376 4212 32428
rect 4988 32419 5040 32428
rect 4988 32385 4997 32419
rect 4997 32385 5031 32419
rect 5031 32385 5040 32419
rect 4988 32376 5040 32385
rect 7840 32376 7892 32428
rect 8944 32376 8996 32428
rect 9864 32376 9916 32428
rect 10508 32419 10560 32428
rect 10508 32385 10542 32419
rect 10542 32385 10560 32419
rect 10508 32376 10560 32385
rect 10692 32419 10744 32428
rect 10692 32385 10701 32419
rect 10701 32385 10735 32419
rect 10735 32385 10744 32419
rect 10692 32376 10744 32385
rect 11612 32376 11664 32428
rect 12072 32419 12124 32428
rect 12072 32385 12106 32419
rect 12106 32385 12124 32419
rect 12072 32376 12124 32385
rect 13820 32419 13872 32428
rect 13820 32385 13829 32419
rect 13829 32385 13863 32419
rect 13863 32385 13872 32419
rect 13820 32376 13872 32385
rect 3700 32351 3752 32360
rect 3700 32317 3709 32351
rect 3709 32317 3743 32351
rect 3743 32317 3752 32351
rect 3700 32308 3752 32317
rect 4252 32351 4304 32360
rect 4252 32317 4261 32351
rect 4261 32317 4295 32351
rect 4295 32317 4304 32351
rect 4252 32308 4304 32317
rect 4620 32308 4672 32360
rect 4528 32240 4580 32292
rect 4068 32172 4120 32224
rect 5448 32308 5500 32360
rect 6368 32351 6420 32360
rect 6368 32317 6377 32351
rect 6377 32317 6411 32351
rect 6411 32317 6420 32351
rect 6368 32308 6420 32317
rect 5724 32240 5776 32292
rect 6644 32172 6696 32224
rect 6736 32172 6788 32224
rect 9220 32240 9272 32292
rect 14924 32419 14976 32428
rect 14924 32385 14958 32419
rect 14958 32385 14976 32419
rect 14924 32376 14976 32385
rect 15108 32419 15160 32428
rect 15108 32385 15117 32419
rect 15117 32385 15151 32419
rect 15151 32385 15160 32419
rect 15108 32376 15160 32385
rect 10140 32283 10192 32292
rect 10140 32249 10149 32283
rect 10149 32249 10183 32283
rect 10183 32249 10192 32283
rect 10140 32240 10192 32249
rect 8208 32172 8260 32224
rect 9956 32172 10008 32224
rect 11152 32172 11204 32224
rect 11336 32215 11388 32224
rect 11336 32181 11345 32215
rect 11345 32181 11379 32215
rect 11379 32181 11388 32215
rect 11336 32172 11388 32181
rect 11796 32351 11848 32360
rect 11796 32317 11805 32351
rect 11805 32317 11839 32351
rect 11839 32317 11848 32351
rect 11796 32308 11848 32317
rect 14096 32351 14148 32360
rect 14096 32317 14105 32351
rect 14105 32317 14139 32351
rect 14139 32317 14148 32351
rect 14096 32308 14148 32317
rect 14188 32308 14240 32360
rect 14648 32308 14700 32360
rect 11796 32172 11848 32224
rect 12532 32172 12584 32224
rect 16396 32376 16448 32428
rect 17224 32376 17276 32428
rect 18512 32419 18564 32428
rect 18512 32385 18521 32419
rect 18521 32385 18555 32419
rect 18555 32385 18564 32419
rect 18512 32376 18564 32385
rect 14280 32172 14332 32224
rect 16028 32215 16080 32224
rect 16028 32181 16037 32215
rect 16037 32181 16071 32215
rect 16071 32181 16080 32215
rect 16028 32172 16080 32181
rect 16396 32172 16448 32224
rect 20812 32555 20864 32564
rect 20812 32521 20821 32555
rect 20821 32521 20855 32555
rect 20855 32521 20864 32555
rect 20812 32512 20864 32521
rect 21456 32512 21508 32564
rect 21548 32512 21600 32564
rect 24584 32512 24636 32564
rect 24768 32555 24820 32564
rect 24768 32521 24777 32555
rect 24777 32521 24811 32555
rect 24811 32521 24820 32555
rect 24768 32512 24820 32521
rect 25412 32555 25464 32564
rect 25412 32521 25421 32555
rect 25421 32521 25455 32555
rect 25455 32521 25464 32555
rect 25412 32512 25464 32521
rect 27988 32512 28040 32564
rect 29184 32512 29236 32564
rect 30380 32555 30432 32564
rect 30380 32521 30389 32555
rect 30389 32521 30423 32555
rect 30423 32521 30432 32555
rect 30380 32512 30432 32521
rect 30748 32555 30800 32564
rect 30748 32521 30757 32555
rect 30757 32521 30791 32555
rect 30791 32521 30800 32555
rect 30748 32512 30800 32521
rect 32128 32555 32180 32564
rect 32128 32521 32137 32555
rect 32137 32521 32171 32555
rect 32171 32521 32180 32555
rect 32128 32512 32180 32521
rect 32496 32555 32548 32564
rect 32496 32521 32505 32555
rect 32505 32521 32539 32555
rect 32539 32521 32548 32555
rect 32496 32512 32548 32521
rect 32680 32512 32732 32564
rect 32956 32512 33008 32564
rect 34244 32512 34296 32564
rect 19064 32376 19116 32428
rect 19156 32419 19208 32428
rect 19156 32385 19165 32419
rect 19165 32385 19199 32419
rect 19199 32385 19208 32419
rect 19156 32376 19208 32385
rect 20904 32419 20956 32428
rect 20904 32385 20913 32419
rect 20913 32385 20947 32419
rect 20947 32385 20956 32419
rect 20904 32376 20956 32385
rect 22744 32444 22796 32496
rect 19892 32351 19944 32360
rect 19892 32317 19901 32351
rect 19901 32317 19935 32351
rect 19935 32317 19944 32351
rect 19892 32308 19944 32317
rect 19984 32351 20036 32360
rect 19984 32317 20018 32351
rect 20018 32317 20036 32351
rect 19984 32308 20036 32317
rect 20168 32351 20220 32360
rect 20168 32317 20177 32351
rect 20177 32317 20211 32351
rect 20211 32317 20220 32351
rect 20168 32308 20220 32317
rect 20720 32308 20772 32360
rect 19708 32240 19760 32292
rect 20812 32240 20864 32292
rect 22192 32419 22244 32428
rect 22192 32385 22201 32419
rect 22201 32385 22235 32419
rect 22235 32385 22244 32419
rect 22192 32376 22244 32385
rect 26792 32444 26844 32496
rect 24676 32308 24728 32360
rect 21456 32240 21508 32292
rect 26332 32376 26384 32428
rect 26700 32376 26752 32428
rect 27988 32419 28040 32428
rect 29552 32444 29604 32496
rect 37372 32512 37424 32564
rect 27988 32385 28022 32419
rect 28022 32385 28040 32419
rect 27988 32376 28040 32385
rect 29184 32419 29236 32428
rect 29184 32385 29218 32419
rect 29218 32385 29236 32419
rect 29184 32376 29236 32385
rect 18144 32215 18196 32224
rect 18144 32181 18153 32215
rect 18153 32181 18187 32215
rect 18187 32181 18196 32215
rect 18144 32172 18196 32181
rect 18880 32172 18932 32224
rect 19248 32172 19300 32224
rect 20352 32172 20404 32224
rect 20904 32172 20956 32224
rect 21364 32215 21416 32224
rect 21364 32181 21373 32215
rect 21373 32181 21407 32215
rect 21407 32181 21416 32215
rect 21364 32172 21416 32181
rect 22100 32172 22152 32224
rect 22468 32172 22520 32224
rect 26608 32308 26660 32360
rect 27160 32351 27212 32360
rect 27160 32317 27169 32351
rect 27169 32317 27203 32351
rect 27203 32317 27212 32351
rect 27160 32308 27212 32317
rect 27528 32308 27580 32360
rect 28172 32351 28224 32360
rect 28172 32317 28181 32351
rect 28181 32317 28215 32351
rect 28215 32317 28224 32351
rect 28172 32308 28224 32317
rect 30656 32308 30708 32360
rect 38016 32444 38068 32496
rect 31024 32351 31076 32360
rect 31024 32317 31033 32351
rect 31033 32317 31067 32351
rect 31067 32317 31076 32351
rect 31024 32308 31076 32317
rect 32680 32351 32732 32360
rect 32680 32317 32689 32351
rect 32689 32317 32723 32351
rect 32723 32317 32732 32351
rect 32680 32308 32732 32317
rect 35348 32308 35400 32360
rect 27620 32283 27672 32292
rect 27620 32249 27629 32283
rect 27629 32249 27663 32283
rect 27663 32249 27672 32283
rect 27620 32240 27672 32249
rect 27160 32172 27212 32224
rect 28632 32172 28684 32224
rect 30196 32240 30248 32292
rect 36820 32240 36872 32292
rect 37096 32308 37148 32360
rect 40500 32376 40552 32428
rect 37556 32351 37608 32360
rect 37556 32317 37565 32351
rect 37565 32317 37599 32351
rect 37599 32317 37608 32351
rect 37556 32308 37608 32317
rect 40224 32351 40276 32360
rect 40224 32317 40233 32351
rect 40233 32317 40267 32351
rect 40267 32317 40276 32351
rect 40224 32308 40276 32317
rect 40776 32308 40828 32360
rect 41236 32419 41288 32428
rect 41236 32385 41245 32419
rect 41245 32385 41279 32419
rect 41279 32385 41288 32419
rect 41236 32376 41288 32385
rect 42064 32512 42116 32564
rect 42432 32555 42484 32564
rect 42432 32521 42441 32555
rect 42441 32521 42475 32555
rect 42475 32521 42484 32555
rect 42432 32512 42484 32521
rect 43904 32512 43956 32564
rect 45468 32512 45520 32564
rect 42708 32444 42760 32496
rect 43168 32487 43220 32496
rect 43168 32453 43177 32487
rect 43177 32453 43211 32487
rect 43211 32453 43220 32487
rect 43168 32444 43220 32453
rect 44180 32444 44232 32496
rect 44916 32444 44968 32496
rect 38568 32240 38620 32292
rect 41328 32240 41380 32292
rect 42156 32419 42208 32428
rect 42156 32385 42165 32419
rect 42165 32385 42199 32419
rect 42199 32385 42208 32419
rect 42156 32376 42208 32385
rect 42616 32376 42668 32428
rect 42340 32308 42392 32360
rect 42892 32351 42944 32360
rect 42892 32317 42901 32351
rect 42901 32317 42935 32351
rect 42935 32317 42944 32351
rect 43444 32419 43496 32428
rect 43444 32385 43453 32419
rect 43453 32385 43487 32419
rect 43487 32385 43496 32419
rect 43444 32376 43496 32385
rect 44364 32376 44416 32428
rect 42892 32308 42944 32317
rect 44640 32351 44692 32360
rect 44640 32317 44649 32351
rect 44649 32317 44683 32351
rect 44683 32317 44692 32351
rect 44640 32308 44692 32317
rect 44824 32351 44876 32360
rect 44824 32317 44833 32351
rect 44833 32317 44867 32351
rect 44867 32317 44876 32351
rect 44824 32308 44876 32317
rect 45008 32419 45060 32428
rect 45008 32385 45017 32419
rect 45017 32385 45051 32419
rect 45051 32385 45060 32419
rect 45008 32376 45060 32385
rect 29644 32172 29696 32224
rect 36544 32172 36596 32224
rect 37648 32215 37700 32224
rect 37648 32181 37657 32215
rect 37657 32181 37691 32215
rect 37691 32181 37700 32215
rect 37648 32172 37700 32181
rect 38476 32172 38528 32224
rect 41512 32172 41564 32224
rect 41604 32172 41656 32224
rect 42524 32172 42576 32224
rect 45376 32240 45428 32292
rect 43076 32215 43128 32224
rect 43076 32181 43085 32215
rect 43085 32181 43119 32215
rect 43119 32181 43128 32215
rect 43076 32172 43128 32181
rect 45100 32215 45152 32224
rect 45100 32181 45109 32215
rect 45109 32181 45143 32215
rect 45143 32181 45152 32215
rect 45100 32172 45152 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 3700 31968 3752 32020
rect 6276 31968 6328 32020
rect 7564 31968 7616 32020
rect 8208 31968 8260 32020
rect 8944 32011 8996 32020
rect 8944 31977 8953 32011
rect 8953 31977 8987 32011
rect 8987 31977 8996 32011
rect 8944 31968 8996 31977
rect 4712 31900 4764 31952
rect 5264 31900 5316 31952
rect 940 31832 992 31884
rect 1676 31875 1728 31884
rect 1676 31841 1685 31875
rect 1685 31841 1719 31875
rect 1719 31841 1728 31875
rect 1676 31832 1728 31841
rect 6368 31875 6420 31884
rect 6368 31841 6377 31875
rect 6377 31841 6411 31875
rect 6411 31841 6420 31875
rect 6368 31832 6420 31841
rect 4712 31764 4764 31816
rect 5356 31764 5408 31816
rect 6644 31807 6696 31816
rect 6644 31773 6678 31807
rect 6678 31773 6696 31807
rect 6644 31764 6696 31773
rect 9588 31900 9640 31952
rect 12532 31968 12584 32020
rect 12808 31968 12860 32020
rect 13636 31968 13688 32020
rect 13912 31968 13964 32020
rect 14004 31900 14056 31952
rect 14188 31968 14240 32020
rect 18512 31968 18564 32020
rect 19984 31968 20036 32020
rect 20260 31968 20312 32020
rect 20352 31968 20404 32020
rect 21364 31968 21416 32020
rect 21732 31968 21784 32020
rect 8668 31875 8720 31884
rect 8668 31841 8677 31875
rect 8677 31841 8711 31875
rect 8711 31841 8720 31875
rect 8668 31832 8720 31841
rect 9220 31875 9272 31884
rect 9220 31841 9229 31875
rect 9229 31841 9263 31875
rect 9263 31841 9272 31875
rect 9220 31832 9272 31841
rect 9772 31832 9824 31884
rect 9956 31832 10008 31884
rect 10600 31832 10652 31884
rect 11336 31832 11388 31884
rect 10416 31807 10468 31816
rect 10416 31773 10425 31807
rect 10425 31773 10459 31807
rect 10459 31773 10468 31807
rect 10416 31764 10468 31773
rect 12532 31875 12584 31884
rect 12532 31841 12541 31875
rect 12541 31841 12575 31875
rect 12575 31841 12584 31875
rect 12532 31832 12584 31841
rect 13176 31832 13228 31884
rect 13268 31875 13320 31884
rect 13268 31841 13277 31875
rect 13277 31841 13311 31875
rect 13311 31841 13320 31875
rect 13268 31832 13320 31841
rect 15292 31900 15344 31952
rect 19156 31900 19208 31952
rect 16396 31875 16448 31884
rect 16396 31841 16405 31875
rect 16405 31841 16439 31875
rect 16439 31841 16448 31875
rect 16396 31832 16448 31841
rect 19064 31832 19116 31884
rect 21088 31900 21140 31952
rect 21456 31900 21508 31952
rect 19524 31832 19576 31884
rect 20168 31875 20220 31884
rect 20168 31841 20177 31875
rect 20177 31841 20211 31875
rect 20211 31841 20220 31875
rect 20168 31832 20220 31841
rect 20260 31875 20312 31884
rect 20260 31841 20294 31875
rect 20294 31841 20312 31875
rect 20260 31832 20312 31841
rect 12808 31764 12860 31816
rect 13360 31764 13412 31816
rect 14280 31764 14332 31816
rect 15936 31807 15988 31816
rect 15936 31773 15945 31807
rect 15945 31773 15979 31807
rect 15979 31773 15988 31807
rect 15936 31764 15988 31773
rect 16028 31764 16080 31816
rect 20444 31807 20496 31816
rect 20444 31773 20453 31807
rect 20453 31773 20487 31807
rect 20487 31773 20496 31807
rect 20444 31764 20496 31773
rect 11520 31696 11572 31748
rect 15752 31696 15804 31748
rect 21180 31764 21232 31816
rect 8484 31671 8536 31680
rect 8484 31637 8493 31671
rect 8493 31637 8527 31671
rect 8527 31637 8536 31671
rect 8484 31628 8536 31637
rect 10140 31628 10192 31680
rect 11612 31628 11664 31680
rect 16028 31671 16080 31680
rect 16028 31637 16037 31671
rect 16037 31637 16071 31671
rect 16071 31637 16080 31671
rect 16028 31628 16080 31637
rect 20996 31628 21048 31680
rect 21180 31671 21232 31680
rect 21180 31637 21189 31671
rect 21189 31637 21223 31671
rect 21223 31637 21232 31671
rect 21180 31628 21232 31637
rect 22008 31968 22060 32020
rect 23204 31968 23256 32020
rect 28172 31968 28224 32020
rect 29184 32011 29236 32020
rect 29184 31977 29193 32011
rect 29193 31977 29227 32011
rect 29227 31977 29236 32011
rect 29184 31968 29236 31977
rect 22836 31900 22888 31952
rect 27344 31900 27396 31952
rect 28908 31900 28960 31952
rect 30656 31968 30708 32020
rect 30748 31968 30800 32020
rect 31024 31968 31076 32020
rect 31300 31900 31352 31952
rect 32036 31900 32088 31952
rect 37556 31968 37608 32020
rect 26608 31875 26660 31884
rect 26608 31841 26617 31875
rect 26617 31841 26651 31875
rect 26651 31841 26660 31875
rect 26608 31832 26660 31841
rect 27160 31832 27212 31884
rect 27528 31875 27580 31884
rect 27528 31841 27537 31875
rect 27537 31841 27571 31875
rect 27571 31841 27580 31875
rect 27528 31832 27580 31841
rect 27988 31832 28040 31884
rect 28356 31832 28408 31884
rect 29276 31832 29328 31884
rect 21548 31807 21600 31816
rect 21548 31773 21557 31807
rect 21557 31773 21591 31807
rect 21591 31773 21600 31807
rect 21548 31764 21600 31773
rect 21640 31807 21692 31816
rect 21640 31773 21649 31807
rect 21649 31773 21683 31807
rect 21683 31773 21692 31807
rect 21640 31764 21692 31773
rect 21732 31764 21784 31816
rect 22100 31807 22152 31816
rect 22100 31773 22134 31807
rect 22134 31773 22152 31807
rect 22100 31764 22152 31773
rect 22376 31764 22428 31816
rect 26700 31764 26752 31816
rect 27804 31807 27856 31816
rect 27804 31773 27813 31807
rect 27813 31773 27847 31807
rect 27847 31773 27856 31807
rect 27804 31764 27856 31773
rect 29368 31807 29420 31816
rect 29368 31773 29377 31807
rect 29377 31773 29411 31807
rect 29411 31773 29420 31807
rect 29368 31764 29420 31773
rect 29552 31807 29604 31816
rect 29552 31773 29561 31807
rect 29561 31773 29595 31807
rect 29595 31773 29604 31807
rect 29552 31764 29604 31773
rect 30840 31832 30892 31884
rect 30380 31764 30432 31816
rect 31484 31764 31536 31816
rect 31852 31764 31904 31816
rect 34612 31764 34664 31816
rect 34888 31807 34940 31816
rect 34888 31773 34895 31807
rect 34895 31773 34940 31807
rect 34888 31764 34940 31773
rect 21824 31628 21876 31680
rect 22376 31628 22428 31680
rect 24584 31628 24636 31680
rect 34520 31696 34572 31748
rect 35256 31764 35308 31816
rect 35348 31764 35400 31816
rect 35992 31764 36044 31816
rect 36084 31807 36136 31816
rect 36084 31773 36093 31807
rect 36093 31773 36127 31807
rect 36127 31773 36136 31807
rect 36084 31764 36136 31773
rect 37464 31764 37516 31816
rect 37648 31875 37700 31884
rect 37648 31841 37657 31875
rect 37657 31841 37691 31875
rect 37691 31841 37700 31875
rect 37648 31832 37700 31841
rect 41972 31968 42024 32020
rect 42340 31968 42392 32020
rect 44640 31968 44692 32020
rect 45008 31900 45060 31952
rect 41512 31832 41564 31884
rect 40224 31764 40276 31816
rect 40592 31764 40644 31816
rect 42248 31764 42300 31816
rect 42708 31764 42760 31816
rect 43720 31764 43772 31816
rect 44916 31764 44968 31816
rect 29000 31671 29052 31680
rect 29000 31637 29009 31671
rect 29009 31637 29043 31671
rect 29043 31637 29052 31671
rect 29000 31628 29052 31637
rect 33968 31671 34020 31680
rect 33968 31637 33977 31671
rect 33977 31637 34011 31671
rect 34011 31637 34020 31671
rect 33968 31628 34020 31637
rect 35164 31628 35216 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 9680 31467 9732 31476
rect 9680 31433 9689 31467
rect 9689 31433 9723 31467
rect 9723 31433 9732 31467
rect 9680 31424 9732 31433
rect 9864 31424 9916 31476
rect 11520 31424 11572 31476
rect 13820 31424 13872 31476
rect 15292 31467 15344 31476
rect 15292 31433 15301 31467
rect 15301 31433 15335 31467
rect 15335 31433 15344 31467
rect 15292 31424 15344 31433
rect 15936 31424 15988 31476
rect 17960 31424 18012 31476
rect 21548 31424 21600 31476
rect 22284 31424 22336 31476
rect 22376 31467 22428 31476
rect 22376 31433 22385 31467
rect 22385 31433 22419 31467
rect 22419 31433 22428 31467
rect 22376 31424 22428 31433
rect 22468 31467 22520 31476
rect 22468 31433 22477 31467
rect 22477 31433 22511 31467
rect 22511 31433 22520 31467
rect 22468 31424 22520 31433
rect 20444 31399 20496 31408
rect 20444 31365 20453 31399
rect 20453 31365 20487 31399
rect 20487 31365 20496 31399
rect 20444 31356 20496 31365
rect 30840 31424 30892 31476
rect 31300 31424 31352 31476
rect 34612 31424 34664 31476
rect 35440 31424 35492 31476
rect 41512 31467 41564 31476
rect 41512 31433 41521 31467
rect 41521 31433 41555 31467
rect 41555 31433 41564 31467
rect 41512 31424 41564 31433
rect 44824 31424 44876 31476
rect 45468 31424 45520 31476
rect 2228 31331 2280 31340
rect 2228 31297 2237 31331
rect 2237 31297 2271 31331
rect 2271 31297 2280 31331
rect 2228 31288 2280 31297
rect 6920 31288 6972 31340
rect 20168 31288 20220 31340
rect 20720 31331 20772 31340
rect 20720 31297 20729 31331
rect 20729 31297 20763 31331
rect 20763 31297 20772 31331
rect 20720 31288 20772 31297
rect 4988 31220 5040 31272
rect 5448 31220 5500 31272
rect 10140 31263 10192 31272
rect 10140 31229 10149 31263
rect 10149 31229 10183 31263
rect 10183 31229 10192 31263
rect 10140 31220 10192 31229
rect 9772 31152 9824 31204
rect 10876 31220 10928 31272
rect 12164 31152 12216 31204
rect 15476 31220 15528 31272
rect 21640 31288 21692 31340
rect 21732 31220 21784 31272
rect 22376 31220 22428 31272
rect 23572 31263 23624 31272
rect 23572 31229 23581 31263
rect 23581 31229 23615 31263
rect 23615 31229 23624 31263
rect 23572 31220 23624 31229
rect 23756 31263 23808 31272
rect 23756 31229 23765 31263
rect 23765 31229 23799 31263
rect 23799 31229 23808 31263
rect 23756 31220 23808 31229
rect 24216 31263 24268 31272
rect 24216 31229 24225 31263
rect 24225 31229 24259 31263
rect 24259 31229 24268 31263
rect 24216 31220 24268 31229
rect 24492 31263 24544 31272
rect 24492 31229 24501 31263
rect 24501 31229 24535 31263
rect 24535 31229 24544 31263
rect 24492 31220 24544 31229
rect 24584 31263 24636 31272
rect 24584 31229 24618 31263
rect 24618 31229 24636 31263
rect 24584 31220 24636 31229
rect 25596 31220 25648 31272
rect 25780 31220 25832 31272
rect 33784 31356 33836 31408
rect 33968 31399 34020 31408
rect 33968 31365 34002 31399
rect 34002 31365 34020 31399
rect 33968 31356 34020 31365
rect 2044 31127 2096 31136
rect 2044 31093 2053 31127
rect 2053 31093 2087 31127
rect 2087 31093 2096 31127
rect 2044 31084 2096 31093
rect 7656 31084 7708 31136
rect 20812 31084 20864 31136
rect 21088 31084 21140 31136
rect 21272 31152 21324 31204
rect 22192 31152 22244 31204
rect 23664 31152 23716 31204
rect 28264 31288 28316 31340
rect 28448 31288 28500 31340
rect 29092 31288 29144 31340
rect 29000 31152 29052 31204
rect 31944 31288 31996 31340
rect 33048 31288 33100 31340
rect 36084 31356 36136 31408
rect 31392 31220 31444 31272
rect 32036 31220 32088 31272
rect 32588 31220 32640 31272
rect 31208 31152 31260 31204
rect 33416 31220 33468 31272
rect 22928 31084 22980 31136
rect 23848 31084 23900 31136
rect 24768 31084 24820 31136
rect 27528 31127 27580 31136
rect 27528 31093 27537 31127
rect 27537 31093 27571 31127
rect 27571 31093 27580 31127
rect 27528 31084 27580 31093
rect 27988 31127 28040 31136
rect 27988 31093 27997 31127
rect 27997 31093 28031 31127
rect 28031 31093 28040 31127
rect 27988 31084 28040 31093
rect 30840 31127 30892 31136
rect 30840 31093 30849 31127
rect 30849 31093 30883 31127
rect 30883 31093 30892 31127
rect 30840 31084 30892 31093
rect 31852 31084 31904 31136
rect 36360 31288 36412 31340
rect 36544 31288 36596 31340
rect 37280 31288 37332 31340
rect 37556 31331 37608 31340
rect 37556 31297 37565 31331
rect 37565 31297 37599 31331
rect 37599 31297 37608 31331
rect 37556 31288 37608 31297
rect 35716 31263 35768 31272
rect 35716 31229 35725 31263
rect 35725 31229 35759 31263
rect 35759 31229 35768 31263
rect 35716 31220 35768 31229
rect 32312 31084 32364 31136
rect 35624 31152 35676 31204
rect 43076 31288 43128 31340
rect 42708 31220 42760 31272
rect 44732 31263 44784 31272
rect 44732 31229 44741 31263
rect 44741 31229 44775 31263
rect 44775 31229 44784 31263
rect 44732 31220 44784 31229
rect 35164 31084 35216 31136
rect 45008 31152 45060 31204
rect 45192 31152 45244 31204
rect 36544 31127 36596 31136
rect 36544 31093 36553 31127
rect 36553 31093 36587 31127
rect 36587 31093 36596 31127
rect 36544 31084 36596 31093
rect 36728 31084 36780 31136
rect 36912 31127 36964 31136
rect 36912 31093 36921 31127
rect 36921 31093 36955 31127
rect 36955 31093 36964 31127
rect 36912 31084 36964 31093
rect 37372 31084 37424 31136
rect 37924 31084 37976 31136
rect 40408 31084 40460 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 4988 30880 5040 30932
rect 12900 30880 12952 30932
rect 13360 30880 13412 30932
rect 17960 30880 18012 30932
rect 21088 30923 21140 30932
rect 21088 30889 21097 30923
rect 21097 30889 21131 30923
rect 21131 30889 21140 30923
rect 21088 30880 21140 30889
rect 21640 30880 21692 30932
rect 23756 30880 23808 30932
rect 1768 30719 1820 30728
rect 1768 30685 1777 30719
rect 1777 30685 1811 30719
rect 1811 30685 1820 30719
rect 1768 30676 1820 30685
rect 2044 30719 2096 30728
rect 2044 30685 2078 30719
rect 2078 30685 2096 30719
rect 2044 30676 2096 30685
rect 10140 30812 10192 30864
rect 10968 30787 11020 30796
rect 10968 30753 10977 30787
rect 10977 30753 11011 30787
rect 11011 30753 11020 30787
rect 10968 30744 11020 30753
rect 13636 30787 13688 30796
rect 13636 30753 13645 30787
rect 13645 30753 13679 30787
rect 13679 30753 13688 30787
rect 13636 30744 13688 30753
rect 20996 30855 21048 30864
rect 20996 30821 21005 30855
rect 21005 30821 21039 30855
rect 21039 30821 21048 30855
rect 20996 30812 21048 30821
rect 22468 30744 22520 30796
rect 22836 30787 22888 30796
rect 22836 30753 22845 30787
rect 22845 30753 22879 30787
rect 22879 30753 22888 30787
rect 22836 30744 22888 30753
rect 4804 30676 4856 30728
rect 2596 30608 2648 30660
rect 4620 30608 4672 30660
rect 3148 30583 3200 30592
rect 3148 30549 3157 30583
rect 3157 30549 3191 30583
rect 3191 30549 3200 30583
rect 3148 30540 3200 30549
rect 3792 30583 3844 30592
rect 3792 30549 3801 30583
rect 3801 30549 3835 30583
rect 3835 30549 3844 30583
rect 3792 30540 3844 30549
rect 4160 30540 4212 30592
rect 16028 30676 16080 30728
rect 16488 30676 16540 30728
rect 21916 30719 21968 30728
rect 21916 30685 21925 30719
rect 21925 30685 21959 30719
rect 21959 30685 21968 30719
rect 21916 30676 21968 30685
rect 24492 30880 24544 30932
rect 24860 30880 24912 30932
rect 27528 30880 27580 30932
rect 31852 30880 31904 30932
rect 31944 30923 31996 30932
rect 31944 30889 31953 30923
rect 31953 30889 31987 30923
rect 31987 30889 31996 30923
rect 31944 30880 31996 30889
rect 33140 30880 33192 30932
rect 33784 30880 33836 30932
rect 34336 30880 34388 30932
rect 35072 30880 35124 30932
rect 35440 30880 35492 30932
rect 24676 30744 24728 30796
rect 24952 30787 25004 30796
rect 24952 30753 24961 30787
rect 24961 30753 24995 30787
rect 24995 30753 25004 30787
rect 24952 30744 25004 30753
rect 27344 30812 27396 30864
rect 27988 30812 28040 30864
rect 31668 30812 31720 30864
rect 27804 30787 27856 30796
rect 27804 30753 27813 30787
rect 27813 30753 27847 30787
rect 27847 30753 27856 30787
rect 27804 30744 27856 30753
rect 30564 30787 30616 30796
rect 30564 30753 30573 30787
rect 30573 30753 30607 30787
rect 30607 30753 30616 30787
rect 30564 30744 30616 30753
rect 32128 30787 32180 30796
rect 32128 30753 32137 30787
rect 32137 30753 32171 30787
rect 32171 30753 32180 30787
rect 32128 30744 32180 30753
rect 32496 30744 32548 30796
rect 32772 30787 32824 30796
rect 32772 30753 32781 30787
rect 32781 30753 32815 30787
rect 32815 30753 32824 30787
rect 32772 30744 32824 30753
rect 34520 30812 34572 30864
rect 28632 30676 28684 30728
rect 30840 30719 30892 30728
rect 30840 30685 30874 30719
rect 30874 30685 30892 30719
rect 5448 30608 5500 30660
rect 8300 30608 8352 30660
rect 13360 30608 13412 30660
rect 15752 30608 15804 30660
rect 21732 30651 21784 30660
rect 21732 30617 21741 30651
rect 21741 30617 21775 30651
rect 21775 30617 21784 30651
rect 21732 30608 21784 30617
rect 6828 30540 6880 30592
rect 10140 30540 10192 30592
rect 13544 30583 13596 30592
rect 13544 30549 13553 30583
rect 13553 30549 13587 30583
rect 13587 30549 13596 30583
rect 13544 30540 13596 30549
rect 19340 30540 19392 30592
rect 20812 30540 20864 30592
rect 21088 30540 21140 30592
rect 21456 30540 21508 30592
rect 26056 30608 26108 30660
rect 29092 30608 29144 30660
rect 30840 30676 30892 30685
rect 32312 30719 32364 30728
rect 32312 30685 32321 30719
rect 32321 30685 32355 30719
rect 32355 30685 32364 30719
rect 32312 30676 32364 30685
rect 33048 30719 33100 30728
rect 33048 30685 33057 30719
rect 33057 30685 33091 30719
rect 33091 30685 33100 30719
rect 33048 30676 33100 30685
rect 33140 30719 33192 30728
rect 33140 30685 33174 30719
rect 33174 30685 33192 30719
rect 33140 30676 33192 30685
rect 33324 30719 33376 30728
rect 33324 30685 33333 30719
rect 33333 30685 33367 30719
rect 33367 30685 33376 30719
rect 33324 30676 33376 30685
rect 34704 30719 34756 30728
rect 34704 30685 34713 30719
rect 34713 30685 34747 30719
rect 34747 30685 34756 30719
rect 34704 30676 34756 30685
rect 31208 30608 31260 30660
rect 25872 30540 25924 30592
rect 29736 30540 29788 30592
rect 30840 30540 30892 30592
rect 32220 30540 32272 30592
rect 35072 30719 35124 30728
rect 35072 30685 35081 30719
rect 35081 30685 35115 30719
rect 35115 30685 35124 30719
rect 35072 30676 35124 30685
rect 35164 30719 35216 30728
rect 35164 30685 35178 30719
rect 35178 30685 35212 30719
rect 35212 30685 35216 30719
rect 35164 30676 35216 30685
rect 35992 30676 36044 30728
rect 36084 30676 36136 30728
rect 40500 30880 40552 30932
rect 46204 30812 46256 30864
rect 36360 30744 36412 30796
rect 36452 30719 36504 30728
rect 36452 30685 36461 30719
rect 36461 30685 36495 30719
rect 36495 30685 36504 30719
rect 36452 30676 36504 30685
rect 39120 30744 39172 30796
rect 40224 30744 40276 30796
rect 37280 30676 37332 30728
rect 37372 30719 37424 30728
rect 37372 30685 37381 30719
rect 37381 30685 37415 30719
rect 37415 30685 37424 30719
rect 37372 30676 37424 30685
rect 37648 30719 37700 30728
rect 37648 30685 37657 30719
rect 37657 30685 37691 30719
rect 37691 30685 37700 30719
rect 37648 30676 37700 30685
rect 40040 30719 40092 30728
rect 40040 30685 40049 30719
rect 40049 30685 40083 30719
rect 40083 30685 40092 30719
rect 40040 30676 40092 30685
rect 35624 30540 35676 30592
rect 36360 30651 36412 30660
rect 36360 30617 36369 30651
rect 36369 30617 36403 30651
rect 36403 30617 36412 30651
rect 36360 30608 36412 30617
rect 40316 30719 40368 30728
rect 40316 30685 40325 30719
rect 40325 30685 40359 30719
rect 40359 30685 40368 30719
rect 40316 30676 40368 30685
rect 40408 30719 40460 30728
rect 40408 30685 40417 30719
rect 40417 30685 40451 30719
rect 40451 30685 40460 30719
rect 40408 30676 40460 30685
rect 45376 30787 45428 30796
rect 45376 30753 45385 30787
rect 45385 30753 45419 30787
rect 45419 30753 45428 30787
rect 45376 30744 45428 30753
rect 45744 30744 45796 30796
rect 45468 30719 45520 30728
rect 45468 30685 45477 30719
rect 45477 30685 45511 30719
rect 45511 30685 45520 30719
rect 45468 30676 45520 30685
rect 46112 30719 46164 30728
rect 46112 30685 46121 30719
rect 46121 30685 46155 30719
rect 46155 30685 46164 30719
rect 46112 30676 46164 30685
rect 36452 30540 36504 30592
rect 37740 30540 37792 30592
rect 39396 30540 39448 30592
rect 40408 30540 40460 30592
rect 40960 30583 41012 30592
rect 40960 30549 40969 30583
rect 40969 30549 41003 30583
rect 41003 30549 41012 30583
rect 40960 30540 41012 30549
rect 45928 30583 45980 30592
rect 45928 30549 45937 30583
rect 45937 30549 45971 30583
rect 45971 30549 45980 30583
rect 45928 30540 45980 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 2228 30336 2280 30388
rect 2412 30311 2464 30320
rect 2412 30277 2421 30311
rect 2421 30277 2455 30311
rect 2455 30277 2464 30311
rect 2412 30268 2464 30277
rect 3148 30336 3200 30388
rect 3792 30268 3844 30320
rect 4620 30336 4672 30388
rect 5448 30379 5500 30388
rect 5448 30345 5457 30379
rect 5457 30345 5491 30379
rect 5491 30345 5500 30379
rect 5448 30336 5500 30345
rect 6828 30379 6880 30388
rect 6828 30345 6837 30379
rect 6837 30345 6871 30379
rect 6871 30345 6880 30379
rect 6828 30336 6880 30345
rect 18328 30336 18380 30388
rect 18696 30336 18748 30388
rect 18788 30379 18840 30388
rect 18788 30345 18797 30379
rect 18797 30345 18831 30379
rect 18831 30345 18840 30379
rect 18788 30336 18840 30345
rect 19340 30336 19392 30388
rect 20352 30336 20404 30388
rect 20536 30336 20588 30388
rect 8300 30268 8352 30320
rect 16028 30311 16080 30320
rect 16028 30277 16037 30311
rect 16037 30277 16071 30311
rect 16071 30277 16080 30311
rect 16028 30268 16080 30277
rect 16120 30268 16172 30320
rect 3056 30200 3108 30252
rect 2412 30132 2464 30184
rect 2596 30132 2648 30184
rect 8576 30200 8628 30252
rect 9956 30200 10008 30252
rect 11980 30243 12032 30252
rect 11980 30209 11989 30243
rect 11989 30209 12023 30243
rect 12023 30209 12032 30243
rect 11980 30200 12032 30209
rect 7656 30132 7708 30184
rect 4804 29996 4856 30048
rect 10508 30132 10560 30184
rect 13728 30175 13780 30184
rect 13728 30141 13737 30175
rect 13737 30141 13771 30175
rect 13771 30141 13780 30175
rect 13728 30132 13780 30141
rect 15936 30243 15988 30252
rect 15936 30209 15945 30243
rect 15945 30209 15979 30243
rect 15979 30209 15988 30243
rect 15936 30200 15988 30209
rect 16488 30268 16540 30320
rect 10692 30064 10744 30116
rect 12716 30064 12768 30116
rect 16120 30132 16172 30184
rect 16304 30200 16356 30252
rect 17040 30243 17092 30252
rect 17040 30209 17049 30243
rect 17049 30209 17083 30243
rect 17083 30209 17092 30243
rect 17040 30200 17092 30209
rect 16396 30132 16448 30184
rect 17684 30132 17736 30184
rect 17960 30132 18012 30184
rect 18512 30132 18564 30184
rect 19984 30268 20036 30320
rect 21732 30268 21784 30320
rect 20904 30243 20956 30252
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 20904 30200 20956 30209
rect 21364 30243 21416 30252
rect 21364 30209 21373 30243
rect 21373 30209 21407 30243
rect 21407 30209 21416 30243
rect 21364 30200 21416 30209
rect 18880 30132 18932 30184
rect 18972 30175 19024 30184
rect 18972 30141 18981 30175
rect 18981 30141 19015 30175
rect 19015 30141 19024 30175
rect 18972 30132 19024 30141
rect 19340 30175 19392 30184
rect 19340 30141 19349 30175
rect 19349 30141 19383 30175
rect 19383 30141 19392 30175
rect 19340 30132 19392 30141
rect 19892 30132 19944 30184
rect 21640 30243 21692 30252
rect 21640 30209 21649 30243
rect 21649 30209 21683 30243
rect 21683 30209 21692 30243
rect 21640 30200 21692 30209
rect 21916 30336 21968 30388
rect 24952 30336 25004 30388
rect 25136 30336 25188 30388
rect 31668 30336 31720 30388
rect 30840 30311 30892 30320
rect 21916 30200 21968 30252
rect 23572 30200 23624 30252
rect 22468 30132 22520 30184
rect 23756 30132 23808 30184
rect 24400 30243 24452 30252
rect 24400 30209 24409 30243
rect 24409 30209 24443 30243
rect 24443 30209 24452 30243
rect 24400 30200 24452 30209
rect 24584 30200 24636 30252
rect 24216 30132 24268 30184
rect 24676 30175 24728 30184
rect 24676 30141 24685 30175
rect 24685 30141 24719 30175
rect 24719 30141 24728 30175
rect 24676 30132 24728 30141
rect 9312 30039 9364 30048
rect 9312 30005 9321 30039
rect 9321 30005 9355 30039
rect 9355 30005 9364 30039
rect 9312 29996 9364 30005
rect 11612 29996 11664 30048
rect 13176 29996 13228 30048
rect 13636 29996 13688 30048
rect 14004 30064 14056 30116
rect 15384 29996 15436 30048
rect 15660 29996 15712 30048
rect 17040 29996 17092 30048
rect 18144 29996 18196 30048
rect 18420 29996 18472 30048
rect 18512 29996 18564 30048
rect 18788 29996 18840 30048
rect 19064 29996 19116 30048
rect 19248 30064 19300 30116
rect 19340 29996 19392 30048
rect 23848 30064 23900 30116
rect 21088 29996 21140 30048
rect 21180 30039 21232 30048
rect 21180 30005 21189 30039
rect 21189 30005 21223 30039
rect 21223 30005 21232 30039
rect 21180 29996 21232 30005
rect 25320 30200 25372 30252
rect 25872 30243 25924 30252
rect 25872 30209 25881 30243
rect 25881 30209 25915 30243
rect 25915 30209 25924 30243
rect 25872 30200 25924 30209
rect 25412 30132 25464 30184
rect 26792 30243 26844 30252
rect 26792 30209 26801 30243
rect 26801 30209 26835 30243
rect 26835 30209 26844 30243
rect 26792 30200 26844 30209
rect 26240 30132 26292 30184
rect 30840 30277 30874 30311
rect 30874 30277 30892 30311
rect 30840 30268 30892 30277
rect 32036 30336 32088 30388
rect 32772 30336 32824 30388
rect 33324 30336 33376 30388
rect 34428 30336 34480 30388
rect 34704 30336 34756 30388
rect 28080 30200 28132 30252
rect 29736 30200 29788 30252
rect 25504 29996 25556 30048
rect 25688 29996 25740 30048
rect 30380 30132 30432 30184
rect 30564 30175 30616 30184
rect 30564 30141 30573 30175
rect 30573 30141 30607 30175
rect 30607 30141 30616 30175
rect 30564 30132 30616 30141
rect 32128 30243 32180 30252
rect 32128 30209 32137 30243
rect 32137 30209 32171 30243
rect 32171 30209 32180 30243
rect 32128 30200 32180 30209
rect 37280 30268 37332 30320
rect 37464 30268 37516 30320
rect 32312 30175 32364 30184
rect 32312 30141 32321 30175
rect 32321 30141 32355 30175
rect 32355 30141 32364 30175
rect 32312 30132 32364 30141
rect 33140 30243 33192 30252
rect 33140 30209 33174 30243
rect 33174 30209 33192 30243
rect 33140 30200 33192 30209
rect 34704 30200 34756 30252
rect 35072 30200 35124 30252
rect 36452 30200 36504 30252
rect 33048 30175 33100 30184
rect 33048 30141 33057 30175
rect 33057 30141 33091 30175
rect 33091 30141 33100 30175
rect 33048 30132 33100 30141
rect 33324 30175 33376 30184
rect 33324 30141 33333 30175
rect 33333 30141 33367 30175
rect 33367 30141 33376 30175
rect 33324 30132 33376 30141
rect 37004 30200 37056 30252
rect 38384 30243 38436 30252
rect 38384 30209 38393 30243
rect 38393 30209 38427 30243
rect 38427 30209 38436 30243
rect 38384 30200 38436 30209
rect 45376 30336 45428 30388
rect 39120 30200 39172 30252
rect 39304 30200 39356 30252
rect 39396 30243 39448 30252
rect 39396 30209 39405 30243
rect 39405 30209 39439 30243
rect 39439 30209 39448 30243
rect 39396 30200 39448 30209
rect 40040 30200 40092 30252
rect 40316 30200 40368 30252
rect 40500 30243 40552 30252
rect 40500 30209 40509 30243
rect 40509 30209 40543 30243
rect 40543 30209 40552 30243
rect 40500 30200 40552 30209
rect 28264 29996 28316 30048
rect 28356 30039 28408 30048
rect 28356 30005 28365 30039
rect 28365 30005 28399 30039
rect 28399 30005 28408 30039
rect 28356 29996 28408 30005
rect 32864 30064 32916 30116
rect 35624 30064 35676 30116
rect 36360 30064 36412 30116
rect 34060 29996 34112 30048
rect 36452 29996 36504 30048
rect 36912 29996 36964 30048
rect 37280 29996 37332 30048
rect 38016 29996 38068 30048
rect 38936 30064 38988 30116
rect 39120 30107 39172 30116
rect 39120 30073 39129 30107
rect 39129 30073 39163 30107
rect 39163 30073 39172 30107
rect 39120 30064 39172 30073
rect 39488 30175 39540 30184
rect 39488 30141 39497 30175
rect 39497 30141 39531 30175
rect 39531 30141 39540 30175
rect 39488 30132 39540 30141
rect 39672 30175 39724 30184
rect 39672 30141 39681 30175
rect 39681 30141 39715 30175
rect 39715 30141 39724 30175
rect 39672 30132 39724 30141
rect 42340 30268 42392 30320
rect 41604 30243 41656 30252
rect 41604 30209 41613 30243
rect 41613 30209 41647 30243
rect 41647 30209 41656 30243
rect 41604 30200 41656 30209
rect 41788 30243 41840 30252
rect 41788 30209 41795 30243
rect 41795 30209 41840 30243
rect 41788 30200 41840 30209
rect 41236 30132 41288 30184
rect 41052 30064 41104 30116
rect 43168 30200 43220 30252
rect 43720 30243 43772 30252
rect 43720 30209 43729 30243
rect 43729 30209 43763 30243
rect 43763 30209 43772 30243
rect 43720 30200 43772 30209
rect 44088 30243 44140 30252
rect 44088 30209 44097 30243
rect 44097 30209 44131 30243
rect 44131 30209 44140 30243
rect 44088 30200 44140 30209
rect 44272 30243 44324 30252
rect 44272 30209 44281 30243
rect 44281 30209 44315 30243
rect 44315 30209 44324 30243
rect 44272 30200 44324 30209
rect 44456 30243 44508 30252
rect 44456 30209 44465 30243
rect 44465 30209 44499 30243
rect 44499 30209 44508 30243
rect 44456 30200 44508 30209
rect 45376 30200 45428 30252
rect 45928 30200 45980 30252
rect 44916 30132 44968 30184
rect 45284 30064 45336 30116
rect 46204 30132 46256 30184
rect 39948 29996 40000 30048
rect 40868 29996 40920 30048
rect 42156 29996 42208 30048
rect 43904 30039 43956 30048
rect 43904 30005 43913 30039
rect 43913 30005 43947 30039
rect 43947 30005 43956 30039
rect 43904 29996 43956 30005
rect 45468 29996 45520 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 8576 29835 8628 29844
rect 8576 29801 8585 29835
rect 8585 29801 8619 29835
rect 8619 29801 8628 29835
rect 8576 29792 8628 29801
rect 17040 29792 17092 29844
rect 5264 29724 5316 29776
rect 9312 29724 9364 29776
rect 1676 29699 1728 29708
rect 1676 29665 1685 29699
rect 1685 29665 1719 29699
rect 1719 29665 1728 29699
rect 1676 29656 1728 29665
rect 6828 29656 6880 29708
rect 7472 29656 7524 29708
rect 19708 29792 19760 29844
rect 20720 29835 20772 29844
rect 20720 29801 20729 29835
rect 20729 29801 20763 29835
rect 20763 29801 20772 29835
rect 20720 29792 20772 29801
rect 21180 29792 21232 29844
rect 25412 29792 25464 29844
rect 25688 29835 25740 29844
rect 25688 29801 25697 29835
rect 25697 29801 25731 29835
rect 25731 29801 25740 29835
rect 25688 29792 25740 29801
rect 26792 29792 26844 29844
rect 27344 29792 27396 29844
rect 27804 29792 27856 29844
rect 28264 29792 28316 29844
rect 31484 29792 31536 29844
rect 38568 29835 38620 29844
rect 38568 29801 38577 29835
rect 38577 29801 38611 29835
rect 38611 29801 38620 29835
rect 38568 29792 38620 29801
rect 39672 29792 39724 29844
rect 39948 29792 40000 29844
rect 40684 29792 40736 29844
rect 25320 29724 25372 29776
rect 25504 29767 25556 29776
rect 25504 29733 25513 29767
rect 25513 29733 25547 29767
rect 25547 29733 25556 29767
rect 25504 29724 25556 29733
rect 26148 29724 26200 29776
rect 10232 29656 10284 29708
rect 10324 29656 10376 29708
rect 10692 29699 10744 29708
rect 10692 29665 10701 29699
rect 10701 29665 10735 29699
rect 10735 29665 10744 29699
rect 10692 29656 10744 29665
rect 15108 29656 15160 29708
rect 940 29588 992 29640
rect 6368 29588 6420 29640
rect 8300 29588 8352 29640
rect 7656 29563 7708 29572
rect 7656 29529 7665 29563
rect 7665 29529 7699 29563
rect 7699 29529 7708 29563
rect 7656 29520 7708 29529
rect 5448 29495 5500 29504
rect 5448 29461 5457 29495
rect 5457 29461 5491 29495
rect 5491 29461 5500 29495
rect 5448 29452 5500 29461
rect 6920 29452 6972 29504
rect 10508 29588 10560 29640
rect 11612 29631 11664 29640
rect 11612 29597 11646 29631
rect 11646 29597 11664 29631
rect 11612 29588 11664 29597
rect 15384 29631 15436 29640
rect 15384 29597 15393 29631
rect 15393 29597 15427 29631
rect 15427 29597 15436 29631
rect 15384 29588 15436 29597
rect 15660 29631 15712 29640
rect 15660 29597 15669 29631
rect 15669 29597 15703 29631
rect 15703 29597 15712 29631
rect 15660 29588 15712 29597
rect 16764 29656 16816 29708
rect 17224 29699 17276 29708
rect 17224 29665 17233 29699
rect 17233 29665 17267 29699
rect 17267 29665 17276 29699
rect 17224 29656 17276 29665
rect 17776 29656 17828 29708
rect 17960 29656 18012 29708
rect 18144 29699 18196 29708
rect 18144 29665 18153 29699
rect 18153 29665 18187 29699
rect 18187 29665 18196 29699
rect 18144 29656 18196 29665
rect 19892 29656 19944 29708
rect 20444 29656 20496 29708
rect 21088 29656 21140 29708
rect 21456 29656 21508 29708
rect 27344 29656 27396 29708
rect 27528 29656 27580 29708
rect 37740 29724 37792 29776
rect 39304 29724 39356 29776
rect 40040 29724 40092 29776
rect 17408 29631 17460 29640
rect 17408 29597 17417 29631
rect 17417 29597 17451 29631
rect 17451 29597 17460 29631
rect 17408 29588 17460 29597
rect 18328 29588 18380 29640
rect 15108 29520 15160 29572
rect 12624 29452 12676 29504
rect 15200 29495 15252 29504
rect 15200 29461 15209 29495
rect 15209 29461 15243 29495
rect 15243 29461 15252 29495
rect 15200 29452 15252 29461
rect 16120 29452 16172 29504
rect 18328 29452 18380 29504
rect 18512 29452 18564 29504
rect 18880 29452 18932 29504
rect 20904 29631 20956 29640
rect 20904 29597 20913 29631
rect 20913 29597 20947 29631
rect 20947 29597 20956 29631
rect 20904 29588 20956 29597
rect 21180 29631 21232 29640
rect 21180 29597 21189 29631
rect 21189 29597 21223 29631
rect 21223 29597 21232 29631
rect 21180 29588 21232 29597
rect 21916 29631 21968 29640
rect 21916 29597 21925 29631
rect 21925 29597 21959 29631
rect 21959 29597 21968 29631
rect 21916 29588 21968 29597
rect 22468 29631 22520 29640
rect 22468 29597 22477 29631
rect 22477 29597 22511 29631
rect 22511 29597 22520 29631
rect 22468 29588 22520 29597
rect 22652 29588 22704 29640
rect 23480 29588 23532 29640
rect 20904 29452 20956 29504
rect 21456 29563 21508 29572
rect 21456 29529 21465 29563
rect 21465 29529 21499 29563
rect 21499 29529 21508 29563
rect 21456 29520 21508 29529
rect 24952 29520 25004 29572
rect 25228 29563 25280 29572
rect 25228 29529 25237 29563
rect 25237 29529 25271 29563
rect 25271 29529 25280 29563
rect 25228 29520 25280 29529
rect 28908 29588 28960 29640
rect 29092 29588 29144 29640
rect 29460 29588 29512 29640
rect 35440 29631 35492 29640
rect 35440 29597 35449 29631
rect 35449 29597 35483 29631
rect 35483 29597 35492 29631
rect 35440 29588 35492 29597
rect 35624 29631 35676 29640
rect 35624 29597 35633 29631
rect 35633 29597 35667 29631
rect 35667 29597 35676 29631
rect 35624 29588 35676 29597
rect 35992 29588 36044 29640
rect 37096 29588 37148 29640
rect 30012 29520 30064 29572
rect 31576 29520 31628 29572
rect 34060 29520 34112 29572
rect 22284 29452 22336 29504
rect 22560 29452 22612 29504
rect 24216 29452 24268 29504
rect 28356 29452 28408 29504
rect 29552 29452 29604 29504
rect 33600 29452 33652 29504
rect 36636 29520 36688 29572
rect 37740 29563 37792 29572
rect 37740 29529 37749 29563
rect 37749 29529 37783 29563
rect 37783 29529 37792 29563
rect 37740 29520 37792 29529
rect 38200 29588 38252 29640
rect 40224 29588 40276 29640
rect 41144 29724 41196 29776
rect 42156 29835 42208 29844
rect 42156 29801 42165 29835
rect 42165 29801 42199 29835
rect 42199 29801 42208 29835
rect 42156 29792 42208 29801
rect 44272 29792 44324 29844
rect 45100 29792 45152 29844
rect 46020 29792 46072 29844
rect 42616 29724 42668 29776
rect 40960 29656 41012 29708
rect 42524 29699 42576 29708
rect 42524 29665 42533 29699
rect 42533 29665 42567 29699
rect 42567 29665 42576 29699
rect 42524 29656 42576 29665
rect 42708 29656 42760 29708
rect 36544 29452 36596 29504
rect 37464 29452 37516 29504
rect 38384 29452 38436 29504
rect 38844 29452 38896 29504
rect 39028 29452 39080 29504
rect 40132 29452 40184 29504
rect 40868 29520 40920 29572
rect 41144 29588 41196 29640
rect 41696 29520 41748 29572
rect 42064 29631 42116 29640
rect 42064 29597 42073 29631
rect 42073 29597 42107 29631
rect 42107 29597 42116 29631
rect 42064 29588 42116 29597
rect 43168 29724 43220 29776
rect 44180 29724 44232 29776
rect 41880 29520 41932 29572
rect 43076 29588 43128 29640
rect 43904 29656 43956 29708
rect 45008 29699 45060 29708
rect 45008 29665 45017 29699
rect 45017 29665 45051 29699
rect 45051 29665 45060 29699
rect 45008 29656 45060 29665
rect 42892 29520 42944 29572
rect 44732 29588 44784 29640
rect 45468 29631 45520 29640
rect 45468 29597 45477 29631
rect 45477 29597 45511 29631
rect 45511 29597 45520 29631
rect 45468 29588 45520 29597
rect 45376 29563 45428 29572
rect 45376 29529 45385 29563
rect 45385 29529 45419 29563
rect 45419 29529 45428 29563
rect 46020 29588 46072 29640
rect 45376 29520 45428 29529
rect 40960 29495 41012 29504
rect 40960 29461 40969 29495
rect 40969 29461 41003 29495
rect 41003 29461 41012 29495
rect 40960 29452 41012 29461
rect 41144 29452 41196 29504
rect 45468 29452 45520 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 2412 29248 2464 29300
rect 5448 29180 5500 29232
rect 6368 29291 6420 29300
rect 6368 29257 6377 29291
rect 6377 29257 6411 29291
rect 6411 29257 6420 29291
rect 6368 29248 6420 29257
rect 9036 29248 9088 29300
rect 9404 29180 9456 29232
rect 6736 29155 6788 29164
rect 6736 29121 6745 29155
rect 6745 29121 6779 29155
rect 6779 29121 6788 29155
rect 6736 29112 6788 29121
rect 4620 29044 4672 29096
rect 4804 29087 4856 29096
rect 4804 29053 4813 29087
rect 4813 29053 4847 29087
rect 4847 29053 4856 29087
rect 4804 29044 4856 29053
rect 7656 29112 7708 29164
rect 7840 29155 7892 29164
rect 7840 29121 7874 29155
rect 7874 29121 7892 29155
rect 7840 29112 7892 29121
rect 9312 29112 9364 29164
rect 9956 29180 10008 29232
rect 15476 29248 15528 29300
rect 15936 29248 15988 29300
rect 17408 29248 17460 29300
rect 11060 29112 11112 29164
rect 13084 29155 13136 29164
rect 13084 29121 13093 29155
rect 13093 29121 13127 29155
rect 13127 29121 13136 29155
rect 13084 29112 13136 29121
rect 7288 28976 7340 29028
rect 9956 29087 10008 29096
rect 9956 29053 9965 29087
rect 9965 29053 9999 29087
rect 9999 29053 10008 29087
rect 9956 29044 10008 29053
rect 10968 29044 11020 29096
rect 14096 29112 14148 29164
rect 15200 29180 15252 29232
rect 17500 29180 17552 29232
rect 17224 29112 17276 29164
rect 19248 29291 19300 29300
rect 19248 29257 19257 29291
rect 19257 29257 19291 29291
rect 19291 29257 19300 29291
rect 19248 29248 19300 29257
rect 19984 29180 20036 29232
rect 18512 29112 18564 29164
rect 19248 29112 19300 29164
rect 20812 29112 20864 29164
rect 29368 29112 29420 29164
rect 29552 29155 29604 29164
rect 29552 29121 29561 29155
rect 29561 29121 29595 29155
rect 29595 29121 29604 29155
rect 29552 29112 29604 29121
rect 29644 29155 29696 29164
rect 29644 29121 29653 29155
rect 29653 29121 29687 29155
rect 29687 29121 29696 29155
rect 29644 29112 29696 29121
rect 34152 29180 34204 29232
rect 37280 29248 37332 29300
rect 32128 29112 32180 29164
rect 33600 29155 33652 29164
rect 33600 29121 33609 29155
rect 33609 29121 33643 29155
rect 33643 29121 33652 29155
rect 33600 29112 33652 29121
rect 33876 29155 33928 29164
rect 33876 29121 33910 29155
rect 33910 29121 33928 29155
rect 33876 29112 33928 29121
rect 36820 29180 36872 29232
rect 9864 28976 9916 29028
rect 9312 28908 9364 28960
rect 9404 28908 9456 28960
rect 11336 28951 11388 28960
rect 11336 28917 11345 28951
rect 11345 28917 11379 28951
rect 11379 28917 11388 28951
rect 11336 28908 11388 28917
rect 13176 28976 13228 29028
rect 12716 28951 12768 28960
rect 12716 28917 12725 28951
rect 12725 28917 12759 28951
rect 12759 28917 12768 28951
rect 12716 28908 12768 28917
rect 15108 29087 15160 29096
rect 15108 29053 15117 29087
rect 15117 29053 15151 29087
rect 15151 29053 15160 29087
rect 15108 29044 15160 29053
rect 17316 29044 17368 29096
rect 16764 28976 16816 29028
rect 17684 28976 17736 29028
rect 17960 29044 18012 29096
rect 18604 29087 18656 29096
rect 18604 29053 18613 29087
rect 18613 29053 18647 29087
rect 18647 29053 18656 29087
rect 18604 29044 18656 29053
rect 18788 29044 18840 29096
rect 29460 29044 29512 29096
rect 18144 28976 18196 29028
rect 21456 28976 21508 29028
rect 32864 29044 32916 29096
rect 33232 29044 33284 29096
rect 34612 29044 34664 29096
rect 30012 29019 30064 29028
rect 30012 28985 30021 29019
rect 30021 28985 30055 29019
rect 30055 28985 30064 29019
rect 30012 28976 30064 28985
rect 15108 28908 15160 28960
rect 18696 28908 18748 28960
rect 32680 28908 32732 28960
rect 33416 28908 33468 28960
rect 35992 29044 36044 29096
rect 36360 29155 36412 29164
rect 36360 29121 36369 29155
rect 36369 29121 36403 29155
rect 36403 29121 36412 29155
rect 36360 29112 36412 29121
rect 36728 29112 36780 29164
rect 37280 29155 37332 29164
rect 37280 29121 37289 29155
rect 37289 29121 37323 29155
rect 37323 29121 37332 29155
rect 37280 29112 37332 29121
rect 38108 29248 38160 29300
rect 38292 29248 38344 29300
rect 38844 29248 38896 29300
rect 39488 29248 39540 29300
rect 41328 29248 41380 29300
rect 38108 29155 38160 29164
rect 38108 29121 38117 29155
rect 38117 29121 38151 29155
rect 38151 29121 38160 29155
rect 38108 29112 38160 29121
rect 38844 29112 38896 29164
rect 39304 29180 39356 29232
rect 40132 29180 40184 29232
rect 41236 29180 41288 29232
rect 39120 29155 39172 29164
rect 39120 29121 39129 29155
rect 39129 29121 39163 29155
rect 39163 29121 39172 29155
rect 39120 29112 39172 29121
rect 40960 29112 41012 29164
rect 41144 29112 41196 29164
rect 41512 29155 41564 29164
rect 41512 29121 41521 29155
rect 41521 29121 41555 29155
rect 41555 29121 41564 29155
rect 41512 29112 41564 29121
rect 41972 29248 42024 29300
rect 37740 28976 37792 29028
rect 39028 28976 39080 29028
rect 40040 29044 40092 29096
rect 41328 29044 41380 29096
rect 41880 29155 41932 29164
rect 41880 29121 41889 29155
rect 41889 29121 41923 29155
rect 41923 29121 41932 29155
rect 41880 29112 41932 29121
rect 42064 29155 42116 29164
rect 42064 29121 42073 29155
rect 42073 29121 42107 29155
rect 42107 29121 42116 29155
rect 42064 29112 42116 29121
rect 42156 29112 42208 29164
rect 42616 29155 42668 29164
rect 42616 29121 42625 29155
rect 42625 29121 42659 29155
rect 42659 29121 42668 29155
rect 42616 29112 42668 29121
rect 43076 29180 43128 29232
rect 43168 29112 43220 29164
rect 46664 29291 46716 29300
rect 46664 29257 46673 29291
rect 46673 29257 46707 29291
rect 46707 29257 46716 29291
rect 46664 29248 46716 29257
rect 43720 29044 43772 29096
rect 44732 29044 44784 29096
rect 45008 29044 45060 29096
rect 42156 28976 42208 29028
rect 37832 28951 37884 28960
rect 37832 28917 37841 28951
rect 37841 28917 37875 28951
rect 37875 28917 37884 28951
rect 37832 28908 37884 28917
rect 41420 28908 41472 28960
rect 41604 28908 41656 28960
rect 41972 28908 42024 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 7840 28704 7892 28756
rect 11060 28704 11112 28756
rect 14096 28747 14148 28756
rect 14096 28713 14105 28747
rect 14105 28713 14139 28747
rect 14139 28713 14148 28747
rect 14096 28704 14148 28713
rect 5908 28679 5960 28688
rect 5908 28645 5917 28679
rect 5917 28645 5951 28679
rect 5951 28645 5960 28679
rect 5908 28636 5960 28645
rect 6736 28636 6788 28688
rect 10968 28636 11020 28688
rect 14004 28636 14056 28688
rect 19248 28704 19300 28756
rect 20260 28704 20312 28756
rect 20812 28704 20864 28756
rect 19800 28636 19852 28688
rect 22192 28636 22244 28688
rect 24400 28636 24452 28688
rect 24676 28636 24728 28688
rect 3240 28611 3292 28620
rect 3240 28577 3249 28611
rect 3249 28577 3283 28611
rect 3283 28577 3292 28611
rect 3240 28568 3292 28577
rect 4436 28543 4488 28552
rect 4436 28509 4445 28543
rect 4445 28509 4479 28543
rect 4479 28509 4488 28543
rect 4436 28500 4488 28509
rect 4528 28543 4580 28552
rect 4528 28509 4537 28543
rect 4537 28509 4571 28543
rect 4571 28509 4580 28543
rect 4528 28500 4580 28509
rect 7104 28568 7156 28620
rect 7288 28611 7340 28620
rect 7288 28577 7297 28611
rect 7297 28577 7331 28611
rect 7331 28577 7340 28611
rect 7288 28568 7340 28577
rect 7472 28611 7524 28620
rect 7472 28577 7481 28611
rect 7481 28577 7515 28611
rect 7515 28577 7524 28611
rect 7472 28568 7524 28577
rect 6460 28500 6512 28552
rect 6736 28500 6788 28552
rect 9404 28568 9456 28620
rect 9864 28568 9916 28620
rect 10876 28568 10928 28620
rect 11336 28568 11388 28620
rect 12624 28611 12676 28620
rect 12624 28577 12633 28611
rect 12633 28577 12667 28611
rect 12667 28577 12676 28611
rect 12624 28568 12676 28577
rect 2320 28364 2372 28416
rect 2964 28407 3016 28416
rect 2964 28373 2973 28407
rect 2973 28373 3007 28407
rect 3007 28373 3016 28407
rect 2964 28364 3016 28373
rect 4068 28364 4120 28416
rect 6828 28407 6880 28416
rect 6828 28373 6837 28407
rect 6837 28373 6871 28407
rect 6871 28373 6880 28407
rect 6828 28364 6880 28373
rect 9404 28475 9456 28484
rect 9404 28441 9413 28475
rect 9413 28441 9447 28475
rect 9447 28441 9456 28475
rect 9404 28432 9456 28441
rect 12900 28543 12952 28552
rect 12900 28509 12909 28543
rect 12909 28509 12943 28543
rect 12943 28509 12952 28543
rect 12900 28500 12952 28509
rect 13636 28500 13688 28552
rect 14280 28543 14332 28552
rect 14280 28509 14289 28543
rect 14289 28509 14323 28543
rect 14323 28509 14332 28543
rect 14280 28500 14332 28509
rect 19340 28568 19392 28620
rect 19432 28568 19484 28620
rect 22376 28568 22428 28620
rect 18420 28543 18472 28552
rect 18420 28509 18429 28543
rect 18429 28509 18463 28543
rect 18463 28509 18472 28543
rect 18420 28500 18472 28509
rect 9312 28407 9364 28416
rect 9312 28373 9321 28407
rect 9321 28373 9355 28407
rect 9355 28373 9364 28407
rect 9312 28364 9364 28373
rect 10600 28407 10652 28416
rect 10600 28373 10609 28407
rect 10609 28373 10643 28407
rect 10643 28373 10652 28407
rect 10600 28364 10652 28373
rect 11060 28407 11112 28416
rect 11060 28373 11069 28407
rect 11069 28373 11103 28407
rect 11103 28373 11112 28407
rect 11060 28364 11112 28373
rect 13820 28432 13872 28484
rect 15108 28432 15160 28484
rect 21272 28543 21324 28552
rect 21272 28509 21281 28543
rect 21281 28509 21315 28543
rect 21315 28509 21324 28543
rect 21272 28500 21324 28509
rect 21824 28500 21876 28552
rect 20168 28475 20220 28484
rect 20168 28441 20177 28475
rect 20177 28441 20211 28475
rect 20211 28441 20220 28475
rect 20168 28432 20220 28441
rect 20720 28432 20772 28484
rect 25964 28568 26016 28620
rect 29460 28704 29512 28756
rect 30196 28704 30248 28756
rect 30564 28704 30616 28756
rect 32496 28704 32548 28756
rect 32680 28704 32732 28756
rect 27252 28636 27304 28688
rect 27528 28568 27580 28620
rect 28540 28679 28592 28688
rect 28540 28645 28549 28679
rect 28549 28645 28583 28679
rect 28583 28645 28592 28679
rect 28540 28636 28592 28645
rect 22560 28500 22612 28552
rect 23296 28500 23348 28552
rect 24860 28500 24912 28552
rect 26148 28543 26200 28552
rect 26148 28509 26157 28543
rect 26157 28509 26191 28543
rect 26191 28509 26200 28543
rect 26148 28500 26200 28509
rect 22928 28432 22980 28484
rect 26608 28432 26660 28484
rect 13452 28364 13504 28416
rect 14004 28364 14056 28416
rect 14464 28407 14516 28416
rect 14464 28373 14473 28407
rect 14473 28373 14507 28407
rect 14507 28373 14516 28407
rect 14464 28364 14516 28373
rect 15384 28407 15436 28416
rect 15384 28373 15393 28407
rect 15393 28373 15427 28407
rect 15427 28373 15436 28407
rect 15384 28364 15436 28373
rect 20352 28364 20404 28416
rect 21548 28407 21600 28416
rect 21548 28373 21557 28407
rect 21557 28373 21591 28407
rect 21591 28373 21600 28407
rect 21548 28364 21600 28373
rect 21732 28364 21784 28416
rect 27252 28364 27304 28416
rect 29092 28500 29144 28552
rect 31576 28568 31628 28620
rect 32588 28611 32640 28620
rect 32588 28577 32597 28611
rect 32597 28577 32631 28611
rect 32631 28577 32640 28611
rect 32588 28568 32640 28577
rect 33324 28568 33376 28620
rect 33508 28611 33560 28620
rect 33508 28577 33517 28611
rect 33517 28577 33551 28611
rect 33551 28577 33560 28611
rect 33508 28568 33560 28577
rect 33876 28747 33928 28756
rect 33876 28713 33885 28747
rect 33885 28713 33919 28747
rect 33919 28713 33928 28747
rect 33876 28704 33928 28713
rect 35808 28704 35860 28756
rect 37648 28704 37700 28756
rect 38660 28704 38712 28756
rect 40776 28704 40828 28756
rect 44548 28704 44600 28756
rect 33876 28500 33928 28552
rect 29000 28475 29052 28484
rect 29000 28441 29009 28475
rect 29009 28441 29043 28475
rect 29043 28441 29052 28475
rect 29000 28432 29052 28441
rect 29184 28432 29236 28484
rect 32680 28432 32732 28484
rect 33416 28475 33468 28484
rect 33416 28441 33425 28475
rect 33425 28441 33459 28475
rect 33459 28441 33468 28475
rect 33416 28432 33468 28441
rect 27620 28407 27672 28416
rect 27620 28373 27629 28407
rect 27629 28373 27663 28407
rect 27663 28373 27672 28407
rect 27620 28364 27672 28373
rect 29644 28364 29696 28416
rect 29920 28364 29972 28416
rect 31944 28364 31996 28416
rect 32864 28364 32916 28416
rect 37832 28500 37884 28552
rect 42064 28611 42116 28620
rect 42064 28577 42073 28611
rect 42073 28577 42107 28611
rect 42107 28577 42116 28611
rect 42064 28568 42116 28577
rect 42432 28568 42484 28620
rect 45468 28568 45520 28620
rect 37004 28432 37056 28484
rect 41788 28543 41840 28552
rect 41788 28509 41797 28543
rect 41797 28509 41831 28543
rect 41831 28509 41840 28543
rect 41788 28500 41840 28509
rect 41972 28500 42024 28552
rect 43720 28543 43772 28552
rect 43720 28509 43729 28543
rect 43729 28509 43763 28543
rect 43763 28509 43772 28543
rect 43720 28500 43772 28509
rect 44180 28500 44232 28552
rect 44916 28500 44968 28552
rect 45008 28543 45060 28552
rect 45008 28509 45017 28543
rect 45017 28509 45051 28543
rect 45051 28509 45060 28543
rect 45008 28500 45060 28509
rect 45100 28500 45152 28552
rect 39028 28432 39080 28484
rect 42616 28364 42668 28416
rect 43996 28364 44048 28416
rect 45192 28407 45244 28416
rect 45192 28373 45201 28407
rect 45201 28373 45235 28407
rect 45235 28373 45244 28407
rect 45192 28364 45244 28373
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 11980 28160 12032 28212
rect 12716 28160 12768 28212
rect 1676 28092 1728 28144
rect 2320 28067 2372 28076
rect 2320 28033 2329 28067
rect 2329 28033 2363 28067
rect 2363 28033 2372 28067
rect 2320 28024 2372 28033
rect 4528 28092 4580 28144
rect 3148 28024 3200 28076
rect 4620 28067 4672 28076
rect 4620 28033 4629 28067
rect 4629 28033 4663 28067
rect 4663 28033 4672 28067
rect 4620 28024 4672 28033
rect 6828 28092 6880 28144
rect 6920 28024 6972 28076
rect 12900 28092 12952 28144
rect 12624 28024 12676 28076
rect 10968 27956 11020 28008
rect 14280 28160 14332 28212
rect 15016 28160 15068 28212
rect 21732 28160 21784 28212
rect 21824 28203 21876 28212
rect 21824 28169 21833 28203
rect 21833 28169 21867 28203
rect 21867 28169 21876 28203
rect 21824 28160 21876 28169
rect 26608 28203 26660 28212
rect 26608 28169 26617 28203
rect 26617 28169 26651 28203
rect 26651 28169 26660 28203
rect 26608 28160 26660 28169
rect 27988 28160 28040 28212
rect 29184 28160 29236 28212
rect 13820 28135 13872 28144
rect 13820 28101 13829 28135
rect 13829 28101 13863 28135
rect 13863 28101 13872 28135
rect 13820 28092 13872 28101
rect 13912 28092 13964 28144
rect 14372 28092 14424 28144
rect 14004 28067 14056 28076
rect 14004 28033 14013 28067
rect 14013 28033 14047 28067
rect 14047 28033 14056 28067
rect 14004 28024 14056 28033
rect 14464 28024 14516 28076
rect 16304 28092 16356 28144
rect 14556 27999 14608 28008
rect 14556 27965 14565 27999
rect 14565 27965 14599 27999
rect 14599 27965 14608 27999
rect 14556 27956 14608 27965
rect 16396 28024 16448 28076
rect 16488 28024 16540 28076
rect 11336 27888 11388 27940
rect 15200 27956 15252 28008
rect 15476 27956 15528 28008
rect 15844 27999 15896 28008
rect 15844 27965 15853 27999
rect 15853 27965 15887 27999
rect 15887 27965 15896 27999
rect 15844 27956 15896 27965
rect 16028 27999 16080 28008
rect 16028 27965 16037 27999
rect 16037 27965 16071 27999
rect 16071 27965 16080 27999
rect 16028 27956 16080 27965
rect 16212 27956 16264 28008
rect 19432 28092 19484 28144
rect 20996 28092 21048 28144
rect 22192 28135 22244 28144
rect 22192 28101 22201 28135
rect 22201 28101 22235 28135
rect 22235 28101 22244 28135
rect 22192 28092 22244 28101
rect 20168 28024 20220 28076
rect 17592 27956 17644 28008
rect 19984 27956 20036 28008
rect 20628 27956 20680 28008
rect 22744 28024 22796 28076
rect 22468 27999 22520 28008
rect 22468 27965 22477 27999
rect 22477 27965 22511 27999
rect 22511 27965 22520 27999
rect 23112 28024 23164 28076
rect 27620 28024 27672 28076
rect 28448 28024 28500 28076
rect 29644 28160 29696 28212
rect 29920 28160 29972 28212
rect 31576 28160 31628 28212
rect 32496 28160 32548 28212
rect 22468 27956 22520 27965
rect 22928 27956 22980 28008
rect 23388 27999 23440 28008
rect 23388 27965 23397 27999
rect 23397 27965 23431 27999
rect 23431 27965 23440 27999
rect 23388 27956 23440 27965
rect 1952 27820 2004 27872
rect 3976 27863 4028 27872
rect 3976 27829 3985 27863
rect 3985 27829 4019 27863
rect 4019 27829 4028 27863
rect 3976 27820 4028 27829
rect 7380 27820 7432 27872
rect 8392 27820 8444 27872
rect 12716 27820 12768 27872
rect 19524 27888 19576 27940
rect 16488 27820 16540 27872
rect 18052 27820 18104 27872
rect 18880 27820 18932 27872
rect 19340 27863 19392 27872
rect 19340 27829 19349 27863
rect 19349 27829 19383 27863
rect 19383 27829 19392 27863
rect 19340 27820 19392 27829
rect 19616 27820 19668 27872
rect 19892 27863 19944 27872
rect 19892 27829 19901 27863
rect 19901 27829 19935 27863
rect 19935 27829 19944 27863
rect 19892 27820 19944 27829
rect 20812 27820 20864 27872
rect 22100 27820 22152 27872
rect 22836 27888 22888 27940
rect 23940 27956 23992 28008
rect 24308 27956 24360 28008
rect 24400 27999 24452 28008
rect 24400 27965 24409 27999
rect 24409 27965 24443 27999
rect 24443 27965 24452 27999
rect 24400 27956 24452 27965
rect 25228 27956 25280 28008
rect 23848 27931 23900 27940
rect 23848 27897 23857 27931
rect 23857 27897 23891 27931
rect 23891 27897 23900 27931
rect 23848 27888 23900 27897
rect 26884 27888 26936 27940
rect 28264 27956 28316 28008
rect 30564 28067 30616 28076
rect 30564 28033 30573 28067
rect 30573 28033 30607 28067
rect 30607 28033 30616 28067
rect 30564 28024 30616 28033
rect 32588 28092 32640 28144
rect 30012 27999 30064 28008
rect 30012 27965 30021 27999
rect 30021 27965 30055 27999
rect 30055 27965 30064 27999
rect 30012 27956 30064 27965
rect 27988 27888 28040 27940
rect 30472 27888 30524 27940
rect 25596 27863 25648 27872
rect 25596 27829 25605 27863
rect 25605 27829 25639 27863
rect 25639 27829 25648 27863
rect 25596 27820 25648 27829
rect 28724 27820 28776 27872
rect 29000 27820 29052 27872
rect 30748 27999 30800 28008
rect 30748 27965 30757 27999
rect 30757 27965 30791 27999
rect 30791 27965 30800 27999
rect 30748 27956 30800 27965
rect 31944 28067 31996 28076
rect 31944 28033 31953 28067
rect 31953 28033 31987 28067
rect 31987 28033 31996 28067
rect 31944 28024 31996 28033
rect 32864 28092 32916 28144
rect 39120 28160 39172 28212
rect 41788 28160 41840 28212
rect 33600 28092 33652 28144
rect 39212 28092 39264 28144
rect 40500 28092 40552 28144
rect 42616 28203 42668 28212
rect 42616 28169 42641 28203
rect 42641 28169 42668 28203
rect 42616 28160 42668 28169
rect 32128 27999 32180 28008
rect 32128 27965 32137 27999
rect 32137 27965 32171 27999
rect 32171 27965 32180 27999
rect 32128 27956 32180 27965
rect 38752 28024 38804 28076
rect 39948 28067 40000 28076
rect 39948 28033 39957 28067
rect 39957 28033 39991 28067
rect 39991 28033 40000 28067
rect 39948 28024 40000 28033
rect 40132 28024 40184 28076
rect 40224 28067 40276 28076
rect 40224 28033 40233 28067
rect 40233 28033 40267 28067
rect 40267 28033 40276 28067
rect 40224 28024 40276 28033
rect 41512 28067 41564 28076
rect 41512 28033 41521 28067
rect 41521 28033 41555 28067
rect 41555 28033 41564 28067
rect 41512 28024 41564 28033
rect 44916 28203 44968 28212
rect 44916 28169 44925 28203
rect 44925 28169 44959 28203
rect 44959 28169 44968 28203
rect 44916 28160 44968 28169
rect 46664 28203 46716 28212
rect 46664 28169 46673 28203
rect 46673 28169 46707 28203
rect 46707 28169 46716 28203
rect 46664 28160 46716 28169
rect 35440 27956 35492 28008
rect 38384 27999 38436 28008
rect 38384 27965 38393 27999
rect 38393 27965 38427 27999
rect 38427 27965 38436 27999
rect 38384 27956 38436 27965
rect 41328 27999 41380 28008
rect 41328 27965 41337 27999
rect 41337 27965 41371 27999
rect 41371 27965 41380 27999
rect 41328 27956 41380 27965
rect 34520 27888 34572 27940
rect 39764 27888 39816 27940
rect 33508 27820 33560 27872
rect 38200 27820 38252 27872
rect 38568 27820 38620 27872
rect 38660 27863 38712 27872
rect 38660 27829 38669 27863
rect 38669 27829 38703 27863
rect 38703 27829 38712 27863
rect 38660 27820 38712 27829
rect 40960 27820 41012 27872
rect 43536 28067 43588 28076
rect 43536 28033 43545 28067
rect 43545 28033 43579 28067
rect 43579 28033 43588 28067
rect 43536 28024 43588 28033
rect 41880 27999 41932 28008
rect 41880 27965 41889 27999
rect 41889 27965 41923 27999
rect 41923 27965 41932 27999
rect 41880 27956 41932 27965
rect 42432 27956 42484 28008
rect 43996 28092 44048 28144
rect 44088 28135 44140 28144
rect 44088 28101 44113 28135
rect 44113 28101 44140 28135
rect 44088 28092 44140 28101
rect 44548 28135 44600 28144
rect 44548 28101 44557 28135
rect 44557 28101 44591 28135
rect 44591 28101 44600 28135
rect 44548 28092 44600 28101
rect 44456 28024 44508 28076
rect 44640 28067 44692 28076
rect 44640 28033 44649 28067
rect 44649 28033 44683 28067
rect 44683 28033 44692 28067
rect 44640 28024 44692 28033
rect 46020 28092 46072 28144
rect 45192 28067 45244 28076
rect 45192 28033 45201 28067
rect 45201 28033 45235 28067
rect 45235 28033 45244 28067
rect 45192 28024 45244 28033
rect 46572 28067 46624 28076
rect 46572 28033 46581 28067
rect 46581 28033 46615 28067
rect 46615 28033 46624 28067
rect 46572 28024 46624 28033
rect 41972 27888 42024 27940
rect 42524 27888 42576 27940
rect 42892 27888 42944 27940
rect 43536 27888 43588 27940
rect 41788 27820 41840 27872
rect 42064 27820 42116 27872
rect 42616 27863 42668 27872
rect 42616 27829 42625 27863
rect 42625 27829 42659 27863
rect 42659 27829 42668 27863
rect 42616 27820 42668 27829
rect 42800 27863 42852 27872
rect 42800 27829 42809 27863
rect 42809 27829 42843 27863
rect 42843 27829 42852 27863
rect 42800 27820 42852 27829
rect 43996 27820 44048 27872
rect 45468 27863 45520 27872
rect 45468 27829 45477 27863
rect 45477 27829 45511 27863
rect 45511 27829 45520 27863
rect 45468 27820 45520 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2964 27616 3016 27668
rect 3148 27659 3200 27668
rect 3148 27625 3157 27659
rect 3157 27625 3191 27659
rect 3191 27625 3200 27659
rect 3148 27616 3200 27625
rect 4620 27616 4672 27668
rect 6460 27659 6512 27668
rect 6460 27625 6469 27659
rect 6469 27625 6503 27659
rect 6503 27625 6512 27659
rect 6460 27616 6512 27625
rect 10968 27616 11020 27668
rect 13820 27616 13872 27668
rect 16304 27616 16356 27668
rect 16580 27616 16632 27668
rect 17592 27659 17644 27668
rect 17592 27625 17601 27659
rect 17601 27625 17635 27659
rect 17635 27625 17644 27659
rect 17592 27616 17644 27625
rect 17684 27616 17736 27668
rect 22468 27616 22520 27668
rect 1676 27523 1728 27532
rect 1676 27489 1685 27523
rect 1685 27489 1719 27523
rect 1719 27489 1728 27523
rect 1676 27480 1728 27489
rect 3056 27480 3108 27532
rect 3608 27480 3660 27532
rect 8668 27548 8720 27600
rect 1952 27455 2004 27464
rect 1952 27421 1986 27455
rect 1986 27421 2004 27455
rect 1952 27412 2004 27421
rect 3976 27412 4028 27464
rect 7472 27480 7524 27532
rect 8024 27480 8076 27532
rect 5908 27412 5960 27464
rect 7012 27412 7064 27464
rect 9128 27480 9180 27532
rect 10140 27523 10192 27532
rect 10140 27489 10149 27523
rect 10149 27489 10183 27523
rect 10183 27489 10192 27523
rect 10140 27480 10192 27489
rect 10600 27480 10652 27532
rect 12624 27548 12676 27600
rect 13912 27548 13964 27600
rect 17040 27548 17092 27600
rect 18696 27548 18748 27600
rect 18972 27591 19024 27600
rect 18972 27557 18981 27591
rect 18981 27557 19015 27591
rect 19015 27557 19024 27591
rect 18972 27548 19024 27557
rect 19800 27548 19852 27600
rect 11980 27480 12032 27532
rect 14280 27480 14332 27532
rect 14648 27480 14700 27532
rect 15108 27480 15160 27532
rect 8208 27455 8260 27464
rect 8208 27421 8217 27455
rect 8217 27421 8251 27455
rect 8251 27421 8260 27455
rect 8208 27412 8260 27421
rect 8300 27344 8352 27396
rect 9312 27344 9364 27396
rect 11336 27344 11388 27396
rect 13268 27412 13320 27464
rect 12900 27344 12952 27396
rect 14648 27344 14700 27396
rect 4068 27276 4120 27328
rect 5908 27319 5960 27328
rect 5908 27285 5917 27319
rect 5917 27285 5951 27319
rect 5951 27285 5960 27319
rect 5908 27276 5960 27285
rect 7196 27276 7248 27328
rect 7932 27276 7984 27328
rect 9956 27276 10008 27328
rect 10048 27319 10100 27328
rect 10048 27285 10057 27319
rect 10057 27285 10091 27319
rect 10091 27285 10100 27319
rect 10048 27276 10100 27285
rect 10784 27276 10836 27328
rect 11796 27276 11848 27328
rect 12532 27276 12584 27328
rect 13268 27276 13320 27328
rect 15200 27412 15252 27464
rect 16948 27455 17000 27464
rect 16948 27421 16957 27455
rect 16957 27421 16991 27455
rect 16991 27421 17000 27455
rect 16948 27412 17000 27421
rect 17040 27455 17092 27464
rect 17040 27421 17049 27455
rect 17049 27421 17083 27455
rect 17083 27421 17092 27455
rect 17040 27412 17092 27421
rect 18420 27412 18472 27464
rect 18696 27412 18748 27464
rect 21548 27455 21600 27464
rect 21548 27421 21582 27455
rect 21582 27421 21600 27455
rect 16396 27344 16448 27396
rect 15844 27276 15896 27328
rect 16672 27276 16724 27328
rect 20352 27344 20404 27396
rect 21548 27412 21600 27421
rect 22100 27412 22152 27464
rect 23204 27616 23256 27668
rect 24032 27616 24084 27668
rect 28448 27659 28500 27668
rect 28448 27625 28457 27659
rect 28457 27625 28491 27659
rect 28491 27625 28500 27659
rect 28448 27616 28500 27625
rect 30012 27616 30064 27668
rect 30564 27616 30616 27668
rect 23388 27480 23440 27532
rect 22836 27412 22888 27464
rect 23112 27344 23164 27396
rect 23204 27387 23256 27396
rect 23204 27353 23213 27387
rect 23213 27353 23247 27387
rect 23247 27353 23256 27387
rect 23204 27344 23256 27353
rect 20168 27276 20220 27328
rect 22192 27276 22244 27328
rect 22468 27276 22520 27328
rect 22744 27276 22796 27328
rect 24032 27412 24084 27464
rect 24216 27412 24268 27464
rect 24768 27344 24820 27396
rect 26332 27480 26384 27532
rect 29644 27548 29696 27600
rect 27620 27412 27672 27464
rect 28540 27412 28592 27464
rect 28724 27455 28776 27464
rect 28724 27421 28733 27455
rect 28733 27421 28767 27455
rect 28767 27421 28776 27455
rect 28724 27412 28776 27421
rect 26516 27276 26568 27328
rect 26608 27319 26660 27328
rect 26608 27285 26617 27319
rect 26617 27285 26651 27319
rect 26651 27285 26660 27319
rect 26608 27276 26660 27285
rect 27988 27276 28040 27328
rect 29092 27480 29144 27532
rect 29920 27480 29972 27532
rect 30196 27523 30248 27532
rect 30196 27489 30205 27523
rect 30205 27489 30239 27523
rect 30239 27489 30248 27523
rect 30196 27480 30248 27489
rect 30932 27480 30984 27532
rect 31300 27480 31352 27532
rect 29552 27455 29604 27464
rect 29552 27421 29561 27455
rect 29561 27421 29595 27455
rect 29595 27421 29604 27455
rect 29552 27412 29604 27421
rect 30472 27455 30524 27464
rect 30472 27421 30481 27455
rect 30481 27421 30515 27455
rect 30515 27421 30524 27455
rect 30472 27412 30524 27421
rect 32680 27523 32732 27532
rect 32680 27489 32689 27523
rect 32689 27489 32723 27523
rect 32723 27489 32732 27523
rect 32680 27480 32732 27489
rect 33232 27480 33284 27532
rect 34520 27591 34572 27600
rect 34520 27557 34529 27591
rect 34529 27557 34563 27591
rect 34563 27557 34572 27591
rect 34520 27548 34572 27557
rect 34060 27480 34112 27532
rect 36636 27616 36688 27668
rect 37648 27659 37700 27668
rect 37648 27625 37657 27659
rect 37657 27625 37691 27659
rect 37691 27625 37700 27659
rect 37648 27616 37700 27625
rect 32864 27455 32916 27464
rect 32864 27421 32873 27455
rect 32873 27421 32907 27455
rect 32907 27421 32916 27455
rect 32864 27412 32916 27421
rect 33600 27455 33652 27464
rect 33600 27421 33609 27455
rect 33609 27421 33643 27455
rect 33643 27421 33652 27455
rect 33600 27412 33652 27421
rect 33876 27455 33928 27464
rect 33876 27421 33885 27455
rect 33885 27421 33919 27455
rect 33919 27421 33928 27455
rect 33876 27412 33928 27421
rect 35164 27455 35216 27464
rect 35164 27421 35173 27455
rect 35173 27421 35207 27455
rect 35207 27421 35216 27455
rect 35164 27412 35216 27421
rect 36084 27412 36136 27464
rect 37096 27548 37148 27600
rect 29184 27344 29236 27396
rect 31576 27344 31628 27396
rect 29920 27276 29972 27328
rect 30472 27276 30524 27328
rect 31852 27319 31904 27328
rect 31852 27285 31861 27319
rect 31861 27285 31895 27319
rect 31895 27285 31904 27319
rect 31852 27276 31904 27285
rect 35624 27344 35676 27396
rect 36912 27387 36964 27396
rect 36912 27353 36921 27387
rect 36921 27353 36955 27387
rect 36955 27353 36964 27387
rect 36912 27344 36964 27353
rect 36636 27319 36688 27328
rect 36636 27285 36645 27319
rect 36645 27285 36679 27319
rect 36679 27285 36688 27319
rect 36636 27276 36688 27285
rect 37464 27480 37516 27532
rect 37096 27412 37148 27464
rect 38200 27616 38252 27668
rect 38660 27616 38712 27668
rect 41788 27616 41840 27668
rect 45652 27616 45704 27668
rect 39120 27548 39172 27600
rect 39212 27548 39264 27600
rect 41420 27548 41472 27600
rect 46112 27548 46164 27600
rect 46204 27591 46256 27600
rect 46204 27557 46213 27591
rect 46213 27557 46247 27591
rect 46247 27557 46256 27591
rect 46204 27548 46256 27557
rect 41788 27480 41840 27532
rect 38292 27276 38344 27328
rect 38568 27344 38620 27396
rect 39120 27412 39172 27464
rect 39396 27344 39448 27396
rect 39948 27344 40000 27396
rect 40316 27412 40368 27464
rect 40040 27276 40092 27328
rect 40776 27344 40828 27396
rect 41052 27344 41104 27396
rect 41144 27387 41196 27396
rect 41144 27353 41153 27387
rect 41153 27353 41187 27387
rect 41187 27353 41196 27387
rect 41144 27344 41196 27353
rect 41512 27412 41564 27464
rect 41972 27480 42024 27532
rect 42800 27480 42852 27532
rect 45468 27523 45520 27532
rect 45468 27489 45477 27523
rect 45477 27489 45511 27523
rect 45511 27489 45520 27523
rect 45468 27480 45520 27489
rect 42248 27412 42300 27464
rect 45652 27455 45704 27464
rect 45652 27421 45661 27455
rect 45661 27421 45695 27455
rect 45695 27421 45704 27455
rect 45652 27412 45704 27421
rect 46204 27412 46256 27464
rect 40684 27276 40736 27328
rect 41972 27344 42024 27396
rect 41880 27276 41932 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 2872 27072 2924 27124
rect 4068 27072 4120 27124
rect 8392 27047 8444 27056
rect 2504 26936 2556 26988
rect 4620 26936 4672 26988
rect 6828 26979 6880 26988
rect 6828 26945 6862 26979
rect 6862 26945 6880 26979
rect 6828 26936 6880 26945
rect 8392 27013 8426 27047
rect 8426 27013 8444 27047
rect 8392 27004 8444 27013
rect 9864 27004 9916 27056
rect 10048 27004 10100 27056
rect 9680 26979 9732 26988
rect 9680 26945 9689 26979
rect 9689 26945 9723 26979
rect 9723 26945 9732 26979
rect 9680 26936 9732 26945
rect 9956 26936 10008 26988
rect 10784 26979 10836 26988
rect 10784 26945 10793 26979
rect 10793 26945 10827 26979
rect 10827 26945 10836 26979
rect 10784 26936 10836 26945
rect 2964 26800 3016 26852
rect 5080 26800 5132 26852
rect 940 26732 992 26784
rect 3976 26732 4028 26784
rect 9128 26868 9180 26920
rect 11796 27115 11848 27124
rect 11796 27081 11805 27115
rect 11805 27081 11839 27115
rect 11839 27081 11848 27115
rect 11796 27072 11848 27081
rect 11980 27115 12032 27124
rect 11980 27081 11989 27115
rect 11989 27081 12023 27115
rect 12023 27081 12032 27115
rect 11980 27072 12032 27081
rect 12900 27115 12952 27124
rect 12900 27081 12909 27115
rect 12909 27081 12943 27115
rect 12943 27081 12952 27115
rect 12900 27072 12952 27081
rect 13452 27072 13504 27124
rect 14556 27072 14608 27124
rect 14740 27072 14792 27124
rect 16764 27072 16816 27124
rect 12256 26936 12308 26988
rect 12532 27047 12584 27056
rect 12532 27013 12541 27047
rect 12541 27013 12575 27047
rect 12575 27013 12584 27047
rect 12532 27004 12584 27013
rect 12716 27047 12768 27056
rect 12716 27013 12725 27047
rect 12725 27013 12759 27047
rect 12759 27013 12768 27047
rect 12716 27004 12768 27013
rect 13452 26979 13504 26988
rect 13452 26945 13461 26979
rect 13461 26945 13495 26979
rect 13495 26945 13504 26979
rect 13452 26936 13504 26945
rect 13636 26979 13688 26988
rect 13636 26945 13645 26979
rect 13645 26945 13679 26979
rect 13679 26945 13688 26979
rect 13636 26936 13688 26945
rect 15384 27004 15436 27056
rect 16580 27004 16632 27056
rect 18420 27072 18472 27124
rect 19064 27115 19116 27124
rect 19064 27081 19073 27115
rect 19073 27081 19107 27115
rect 19107 27081 19116 27115
rect 19064 27072 19116 27081
rect 21272 27072 21324 27124
rect 16948 27004 17000 27056
rect 18236 27047 18288 27056
rect 18236 27013 18245 27047
rect 18245 27013 18279 27047
rect 18279 27013 18288 27047
rect 18236 27004 18288 27013
rect 18788 27047 18840 27056
rect 18788 27013 18797 27047
rect 18797 27013 18831 27047
rect 18831 27013 18840 27047
rect 18788 27004 18840 27013
rect 22468 27004 22520 27056
rect 25320 27004 25372 27056
rect 14464 26936 14516 26988
rect 14740 26936 14792 26988
rect 7932 26843 7984 26852
rect 7932 26809 7941 26843
rect 7941 26809 7975 26843
rect 7975 26809 7984 26843
rect 7932 26800 7984 26809
rect 10968 26800 11020 26852
rect 11796 26868 11848 26920
rect 12348 26911 12400 26920
rect 12348 26877 12357 26911
rect 12357 26877 12391 26911
rect 12391 26877 12400 26911
rect 12348 26868 12400 26877
rect 12900 26868 12952 26920
rect 13820 26868 13872 26920
rect 15200 26868 15252 26920
rect 16396 26936 16448 26988
rect 17224 26979 17276 26988
rect 17224 26945 17233 26979
rect 17233 26945 17267 26979
rect 17267 26945 17276 26979
rect 17224 26936 17276 26945
rect 17408 26979 17460 26988
rect 17408 26945 17417 26979
rect 17417 26945 17451 26979
rect 17451 26945 17460 26979
rect 17408 26936 17460 26945
rect 16764 26911 16816 26920
rect 16764 26877 16773 26911
rect 16773 26877 16807 26911
rect 16807 26877 16816 26911
rect 16764 26868 16816 26877
rect 16948 26868 17000 26920
rect 18604 26936 18656 26988
rect 21364 26936 21416 26988
rect 21456 26979 21508 26988
rect 21456 26945 21465 26979
rect 21465 26945 21499 26979
rect 21499 26945 21508 26979
rect 21456 26936 21508 26945
rect 21732 26936 21784 26988
rect 22192 26979 22244 26988
rect 22192 26945 22201 26979
rect 22201 26945 22235 26979
rect 22235 26945 22244 26979
rect 22192 26936 22244 26945
rect 20996 26868 21048 26920
rect 21088 26868 21140 26920
rect 22376 26911 22428 26920
rect 22376 26877 22385 26911
rect 22385 26877 22419 26911
rect 22419 26877 22428 26911
rect 22376 26868 22428 26877
rect 9772 26732 9824 26784
rect 10048 26775 10100 26784
rect 10048 26741 10057 26775
rect 10057 26741 10091 26775
rect 10091 26741 10100 26775
rect 10048 26732 10100 26741
rect 10784 26732 10836 26784
rect 12256 26800 12308 26852
rect 22468 26800 22520 26852
rect 13636 26732 13688 26784
rect 14280 26732 14332 26784
rect 16028 26732 16080 26784
rect 19708 26732 19760 26784
rect 20812 26732 20864 26784
rect 20996 26732 21048 26784
rect 23296 26936 23348 26988
rect 24032 26936 24084 26988
rect 25044 26936 25096 26988
rect 26608 27072 26660 27124
rect 26516 27004 26568 27056
rect 22928 26911 22980 26920
rect 22928 26877 22937 26911
rect 22937 26877 22971 26911
rect 22971 26877 22980 26911
rect 22928 26868 22980 26877
rect 23848 26911 23900 26920
rect 23848 26877 23857 26911
rect 23857 26877 23891 26911
rect 23891 26877 23900 26911
rect 23848 26868 23900 26877
rect 24124 26911 24176 26920
rect 24124 26877 24133 26911
rect 24133 26877 24167 26911
rect 24167 26877 24176 26911
rect 24124 26868 24176 26877
rect 23572 26843 23624 26852
rect 23572 26809 23581 26843
rect 23581 26809 23615 26843
rect 23615 26809 23624 26843
rect 23572 26800 23624 26809
rect 25964 26979 26016 26988
rect 25964 26945 25973 26979
rect 25973 26945 26007 26979
rect 26007 26945 26016 26979
rect 25964 26936 26016 26945
rect 26884 26936 26936 26988
rect 27620 26936 27672 26988
rect 25596 26868 25648 26920
rect 29276 27072 29328 27124
rect 29736 27072 29788 27124
rect 30196 27072 30248 27124
rect 32864 27072 32916 27124
rect 29092 26979 29144 26988
rect 29092 26945 29101 26979
rect 29101 26945 29135 26979
rect 29135 26945 29144 26979
rect 29092 26936 29144 26945
rect 29828 26979 29880 26988
rect 29828 26945 29837 26979
rect 29837 26945 29871 26979
rect 29871 26945 29880 26979
rect 29828 26936 29880 26945
rect 31852 26936 31904 26988
rect 32680 26936 32732 26988
rect 35164 27072 35216 27124
rect 36636 27072 36688 27124
rect 38384 27072 38436 27124
rect 38752 27115 38804 27124
rect 38752 27081 38761 27115
rect 38761 27081 38795 27115
rect 38795 27081 38804 27115
rect 38752 27072 38804 27081
rect 34060 26979 34112 26988
rect 34060 26945 34094 26979
rect 34094 26945 34112 26979
rect 34060 26936 34112 26945
rect 35440 26936 35492 26988
rect 36360 26979 36412 26988
rect 36360 26945 36369 26979
rect 36369 26945 36403 26979
rect 36403 26945 36412 26979
rect 36360 26936 36412 26945
rect 36912 27004 36964 27056
rect 41144 27072 41196 27124
rect 37372 26936 37424 26988
rect 38108 26936 38160 26988
rect 38292 26979 38344 26988
rect 38292 26945 38301 26979
rect 38301 26945 38335 26979
rect 38335 26945 38344 26979
rect 38292 26936 38344 26945
rect 40684 27004 40736 27056
rect 39396 26979 39448 26988
rect 39396 26945 39405 26979
rect 39405 26945 39439 26979
rect 39439 26945 39448 26979
rect 39396 26936 39448 26945
rect 39764 26979 39816 26988
rect 39764 26945 39773 26979
rect 39773 26945 39807 26979
rect 39807 26945 39816 26979
rect 39764 26936 39816 26945
rect 39948 26936 40000 26988
rect 42064 27072 42116 27124
rect 45652 27072 45704 27124
rect 41788 27004 41840 27056
rect 42432 27004 42484 27056
rect 42248 26936 42300 26988
rect 42616 26979 42668 26988
rect 42616 26945 42625 26979
rect 42625 26945 42659 26979
rect 42659 26945 42668 26979
rect 42616 26936 42668 26945
rect 43352 27004 43404 27056
rect 29644 26868 29696 26920
rect 30840 26868 30892 26920
rect 33600 26868 33652 26920
rect 34244 26911 34296 26920
rect 34244 26877 34253 26911
rect 34253 26877 34287 26911
rect 34287 26877 34296 26911
rect 34244 26868 34296 26877
rect 35348 26868 35400 26920
rect 38568 26868 38620 26920
rect 41604 26868 41656 26920
rect 42432 26868 42484 26920
rect 42984 26911 43036 26920
rect 42984 26877 42993 26911
rect 42993 26877 43027 26911
rect 43027 26877 43036 26911
rect 43260 26979 43312 26988
rect 43260 26945 43269 26979
rect 43269 26945 43303 26979
rect 43303 26945 43312 26979
rect 43260 26936 43312 26945
rect 45560 26979 45612 26988
rect 45560 26945 45569 26979
rect 45569 26945 45603 26979
rect 45603 26945 45612 26979
rect 45560 26936 45612 26945
rect 45744 26936 45796 26988
rect 46756 26936 46808 26988
rect 42984 26868 43036 26877
rect 24032 26732 24084 26784
rect 24308 26732 24360 26784
rect 24768 26775 24820 26784
rect 24768 26741 24777 26775
rect 24777 26741 24811 26775
rect 24811 26741 24820 26775
rect 24768 26732 24820 26741
rect 25228 26775 25280 26784
rect 25228 26741 25237 26775
rect 25237 26741 25271 26775
rect 25271 26741 25280 26775
rect 25228 26732 25280 26741
rect 29460 26800 29512 26852
rect 29000 26732 29052 26784
rect 33692 26843 33744 26852
rect 33692 26809 33701 26843
rect 33701 26809 33735 26843
rect 33735 26809 33744 26843
rect 33692 26800 33744 26809
rect 40316 26800 40368 26852
rect 41880 26843 41932 26852
rect 41880 26809 41889 26843
rect 41889 26809 41923 26843
rect 41923 26809 41932 26843
rect 41880 26800 41932 26809
rect 42064 26800 42116 26852
rect 46020 26843 46072 26852
rect 46020 26809 46029 26843
rect 46029 26809 46063 26843
rect 46063 26809 46072 26843
rect 46020 26800 46072 26809
rect 30288 26732 30340 26784
rect 30564 26732 30616 26784
rect 32036 26732 32088 26784
rect 33324 26732 33376 26784
rect 37096 26775 37148 26784
rect 37096 26741 37105 26775
rect 37105 26741 37139 26775
rect 37139 26741 37148 26775
rect 37096 26732 37148 26741
rect 38752 26732 38804 26784
rect 39120 26732 39172 26784
rect 41236 26732 41288 26784
rect 44640 26732 44692 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2780 26528 2832 26580
rect 4528 26528 4580 26580
rect 4068 26435 4120 26444
rect 4068 26401 4077 26435
rect 4077 26401 4111 26435
rect 4111 26401 4120 26435
rect 4068 26392 4120 26401
rect 4620 26392 4672 26444
rect 4712 26435 4764 26444
rect 4712 26401 4721 26435
rect 4721 26401 4755 26435
rect 4755 26401 4764 26435
rect 4712 26392 4764 26401
rect 5632 26528 5684 26580
rect 6092 26528 6144 26580
rect 6276 26528 6328 26580
rect 6828 26528 6880 26580
rect 5724 26460 5776 26512
rect 8576 26460 8628 26512
rect 5080 26435 5132 26444
rect 5080 26401 5114 26435
rect 5114 26401 5132 26435
rect 5080 26392 5132 26401
rect 1676 26324 1728 26376
rect 3976 26367 4028 26376
rect 3976 26333 3985 26367
rect 3985 26333 4019 26367
rect 4019 26333 4028 26367
rect 3976 26324 4028 26333
rect 4252 26367 4304 26376
rect 4252 26333 4261 26367
rect 4261 26333 4295 26367
rect 4295 26333 4304 26367
rect 4252 26324 4304 26333
rect 6184 26367 6236 26376
rect 6184 26333 6193 26367
rect 6193 26333 6227 26367
rect 6227 26333 6236 26367
rect 6184 26324 6236 26333
rect 7196 26367 7248 26376
rect 7196 26333 7205 26367
rect 7205 26333 7239 26367
rect 7239 26333 7248 26367
rect 7196 26324 7248 26333
rect 2044 26256 2096 26308
rect 6828 26256 6880 26308
rect 7932 26392 7984 26444
rect 9864 26528 9916 26580
rect 12992 26571 13044 26580
rect 12992 26537 13001 26571
rect 13001 26537 13035 26571
rect 13035 26537 13044 26571
rect 12992 26528 13044 26537
rect 8024 26324 8076 26376
rect 12348 26392 12400 26444
rect 10048 26324 10100 26376
rect 10784 26324 10836 26376
rect 3884 26188 3936 26240
rect 4620 26188 4672 26240
rect 4988 26188 5040 26240
rect 8300 26256 8352 26308
rect 10416 26256 10468 26308
rect 12532 26324 12584 26376
rect 12716 26324 12768 26376
rect 13820 26503 13872 26512
rect 13820 26469 13829 26503
rect 13829 26469 13863 26503
rect 13863 26469 13872 26503
rect 13820 26460 13872 26469
rect 14556 26528 14608 26580
rect 15108 26528 15160 26580
rect 25228 26528 25280 26580
rect 15200 26460 15252 26512
rect 15476 26460 15528 26512
rect 13544 26324 13596 26376
rect 10600 26231 10652 26240
rect 10600 26197 10609 26231
rect 10609 26197 10643 26231
rect 10643 26197 10652 26231
rect 12900 26256 12952 26308
rect 13636 26299 13688 26308
rect 13636 26265 13645 26299
rect 13645 26265 13679 26299
rect 13679 26265 13688 26299
rect 15752 26435 15804 26444
rect 15752 26401 15761 26435
rect 15761 26401 15795 26435
rect 15795 26401 15804 26435
rect 15752 26392 15804 26401
rect 16120 26392 16172 26444
rect 17040 26460 17092 26512
rect 20352 26503 20404 26512
rect 20352 26469 20361 26503
rect 20361 26469 20395 26503
rect 20395 26469 20404 26503
rect 20352 26460 20404 26469
rect 20812 26503 20864 26512
rect 20812 26469 20821 26503
rect 20821 26469 20855 26503
rect 20855 26469 20864 26503
rect 20812 26460 20864 26469
rect 16764 26392 16816 26444
rect 14648 26324 14700 26376
rect 14740 26324 14792 26376
rect 13636 26256 13688 26265
rect 10600 26188 10652 26197
rect 12256 26188 12308 26240
rect 13268 26188 13320 26240
rect 13912 26188 13964 26240
rect 16212 26324 16264 26376
rect 17040 26367 17092 26376
rect 17040 26333 17049 26367
rect 17049 26333 17083 26367
rect 17083 26333 17092 26367
rect 17040 26324 17092 26333
rect 17408 26392 17460 26444
rect 20536 26392 20588 26444
rect 18604 26367 18656 26376
rect 18604 26333 18613 26367
rect 18613 26333 18647 26367
rect 18647 26333 18656 26367
rect 18604 26324 18656 26333
rect 20628 26367 20680 26376
rect 20628 26333 20637 26367
rect 20637 26333 20671 26367
rect 20671 26333 20680 26367
rect 20628 26324 20680 26333
rect 21180 26324 21232 26376
rect 16028 26256 16080 26308
rect 16856 26256 16908 26308
rect 17592 26299 17644 26308
rect 17592 26265 17601 26299
rect 17601 26265 17635 26299
rect 17635 26265 17644 26299
rect 17592 26256 17644 26265
rect 19616 26256 19668 26308
rect 19984 26256 20036 26308
rect 24768 26460 24820 26512
rect 26332 26460 26384 26512
rect 34060 26528 34112 26580
rect 35348 26528 35400 26580
rect 37648 26528 37700 26580
rect 42616 26528 42668 26580
rect 43168 26528 43220 26580
rect 46020 26571 46072 26580
rect 46020 26537 46029 26571
rect 46029 26537 46063 26571
rect 46063 26537 46072 26571
rect 46020 26528 46072 26537
rect 46204 26571 46256 26580
rect 46204 26537 46213 26571
rect 46213 26537 46247 26571
rect 46247 26537 46256 26571
rect 46204 26528 46256 26537
rect 23480 26392 23532 26444
rect 36360 26460 36412 26512
rect 38384 26460 38436 26512
rect 40960 26460 41012 26512
rect 42800 26460 42852 26512
rect 46756 26571 46808 26580
rect 46756 26537 46765 26571
rect 46765 26537 46799 26571
rect 46799 26537 46808 26571
rect 46756 26528 46808 26537
rect 31576 26392 31628 26444
rect 38568 26392 38620 26444
rect 22928 26256 22980 26308
rect 23940 26324 23992 26376
rect 26056 26324 26108 26376
rect 26148 26324 26200 26376
rect 28540 26324 28592 26376
rect 30564 26367 30616 26376
rect 30564 26333 30573 26367
rect 30573 26333 30607 26367
rect 30607 26333 30616 26367
rect 30564 26324 30616 26333
rect 31852 26324 31904 26376
rect 32036 26367 32088 26376
rect 32036 26333 32070 26367
rect 32070 26333 32088 26367
rect 32036 26324 32088 26333
rect 32772 26324 32824 26376
rect 33968 26324 34020 26376
rect 34152 26324 34204 26376
rect 37372 26324 37424 26376
rect 38200 26367 38252 26376
rect 38200 26333 38209 26367
rect 38209 26333 38243 26367
rect 38243 26333 38252 26367
rect 42616 26392 42668 26444
rect 38200 26324 38252 26333
rect 41696 26324 41748 26376
rect 41972 26367 42024 26376
rect 41972 26333 41981 26367
rect 41981 26333 42015 26367
rect 42015 26333 42024 26367
rect 41972 26324 42024 26333
rect 42248 26367 42300 26376
rect 42248 26333 42257 26367
rect 42257 26333 42291 26367
rect 42291 26333 42300 26367
rect 42248 26324 42300 26333
rect 42432 26324 42484 26376
rect 17040 26188 17092 26240
rect 17224 26188 17276 26240
rect 23756 26188 23808 26240
rect 26240 26299 26292 26308
rect 26240 26265 26249 26299
rect 26249 26265 26283 26299
rect 26283 26265 26292 26299
rect 26240 26256 26292 26265
rect 33324 26256 33376 26308
rect 37096 26256 37148 26308
rect 43260 26392 43312 26444
rect 42984 26367 43036 26376
rect 42984 26333 42993 26367
rect 42993 26333 43027 26367
rect 43027 26333 43036 26367
rect 42984 26324 43036 26333
rect 43168 26367 43220 26376
rect 43168 26333 43177 26367
rect 43177 26333 43211 26367
rect 43211 26333 43220 26367
rect 43168 26324 43220 26333
rect 43352 26367 43404 26376
rect 43352 26333 43361 26367
rect 43361 26333 43395 26367
rect 43395 26333 43404 26367
rect 43352 26324 43404 26333
rect 45744 26367 45796 26376
rect 45744 26333 45753 26367
rect 45753 26333 45787 26367
rect 45787 26333 45796 26367
rect 45744 26324 45796 26333
rect 26056 26188 26108 26240
rect 39120 26188 39172 26240
rect 39672 26188 39724 26240
rect 43996 26256 44048 26308
rect 43260 26188 43312 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 2044 26027 2096 26036
rect 2044 25993 2053 26027
rect 2053 25993 2087 26027
rect 2087 25993 2096 26027
rect 2044 25984 2096 25993
rect 2780 26027 2832 26036
rect 2780 25993 2789 26027
rect 2789 25993 2823 26027
rect 2823 25993 2832 26027
rect 2780 25984 2832 25993
rect 2872 26027 2924 26036
rect 2872 25993 2881 26027
rect 2881 25993 2915 26027
rect 2915 25993 2924 26027
rect 2872 25984 2924 25993
rect 6276 25984 6328 26036
rect 12532 25984 12584 26036
rect 14832 25984 14884 26036
rect 15752 25984 15804 26036
rect 22008 25984 22060 26036
rect 23112 25984 23164 26036
rect 25872 25984 25924 26036
rect 29460 25984 29512 26036
rect 9864 25916 9916 25968
rect 4068 25848 4120 25900
rect 4896 25891 4948 25900
rect 4896 25857 4905 25891
rect 4905 25857 4939 25891
rect 4939 25857 4948 25891
rect 4896 25848 4948 25857
rect 5080 25848 5132 25900
rect 7656 25848 7708 25900
rect 8576 25891 8628 25900
rect 8576 25857 8585 25891
rect 8585 25857 8619 25891
rect 8619 25857 8628 25891
rect 8576 25848 8628 25857
rect 9404 25848 9456 25900
rect 13268 25916 13320 25968
rect 13452 25916 13504 25968
rect 10600 25848 10652 25900
rect 14740 25916 14792 25968
rect 16304 25916 16356 25968
rect 17592 25916 17644 25968
rect 4252 25780 4304 25832
rect 5356 25780 5408 25832
rect 7472 25823 7524 25832
rect 7472 25789 7481 25823
rect 7481 25789 7515 25823
rect 7515 25789 7524 25823
rect 7472 25780 7524 25789
rect 8024 25780 8076 25832
rect 9128 25780 9180 25832
rect 9772 25780 9824 25832
rect 4712 25712 4764 25764
rect 6184 25712 6236 25764
rect 6460 25712 6512 25764
rect 14280 25891 14332 25900
rect 14280 25857 14289 25891
rect 14289 25857 14323 25891
rect 14323 25857 14332 25891
rect 14280 25848 14332 25857
rect 14372 25891 14424 25900
rect 14372 25857 14381 25891
rect 14381 25857 14415 25891
rect 14415 25857 14424 25891
rect 14372 25848 14424 25857
rect 15476 25891 15528 25900
rect 15476 25857 15485 25891
rect 15485 25857 15519 25891
rect 15519 25857 15528 25891
rect 15476 25848 15528 25857
rect 20720 25916 20772 25968
rect 20812 25916 20864 25968
rect 34152 25916 34204 25968
rect 41144 25916 41196 25968
rect 11796 25823 11848 25832
rect 11796 25789 11805 25823
rect 11805 25789 11839 25823
rect 11839 25789 11848 25823
rect 11796 25780 11848 25789
rect 12624 25780 12676 25832
rect 12992 25780 13044 25832
rect 14096 25780 14148 25832
rect 23020 25848 23072 25900
rect 23296 25891 23348 25900
rect 23296 25857 23305 25891
rect 23305 25857 23339 25891
rect 23339 25857 23348 25891
rect 23296 25848 23348 25857
rect 23388 25891 23440 25900
rect 23388 25857 23397 25891
rect 23397 25857 23431 25891
rect 23431 25857 23440 25891
rect 23388 25848 23440 25857
rect 22008 25780 22060 25832
rect 22836 25780 22888 25832
rect 5172 25644 5224 25696
rect 6828 25644 6880 25696
rect 8392 25687 8444 25696
rect 8392 25653 8401 25687
rect 8401 25653 8435 25687
rect 8435 25653 8444 25687
rect 8392 25644 8444 25653
rect 10968 25644 11020 25696
rect 17316 25712 17368 25764
rect 23756 25780 23808 25832
rect 25688 25848 25740 25900
rect 25964 25891 26016 25900
rect 25964 25857 25973 25891
rect 25973 25857 26007 25891
rect 26007 25857 26016 25891
rect 25964 25848 26016 25857
rect 33048 25848 33100 25900
rect 36544 25891 36596 25900
rect 36544 25857 36553 25891
rect 36553 25857 36587 25891
rect 36587 25857 36596 25891
rect 36544 25848 36596 25857
rect 37004 25848 37056 25900
rect 37924 25848 37976 25900
rect 39672 25891 39724 25900
rect 39672 25857 39681 25891
rect 39681 25857 39715 25891
rect 39715 25857 39724 25891
rect 39672 25848 39724 25857
rect 42892 25984 42944 26036
rect 44088 25984 44140 26036
rect 45560 25984 45612 26036
rect 43996 25916 44048 25968
rect 42524 25848 42576 25900
rect 43260 25891 43312 25900
rect 43260 25857 43269 25891
rect 43269 25857 43303 25891
rect 43303 25857 43312 25891
rect 43260 25848 43312 25857
rect 30564 25780 30616 25832
rect 33508 25823 33560 25832
rect 33508 25789 33517 25823
rect 33517 25789 33551 25823
rect 33551 25789 33560 25823
rect 33508 25780 33560 25789
rect 34428 25780 34480 25832
rect 34704 25780 34756 25832
rect 42064 25780 42116 25832
rect 42616 25780 42668 25832
rect 42800 25823 42852 25832
rect 42800 25789 42809 25823
rect 42809 25789 42843 25823
rect 42843 25789 42852 25823
rect 42800 25780 42852 25789
rect 43168 25823 43220 25832
rect 43168 25789 43177 25823
rect 43177 25789 43211 25823
rect 43211 25789 43220 25823
rect 43168 25780 43220 25789
rect 36084 25712 36136 25764
rect 13544 25687 13596 25696
rect 13544 25653 13553 25687
rect 13553 25653 13587 25687
rect 13587 25653 13596 25687
rect 13544 25644 13596 25653
rect 14188 25644 14240 25696
rect 17500 25644 17552 25696
rect 18052 25644 18104 25696
rect 19800 25644 19852 25696
rect 23388 25644 23440 25696
rect 31116 25644 31168 25696
rect 33600 25644 33652 25696
rect 36176 25644 36228 25696
rect 40316 25644 40368 25696
rect 42524 25687 42576 25696
rect 42524 25653 42533 25687
rect 42533 25653 42567 25687
rect 42567 25653 42576 25687
rect 42524 25644 42576 25653
rect 43260 25644 43312 25696
rect 43904 25644 43956 25696
rect 44088 25712 44140 25764
rect 45744 25891 45796 25900
rect 45744 25857 45753 25891
rect 45753 25857 45787 25891
rect 45787 25857 45796 25891
rect 45744 25848 45796 25857
rect 46204 25848 46256 25900
rect 45284 25644 45336 25696
rect 46020 25687 46072 25696
rect 46020 25653 46029 25687
rect 46029 25653 46063 25687
rect 46063 25653 46072 25687
rect 46020 25644 46072 25653
rect 46296 25644 46348 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 5172 25483 5224 25492
rect 5172 25449 5181 25483
rect 5181 25449 5215 25483
rect 5215 25449 5224 25483
rect 5172 25440 5224 25449
rect 7472 25304 7524 25356
rect 8024 25304 8076 25356
rect 1676 25236 1728 25288
rect 3884 25236 3936 25288
rect 6828 25279 6880 25288
rect 6828 25245 6837 25279
rect 6837 25245 6871 25279
rect 6871 25245 6880 25279
rect 6828 25236 6880 25245
rect 7656 25279 7708 25288
rect 7656 25245 7665 25279
rect 7665 25245 7699 25279
rect 7699 25245 7708 25279
rect 13084 25440 13136 25492
rect 14372 25440 14424 25492
rect 12716 25415 12768 25424
rect 12716 25381 12725 25415
rect 12725 25381 12759 25415
rect 12759 25381 12768 25415
rect 12716 25372 12768 25381
rect 9772 25304 9824 25356
rect 9864 25304 9916 25356
rect 12808 25304 12860 25356
rect 18696 25440 18748 25492
rect 28908 25440 28960 25492
rect 16212 25372 16264 25424
rect 17316 25372 17368 25424
rect 17500 25372 17552 25424
rect 7656 25236 7708 25245
rect 9404 25279 9456 25288
rect 9404 25245 9413 25279
rect 9413 25245 9447 25279
rect 9447 25245 9456 25279
rect 9404 25236 9456 25245
rect 12164 25236 12216 25288
rect 12624 25236 12676 25288
rect 14096 25279 14148 25288
rect 14096 25245 14105 25279
rect 14105 25245 14139 25279
rect 14139 25245 14148 25279
rect 14096 25236 14148 25245
rect 2780 25168 2832 25220
rect 8944 25168 8996 25220
rect 3240 25143 3292 25152
rect 3240 25109 3249 25143
rect 3249 25109 3283 25143
rect 3283 25109 3292 25143
rect 3240 25100 3292 25109
rect 6552 25100 6604 25152
rect 7288 25143 7340 25152
rect 7288 25109 7297 25143
rect 7297 25109 7331 25143
rect 7331 25109 7340 25143
rect 7288 25100 7340 25109
rect 12072 25143 12124 25152
rect 12072 25109 12081 25143
rect 12081 25109 12115 25143
rect 12115 25109 12124 25143
rect 12072 25100 12124 25109
rect 16764 25347 16816 25356
rect 16304 25279 16356 25288
rect 16304 25245 16313 25279
rect 16313 25245 16347 25279
rect 16347 25245 16356 25279
rect 16304 25236 16356 25245
rect 16764 25313 16773 25347
rect 16773 25313 16807 25347
rect 16807 25313 16816 25347
rect 16764 25304 16816 25313
rect 20812 25304 20864 25356
rect 21272 25347 21324 25356
rect 21272 25313 21281 25347
rect 21281 25313 21315 25347
rect 21315 25313 21324 25347
rect 21272 25304 21324 25313
rect 17040 25236 17092 25288
rect 17316 25279 17368 25288
rect 17316 25245 17325 25279
rect 17325 25245 17359 25279
rect 17359 25245 17368 25279
rect 17316 25236 17368 25245
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 18052 25279 18104 25288
rect 18052 25245 18061 25279
rect 18061 25245 18095 25279
rect 18095 25245 18104 25279
rect 18052 25236 18104 25245
rect 18236 25236 18288 25288
rect 21548 25415 21600 25424
rect 21548 25381 21557 25415
rect 21557 25381 21591 25415
rect 21591 25381 21600 25415
rect 21548 25372 21600 25381
rect 24124 25415 24176 25424
rect 24124 25381 24133 25415
rect 24133 25381 24167 25415
rect 24167 25381 24176 25415
rect 24124 25372 24176 25381
rect 30656 25372 30708 25424
rect 33876 25440 33928 25492
rect 38384 25440 38436 25492
rect 36268 25347 36320 25356
rect 22100 25236 22152 25288
rect 23112 25279 23164 25288
rect 23112 25245 23121 25279
rect 23121 25245 23155 25279
rect 23155 25245 23164 25279
rect 23112 25236 23164 25245
rect 23388 25279 23440 25288
rect 23388 25245 23397 25279
rect 23397 25245 23431 25279
rect 23431 25245 23440 25279
rect 23388 25236 23440 25245
rect 26240 25236 26292 25288
rect 29920 25236 29972 25288
rect 30840 25236 30892 25288
rect 31024 25279 31076 25288
rect 31024 25245 31033 25279
rect 31033 25245 31067 25279
rect 31067 25245 31076 25279
rect 31024 25236 31076 25245
rect 31760 25236 31812 25288
rect 33048 25236 33100 25288
rect 36268 25313 36277 25347
rect 36277 25313 36311 25347
rect 36311 25313 36320 25347
rect 36268 25304 36320 25313
rect 37280 25347 37332 25356
rect 37280 25313 37289 25347
rect 37289 25313 37323 25347
rect 37323 25313 37332 25347
rect 37280 25304 37332 25313
rect 38844 25372 38896 25424
rect 45284 25415 45336 25424
rect 45284 25381 45293 25415
rect 45293 25381 45327 25415
rect 45327 25381 45336 25415
rect 45284 25372 45336 25381
rect 35348 25236 35400 25288
rect 36544 25279 36596 25288
rect 36544 25245 36553 25279
rect 36553 25245 36587 25279
rect 36587 25245 36596 25279
rect 36544 25236 36596 25245
rect 37096 25236 37148 25288
rect 26056 25211 26108 25220
rect 26056 25177 26065 25211
rect 26065 25177 26099 25211
rect 26099 25177 26108 25211
rect 26056 25168 26108 25177
rect 17776 25143 17828 25152
rect 17776 25109 17785 25143
rect 17785 25109 17819 25143
rect 17819 25109 17828 25143
rect 17776 25100 17828 25109
rect 25228 25100 25280 25152
rect 28172 25168 28224 25220
rect 33232 25168 33284 25220
rect 26976 25143 27028 25152
rect 26976 25109 26985 25143
rect 26985 25109 27019 25143
rect 27019 25109 27028 25143
rect 26976 25100 27028 25109
rect 30840 25143 30892 25152
rect 30840 25109 30849 25143
rect 30849 25109 30883 25143
rect 30883 25109 30892 25143
rect 30840 25100 30892 25109
rect 34336 25100 34388 25152
rect 34520 25143 34572 25152
rect 34520 25109 34529 25143
rect 34529 25109 34563 25143
rect 34563 25109 34572 25143
rect 34520 25100 34572 25109
rect 35440 25100 35492 25152
rect 38476 25279 38528 25288
rect 38476 25245 38485 25279
rect 38485 25245 38519 25279
rect 38519 25245 38528 25279
rect 38476 25236 38528 25245
rect 43720 25304 43772 25356
rect 43904 25347 43956 25356
rect 43904 25313 43913 25347
rect 43913 25313 43947 25347
rect 43947 25313 43956 25347
rect 43904 25304 43956 25313
rect 45836 25304 45888 25356
rect 39120 25236 39172 25288
rect 40316 25279 40368 25288
rect 40316 25245 40325 25279
rect 40325 25245 40359 25279
rect 40359 25245 40368 25279
rect 40316 25236 40368 25245
rect 43996 25279 44048 25288
rect 43996 25245 44005 25279
rect 44005 25245 44039 25279
rect 44039 25245 44048 25279
rect 43996 25236 44048 25245
rect 44456 25279 44508 25288
rect 44456 25245 44465 25279
rect 44465 25245 44499 25279
rect 44499 25245 44508 25279
rect 44456 25236 44508 25245
rect 44548 25236 44600 25288
rect 45928 25279 45980 25288
rect 45928 25245 45937 25279
rect 45937 25245 45971 25279
rect 45971 25245 45980 25279
rect 45928 25236 45980 25245
rect 38752 25168 38804 25220
rect 39304 25211 39356 25220
rect 39304 25177 39313 25211
rect 39313 25177 39347 25211
rect 39347 25177 39356 25211
rect 39304 25168 39356 25177
rect 45744 25168 45796 25220
rect 38844 25100 38896 25152
rect 38936 25100 38988 25152
rect 40040 25100 40092 25152
rect 40868 25100 40920 25152
rect 44732 25100 44784 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 2780 24939 2832 24948
rect 2780 24905 2789 24939
rect 2789 24905 2823 24939
rect 2823 24905 2832 24939
rect 2780 24896 2832 24905
rect 5264 24896 5316 24948
rect 5632 24896 5684 24948
rect 13268 24896 13320 24948
rect 18052 24896 18104 24948
rect 18604 24896 18656 24948
rect 5540 24828 5592 24880
rect 6000 24828 6052 24880
rect 8392 24828 8444 24880
rect 940 24760 992 24812
rect 2412 24735 2464 24744
rect 2412 24701 2421 24735
rect 2421 24701 2455 24735
rect 2455 24701 2464 24735
rect 2412 24692 2464 24701
rect 2504 24735 2556 24744
rect 2504 24701 2513 24735
rect 2513 24701 2547 24735
rect 2547 24701 2556 24735
rect 2504 24692 2556 24701
rect 7380 24760 7432 24812
rect 7196 24692 7248 24744
rect 9128 24760 9180 24812
rect 9680 24760 9732 24812
rect 12440 24760 12492 24812
rect 18236 24828 18288 24880
rect 19892 24896 19944 24948
rect 25228 24896 25280 24948
rect 1584 24599 1636 24608
rect 1584 24565 1593 24599
rect 1593 24565 1627 24599
rect 1627 24565 1636 24599
rect 1584 24556 1636 24565
rect 11520 24692 11572 24744
rect 16028 24692 16080 24744
rect 17776 24735 17828 24744
rect 17776 24701 17785 24735
rect 17785 24701 17819 24735
rect 17819 24701 17828 24735
rect 17776 24692 17828 24701
rect 18972 24692 19024 24744
rect 19432 24803 19484 24812
rect 19432 24769 19441 24803
rect 19441 24769 19475 24803
rect 19475 24769 19484 24803
rect 19432 24760 19484 24769
rect 21272 24828 21324 24880
rect 24492 24828 24544 24880
rect 19524 24735 19576 24744
rect 19524 24701 19533 24735
rect 19533 24701 19567 24735
rect 19567 24701 19576 24735
rect 19524 24692 19576 24701
rect 14096 24624 14148 24676
rect 10600 24556 10652 24608
rect 19616 24624 19668 24676
rect 19156 24599 19208 24608
rect 19156 24565 19165 24599
rect 19165 24565 19199 24599
rect 19199 24565 19208 24599
rect 22376 24803 22428 24812
rect 22376 24769 22385 24803
rect 22385 24769 22419 24803
rect 22419 24769 22428 24803
rect 22376 24760 22428 24769
rect 25228 24760 25280 24812
rect 26976 24896 27028 24948
rect 33232 24896 33284 24948
rect 36176 24896 36228 24948
rect 36268 24896 36320 24948
rect 36912 24896 36964 24948
rect 41144 24939 41196 24948
rect 41144 24905 41153 24939
rect 41153 24905 41187 24939
rect 41187 24905 41196 24939
rect 41144 24896 41196 24905
rect 25504 24760 25556 24812
rect 26056 24760 26108 24812
rect 27252 24803 27304 24812
rect 27252 24769 27286 24803
rect 27286 24769 27304 24803
rect 27252 24760 27304 24769
rect 30656 24828 30708 24880
rect 30840 24871 30892 24880
rect 30840 24837 30874 24871
rect 30874 24837 30892 24871
rect 30840 24828 30892 24837
rect 28724 24760 28776 24812
rect 30196 24803 30248 24812
rect 30196 24769 30205 24803
rect 30205 24769 30239 24803
rect 30239 24769 30248 24803
rect 30196 24760 30248 24769
rect 30472 24803 30524 24812
rect 30472 24769 30481 24803
rect 30481 24769 30515 24803
rect 30515 24769 30524 24803
rect 30472 24760 30524 24769
rect 32404 24803 32456 24812
rect 32404 24769 32413 24803
rect 32413 24769 32447 24803
rect 32447 24769 32456 24803
rect 32404 24760 32456 24769
rect 33324 24803 33376 24812
rect 33324 24769 33333 24803
rect 33333 24769 33367 24803
rect 33367 24769 33376 24803
rect 33324 24760 33376 24769
rect 34336 24803 34388 24812
rect 34336 24769 34345 24803
rect 34345 24769 34379 24803
rect 34379 24769 34388 24803
rect 34336 24760 34388 24769
rect 34612 24803 34664 24812
rect 34612 24769 34621 24803
rect 34621 24769 34655 24803
rect 34655 24769 34664 24803
rect 34612 24760 34664 24769
rect 37280 24828 37332 24880
rect 38844 24828 38896 24880
rect 41696 24896 41748 24948
rect 44180 24896 44232 24948
rect 36360 24760 36412 24812
rect 38568 24803 38620 24812
rect 38568 24769 38577 24803
rect 38577 24769 38611 24803
rect 38611 24769 38620 24803
rect 38568 24760 38620 24769
rect 20444 24735 20496 24744
rect 20444 24701 20453 24735
rect 20453 24701 20487 24735
rect 20487 24701 20496 24735
rect 20444 24692 20496 24701
rect 20536 24735 20588 24744
rect 20536 24701 20570 24735
rect 20570 24701 20588 24735
rect 20536 24692 20588 24701
rect 21456 24692 21508 24744
rect 22100 24735 22152 24744
rect 22100 24701 22109 24735
rect 22109 24701 22143 24735
rect 22143 24701 22152 24735
rect 22100 24692 22152 24701
rect 26976 24735 27028 24744
rect 26976 24701 26985 24735
rect 26985 24701 27019 24735
rect 27019 24701 27028 24735
rect 26976 24692 27028 24701
rect 29092 24735 29144 24744
rect 29092 24701 29101 24735
rect 29101 24701 29135 24735
rect 29135 24701 29144 24735
rect 29092 24692 29144 24701
rect 20260 24624 20312 24676
rect 19156 24556 19208 24565
rect 20720 24556 20772 24608
rect 21916 24556 21968 24608
rect 22468 24556 22520 24608
rect 23112 24599 23164 24608
rect 23112 24565 23121 24599
rect 23121 24565 23155 24599
rect 23155 24565 23164 24599
rect 23112 24556 23164 24565
rect 24676 24556 24728 24608
rect 26608 24556 26660 24608
rect 26700 24556 26752 24608
rect 26976 24556 27028 24608
rect 29368 24624 29420 24676
rect 29644 24624 29696 24676
rect 30012 24692 30064 24744
rect 30564 24735 30616 24744
rect 30564 24701 30573 24735
rect 30573 24701 30607 24735
rect 30607 24701 30616 24735
rect 30564 24692 30616 24701
rect 33416 24735 33468 24744
rect 33416 24701 33425 24735
rect 33425 24701 33459 24735
rect 33459 24701 33468 24735
rect 33416 24692 33468 24701
rect 33784 24692 33836 24744
rect 33968 24692 34020 24744
rect 34152 24692 34204 24744
rect 36176 24692 36228 24744
rect 39212 24760 39264 24812
rect 39580 24803 39632 24812
rect 39580 24769 39589 24803
rect 39589 24769 39623 24803
rect 39623 24769 39632 24803
rect 39580 24760 39632 24769
rect 40684 24803 40736 24812
rect 40684 24769 40693 24803
rect 40693 24769 40727 24803
rect 40727 24769 40736 24803
rect 40684 24760 40736 24769
rect 39396 24692 39448 24744
rect 40868 24803 40920 24812
rect 40868 24769 40877 24803
rect 40877 24769 40911 24803
rect 40911 24769 40920 24803
rect 40868 24760 40920 24769
rect 41788 24828 41840 24880
rect 41420 24803 41472 24812
rect 41420 24769 41429 24803
rect 41429 24769 41463 24803
rect 41463 24769 41472 24803
rect 41420 24760 41472 24769
rect 42524 24760 42576 24812
rect 44548 24828 44600 24880
rect 43996 24760 44048 24812
rect 44456 24760 44508 24812
rect 44732 24803 44784 24812
rect 44732 24769 44741 24803
rect 44741 24769 44775 24803
rect 44775 24769 44784 24803
rect 44732 24760 44784 24769
rect 46388 24760 46440 24812
rect 41236 24692 41288 24744
rect 41512 24735 41564 24744
rect 41512 24701 41521 24735
rect 41521 24701 41555 24735
rect 41555 24701 41564 24735
rect 41512 24692 41564 24701
rect 30380 24624 30432 24676
rect 32956 24624 33008 24676
rect 40132 24624 40184 24676
rect 43720 24624 43772 24676
rect 28356 24599 28408 24608
rect 28356 24565 28365 24599
rect 28365 24565 28399 24599
rect 28399 24565 28408 24599
rect 28356 24556 28408 24565
rect 29736 24556 29788 24608
rect 29828 24556 29880 24608
rect 31668 24556 31720 24608
rect 32220 24599 32272 24608
rect 32220 24565 32229 24599
rect 32229 24565 32263 24599
rect 32263 24565 32272 24599
rect 32220 24556 32272 24565
rect 33232 24556 33284 24608
rect 39212 24556 39264 24608
rect 39488 24556 39540 24608
rect 46572 24599 46624 24608
rect 46572 24565 46581 24599
rect 46581 24565 46615 24599
rect 46615 24565 46624 24599
rect 46572 24556 46624 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 7472 24352 7524 24404
rect 8944 24284 8996 24336
rect 4528 24148 4580 24200
rect 4804 24148 4856 24200
rect 3700 24080 3752 24132
rect 4620 24012 4672 24064
rect 4804 24012 4856 24064
rect 6276 24259 6328 24268
rect 6276 24225 6285 24259
rect 6285 24225 6319 24259
rect 6319 24225 6328 24259
rect 6276 24216 6328 24225
rect 6552 24191 6604 24200
rect 6552 24157 6586 24191
rect 6586 24157 6604 24191
rect 6552 24148 6604 24157
rect 7288 24148 7340 24200
rect 14372 24352 14424 24404
rect 13084 24284 13136 24336
rect 13636 24284 13688 24336
rect 13176 24216 13228 24268
rect 9312 24080 9364 24132
rect 7380 24012 7432 24064
rect 8300 24012 8352 24064
rect 14096 24191 14148 24200
rect 14096 24157 14105 24191
rect 14105 24157 14139 24191
rect 14139 24157 14148 24191
rect 14096 24148 14148 24157
rect 16028 24259 16080 24268
rect 16028 24225 16037 24259
rect 16037 24225 16071 24259
rect 16071 24225 16080 24259
rect 16028 24216 16080 24225
rect 12808 24080 12860 24132
rect 13636 24080 13688 24132
rect 13268 24012 13320 24064
rect 13360 24012 13412 24064
rect 15936 24191 15988 24200
rect 15936 24157 15945 24191
rect 15945 24157 15979 24191
rect 15979 24157 15988 24191
rect 15936 24148 15988 24157
rect 14556 24012 14608 24064
rect 15016 24012 15068 24064
rect 15476 24012 15528 24064
rect 17592 24352 17644 24404
rect 19432 24352 19484 24404
rect 19616 24352 19668 24404
rect 18880 24216 18932 24268
rect 19156 24148 19208 24200
rect 20168 24259 20220 24268
rect 20168 24225 20177 24259
rect 20177 24225 20211 24259
rect 20211 24225 20220 24259
rect 20168 24216 20220 24225
rect 20536 24259 20588 24268
rect 20536 24225 20570 24259
rect 20570 24225 20588 24259
rect 20536 24216 20588 24225
rect 20720 24259 20772 24268
rect 20720 24225 20729 24259
rect 20729 24225 20763 24259
rect 20763 24225 20772 24259
rect 20720 24216 20772 24225
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 20444 24191 20496 24200
rect 20444 24157 20453 24191
rect 20453 24157 20487 24191
rect 20487 24157 20496 24191
rect 20444 24148 20496 24157
rect 19708 24080 19760 24132
rect 17408 24055 17460 24064
rect 17408 24021 17417 24055
rect 17417 24021 17451 24055
rect 17451 24021 17460 24055
rect 17408 24012 17460 24021
rect 17592 24012 17644 24064
rect 20168 24012 20220 24064
rect 21548 24352 21600 24404
rect 22376 24352 22428 24404
rect 23112 24352 23164 24404
rect 21916 24327 21968 24336
rect 21916 24293 21925 24327
rect 21925 24293 21959 24327
rect 21959 24293 21968 24327
rect 21916 24284 21968 24293
rect 22836 24284 22888 24336
rect 26056 24395 26108 24404
rect 26056 24361 26065 24395
rect 26065 24361 26099 24395
rect 26099 24361 26108 24395
rect 26056 24352 26108 24361
rect 26976 24352 27028 24404
rect 27252 24352 27304 24404
rect 27896 24352 27948 24404
rect 28632 24352 28684 24404
rect 28724 24352 28776 24404
rect 31024 24352 31076 24404
rect 22376 24191 22428 24200
rect 22376 24157 22385 24191
rect 22385 24157 22419 24191
rect 22419 24157 22428 24191
rect 22376 24148 22428 24157
rect 26700 24284 26752 24336
rect 21640 24123 21692 24132
rect 21640 24089 21649 24123
rect 21649 24089 21683 24123
rect 21683 24089 21692 24123
rect 21640 24080 21692 24089
rect 23388 24216 23440 24268
rect 26976 24259 27028 24268
rect 26976 24225 26985 24259
rect 26985 24225 27019 24259
rect 27019 24225 27028 24259
rect 26976 24216 27028 24225
rect 27528 24216 27580 24268
rect 28080 24259 28132 24268
rect 28080 24225 28089 24259
rect 28089 24225 28123 24259
rect 28123 24225 28132 24259
rect 28080 24216 28132 24225
rect 29092 24284 29144 24336
rect 33232 24352 33284 24404
rect 33324 24352 33376 24404
rect 33784 24352 33836 24404
rect 36820 24352 36872 24404
rect 37004 24352 37056 24404
rect 33508 24284 33560 24336
rect 29000 24216 29052 24268
rect 29184 24216 29236 24268
rect 23204 24148 23256 24200
rect 23756 24148 23808 24200
rect 23940 24148 23992 24200
rect 24308 24148 24360 24200
rect 24676 24191 24728 24200
rect 24676 24157 24710 24191
rect 24710 24157 24728 24191
rect 24676 24148 24728 24157
rect 24032 24123 24084 24132
rect 24032 24089 24041 24123
rect 24041 24089 24075 24123
rect 24075 24089 24084 24123
rect 24032 24080 24084 24089
rect 23204 24055 23256 24064
rect 23204 24021 23213 24055
rect 23213 24021 23247 24055
rect 23247 24021 23256 24055
rect 23204 24012 23256 24021
rect 23940 24012 23992 24064
rect 25780 24148 25832 24200
rect 26056 24012 26108 24064
rect 26700 24191 26752 24200
rect 26700 24157 26709 24191
rect 26709 24157 26743 24191
rect 26743 24157 26752 24191
rect 26700 24148 26752 24157
rect 26608 24080 26660 24132
rect 27068 24148 27120 24200
rect 27804 24148 27856 24200
rect 28356 24191 28408 24200
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 28632 24191 28684 24200
rect 28632 24157 28641 24191
rect 28641 24157 28675 24191
rect 28675 24157 28684 24191
rect 28632 24148 28684 24157
rect 29736 24191 29788 24200
rect 29736 24157 29745 24191
rect 29745 24157 29779 24191
rect 29779 24157 29788 24191
rect 29736 24148 29788 24157
rect 29828 24191 29880 24200
rect 29828 24157 29837 24191
rect 29837 24157 29871 24191
rect 29871 24157 29880 24191
rect 29828 24148 29880 24157
rect 30472 24216 30524 24268
rect 30840 24216 30892 24268
rect 31392 24259 31444 24268
rect 31392 24225 31401 24259
rect 31401 24225 31435 24259
rect 31435 24225 31444 24259
rect 31392 24216 31444 24225
rect 34244 24259 34296 24268
rect 34244 24225 34253 24259
rect 34253 24225 34287 24259
rect 34287 24225 34296 24259
rect 34244 24216 34296 24225
rect 37832 24284 37884 24336
rect 38568 24284 38620 24336
rect 31208 24148 31260 24200
rect 31760 24148 31812 24200
rect 32220 24191 32272 24200
rect 32220 24157 32254 24191
rect 32254 24157 32272 24191
rect 32220 24148 32272 24157
rect 33508 24148 33560 24200
rect 33876 24148 33928 24200
rect 27528 24080 27580 24132
rect 29552 24123 29604 24132
rect 29552 24089 29561 24123
rect 29561 24089 29595 24123
rect 29595 24089 29604 24123
rect 29552 24080 29604 24089
rect 34520 24148 34572 24200
rect 29368 24012 29420 24064
rect 31668 24012 31720 24064
rect 32772 24012 32824 24064
rect 34152 24080 34204 24132
rect 34336 24080 34388 24132
rect 36452 24216 36504 24268
rect 36728 24216 36780 24268
rect 35440 24148 35492 24200
rect 36360 24080 36412 24132
rect 36636 24080 36688 24132
rect 38292 24191 38344 24200
rect 38292 24157 38301 24191
rect 38301 24157 38335 24191
rect 38335 24157 38344 24191
rect 38292 24148 38344 24157
rect 38476 24191 38528 24200
rect 38476 24157 38483 24191
rect 38483 24157 38528 24191
rect 38476 24148 38528 24157
rect 41512 24352 41564 24404
rect 42156 24284 42208 24336
rect 42432 24259 42484 24268
rect 42432 24225 42441 24259
rect 42441 24225 42475 24259
rect 42475 24225 42484 24259
rect 42432 24216 42484 24225
rect 42524 24259 42576 24268
rect 42524 24225 42533 24259
rect 42533 24225 42567 24259
rect 42567 24225 42576 24259
rect 42524 24216 42576 24225
rect 39304 24148 39356 24200
rect 40040 24191 40092 24200
rect 40040 24157 40049 24191
rect 40049 24157 40083 24191
rect 40083 24157 40092 24191
rect 40040 24148 40092 24157
rect 41604 24148 41656 24200
rect 41880 24148 41932 24200
rect 41972 24191 42024 24200
rect 41972 24157 41981 24191
rect 41981 24157 42015 24191
rect 42015 24157 42024 24191
rect 41972 24148 42024 24157
rect 43076 24191 43128 24200
rect 43076 24157 43085 24191
rect 43085 24157 43119 24191
rect 43119 24157 43128 24191
rect 43076 24148 43128 24157
rect 44456 24284 44508 24336
rect 43352 24259 43404 24268
rect 43352 24225 43361 24259
rect 43361 24225 43395 24259
rect 43395 24225 43404 24259
rect 43352 24216 43404 24225
rect 45928 24216 45980 24268
rect 43260 24191 43312 24200
rect 43260 24157 43269 24191
rect 43269 24157 43303 24191
rect 43303 24157 43312 24191
rect 43260 24148 43312 24157
rect 44916 24148 44968 24200
rect 45192 24191 45244 24200
rect 45192 24157 45201 24191
rect 45201 24157 45235 24191
rect 45235 24157 45244 24191
rect 45192 24148 45244 24157
rect 45560 24148 45612 24200
rect 43536 24080 43588 24132
rect 45468 24123 45520 24132
rect 45468 24089 45477 24123
rect 45477 24089 45511 24123
rect 45511 24089 45520 24123
rect 45468 24080 45520 24089
rect 45652 24080 45704 24132
rect 46020 24191 46072 24200
rect 46020 24157 46029 24191
rect 46029 24157 46063 24191
rect 46063 24157 46072 24191
rect 46020 24148 46072 24157
rect 46664 24216 46716 24268
rect 45928 24080 45980 24132
rect 34704 24012 34756 24064
rect 35440 24012 35492 24064
rect 36084 24012 36136 24064
rect 36820 24012 36872 24064
rect 38384 24012 38436 24064
rect 39764 24012 39816 24064
rect 40592 24012 40644 24064
rect 42156 24012 42208 24064
rect 46572 24191 46624 24200
rect 46572 24157 46581 24191
rect 46581 24157 46615 24191
rect 46615 24157 46624 24191
rect 46572 24148 46624 24157
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 11520 23808 11572 23860
rect 12900 23808 12952 23860
rect 15936 23808 15988 23860
rect 17408 23808 17460 23860
rect 18788 23808 18840 23860
rect 19524 23808 19576 23860
rect 23112 23808 23164 23860
rect 23204 23808 23256 23860
rect 3240 23672 3292 23724
rect 5540 23715 5592 23724
rect 5540 23681 5549 23715
rect 5549 23681 5583 23715
rect 5583 23681 5592 23715
rect 5540 23672 5592 23681
rect 9128 23715 9180 23724
rect 9128 23681 9137 23715
rect 9137 23681 9171 23715
rect 9171 23681 9180 23715
rect 9128 23672 9180 23681
rect 10968 23672 11020 23724
rect 12164 23672 12216 23724
rect 12440 23672 12492 23724
rect 12992 23715 13044 23724
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 13360 23715 13412 23724
rect 13360 23681 13369 23715
rect 13369 23681 13403 23715
rect 13403 23681 13412 23715
rect 13360 23672 13412 23681
rect 13636 23672 13688 23724
rect 5080 23604 5132 23656
rect 5264 23647 5316 23656
rect 5264 23613 5273 23647
rect 5273 23613 5307 23647
rect 5307 23613 5316 23647
rect 5264 23604 5316 23613
rect 5724 23604 5776 23656
rect 6184 23647 6236 23656
rect 6184 23613 6193 23647
rect 6193 23613 6227 23647
rect 6227 23613 6236 23647
rect 6184 23604 6236 23613
rect 9220 23647 9272 23656
rect 9220 23613 9229 23647
rect 9229 23613 9263 23647
rect 9263 23613 9272 23647
rect 9220 23604 9272 23613
rect 9312 23647 9364 23656
rect 9312 23613 9321 23647
rect 9321 23613 9355 23647
rect 9355 23613 9364 23647
rect 9312 23604 9364 23613
rect 12900 23647 12952 23656
rect 12900 23613 12909 23647
rect 12909 23613 12943 23647
rect 12943 23613 12952 23647
rect 12900 23604 12952 23613
rect 17592 23783 17644 23792
rect 17592 23749 17601 23783
rect 17601 23749 17635 23783
rect 17635 23749 17644 23783
rect 17592 23740 17644 23749
rect 19432 23740 19484 23792
rect 19800 23740 19852 23792
rect 15016 23672 15068 23724
rect 15384 23715 15436 23724
rect 15384 23681 15393 23715
rect 15393 23681 15427 23715
rect 15427 23681 15436 23715
rect 15384 23672 15436 23681
rect 15476 23672 15528 23724
rect 20812 23740 20864 23792
rect 20904 23740 20956 23792
rect 19984 23715 20036 23724
rect 19984 23681 19993 23715
rect 19993 23681 20027 23715
rect 20027 23681 20036 23715
rect 19984 23672 20036 23681
rect 21088 23715 21140 23724
rect 21088 23681 21097 23715
rect 21097 23681 21131 23715
rect 21131 23681 21140 23715
rect 21088 23672 21140 23681
rect 21272 23715 21324 23724
rect 21272 23681 21281 23715
rect 21281 23681 21315 23715
rect 21315 23681 21324 23715
rect 21272 23672 21324 23681
rect 21456 23740 21508 23792
rect 24032 23740 24084 23792
rect 25228 23851 25280 23860
rect 25228 23817 25237 23851
rect 25237 23817 25271 23851
rect 25271 23817 25280 23851
rect 25228 23808 25280 23817
rect 27068 23851 27120 23860
rect 27068 23817 27077 23851
rect 27077 23817 27111 23851
rect 27111 23817 27120 23851
rect 27068 23808 27120 23817
rect 29092 23808 29144 23860
rect 29644 23808 29696 23860
rect 32404 23851 32456 23860
rect 32404 23817 32413 23851
rect 32413 23817 32447 23851
rect 32447 23817 32456 23851
rect 32404 23808 32456 23817
rect 32772 23851 32824 23860
rect 32772 23817 32781 23851
rect 32781 23817 32815 23851
rect 32815 23817 32824 23851
rect 32772 23808 32824 23817
rect 33600 23808 33652 23860
rect 34612 23808 34664 23860
rect 35256 23851 35308 23860
rect 35256 23817 35265 23851
rect 35265 23817 35299 23851
rect 35299 23817 35308 23851
rect 35256 23808 35308 23817
rect 35348 23851 35400 23860
rect 35348 23817 35357 23851
rect 35357 23817 35391 23851
rect 35391 23817 35400 23851
rect 35348 23808 35400 23817
rect 35440 23808 35492 23860
rect 38292 23808 38344 23860
rect 42156 23808 42208 23860
rect 42340 23808 42392 23860
rect 43076 23808 43128 23860
rect 43996 23851 44048 23860
rect 43996 23817 44005 23851
rect 44005 23817 44039 23851
rect 44039 23817 44048 23851
rect 43996 23808 44048 23817
rect 44456 23808 44508 23860
rect 45192 23808 45244 23860
rect 46664 23808 46716 23860
rect 27620 23740 27672 23792
rect 31300 23740 31352 23792
rect 33324 23740 33376 23792
rect 4896 23536 4948 23588
rect 17224 23647 17276 23656
rect 17224 23613 17233 23647
rect 17233 23613 17267 23647
rect 17267 23613 17276 23647
rect 17224 23604 17276 23613
rect 2044 23468 2096 23520
rect 4528 23468 4580 23520
rect 5540 23468 5592 23520
rect 8024 23468 8076 23520
rect 8760 23511 8812 23520
rect 8760 23477 8769 23511
rect 8769 23477 8803 23511
rect 8803 23477 8812 23511
rect 8760 23468 8812 23477
rect 13176 23511 13228 23520
rect 13176 23477 13185 23511
rect 13185 23477 13219 23511
rect 13219 23477 13228 23511
rect 13176 23468 13228 23477
rect 15108 23511 15160 23520
rect 15108 23477 15117 23511
rect 15117 23477 15151 23511
rect 15151 23477 15160 23511
rect 20444 23604 20496 23656
rect 21456 23604 21508 23656
rect 21640 23672 21692 23724
rect 23940 23672 23992 23724
rect 26056 23672 26108 23724
rect 28264 23672 28316 23724
rect 28908 23715 28960 23724
rect 28908 23681 28942 23715
rect 28942 23681 28960 23715
rect 28908 23672 28960 23681
rect 30472 23715 30524 23724
rect 30472 23681 30481 23715
rect 30481 23681 30515 23715
rect 30515 23681 30524 23715
rect 30472 23672 30524 23681
rect 34336 23715 34388 23724
rect 34336 23681 34345 23715
rect 34345 23681 34379 23715
rect 34379 23681 34388 23715
rect 34336 23672 34388 23681
rect 21916 23604 21968 23656
rect 19248 23536 19300 23588
rect 19708 23536 19760 23588
rect 19800 23536 19852 23588
rect 20628 23536 20680 23588
rect 25504 23604 25556 23656
rect 15108 23468 15160 23477
rect 19524 23468 19576 23520
rect 19984 23468 20036 23520
rect 20168 23468 20220 23520
rect 25228 23536 25280 23588
rect 25596 23536 25648 23588
rect 27712 23604 27764 23656
rect 27988 23604 28040 23656
rect 27804 23536 27856 23588
rect 29092 23647 29144 23656
rect 29092 23613 29101 23647
rect 29101 23613 29135 23647
rect 29135 23613 29144 23647
rect 29092 23604 29144 23613
rect 29460 23604 29512 23656
rect 29828 23604 29880 23656
rect 31392 23604 31444 23656
rect 33048 23647 33100 23656
rect 33048 23613 33057 23647
rect 33057 23613 33091 23647
rect 33091 23613 33100 23647
rect 33048 23604 33100 23613
rect 33416 23647 33468 23656
rect 33416 23613 33425 23647
rect 33425 23613 33459 23647
rect 33459 23613 33468 23647
rect 33416 23604 33468 23613
rect 27436 23468 27488 23520
rect 27528 23468 27580 23520
rect 28540 23579 28592 23588
rect 28540 23545 28549 23579
rect 28549 23545 28583 23579
rect 28583 23545 28592 23579
rect 28540 23536 28592 23545
rect 31208 23536 31260 23588
rect 30196 23468 30248 23520
rect 34152 23604 34204 23656
rect 34612 23647 34664 23656
rect 34612 23613 34621 23647
rect 34621 23613 34655 23647
rect 34655 23613 34664 23647
rect 34612 23604 34664 23613
rect 36084 23672 36136 23724
rect 36544 23672 36596 23724
rect 38108 23715 38160 23724
rect 38108 23681 38117 23715
rect 38117 23681 38151 23715
rect 38151 23681 38160 23715
rect 38108 23672 38160 23681
rect 38292 23672 38344 23724
rect 39488 23715 39540 23724
rect 39488 23681 39497 23715
rect 39497 23681 39531 23715
rect 39531 23681 39540 23715
rect 39488 23672 39540 23681
rect 39764 23715 39816 23724
rect 39764 23681 39773 23715
rect 39773 23681 39807 23715
rect 39807 23681 39816 23715
rect 39764 23672 39816 23681
rect 39948 23715 40000 23724
rect 39948 23681 39957 23715
rect 39957 23681 39991 23715
rect 39991 23681 40000 23715
rect 39948 23672 40000 23681
rect 40500 23672 40552 23724
rect 40592 23715 40644 23724
rect 40592 23681 40601 23715
rect 40601 23681 40635 23715
rect 40635 23681 40644 23715
rect 40592 23672 40644 23681
rect 41880 23740 41932 23792
rect 42800 23740 42852 23792
rect 43352 23740 43404 23792
rect 45468 23740 45520 23792
rect 41420 23672 41472 23724
rect 41604 23715 41656 23724
rect 41604 23681 41613 23715
rect 41613 23681 41647 23715
rect 41647 23681 41656 23715
rect 41604 23672 41656 23681
rect 41696 23672 41748 23724
rect 33784 23536 33836 23588
rect 33876 23536 33928 23588
rect 35348 23536 35400 23588
rect 36360 23604 36412 23656
rect 43720 23715 43772 23724
rect 43720 23681 43729 23715
rect 43729 23681 43763 23715
rect 43763 23681 43772 23715
rect 43720 23672 43772 23681
rect 36544 23536 36596 23588
rect 37372 23536 37424 23588
rect 39396 23536 39448 23588
rect 39764 23536 39816 23588
rect 39304 23468 39356 23520
rect 39948 23468 40000 23520
rect 42248 23536 42300 23588
rect 43076 23604 43128 23656
rect 44272 23672 44324 23724
rect 44456 23604 44508 23656
rect 45376 23604 45428 23656
rect 45652 23740 45704 23792
rect 45928 23672 45980 23724
rect 45744 23647 45796 23656
rect 45744 23613 45753 23647
rect 45753 23613 45787 23647
rect 45787 23613 45796 23647
rect 45744 23604 45796 23613
rect 46388 23579 46440 23588
rect 46388 23545 46397 23579
rect 46397 23545 46431 23579
rect 46431 23545 46440 23579
rect 46388 23536 46440 23545
rect 43720 23468 43772 23520
rect 44180 23468 44232 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2136 23264 2188 23316
rect 3792 23196 3844 23248
rect 12992 23264 13044 23316
rect 15384 23264 15436 23316
rect 17408 23239 17460 23248
rect 17408 23205 17417 23239
rect 17417 23205 17451 23239
rect 17451 23205 17460 23239
rect 17408 23196 17460 23205
rect 1676 23060 1728 23112
rect 2044 23103 2096 23112
rect 2044 23069 2078 23103
rect 2078 23069 2096 23103
rect 2044 23060 2096 23069
rect 4620 23128 4672 23180
rect 5080 23128 5132 23180
rect 5172 23171 5224 23180
rect 5172 23137 5181 23171
rect 5181 23137 5215 23171
rect 5215 23137 5224 23171
rect 5172 23128 5224 23137
rect 5632 23128 5684 23180
rect 4528 23103 4580 23112
rect 4528 23069 4537 23103
rect 4537 23069 4571 23103
rect 4571 23069 4580 23103
rect 4528 23060 4580 23069
rect 4896 23060 4948 23112
rect 5448 23103 5500 23112
rect 5448 23069 5457 23103
rect 5457 23069 5491 23103
rect 5491 23069 5500 23103
rect 5448 23060 5500 23069
rect 5724 23103 5776 23112
rect 5724 23069 5733 23103
rect 5733 23069 5767 23103
rect 5767 23069 5776 23103
rect 5724 23060 5776 23069
rect 8760 23103 8812 23112
rect 8760 23069 8769 23103
rect 8769 23069 8803 23103
rect 8803 23069 8812 23103
rect 8760 23060 8812 23069
rect 8944 23103 8996 23112
rect 8944 23069 8953 23103
rect 8953 23069 8987 23103
rect 8987 23069 8996 23103
rect 8944 23060 8996 23069
rect 14740 23171 14792 23180
rect 14740 23137 14749 23171
rect 14749 23137 14783 23171
rect 14783 23137 14792 23171
rect 14740 23128 14792 23137
rect 9680 23060 9732 23112
rect 15568 23103 15620 23112
rect 15568 23069 15577 23103
rect 15577 23069 15611 23103
rect 15611 23069 15620 23103
rect 15568 23060 15620 23069
rect 15660 23103 15712 23112
rect 15660 23069 15669 23103
rect 15669 23069 15703 23103
rect 15703 23069 15712 23103
rect 15660 23060 15712 23069
rect 4620 22924 4672 22976
rect 5632 22924 5684 22976
rect 6276 22924 6328 22976
rect 9404 22992 9456 23044
rect 9496 22924 9548 22976
rect 11888 22992 11940 23044
rect 13360 22992 13412 23044
rect 15108 22992 15160 23044
rect 14556 22967 14608 22976
rect 14556 22933 14565 22967
rect 14565 22933 14599 22967
rect 14599 22933 14608 22967
rect 14556 22924 14608 22933
rect 17592 23103 17644 23112
rect 17592 23069 17601 23103
rect 17601 23069 17635 23103
rect 17635 23069 17644 23103
rect 17592 23060 17644 23069
rect 17684 23103 17736 23112
rect 17684 23069 17693 23103
rect 17693 23069 17727 23103
rect 17727 23069 17736 23103
rect 17684 23060 17736 23069
rect 18788 23264 18840 23316
rect 21548 23196 21600 23248
rect 21640 23128 21692 23180
rect 22008 23128 22060 23180
rect 17408 22992 17460 23044
rect 18052 22992 18104 23044
rect 22744 23103 22796 23112
rect 22744 23069 22753 23103
rect 22753 23069 22787 23103
rect 22787 23069 22796 23103
rect 22744 23060 22796 23069
rect 24492 23196 24544 23248
rect 25596 23196 25648 23248
rect 26240 23196 26292 23248
rect 27712 23196 27764 23248
rect 23204 23128 23256 23180
rect 24676 23128 24728 23180
rect 29828 23128 29880 23180
rect 23388 23103 23440 23112
rect 23388 23069 23397 23103
rect 23397 23069 23431 23103
rect 23431 23069 23440 23103
rect 23388 23060 23440 23069
rect 23756 23060 23808 23112
rect 25596 23060 25648 23112
rect 29644 23060 29696 23112
rect 30012 23060 30064 23112
rect 30196 23103 30248 23112
rect 30196 23069 30230 23103
rect 30230 23069 30248 23103
rect 30196 23060 30248 23069
rect 31208 23264 31260 23316
rect 31392 23264 31444 23316
rect 32036 23264 32088 23316
rect 36636 23264 36688 23316
rect 38844 23264 38896 23316
rect 41880 23264 41932 23316
rect 42432 23264 42484 23316
rect 32956 23196 33008 23248
rect 34060 23196 34112 23248
rect 31024 23128 31076 23180
rect 32956 23060 33008 23112
rect 33324 23171 33376 23180
rect 33324 23137 33333 23171
rect 33333 23137 33367 23171
rect 33367 23137 33376 23171
rect 33324 23128 33376 23137
rect 34704 23128 34756 23180
rect 42064 23196 42116 23248
rect 36912 23171 36964 23180
rect 36912 23137 36921 23171
rect 36921 23137 36955 23171
rect 36955 23137 36964 23171
rect 36912 23128 36964 23137
rect 38660 23128 38712 23180
rect 39028 23128 39080 23180
rect 42524 23171 42576 23180
rect 42524 23137 42533 23171
rect 42533 23137 42567 23171
rect 42567 23137 42576 23171
rect 42524 23128 42576 23137
rect 43076 23196 43128 23248
rect 44640 23196 44692 23248
rect 46388 23196 46440 23248
rect 46940 23196 46992 23248
rect 17040 22967 17092 22976
rect 17040 22933 17049 22967
rect 17049 22933 17083 22967
rect 17083 22933 17092 22967
rect 17040 22924 17092 22933
rect 19892 22924 19944 22976
rect 22008 22924 22060 22976
rect 22560 22967 22612 22976
rect 22560 22933 22569 22967
rect 22569 22933 22603 22967
rect 22603 22933 22612 22967
rect 22560 22924 22612 22933
rect 32864 22992 32916 23044
rect 24952 22924 25004 22976
rect 27620 22924 27672 22976
rect 31024 22924 31076 22976
rect 36820 23060 36872 23112
rect 39672 23060 39724 23112
rect 42432 23060 42484 23112
rect 42892 23060 42944 23112
rect 43720 23171 43772 23180
rect 43720 23137 43729 23171
rect 43729 23137 43763 23171
rect 43763 23137 43772 23171
rect 43720 23128 43772 23137
rect 43536 23103 43588 23112
rect 43536 23069 43545 23103
rect 43545 23069 43579 23103
rect 43579 23069 43588 23103
rect 43536 23060 43588 23069
rect 43628 23060 43680 23112
rect 44180 23103 44232 23112
rect 44180 23069 44189 23103
rect 44189 23069 44223 23103
rect 44223 23069 44232 23103
rect 44180 23060 44232 23069
rect 44272 23103 44324 23112
rect 44272 23069 44281 23103
rect 44281 23069 44315 23103
rect 44315 23069 44324 23103
rect 44272 23060 44324 23069
rect 44916 23128 44968 23180
rect 43720 22992 43772 23044
rect 45192 22992 45244 23044
rect 45928 23060 45980 23112
rect 45744 22992 45796 23044
rect 46572 23103 46624 23112
rect 46572 23069 46581 23103
rect 46581 23069 46615 23103
rect 46615 23069 46624 23103
rect 46572 23060 46624 23069
rect 38384 22924 38436 22976
rect 42616 22924 42668 22976
rect 42892 22967 42944 22976
rect 42892 22933 42901 22967
rect 42901 22933 42935 22967
rect 42935 22933 42944 22967
rect 42892 22924 42944 22933
rect 43260 22967 43312 22976
rect 43260 22933 43269 22967
rect 43269 22933 43303 22967
rect 43303 22933 43312 22967
rect 43260 22924 43312 22933
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 3240 22763 3292 22772
rect 3240 22729 3249 22763
rect 3249 22729 3283 22763
rect 3283 22729 3292 22763
rect 3240 22720 3292 22729
rect 3792 22720 3844 22772
rect 3700 22695 3752 22704
rect 3700 22661 3709 22695
rect 3709 22661 3743 22695
rect 3743 22661 3752 22695
rect 3700 22652 3752 22661
rect 4804 22720 4856 22772
rect 5356 22720 5408 22772
rect 5724 22720 5776 22772
rect 8392 22720 8444 22772
rect 5632 22652 5684 22704
rect 2044 22627 2096 22636
rect 2044 22593 2078 22627
rect 2078 22593 2096 22627
rect 2044 22584 2096 22593
rect 5356 22584 5408 22636
rect 8392 22584 8444 22636
rect 8576 22720 8628 22772
rect 9220 22720 9272 22772
rect 10784 22720 10836 22772
rect 11152 22720 11204 22772
rect 12900 22720 12952 22772
rect 12992 22720 13044 22772
rect 15292 22720 15344 22772
rect 15568 22720 15620 22772
rect 17592 22720 17644 22772
rect 9404 22652 9456 22704
rect 8852 22627 8904 22636
rect 8852 22593 8861 22627
rect 8861 22593 8895 22627
rect 8895 22593 8904 22627
rect 8852 22584 8904 22593
rect 9128 22584 9180 22636
rect 9496 22627 9548 22636
rect 9496 22593 9505 22627
rect 9505 22593 9539 22627
rect 9539 22593 9548 22627
rect 9496 22584 9548 22593
rect 1676 22516 1728 22568
rect 3792 22559 3844 22568
rect 3792 22525 3801 22559
rect 3801 22525 3835 22559
rect 3835 22525 3844 22559
rect 3792 22516 3844 22525
rect 4804 22559 4856 22568
rect 4804 22525 4813 22559
rect 4813 22525 4847 22559
rect 4847 22525 4856 22559
rect 4804 22516 4856 22525
rect 8208 22559 8260 22568
rect 8208 22525 8217 22559
rect 8217 22525 8251 22559
rect 8251 22525 8260 22559
rect 8208 22516 8260 22525
rect 8484 22516 8536 22568
rect 6184 22448 6236 22500
rect 2964 22380 3016 22432
rect 5540 22380 5592 22432
rect 7104 22380 7156 22432
rect 7840 22448 7892 22500
rect 9680 22559 9732 22568
rect 9680 22525 9689 22559
rect 9689 22525 9723 22559
rect 9723 22525 9732 22559
rect 9680 22516 9732 22525
rect 11888 22584 11940 22636
rect 11980 22584 12032 22636
rect 12532 22584 12584 22636
rect 12808 22584 12860 22636
rect 13176 22627 13228 22636
rect 13176 22593 13210 22627
rect 13210 22593 13228 22627
rect 13176 22584 13228 22593
rect 10416 22559 10468 22568
rect 10416 22525 10425 22559
rect 10425 22525 10459 22559
rect 10459 22525 10468 22559
rect 10416 22516 10468 22525
rect 10508 22559 10560 22568
rect 10508 22525 10542 22559
rect 10542 22525 10560 22559
rect 10508 22516 10560 22525
rect 13912 22448 13964 22500
rect 17500 22652 17552 22704
rect 20720 22720 20772 22772
rect 21548 22763 21600 22772
rect 21548 22729 21557 22763
rect 21557 22729 21591 22763
rect 21591 22729 21600 22763
rect 21548 22720 21600 22729
rect 16488 22584 16540 22636
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 17040 22584 17092 22593
rect 22744 22720 22796 22772
rect 23940 22720 23992 22772
rect 22560 22652 22612 22704
rect 28540 22652 28592 22704
rect 30472 22763 30524 22772
rect 30472 22729 30481 22763
rect 30481 22729 30515 22763
rect 30515 22729 30524 22763
rect 30472 22720 30524 22729
rect 31208 22720 31260 22772
rect 32956 22720 33008 22772
rect 38752 22763 38804 22772
rect 38752 22729 38761 22763
rect 38761 22729 38795 22763
rect 38795 22729 38804 22763
rect 38752 22720 38804 22729
rect 39672 22720 39724 22772
rect 44456 22720 44508 22772
rect 38200 22652 38252 22704
rect 14832 22559 14884 22568
rect 14832 22525 14841 22559
rect 14841 22525 14875 22559
rect 14875 22525 14884 22559
rect 14832 22516 14884 22525
rect 14924 22559 14976 22568
rect 14924 22525 14933 22559
rect 14933 22525 14967 22559
rect 14967 22525 14976 22559
rect 14924 22516 14976 22525
rect 16212 22516 16264 22568
rect 17224 22559 17276 22568
rect 17224 22525 17233 22559
rect 17233 22525 17267 22559
rect 17267 22525 17276 22559
rect 17224 22516 17276 22525
rect 18788 22559 18840 22568
rect 18788 22525 18797 22559
rect 18797 22525 18831 22559
rect 18831 22525 18840 22559
rect 18788 22516 18840 22525
rect 18880 22559 18932 22568
rect 18880 22525 18889 22559
rect 18889 22525 18923 22559
rect 18923 22525 18932 22559
rect 18880 22516 18932 22525
rect 19708 22559 19760 22568
rect 19708 22525 19717 22559
rect 19717 22525 19751 22559
rect 19751 22525 19760 22559
rect 19708 22516 19760 22525
rect 19892 22559 19944 22568
rect 19892 22525 19901 22559
rect 19901 22525 19935 22559
rect 19935 22525 19944 22559
rect 19892 22516 19944 22525
rect 20260 22516 20312 22568
rect 20628 22559 20680 22568
rect 20628 22525 20637 22559
rect 20637 22525 20671 22559
rect 20671 22525 20680 22559
rect 20628 22516 20680 22525
rect 20720 22559 20772 22568
rect 20720 22525 20754 22559
rect 20754 22525 20772 22559
rect 20720 22516 20772 22525
rect 20904 22559 20956 22568
rect 20904 22525 20913 22559
rect 20913 22525 20947 22559
rect 20947 22525 20956 22559
rect 20904 22516 20956 22525
rect 21272 22516 21324 22568
rect 21548 22516 21600 22568
rect 22468 22516 22520 22568
rect 23480 22584 23532 22636
rect 22744 22516 22796 22568
rect 22928 22559 22980 22568
rect 22928 22525 22937 22559
rect 22937 22525 22971 22559
rect 22971 22525 22980 22559
rect 22928 22516 22980 22525
rect 22008 22448 22060 22500
rect 23664 22516 23716 22568
rect 24400 22584 24452 22636
rect 24584 22627 24636 22636
rect 24584 22593 24618 22627
rect 24618 22593 24636 22627
rect 24584 22584 24636 22593
rect 25412 22584 25464 22636
rect 27620 22627 27672 22636
rect 27620 22593 27629 22627
rect 27629 22593 27663 22627
rect 27663 22593 27672 22627
rect 27620 22584 27672 22593
rect 16212 22423 16264 22432
rect 16212 22389 16221 22423
rect 16221 22389 16255 22423
rect 16255 22389 16264 22423
rect 16212 22380 16264 22389
rect 20260 22380 20312 22432
rect 24032 22448 24084 22500
rect 22468 22423 22520 22432
rect 22468 22389 22477 22423
rect 22477 22389 22511 22423
rect 22511 22389 22520 22423
rect 22468 22380 22520 22389
rect 24308 22380 24360 22432
rect 27068 22516 27120 22568
rect 25596 22448 25648 22500
rect 26976 22448 27028 22500
rect 27160 22448 27212 22500
rect 29092 22584 29144 22636
rect 30656 22584 30708 22636
rect 31300 22584 31352 22636
rect 36268 22584 36320 22636
rect 38476 22627 38528 22636
rect 38476 22593 38485 22627
rect 38485 22593 38519 22627
rect 38519 22593 38528 22627
rect 38476 22584 38528 22593
rect 38752 22627 38804 22636
rect 38752 22593 38761 22627
rect 38761 22593 38795 22627
rect 38795 22593 38804 22627
rect 38752 22584 38804 22593
rect 39120 22627 39172 22636
rect 39120 22593 39129 22627
rect 39129 22593 39163 22627
rect 39163 22593 39172 22627
rect 39120 22584 39172 22593
rect 42708 22627 42760 22636
rect 42708 22593 42717 22627
rect 42717 22593 42751 22627
rect 42751 22593 42760 22627
rect 42708 22584 42760 22593
rect 42892 22627 42944 22636
rect 42892 22593 42901 22627
rect 42901 22593 42935 22627
rect 42935 22593 42944 22627
rect 42892 22584 42944 22593
rect 28356 22559 28408 22568
rect 28356 22525 28365 22559
rect 28365 22525 28399 22559
rect 28399 22525 28408 22559
rect 28356 22516 28408 22525
rect 29460 22559 29512 22568
rect 29460 22525 29469 22559
rect 29469 22525 29503 22559
rect 29503 22525 29512 22559
rect 29460 22516 29512 22525
rect 28172 22448 28224 22500
rect 29368 22448 29420 22500
rect 37372 22516 37424 22568
rect 42616 22516 42668 22568
rect 43260 22516 43312 22568
rect 39856 22448 39908 22500
rect 43812 22448 43864 22500
rect 25780 22380 25832 22432
rect 27988 22380 28040 22432
rect 28908 22380 28960 22432
rect 30012 22380 30064 22432
rect 30656 22380 30708 22432
rect 31208 22380 31260 22432
rect 32864 22380 32916 22432
rect 38752 22380 38804 22432
rect 43260 22380 43312 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 2044 22176 2096 22228
rect 3240 22083 3292 22092
rect 3240 22049 3249 22083
rect 3249 22049 3283 22083
rect 3283 22049 3292 22083
rect 3240 22040 3292 22049
rect 940 21972 992 22024
rect 2412 21836 2464 21888
rect 2964 22015 3016 22024
rect 2964 21981 2973 22015
rect 2973 21981 3007 22015
rect 3007 21981 3016 22015
rect 2964 21972 3016 21981
rect 4804 22176 4856 22228
rect 5264 22219 5316 22228
rect 5264 22185 5273 22219
rect 5273 22185 5307 22219
rect 5307 22185 5316 22219
rect 5264 22176 5316 22185
rect 5356 22219 5408 22228
rect 5356 22185 5365 22219
rect 5365 22185 5399 22219
rect 5399 22185 5408 22219
rect 5356 22176 5408 22185
rect 8208 22176 8260 22228
rect 8392 22176 8444 22228
rect 10508 22176 10560 22228
rect 10784 22176 10836 22228
rect 6276 22108 6328 22160
rect 8852 22108 8904 22160
rect 13176 22176 13228 22228
rect 15660 22176 15712 22228
rect 4620 21972 4672 22024
rect 7196 22083 7248 22092
rect 7196 22049 7205 22083
rect 7205 22049 7239 22083
rect 7239 22049 7248 22083
rect 7196 22040 7248 22049
rect 9496 22083 9548 22092
rect 9496 22049 9505 22083
rect 9505 22049 9539 22083
rect 9539 22049 9548 22083
rect 9496 22040 9548 22049
rect 10140 22083 10192 22092
rect 10140 22049 10149 22083
rect 10149 22049 10183 22083
rect 10183 22049 10192 22083
rect 10140 22040 10192 22049
rect 14832 22108 14884 22160
rect 17500 22219 17552 22228
rect 17500 22185 17509 22219
rect 17509 22185 17543 22219
rect 17543 22185 17552 22219
rect 17500 22176 17552 22185
rect 18788 22176 18840 22228
rect 17684 22108 17736 22160
rect 20168 22108 20220 22160
rect 21824 22108 21876 22160
rect 22008 22108 22060 22160
rect 23480 22219 23532 22228
rect 23480 22185 23489 22219
rect 23489 22185 23523 22219
rect 23523 22185 23532 22219
rect 23480 22176 23532 22185
rect 24860 22176 24912 22228
rect 25780 22176 25832 22228
rect 26332 22176 26384 22228
rect 28172 22176 28224 22228
rect 24492 22108 24544 22160
rect 10416 22083 10468 22092
rect 10416 22049 10425 22083
rect 10425 22049 10459 22083
rect 10459 22049 10468 22083
rect 10416 22040 10468 22049
rect 10508 22083 10560 22092
rect 10508 22049 10542 22083
rect 10542 22049 10560 22083
rect 10508 22040 10560 22049
rect 5724 22015 5776 22024
rect 5724 21981 5733 22015
rect 5733 21981 5767 22015
rect 5767 21981 5776 22015
rect 5724 21972 5776 21981
rect 5816 21972 5868 22024
rect 6092 21972 6144 22024
rect 7104 22015 7156 22024
rect 7104 21981 7113 22015
rect 7113 21981 7147 22015
rect 7147 21981 7156 22015
rect 7104 21972 7156 21981
rect 9680 22015 9732 22024
rect 9680 21981 9689 22015
rect 9689 21981 9723 22015
rect 9723 21981 9732 22015
rect 9680 21972 9732 21981
rect 10692 22015 10744 22024
rect 10692 21981 10701 22015
rect 10701 21981 10735 22015
rect 10735 21981 10744 22015
rect 10692 21972 10744 21981
rect 11980 22040 12032 22092
rect 13912 21972 13964 22024
rect 14648 21972 14700 22024
rect 18696 22040 18748 22092
rect 19156 22040 19208 22092
rect 19892 22083 19944 22092
rect 19892 22049 19901 22083
rect 19901 22049 19935 22083
rect 19935 22049 19944 22083
rect 19892 22040 19944 22049
rect 20628 22083 20680 22092
rect 20628 22049 20637 22083
rect 20637 22049 20671 22083
rect 20671 22049 20680 22083
rect 20628 22040 20680 22049
rect 20720 22083 20772 22092
rect 20720 22049 20754 22083
rect 20754 22049 20772 22083
rect 20720 22040 20772 22049
rect 21088 22040 21140 22092
rect 21272 22040 21324 22092
rect 23940 22083 23992 22092
rect 23940 22049 23949 22083
rect 23949 22049 23983 22083
rect 23983 22049 23992 22083
rect 23940 22040 23992 22049
rect 24676 22040 24728 22092
rect 24768 22040 24820 22092
rect 25596 22108 25648 22160
rect 31208 22219 31260 22228
rect 31208 22185 31217 22219
rect 31217 22185 31251 22219
rect 31251 22185 31260 22219
rect 31208 22176 31260 22185
rect 35716 22176 35768 22228
rect 38476 22176 38528 22228
rect 38752 22176 38804 22228
rect 43352 22176 43404 22228
rect 16764 21972 16816 22024
rect 18788 21972 18840 22024
rect 19708 22015 19760 22024
rect 19708 21981 19717 22015
rect 19717 21981 19751 22015
rect 19751 21981 19760 22015
rect 19708 21972 19760 21981
rect 22836 21972 22888 22024
rect 24308 21972 24360 22024
rect 25964 22083 26016 22092
rect 25964 22049 25973 22083
rect 25973 22049 26007 22083
rect 26007 22049 26016 22083
rect 25964 22040 26016 22049
rect 26056 22040 26108 22092
rect 27068 22040 27120 22092
rect 31300 22040 31352 22092
rect 34612 22108 34664 22160
rect 35072 22108 35124 22160
rect 36268 22108 36320 22160
rect 36912 22108 36964 22160
rect 3700 21836 3752 21888
rect 5816 21879 5868 21888
rect 5816 21845 5825 21879
rect 5825 21845 5859 21879
rect 5859 21845 5868 21879
rect 5816 21836 5868 21845
rect 11888 21904 11940 21956
rect 17316 21904 17368 21956
rect 10692 21836 10744 21888
rect 11336 21879 11388 21888
rect 11336 21845 11345 21879
rect 11345 21845 11379 21879
rect 11379 21845 11388 21879
rect 11336 21836 11388 21845
rect 11796 21879 11848 21888
rect 11796 21845 11805 21879
rect 11805 21845 11839 21879
rect 11839 21845 11848 21879
rect 11796 21836 11848 21845
rect 13636 21836 13688 21888
rect 14924 21836 14976 21888
rect 18328 21904 18380 21956
rect 17960 21836 18012 21888
rect 18144 21836 18196 21888
rect 18696 21836 18748 21888
rect 22468 21904 22520 21956
rect 23572 21904 23624 21956
rect 23940 21904 23992 21956
rect 24032 21904 24084 21956
rect 24768 21904 24820 21956
rect 25412 21972 25464 22024
rect 24492 21879 24544 21888
rect 24492 21845 24501 21879
rect 24501 21845 24535 21879
rect 24535 21845 24544 21879
rect 24492 21836 24544 21845
rect 24676 21836 24728 21888
rect 24952 21836 25004 21888
rect 26332 22015 26384 22024
rect 26332 21981 26366 22015
rect 26366 21981 26384 22015
rect 26332 21972 26384 21981
rect 26516 22015 26568 22024
rect 26516 21981 26525 22015
rect 26525 21981 26559 22015
rect 26559 21981 26568 22015
rect 26516 21972 26568 21981
rect 28080 21972 28132 22024
rect 28356 21972 28408 22024
rect 28908 22015 28960 22024
rect 28908 21981 28917 22015
rect 28917 21981 28951 22015
rect 28951 21981 28960 22015
rect 28908 21972 28960 21981
rect 29736 22015 29788 22024
rect 29736 21981 29745 22015
rect 29745 21981 29779 22015
rect 29779 21981 29788 22015
rect 29736 21972 29788 21981
rect 30012 22015 30064 22024
rect 30012 21981 30046 22015
rect 30046 21981 30064 22015
rect 30012 21972 30064 21981
rect 27804 21904 27856 21956
rect 28540 21904 28592 21956
rect 33784 21972 33836 22024
rect 33968 21972 34020 22024
rect 35256 22083 35308 22092
rect 35256 22049 35265 22083
rect 35265 22049 35299 22083
rect 35299 22049 35308 22083
rect 35256 22040 35308 22049
rect 35348 22040 35400 22092
rect 36360 22040 36412 22092
rect 39856 22108 39908 22160
rect 42524 22108 42576 22160
rect 32404 21904 32456 21956
rect 34612 21904 34664 21956
rect 35164 21972 35216 22024
rect 35440 21972 35492 22024
rect 35716 22015 35768 22024
rect 35716 21981 35725 22015
rect 35725 21981 35759 22015
rect 35759 21981 35768 22015
rect 35716 21972 35768 21981
rect 36912 21972 36964 22024
rect 37372 21972 37424 22024
rect 37556 21972 37608 22024
rect 38752 21972 38804 22024
rect 39488 22040 39540 22092
rect 42892 22108 42944 22160
rect 26148 21836 26200 21888
rect 27344 21836 27396 21888
rect 27620 21836 27672 21888
rect 28724 21879 28776 21888
rect 28724 21845 28733 21879
rect 28733 21845 28767 21879
rect 28767 21845 28776 21879
rect 28724 21836 28776 21845
rect 30380 21836 30432 21888
rect 33968 21836 34020 21888
rect 36084 21836 36136 21888
rect 36360 21879 36412 21888
rect 36360 21845 36369 21879
rect 36369 21845 36403 21879
rect 36403 21845 36412 21879
rect 36360 21836 36412 21845
rect 36636 21836 36688 21888
rect 38844 21904 38896 21956
rect 38568 21836 38620 21888
rect 40040 21972 40092 22024
rect 42432 22015 42484 22024
rect 42432 21981 42441 22015
rect 42441 21981 42475 22015
rect 42475 21981 42484 22015
rect 42432 21972 42484 21981
rect 42616 22015 42668 22024
rect 42616 21981 42625 22015
rect 42625 21981 42659 22015
rect 42659 21981 42668 22015
rect 42616 21972 42668 21981
rect 42708 22015 42760 22024
rect 42708 21981 42717 22015
rect 42717 21981 42751 22015
rect 42751 21981 42760 22015
rect 42708 21972 42760 21981
rect 42800 22015 42852 22024
rect 42800 21981 42813 22015
rect 42813 21981 42847 22015
rect 42847 21981 42852 22015
rect 42800 21972 42852 21981
rect 39948 21836 40000 21888
rect 41604 21836 41656 21888
rect 42156 21879 42208 21888
rect 42156 21845 42165 21879
rect 42165 21845 42199 21879
rect 42199 21845 42208 21879
rect 42156 21836 42208 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 5816 21632 5868 21684
rect 8852 21632 8904 21684
rect 7196 21539 7248 21548
rect 7196 21505 7205 21539
rect 7205 21505 7239 21539
rect 7239 21505 7248 21539
rect 7196 21496 7248 21505
rect 7472 21539 7524 21548
rect 7472 21505 7506 21539
rect 7506 21505 7524 21539
rect 7472 21496 7524 21505
rect 10784 21675 10836 21684
rect 10784 21641 10793 21675
rect 10793 21641 10827 21675
rect 10827 21641 10836 21675
rect 10784 21632 10836 21641
rect 11336 21632 11388 21684
rect 19248 21607 19300 21616
rect 19248 21573 19257 21607
rect 19257 21573 19291 21607
rect 19291 21573 19300 21607
rect 19248 21564 19300 21573
rect 23848 21632 23900 21684
rect 24584 21632 24636 21684
rect 24768 21632 24820 21684
rect 27344 21675 27396 21684
rect 27344 21641 27353 21675
rect 27353 21641 27387 21675
rect 27387 21641 27396 21675
rect 27344 21632 27396 21641
rect 27804 21675 27856 21684
rect 27804 21641 27813 21675
rect 27813 21641 27847 21675
rect 27847 21641 27856 21675
rect 27804 21632 27856 21641
rect 10692 21539 10744 21548
rect 10692 21505 10701 21539
rect 10701 21505 10735 21539
rect 10735 21505 10744 21539
rect 10692 21496 10744 21505
rect 14556 21496 14608 21548
rect 16120 21496 16172 21548
rect 10416 21360 10468 21412
rect 15752 21428 15804 21480
rect 17132 21471 17184 21480
rect 17132 21437 17141 21471
rect 17141 21437 17175 21471
rect 17175 21437 17184 21471
rect 17132 21428 17184 21437
rect 17224 21428 17276 21480
rect 18052 21539 18104 21548
rect 18052 21505 18061 21539
rect 18061 21505 18095 21539
rect 18095 21505 18104 21539
rect 18052 21496 18104 21505
rect 18144 21539 18196 21548
rect 18144 21505 18178 21539
rect 18178 21505 18196 21539
rect 18144 21496 18196 21505
rect 18328 21539 18380 21548
rect 18328 21505 18337 21539
rect 18337 21505 18371 21539
rect 18371 21505 18380 21539
rect 18328 21496 18380 21505
rect 19064 21496 19116 21548
rect 19892 21496 19944 21548
rect 21456 21496 21508 21548
rect 21640 21539 21692 21548
rect 21640 21505 21649 21539
rect 21649 21505 21683 21539
rect 21683 21505 21692 21539
rect 21640 21496 21692 21505
rect 21824 21496 21876 21548
rect 22560 21539 22612 21548
rect 22560 21505 22571 21539
rect 22571 21505 22612 21539
rect 22560 21496 22612 21505
rect 17868 21360 17920 21412
rect 10140 21292 10192 21344
rect 15844 21292 15896 21344
rect 18144 21292 18196 21344
rect 20812 21292 20864 21344
rect 22100 21428 22152 21480
rect 22192 21471 22244 21480
rect 22192 21437 22201 21471
rect 22201 21437 22235 21471
rect 22235 21437 22244 21471
rect 22192 21428 22244 21437
rect 24400 21564 24452 21616
rect 32404 21632 32456 21684
rect 28724 21564 28776 21616
rect 29736 21564 29788 21616
rect 31760 21564 31812 21616
rect 22928 21496 22980 21548
rect 24308 21496 24360 21548
rect 24492 21496 24544 21548
rect 24768 21539 24820 21548
rect 24768 21505 24777 21539
rect 24777 21505 24811 21539
rect 24811 21505 24820 21539
rect 24768 21496 24820 21505
rect 25688 21539 25740 21548
rect 25688 21505 25697 21539
rect 25697 21505 25731 21539
rect 25731 21505 25740 21539
rect 25688 21496 25740 21505
rect 25780 21539 25832 21548
rect 25780 21505 25814 21539
rect 25814 21505 25832 21539
rect 25780 21496 25832 21505
rect 25964 21539 26016 21548
rect 25964 21505 25973 21539
rect 25973 21505 26007 21539
rect 26007 21505 26016 21539
rect 25964 21496 26016 21505
rect 27988 21539 28040 21548
rect 27988 21505 27997 21539
rect 27997 21505 28031 21539
rect 28031 21505 28040 21539
rect 27988 21496 28040 21505
rect 28080 21539 28132 21548
rect 28080 21505 28089 21539
rect 28089 21505 28123 21539
rect 28123 21505 28132 21539
rect 28080 21496 28132 21505
rect 24952 21471 25004 21480
rect 24952 21437 24961 21471
rect 24961 21437 24995 21471
rect 24995 21437 25004 21471
rect 24952 21428 25004 21437
rect 25044 21428 25096 21480
rect 30748 21496 30800 21548
rect 32956 21675 33008 21684
rect 32956 21641 32965 21675
rect 32965 21641 32999 21675
rect 32999 21641 33008 21675
rect 32956 21632 33008 21641
rect 33324 21496 33376 21548
rect 33600 21632 33652 21684
rect 35256 21632 35308 21684
rect 36084 21564 36136 21616
rect 36912 21632 36964 21684
rect 38844 21632 38896 21684
rect 40316 21632 40368 21684
rect 38752 21564 38804 21616
rect 39948 21564 40000 21616
rect 42708 21564 42760 21616
rect 35348 21539 35400 21548
rect 35348 21505 35357 21539
rect 35357 21505 35391 21539
rect 35391 21505 35400 21539
rect 35348 21496 35400 21505
rect 36360 21496 36412 21548
rect 39764 21496 39816 21548
rect 22468 21360 22520 21412
rect 22744 21360 22796 21412
rect 23940 21360 23992 21412
rect 22284 21292 22336 21344
rect 22560 21292 22612 21344
rect 27160 21360 27212 21412
rect 33048 21471 33100 21480
rect 33048 21437 33057 21471
rect 33057 21437 33091 21471
rect 33091 21437 33100 21471
rect 33048 21428 33100 21437
rect 33232 21428 33284 21480
rect 33692 21428 33744 21480
rect 34060 21471 34112 21480
rect 34060 21437 34069 21471
rect 34069 21437 34103 21471
rect 34103 21437 34112 21471
rect 34060 21428 34112 21437
rect 34336 21471 34388 21480
rect 34336 21437 34345 21471
rect 34345 21437 34379 21471
rect 34379 21437 34388 21471
rect 34336 21428 34388 21437
rect 34520 21428 34572 21480
rect 34980 21428 35032 21480
rect 36452 21428 36504 21480
rect 36820 21428 36872 21480
rect 29460 21403 29512 21412
rect 29460 21369 29469 21403
rect 29469 21369 29503 21403
rect 29503 21369 29512 21403
rect 29460 21360 29512 21369
rect 32956 21360 33008 21412
rect 33968 21360 34020 21412
rect 26516 21292 26568 21344
rect 31024 21292 31076 21344
rect 32220 21335 32272 21344
rect 32220 21301 32229 21335
rect 32229 21301 32263 21335
rect 32263 21301 32272 21335
rect 32220 21292 32272 21301
rect 33508 21292 33560 21344
rect 36636 21292 36688 21344
rect 38844 21428 38896 21480
rect 41604 21496 41656 21548
rect 42156 21496 42208 21548
rect 43168 21539 43220 21548
rect 43168 21505 43177 21539
rect 43177 21505 43211 21539
rect 43211 21505 43220 21539
rect 43168 21496 43220 21505
rect 43260 21539 43312 21548
rect 43260 21505 43269 21539
rect 43269 21505 43303 21539
rect 43303 21505 43312 21539
rect 43260 21496 43312 21505
rect 46756 21496 46808 21548
rect 41696 21428 41748 21480
rect 42616 21360 42668 21412
rect 43904 21428 43956 21480
rect 39580 21292 39632 21344
rect 40408 21292 40460 21344
rect 40960 21292 41012 21344
rect 41880 21292 41932 21344
rect 45744 21292 45796 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 7472 21131 7524 21140
rect 7472 21097 7481 21131
rect 7481 21097 7515 21131
rect 7515 21097 7524 21131
rect 7472 21088 7524 21097
rect 10692 21088 10744 21140
rect 13912 21131 13964 21140
rect 13912 21097 13921 21131
rect 13921 21097 13955 21131
rect 13955 21097 13964 21131
rect 13912 21088 13964 21097
rect 18052 21088 18104 21140
rect 20812 21131 20864 21140
rect 20812 21097 20821 21131
rect 20821 21097 20855 21131
rect 20855 21097 20864 21131
rect 20812 21088 20864 21097
rect 20904 21088 20956 21140
rect 22468 21088 22520 21140
rect 22928 21088 22980 21140
rect 23848 21088 23900 21140
rect 25964 21088 26016 21140
rect 26056 21088 26108 21140
rect 33508 21088 33560 21140
rect 33968 21088 34020 21140
rect 35256 21088 35308 21140
rect 35532 21088 35584 21140
rect 39672 21088 39724 21140
rect 43904 21131 43956 21140
rect 43904 21097 43913 21131
rect 43913 21097 43947 21131
rect 43947 21097 43956 21131
rect 43904 21088 43956 21097
rect 46020 21088 46072 21140
rect 46296 21088 46348 21140
rect 46756 21131 46808 21140
rect 46756 21097 46765 21131
rect 46765 21097 46799 21131
rect 46799 21097 46808 21131
rect 46756 21088 46808 21097
rect 11888 21063 11940 21072
rect 11888 21029 11897 21063
rect 11897 21029 11931 21063
rect 11931 21029 11940 21063
rect 11888 21020 11940 21029
rect 18696 21020 18748 21072
rect 23940 21020 23992 21072
rect 26148 21020 26200 21072
rect 29460 21020 29512 21072
rect 33324 21063 33376 21072
rect 33324 21029 33333 21063
rect 33333 21029 33367 21063
rect 33367 21029 33376 21063
rect 33324 21020 33376 21029
rect 34520 21020 34572 21072
rect 3792 20952 3844 21004
rect 7196 20952 7248 21004
rect 11428 20952 11480 21004
rect 12256 20952 12308 21004
rect 17224 20995 17276 21004
rect 17224 20961 17233 20995
rect 17233 20961 17267 20995
rect 17267 20961 17276 20995
rect 17224 20952 17276 20961
rect 17592 20952 17644 21004
rect 18972 20952 19024 21004
rect 2136 20791 2188 20800
rect 2136 20757 2145 20791
rect 2145 20757 2179 20791
rect 2179 20757 2188 20791
rect 2136 20748 2188 20757
rect 4804 20884 4856 20936
rect 8484 20884 8536 20936
rect 10140 20884 10192 20936
rect 10600 20884 10652 20936
rect 5356 20816 5408 20868
rect 10968 20816 11020 20868
rect 2964 20791 3016 20800
rect 2964 20757 2973 20791
rect 2973 20757 3007 20791
rect 3007 20757 3016 20791
rect 2964 20748 3016 20757
rect 3056 20791 3108 20800
rect 3056 20757 3065 20791
rect 3065 20757 3099 20791
rect 3099 20757 3108 20791
rect 3056 20748 3108 20757
rect 3976 20748 4028 20800
rect 6368 20791 6420 20800
rect 6368 20757 6377 20791
rect 6377 20757 6411 20791
rect 6411 20757 6420 20791
rect 6368 20748 6420 20757
rect 11888 20884 11940 20936
rect 12532 20927 12584 20936
rect 12532 20893 12541 20927
rect 12541 20893 12575 20927
rect 12575 20893 12584 20927
rect 12532 20884 12584 20893
rect 12992 20816 13044 20868
rect 15292 20884 15344 20936
rect 17132 20884 17184 20936
rect 14740 20859 14792 20868
rect 14740 20825 14774 20859
rect 14774 20825 14792 20859
rect 14740 20816 14792 20825
rect 15200 20748 15252 20800
rect 15752 20748 15804 20800
rect 15844 20791 15896 20800
rect 15844 20757 15853 20791
rect 15853 20757 15887 20791
rect 15887 20757 15896 20791
rect 15844 20748 15896 20757
rect 16120 20791 16172 20800
rect 16120 20757 16129 20791
rect 16129 20757 16163 20791
rect 16163 20757 16172 20791
rect 16120 20748 16172 20757
rect 17960 20927 18012 20936
rect 17960 20893 17969 20927
rect 17969 20893 18003 20927
rect 18003 20893 18012 20927
rect 17960 20884 18012 20893
rect 18144 20884 18196 20936
rect 18512 20748 18564 20800
rect 19248 20748 19300 20800
rect 20720 20884 20772 20936
rect 20996 20927 21048 20936
rect 20996 20893 21005 20927
rect 21005 20893 21039 20927
rect 21039 20893 21048 20927
rect 20996 20884 21048 20893
rect 22284 20884 22336 20936
rect 24308 20884 24360 20936
rect 24860 20884 24912 20936
rect 26056 20884 26108 20936
rect 24768 20816 24820 20868
rect 31944 20927 31996 20936
rect 31944 20893 31953 20927
rect 31953 20893 31987 20927
rect 31987 20893 31996 20927
rect 31944 20884 31996 20893
rect 32220 20927 32272 20936
rect 32220 20893 32254 20927
rect 32254 20893 32272 20927
rect 32220 20884 32272 20893
rect 33968 20952 34020 21004
rect 34244 20995 34296 21004
rect 34244 20961 34253 20995
rect 34253 20961 34287 20995
rect 34287 20961 34296 20995
rect 34244 20952 34296 20961
rect 34336 20952 34388 21004
rect 36912 20952 36964 21004
rect 42524 20952 42576 21004
rect 42892 20952 42944 21004
rect 20628 20748 20680 20800
rect 23296 20748 23348 20800
rect 33416 20791 33468 20800
rect 33416 20757 33425 20791
rect 33425 20757 33459 20791
rect 33459 20757 33468 20791
rect 33416 20748 33468 20757
rect 34428 20816 34480 20868
rect 37280 20884 37332 20936
rect 38016 20884 38068 20936
rect 38568 20884 38620 20936
rect 40132 20927 40184 20936
rect 40132 20893 40141 20927
rect 40141 20893 40175 20927
rect 40175 20893 40184 20927
rect 40132 20884 40184 20893
rect 43352 20927 43404 20936
rect 43352 20893 43361 20927
rect 43361 20893 43395 20927
rect 43395 20893 43404 20927
rect 43352 20884 43404 20893
rect 44640 20952 44692 21004
rect 45744 20995 45796 21004
rect 45744 20961 45753 20995
rect 45753 20961 45787 20995
rect 45787 20961 45796 20995
rect 45744 20952 45796 20961
rect 34152 20748 34204 20800
rect 40684 20816 40736 20868
rect 42892 20816 42944 20868
rect 43628 20859 43680 20868
rect 43628 20825 43637 20859
rect 43637 20825 43671 20859
rect 43671 20825 43680 20859
rect 43628 20816 43680 20825
rect 46204 20884 46256 20936
rect 44548 20816 44600 20868
rect 45560 20816 45612 20868
rect 36636 20748 36688 20800
rect 41052 20748 41104 20800
rect 42984 20748 43036 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 2964 20544 3016 20596
rect 3884 20544 3936 20596
rect 2136 20476 2188 20528
rect 3976 20519 4028 20528
rect 3976 20485 3985 20519
rect 3985 20485 4019 20519
rect 4019 20485 4028 20519
rect 6920 20544 6972 20596
rect 8300 20519 8352 20528
rect 3976 20476 4028 20485
rect 8300 20485 8334 20519
rect 8334 20485 8352 20519
rect 8300 20476 8352 20485
rect 2504 20408 2556 20460
rect 1676 20383 1728 20392
rect 1676 20349 1685 20383
rect 1685 20349 1719 20383
rect 1719 20349 1728 20383
rect 1676 20340 1728 20349
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 5540 20451 5592 20460
rect 5540 20417 5549 20451
rect 5549 20417 5583 20451
rect 5583 20417 5592 20451
rect 5540 20408 5592 20417
rect 7656 20451 7708 20460
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 8116 20408 8168 20460
rect 9864 20408 9916 20460
rect 4436 20340 4488 20392
rect 3332 20272 3384 20324
rect 4160 20272 4212 20324
rect 1952 20204 2004 20256
rect 3516 20247 3568 20256
rect 3516 20213 3525 20247
rect 3525 20213 3559 20247
rect 3559 20213 3568 20247
rect 3516 20204 3568 20213
rect 4712 20340 4764 20392
rect 5264 20383 5316 20392
rect 5264 20349 5273 20383
rect 5273 20349 5307 20383
rect 5307 20349 5316 20383
rect 5264 20340 5316 20349
rect 5448 20340 5500 20392
rect 5724 20340 5776 20392
rect 7196 20340 7248 20392
rect 11152 20408 11204 20460
rect 12072 20544 12124 20596
rect 12992 20587 13044 20596
rect 12992 20553 13001 20587
rect 13001 20553 13035 20587
rect 13035 20553 13044 20587
rect 12992 20544 13044 20553
rect 11888 20340 11940 20392
rect 12532 20383 12584 20392
rect 12532 20349 12541 20383
rect 12541 20349 12575 20383
rect 12575 20349 12584 20383
rect 12532 20340 12584 20349
rect 12624 20383 12676 20392
rect 12624 20349 12633 20383
rect 12633 20349 12667 20383
rect 12667 20349 12676 20383
rect 12624 20340 12676 20349
rect 13912 20544 13964 20596
rect 14740 20587 14792 20596
rect 14740 20553 14749 20587
rect 14749 20553 14783 20587
rect 14783 20553 14792 20587
rect 14740 20544 14792 20553
rect 13636 20408 13688 20460
rect 15844 20544 15896 20596
rect 18512 20587 18564 20596
rect 18512 20553 18521 20587
rect 18521 20553 18555 20587
rect 18555 20553 18564 20587
rect 18512 20544 18564 20553
rect 15936 20451 15988 20460
rect 15936 20417 15945 20451
rect 15945 20417 15979 20451
rect 15979 20417 15988 20451
rect 15936 20408 15988 20417
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 17684 20408 17736 20460
rect 19984 20408 20036 20460
rect 20260 20476 20312 20528
rect 21272 20476 21324 20528
rect 4712 20204 4764 20256
rect 4896 20204 4948 20256
rect 9220 20272 9272 20324
rect 16212 20340 16264 20392
rect 19064 20340 19116 20392
rect 20444 20451 20496 20460
rect 20444 20417 20453 20451
rect 20453 20417 20487 20451
rect 20487 20417 20496 20451
rect 20444 20408 20496 20417
rect 21456 20408 21508 20460
rect 24400 20408 24452 20460
rect 29736 20451 29788 20460
rect 29736 20417 29745 20451
rect 29745 20417 29779 20451
rect 29779 20417 29788 20451
rect 29736 20408 29788 20417
rect 19248 20315 19300 20324
rect 19248 20281 19257 20315
rect 19257 20281 19291 20315
rect 19291 20281 19300 20315
rect 19248 20272 19300 20281
rect 23296 20272 23348 20324
rect 24308 20272 24360 20324
rect 26240 20272 26292 20324
rect 6184 20247 6236 20256
rect 6184 20213 6193 20247
rect 6193 20213 6227 20247
rect 6227 20213 6236 20247
rect 6184 20204 6236 20213
rect 8300 20204 8352 20256
rect 9312 20204 9364 20256
rect 9404 20247 9456 20256
rect 9404 20213 9413 20247
rect 9413 20213 9447 20247
rect 9447 20213 9456 20247
rect 9404 20204 9456 20213
rect 9956 20247 10008 20256
rect 9956 20213 9965 20247
rect 9965 20213 9999 20247
rect 9999 20213 10008 20247
rect 9956 20204 10008 20213
rect 10508 20204 10560 20256
rect 20720 20204 20772 20256
rect 23388 20247 23440 20256
rect 23388 20213 23397 20247
rect 23397 20213 23431 20247
rect 23431 20213 23440 20247
rect 23388 20204 23440 20213
rect 24676 20204 24728 20256
rect 27896 20204 27948 20256
rect 31668 20544 31720 20596
rect 33692 20544 33744 20596
rect 34336 20544 34388 20596
rect 34704 20544 34756 20596
rect 37464 20544 37516 20596
rect 38384 20544 38436 20596
rect 31392 20408 31444 20460
rect 33600 20408 33652 20460
rect 43444 20544 43496 20596
rect 44548 20544 44600 20596
rect 46664 20587 46716 20596
rect 46664 20553 46673 20587
rect 46673 20553 46707 20587
rect 46707 20553 46716 20587
rect 46664 20544 46716 20553
rect 34520 20451 34572 20460
rect 34520 20417 34554 20451
rect 34554 20417 34572 20451
rect 34520 20408 34572 20417
rect 34704 20451 34756 20460
rect 34704 20417 34713 20451
rect 34713 20417 34747 20451
rect 34747 20417 34756 20451
rect 34704 20408 34756 20417
rect 37464 20408 37516 20460
rect 37924 20408 37976 20460
rect 30012 20383 30064 20392
rect 30012 20349 30021 20383
rect 30021 20349 30055 20383
rect 30055 20349 30064 20383
rect 30012 20340 30064 20349
rect 33140 20340 33192 20392
rect 34428 20383 34480 20392
rect 34428 20349 34437 20383
rect 34437 20349 34471 20383
rect 34471 20349 34480 20383
rect 34428 20340 34480 20349
rect 38660 20340 38712 20392
rect 30472 20204 30524 20256
rect 31852 20204 31904 20256
rect 33968 20272 34020 20324
rect 37924 20272 37976 20324
rect 40684 20408 40736 20460
rect 40960 20408 41012 20460
rect 41328 20451 41380 20460
rect 41328 20417 41337 20451
rect 41337 20417 41371 20451
rect 41371 20417 41380 20451
rect 41328 20408 41380 20417
rect 41420 20451 41472 20460
rect 41420 20417 41429 20451
rect 41429 20417 41463 20451
rect 41463 20417 41472 20451
rect 41420 20408 41472 20417
rect 41604 20408 41656 20460
rect 42340 20408 42392 20460
rect 40224 20340 40276 20392
rect 42708 20451 42760 20460
rect 42708 20417 42717 20451
rect 42717 20417 42751 20451
rect 42751 20417 42760 20451
rect 42708 20408 42760 20417
rect 42984 20451 43036 20460
rect 42984 20417 42993 20451
rect 42993 20417 43027 20451
rect 43027 20417 43036 20451
rect 42984 20408 43036 20417
rect 43536 20451 43588 20460
rect 43536 20417 43545 20451
rect 43545 20417 43579 20451
rect 43579 20417 43588 20451
rect 43536 20408 43588 20417
rect 46204 20451 46256 20460
rect 46204 20417 46213 20451
rect 46213 20417 46247 20451
rect 46247 20417 46256 20451
rect 46204 20408 46256 20417
rect 46480 20451 46532 20460
rect 46480 20417 46489 20451
rect 46489 20417 46523 20451
rect 46523 20417 46532 20451
rect 46480 20408 46532 20417
rect 38844 20272 38896 20324
rect 41604 20272 41656 20324
rect 42340 20272 42392 20324
rect 45284 20383 45336 20392
rect 45284 20349 45293 20383
rect 45293 20349 45327 20383
rect 45327 20349 45336 20383
rect 45284 20340 45336 20349
rect 40040 20204 40092 20256
rect 40868 20247 40920 20256
rect 40868 20213 40877 20247
rect 40877 20213 40911 20247
rect 40911 20213 40920 20247
rect 40868 20204 40920 20213
rect 41512 20204 41564 20256
rect 42432 20247 42484 20256
rect 42432 20213 42441 20247
rect 42441 20213 42475 20247
rect 42475 20213 42484 20247
rect 42432 20204 42484 20213
rect 43168 20247 43220 20256
rect 43168 20213 43177 20247
rect 43177 20213 43211 20247
rect 43211 20213 43220 20247
rect 43168 20204 43220 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2964 20000 3016 20052
rect 5448 20000 5500 20052
rect 6184 20000 6236 20052
rect 12532 20000 12584 20052
rect 17040 20000 17092 20052
rect 4160 19932 4212 19984
rect 4896 19932 4948 19984
rect 5172 19975 5224 19984
rect 5172 19941 5181 19975
rect 5181 19941 5215 19975
rect 5215 19941 5224 19975
rect 5172 19932 5224 19941
rect 6276 19932 6328 19984
rect 3884 19864 3936 19916
rect 5264 19864 5316 19916
rect 5540 19907 5592 19916
rect 5540 19873 5574 19907
rect 5574 19873 5592 19907
rect 5540 19864 5592 19873
rect 6092 19864 6144 19916
rect 6644 19864 6696 19916
rect 6920 19907 6972 19916
rect 6920 19873 6929 19907
rect 6929 19873 6963 19907
rect 6963 19873 6972 19907
rect 6920 19864 6972 19873
rect 10416 19932 10468 19984
rect 15936 19932 15988 19984
rect 24400 20043 24452 20052
rect 24400 20009 24409 20043
rect 24409 20009 24443 20043
rect 24443 20009 24452 20043
rect 24400 20000 24452 20009
rect 24768 20000 24820 20052
rect 13820 19864 13872 19916
rect 14004 19864 14056 19916
rect 26148 19932 26200 19984
rect 26240 19975 26292 19984
rect 26240 19941 26249 19975
rect 26249 19941 26283 19975
rect 26283 19941 26292 19975
rect 26240 19932 26292 19941
rect 28908 19932 28960 19984
rect 29368 19932 29420 19984
rect 29736 20000 29788 20052
rect 31392 20043 31444 20052
rect 31392 20009 31401 20043
rect 31401 20009 31435 20043
rect 31435 20009 31444 20043
rect 31392 20000 31444 20009
rect 34428 20000 34480 20052
rect 36912 20000 36964 20052
rect 38568 20000 38620 20052
rect 41420 20000 41472 20052
rect 41604 20000 41656 20052
rect 42616 20000 42668 20052
rect 42984 20000 43036 20052
rect 43536 20000 43588 20052
rect 45928 20043 45980 20052
rect 45928 20009 45937 20043
rect 45937 20009 45971 20043
rect 45971 20009 45980 20043
rect 45928 20000 45980 20009
rect 46204 20043 46256 20052
rect 46204 20009 46213 20043
rect 46213 20009 46247 20043
rect 46247 20009 46256 20043
rect 46204 20000 46256 20009
rect 18328 19864 18380 19916
rect 18788 19864 18840 19916
rect 19892 19864 19944 19916
rect 21180 19864 21232 19916
rect 22836 19907 22888 19916
rect 22836 19873 22845 19907
rect 22845 19873 22879 19907
rect 22879 19873 22888 19907
rect 22836 19864 22888 19873
rect 24676 19864 24728 19916
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 1952 19839 2004 19848
rect 1952 19805 1986 19839
rect 1986 19805 2004 19839
rect 1952 19796 2004 19805
rect 3516 19796 3568 19848
rect 4528 19839 4580 19848
rect 4528 19805 4537 19839
rect 4537 19805 4571 19839
rect 4571 19805 4580 19839
rect 4528 19796 4580 19805
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 6368 19796 6420 19848
rect 8484 19839 8536 19848
rect 8484 19805 8493 19839
rect 8493 19805 8527 19839
rect 8527 19805 8536 19839
rect 8484 19796 8536 19805
rect 11612 19796 11664 19848
rect 15660 19796 15712 19848
rect 17316 19796 17368 19848
rect 18512 19796 18564 19848
rect 20076 19839 20128 19848
rect 20076 19805 20085 19839
rect 20085 19805 20119 19839
rect 20119 19805 20128 19839
rect 20076 19796 20128 19805
rect 3976 19703 4028 19712
rect 3976 19669 3985 19703
rect 3985 19669 4019 19703
rect 4019 19669 4028 19703
rect 3976 19660 4028 19669
rect 6644 19728 6696 19780
rect 11704 19728 11756 19780
rect 11980 19728 12032 19780
rect 12900 19771 12952 19780
rect 12900 19737 12909 19771
rect 12909 19737 12943 19771
rect 12943 19737 12952 19771
rect 12900 19728 12952 19737
rect 15200 19728 15252 19780
rect 19064 19728 19116 19780
rect 20720 19796 20772 19848
rect 23388 19796 23440 19848
rect 23480 19796 23532 19848
rect 24768 19796 24820 19848
rect 26332 19864 26384 19916
rect 29000 19864 29052 19916
rect 29092 19864 29144 19916
rect 30564 19864 30616 19916
rect 31116 19932 31168 19984
rect 37740 19932 37792 19984
rect 31024 19864 31076 19916
rect 32036 19907 32088 19916
rect 32036 19873 32045 19907
rect 32045 19873 32079 19907
rect 32079 19873 32088 19907
rect 32036 19864 32088 19873
rect 25596 19839 25648 19848
rect 25596 19805 25605 19839
rect 25605 19805 25639 19839
rect 25639 19805 25648 19839
rect 25596 19796 25648 19805
rect 25688 19796 25740 19848
rect 6368 19703 6420 19712
rect 6368 19669 6377 19703
rect 6377 19669 6411 19703
rect 6411 19669 6420 19703
rect 6368 19660 6420 19669
rect 6460 19703 6512 19712
rect 6460 19669 6469 19703
rect 6469 19669 6503 19703
rect 6503 19669 6512 19703
rect 6460 19660 6512 19669
rect 9864 19660 9916 19712
rect 10508 19660 10560 19712
rect 15384 19660 15436 19712
rect 17960 19660 18012 19712
rect 20996 19728 21048 19780
rect 24676 19728 24728 19780
rect 19984 19660 20036 19712
rect 20720 19660 20772 19712
rect 21180 19703 21232 19712
rect 21180 19669 21189 19703
rect 21189 19669 21223 19703
rect 21223 19669 21232 19703
rect 21180 19660 21232 19669
rect 23020 19660 23072 19712
rect 26516 19839 26568 19848
rect 26516 19805 26525 19839
rect 26525 19805 26559 19839
rect 26559 19805 26568 19839
rect 26516 19796 26568 19805
rect 26792 19839 26844 19848
rect 26792 19805 26801 19839
rect 26801 19805 26835 19839
rect 26835 19805 26844 19839
rect 26792 19796 26844 19805
rect 28540 19796 28592 19848
rect 31852 19796 31904 19848
rect 31944 19796 31996 19848
rect 33416 19839 33468 19848
rect 33416 19805 33450 19839
rect 33450 19805 33468 19839
rect 33416 19796 33468 19805
rect 37556 19839 37608 19848
rect 37556 19805 37565 19839
rect 37565 19805 37599 19839
rect 37599 19805 37608 19839
rect 37556 19796 37608 19805
rect 40868 19864 40920 19916
rect 37832 19839 37884 19848
rect 37832 19805 37841 19839
rect 37841 19805 37875 19839
rect 37875 19805 37884 19839
rect 37832 19796 37884 19805
rect 37924 19839 37976 19848
rect 37924 19805 37938 19839
rect 37938 19805 37972 19839
rect 37972 19805 37976 19839
rect 37924 19796 37976 19805
rect 38752 19796 38804 19848
rect 41512 19839 41564 19848
rect 41512 19805 41521 19839
rect 41521 19805 41555 19839
rect 41555 19805 41564 19839
rect 41512 19796 41564 19805
rect 42432 19796 42484 19848
rect 43352 19796 43404 19848
rect 44548 19839 44600 19848
rect 44548 19805 44557 19839
rect 44557 19805 44591 19839
rect 44591 19805 44600 19839
rect 44548 19796 44600 19805
rect 44640 19839 44692 19848
rect 44640 19805 44649 19839
rect 44649 19805 44683 19839
rect 44683 19805 44692 19839
rect 44640 19796 44692 19805
rect 45560 19796 45612 19848
rect 28632 19728 28684 19780
rect 29368 19728 29420 19780
rect 42800 19771 42852 19780
rect 42800 19737 42809 19771
rect 42809 19737 42843 19771
rect 42843 19737 42852 19771
rect 42800 19728 42852 19737
rect 27436 19703 27488 19712
rect 27436 19669 27445 19703
rect 27445 19669 27479 19703
rect 27479 19669 27488 19703
rect 27436 19660 27488 19669
rect 27896 19703 27948 19712
rect 27896 19669 27905 19703
rect 27905 19669 27939 19703
rect 27939 19669 27948 19703
rect 27896 19660 27948 19669
rect 29276 19703 29328 19712
rect 29276 19669 29285 19703
rect 29285 19669 29319 19703
rect 29319 19669 29328 19703
rect 29276 19660 29328 19669
rect 32496 19660 32548 19712
rect 37832 19660 37884 19712
rect 44180 19703 44232 19712
rect 44180 19669 44189 19703
rect 44189 19669 44223 19703
rect 44223 19669 44232 19703
rect 44180 19660 44232 19669
rect 44364 19660 44416 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 1308 19456 1360 19508
rect 2504 19456 2556 19508
rect 2964 19499 3016 19508
rect 2964 19465 2973 19499
rect 2973 19465 3007 19499
rect 3007 19465 3016 19499
rect 2964 19456 3016 19465
rect 3056 19499 3108 19508
rect 3056 19465 3065 19499
rect 3065 19465 3099 19499
rect 3099 19465 3108 19499
rect 3056 19456 3108 19465
rect 4528 19456 4580 19508
rect 5356 19499 5408 19508
rect 5356 19465 5365 19499
rect 5365 19465 5399 19499
rect 5399 19465 5408 19499
rect 5356 19456 5408 19465
rect 3332 19388 3384 19440
rect 3976 19388 4028 19440
rect 4068 19388 4120 19440
rect 8300 19456 8352 19508
rect 10508 19499 10560 19508
rect 10508 19465 10517 19499
rect 10517 19465 10551 19499
rect 10551 19465 10560 19499
rect 10508 19456 10560 19465
rect 11704 19499 11756 19508
rect 11704 19465 11713 19499
rect 11713 19465 11747 19499
rect 11747 19465 11756 19499
rect 11704 19456 11756 19465
rect 6368 19388 6420 19440
rect 15200 19388 15252 19440
rect 17684 19456 17736 19508
rect 20076 19456 20128 19508
rect 24124 19456 24176 19508
rect 23296 19388 23348 19440
rect 1676 19320 1728 19372
rect 4160 19320 4212 19372
rect 4804 19320 4856 19372
rect 5356 19320 5408 19372
rect 6460 19320 6512 19372
rect 9404 19320 9456 19372
rect 11428 19320 11480 19372
rect 3240 19295 3292 19304
rect 3240 19261 3249 19295
rect 3249 19261 3283 19295
rect 3283 19261 3292 19295
rect 3240 19252 3292 19261
rect 13084 19363 13136 19372
rect 13084 19329 13093 19363
rect 13093 19329 13127 19363
rect 13127 19329 13136 19363
rect 13084 19320 13136 19329
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 15752 19320 15804 19329
rect 15844 19363 15896 19372
rect 15844 19329 15853 19363
rect 15853 19329 15887 19363
rect 15887 19329 15896 19363
rect 15844 19320 15896 19329
rect 15568 19252 15620 19304
rect 18236 19320 18288 19372
rect 23480 19320 23532 19372
rect 26792 19320 26844 19372
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27160 19320 27212 19329
rect 19984 19252 20036 19304
rect 11704 19184 11756 19236
rect 12808 19116 12860 19168
rect 14832 19184 14884 19236
rect 19064 19184 19116 19236
rect 22928 19295 22980 19304
rect 22928 19261 22937 19295
rect 22937 19261 22971 19295
rect 22971 19261 22980 19295
rect 22928 19252 22980 19261
rect 23020 19252 23072 19304
rect 23296 19295 23348 19304
rect 23296 19261 23305 19295
rect 23305 19261 23339 19295
rect 23339 19261 23348 19295
rect 23296 19252 23348 19261
rect 23204 19184 23256 19236
rect 23664 19184 23716 19236
rect 16028 19116 16080 19168
rect 21180 19116 21232 19168
rect 21456 19116 21508 19168
rect 22100 19116 22152 19168
rect 24032 19295 24084 19304
rect 24032 19261 24041 19295
rect 24041 19261 24075 19295
rect 24075 19261 24084 19295
rect 24032 19252 24084 19261
rect 24124 19295 24176 19304
rect 24124 19261 24158 19295
rect 24158 19261 24176 19295
rect 24124 19252 24176 19261
rect 24676 19252 24728 19304
rect 28632 19227 28684 19236
rect 28632 19193 28641 19227
rect 28641 19193 28675 19227
rect 28675 19193 28684 19227
rect 28632 19184 28684 19193
rect 28908 19363 28960 19372
rect 28908 19329 28917 19363
rect 28917 19329 28951 19363
rect 28951 19329 28960 19363
rect 28908 19320 28960 19329
rect 29276 19456 29328 19508
rect 34060 19456 34112 19508
rect 35992 19456 36044 19508
rect 36360 19456 36412 19508
rect 37556 19456 37608 19508
rect 38752 19456 38804 19508
rect 29276 19363 29328 19372
rect 29276 19329 29310 19363
rect 29310 19329 29328 19363
rect 29276 19320 29328 19329
rect 30196 19320 30248 19372
rect 30840 19320 30892 19372
rect 31300 19320 31352 19372
rect 31668 19320 31720 19372
rect 30472 19295 30524 19304
rect 30472 19261 30481 19295
rect 30481 19261 30515 19295
rect 30515 19261 30524 19295
rect 30472 19252 30524 19261
rect 31576 19295 31628 19304
rect 31576 19261 31585 19295
rect 31585 19261 31619 19295
rect 31619 19261 31628 19295
rect 31576 19252 31628 19261
rect 31852 19252 31904 19304
rect 33508 19295 33560 19304
rect 33508 19261 33517 19295
rect 33517 19261 33551 19295
rect 33551 19261 33560 19295
rect 33508 19252 33560 19261
rect 31024 19227 31076 19236
rect 31024 19193 31033 19227
rect 31033 19193 31067 19227
rect 31067 19193 31076 19227
rect 31024 19184 31076 19193
rect 24216 19116 24268 19168
rect 24860 19116 24912 19168
rect 25596 19116 25648 19168
rect 27620 19116 27672 19168
rect 28172 19116 28224 19168
rect 29644 19116 29696 19168
rect 30564 19116 30616 19168
rect 35992 19320 36044 19372
rect 33692 19295 33744 19304
rect 33692 19261 33701 19295
rect 33701 19261 33735 19295
rect 33735 19261 33744 19295
rect 33692 19252 33744 19261
rect 33876 19252 33928 19304
rect 34244 19252 34296 19304
rect 34520 19295 34572 19304
rect 34520 19261 34554 19295
rect 34554 19261 34572 19295
rect 34520 19252 34572 19261
rect 34888 19252 34940 19304
rect 37832 19363 37884 19372
rect 37832 19329 37841 19363
rect 37841 19329 37875 19363
rect 37875 19329 37884 19363
rect 37832 19320 37884 19329
rect 38384 19363 38436 19372
rect 38384 19329 38393 19363
rect 38393 19329 38427 19363
rect 38427 19329 38436 19363
rect 38384 19320 38436 19329
rect 38752 19320 38804 19372
rect 43812 19456 43864 19508
rect 44180 19456 44232 19508
rect 38568 19295 38620 19304
rect 38568 19261 38577 19295
rect 38577 19261 38611 19295
rect 38611 19261 38620 19295
rect 38568 19252 38620 19261
rect 40500 19363 40552 19372
rect 40500 19329 40509 19363
rect 40509 19329 40543 19363
rect 40543 19329 40552 19363
rect 40500 19320 40552 19329
rect 40592 19320 40644 19372
rect 42800 19388 42852 19440
rect 41328 19252 41380 19304
rect 43352 19320 43404 19372
rect 44272 19363 44324 19372
rect 44272 19329 44281 19363
rect 44281 19329 44315 19363
rect 44315 19329 44324 19363
rect 44272 19320 44324 19329
rect 37832 19184 37884 19236
rect 35716 19159 35768 19168
rect 35716 19125 35725 19159
rect 35725 19125 35759 19159
rect 35759 19125 35768 19159
rect 35716 19116 35768 19125
rect 40592 19227 40644 19236
rect 40592 19193 40601 19227
rect 40601 19193 40635 19227
rect 40635 19193 40644 19227
rect 40592 19184 40644 19193
rect 41420 19184 41472 19236
rect 42340 19252 42392 19304
rect 44364 19295 44416 19304
rect 44364 19261 44373 19295
rect 44373 19261 44407 19295
rect 44407 19261 44416 19295
rect 44364 19252 44416 19261
rect 45284 19252 45336 19304
rect 39212 19116 39264 19168
rect 42800 19116 42852 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3240 18912 3292 18964
rect 3976 18912 4028 18964
rect 10324 18887 10376 18896
rect 10324 18853 10333 18887
rect 10333 18853 10367 18887
rect 10367 18853 10376 18887
rect 10324 18844 10376 18853
rect 11152 18887 11204 18896
rect 11152 18853 11161 18887
rect 11161 18853 11195 18887
rect 11195 18853 11204 18887
rect 11152 18844 11204 18853
rect 11244 18776 11296 18828
rect 11704 18819 11756 18828
rect 11704 18785 11713 18819
rect 11713 18785 11747 18819
rect 11747 18785 11756 18819
rect 11704 18776 11756 18785
rect 14464 18776 14516 18828
rect 14832 18819 14884 18828
rect 14832 18785 14841 18819
rect 14841 18785 14875 18819
rect 14875 18785 14884 18819
rect 14832 18776 14884 18785
rect 15108 18776 15160 18828
rect 6920 18751 6972 18760
rect 6920 18717 6929 18751
rect 6929 18717 6963 18751
rect 6963 18717 6972 18751
rect 6920 18708 6972 18717
rect 8208 18708 8260 18760
rect 10324 18708 10376 18760
rect 10692 18751 10744 18760
rect 10692 18717 10701 18751
rect 10701 18717 10735 18751
rect 10735 18717 10744 18751
rect 10692 18708 10744 18717
rect 11520 18751 11572 18760
rect 11520 18717 11554 18751
rect 11554 18717 11572 18751
rect 11520 18708 11572 18717
rect 12532 18751 12584 18760
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 12808 18751 12860 18760
rect 12808 18717 12842 18751
rect 12842 18717 12860 18751
rect 12808 18708 12860 18717
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 14740 18708 14792 18760
rect 15936 18708 15988 18760
rect 16028 18751 16080 18760
rect 16028 18717 16037 18751
rect 16037 18717 16071 18751
rect 16071 18717 16080 18751
rect 16028 18708 16080 18717
rect 16764 18844 16816 18896
rect 17316 18844 17368 18896
rect 19064 18887 19116 18896
rect 19064 18853 19073 18887
rect 19073 18853 19107 18887
rect 19107 18853 19116 18887
rect 19064 18844 19116 18853
rect 16672 18776 16724 18828
rect 17684 18819 17736 18828
rect 17684 18785 17693 18819
rect 17693 18785 17727 18819
rect 17727 18785 17736 18819
rect 17684 18776 17736 18785
rect 6644 18640 6696 18692
rect 8576 18640 8628 18692
rect 8392 18572 8444 18624
rect 11336 18572 11388 18624
rect 13912 18615 13964 18624
rect 13912 18581 13921 18615
rect 13921 18581 13955 18615
rect 13955 18581 13964 18615
rect 13912 18572 13964 18581
rect 14096 18615 14148 18624
rect 14096 18581 14105 18615
rect 14105 18581 14139 18615
rect 14139 18581 14148 18615
rect 14096 18572 14148 18581
rect 17316 18683 17368 18692
rect 17316 18649 17325 18683
rect 17325 18649 17359 18683
rect 17359 18649 17368 18683
rect 17316 18640 17368 18649
rect 19064 18708 19116 18760
rect 19800 18819 19852 18828
rect 19800 18785 19809 18819
rect 19809 18785 19843 18819
rect 19843 18785 19852 18819
rect 19800 18776 19852 18785
rect 20352 18912 20404 18964
rect 21088 18844 21140 18896
rect 21180 18844 21232 18896
rect 20260 18751 20312 18760
rect 20260 18717 20269 18751
rect 20269 18717 20303 18751
rect 20303 18717 20312 18751
rect 20260 18708 20312 18717
rect 20444 18708 20496 18760
rect 20996 18776 21048 18828
rect 24124 18912 24176 18964
rect 24216 18912 24268 18964
rect 27160 18912 27212 18964
rect 29276 18912 29328 18964
rect 30104 18912 30156 18964
rect 30288 18912 30340 18964
rect 37648 18912 37700 18964
rect 38660 18912 38712 18964
rect 41328 18955 41380 18964
rect 41328 18921 41337 18955
rect 41337 18921 41371 18955
rect 41371 18921 41380 18955
rect 41328 18912 41380 18921
rect 38752 18844 38804 18896
rect 21916 18819 21968 18828
rect 21916 18785 21925 18819
rect 21925 18785 21959 18819
rect 21959 18785 21968 18819
rect 21916 18776 21968 18785
rect 23664 18776 23716 18828
rect 24308 18776 24360 18828
rect 24860 18819 24912 18828
rect 24860 18785 24869 18819
rect 24869 18785 24903 18819
rect 24903 18785 24912 18819
rect 24860 18776 24912 18785
rect 21640 18751 21692 18760
rect 21640 18717 21649 18751
rect 21649 18717 21683 18751
rect 21683 18717 21692 18751
rect 21640 18708 21692 18717
rect 22560 18708 22612 18760
rect 22744 18708 22796 18760
rect 25596 18776 25648 18828
rect 25688 18819 25740 18828
rect 25688 18785 25697 18819
rect 25697 18785 25731 18819
rect 25731 18785 25740 18819
rect 25688 18776 25740 18785
rect 25872 18776 25924 18828
rect 26424 18819 26476 18828
rect 26424 18785 26433 18819
rect 26433 18785 26467 18819
rect 26467 18785 26476 18819
rect 26424 18776 26476 18785
rect 27344 18819 27396 18828
rect 27344 18785 27353 18819
rect 27353 18785 27387 18819
rect 27387 18785 27396 18819
rect 27344 18776 27396 18785
rect 27896 18819 27948 18828
rect 27896 18785 27905 18819
rect 27905 18785 27939 18819
rect 27939 18785 27948 18819
rect 27896 18776 27948 18785
rect 28172 18776 28224 18828
rect 26608 18708 26660 18760
rect 26700 18751 26752 18760
rect 26700 18717 26709 18751
rect 26709 18717 26743 18751
rect 26743 18717 26752 18751
rect 26700 18708 26752 18717
rect 27620 18708 27672 18760
rect 31576 18776 31628 18828
rect 40408 18776 40460 18828
rect 41420 18819 41472 18828
rect 41420 18785 41429 18819
rect 41429 18785 41463 18819
rect 41463 18785 41472 18819
rect 41420 18776 41472 18785
rect 41788 18776 41840 18828
rect 44272 18776 44324 18828
rect 17684 18640 17736 18692
rect 18696 18640 18748 18692
rect 20352 18640 20404 18692
rect 22468 18640 22520 18692
rect 19248 18615 19300 18624
rect 19248 18581 19257 18615
rect 19257 18581 19291 18615
rect 19291 18581 19300 18615
rect 19248 18572 19300 18581
rect 19708 18615 19760 18624
rect 19708 18581 19717 18615
rect 19717 18581 19751 18615
rect 19751 18581 19760 18615
rect 19708 18572 19760 18581
rect 20444 18615 20496 18624
rect 20444 18581 20453 18615
rect 20453 18581 20487 18615
rect 20487 18581 20496 18615
rect 20444 18572 20496 18581
rect 24952 18640 25004 18692
rect 27528 18640 27580 18692
rect 28448 18640 28500 18692
rect 23480 18572 23532 18624
rect 27436 18572 27488 18624
rect 29736 18708 29788 18760
rect 30012 18751 30064 18760
rect 30012 18717 30021 18751
rect 30021 18717 30055 18751
rect 30055 18717 30064 18751
rect 30012 18708 30064 18717
rect 31760 18751 31812 18760
rect 31760 18717 31769 18751
rect 31769 18717 31803 18751
rect 31803 18717 31812 18751
rect 31760 18708 31812 18717
rect 33784 18708 33836 18760
rect 30564 18640 30616 18692
rect 32496 18640 32548 18692
rect 34152 18708 34204 18760
rect 34336 18708 34388 18760
rect 35716 18751 35768 18760
rect 35716 18717 35750 18751
rect 35750 18717 35768 18751
rect 35716 18708 35768 18717
rect 36820 18708 36872 18760
rect 38108 18708 38160 18760
rect 38384 18751 38436 18760
rect 38384 18717 38393 18751
rect 38393 18717 38427 18751
rect 38427 18717 38436 18751
rect 38384 18708 38436 18717
rect 38660 18708 38712 18760
rect 40040 18751 40092 18760
rect 40040 18717 40049 18751
rect 40049 18717 40083 18751
rect 40083 18717 40092 18751
rect 40040 18708 40092 18717
rect 36636 18640 36688 18692
rect 37832 18640 37884 18692
rect 39120 18640 39172 18692
rect 40500 18751 40552 18760
rect 40500 18717 40509 18751
rect 40509 18717 40543 18751
rect 40543 18717 40552 18751
rect 40500 18708 40552 18717
rect 40592 18708 40644 18760
rect 41144 18708 41196 18760
rect 42064 18708 42116 18760
rect 44548 18751 44600 18760
rect 44548 18717 44557 18751
rect 44557 18717 44591 18751
rect 44591 18717 44600 18751
rect 44548 18708 44600 18717
rect 44732 18751 44784 18760
rect 44732 18717 44741 18751
rect 44741 18717 44775 18751
rect 44775 18717 44784 18751
rect 44732 18708 44784 18717
rect 46112 18751 46164 18760
rect 46112 18717 46121 18751
rect 46121 18717 46155 18751
rect 46155 18717 46164 18751
rect 46112 18708 46164 18717
rect 32588 18572 32640 18624
rect 36084 18572 36136 18624
rect 37924 18572 37976 18624
rect 40592 18572 40644 18624
rect 44272 18640 44324 18692
rect 44640 18640 44692 18692
rect 41512 18572 41564 18624
rect 44824 18615 44876 18624
rect 44824 18581 44833 18615
rect 44833 18581 44867 18615
rect 44867 18581 44876 18615
rect 44824 18572 44876 18581
rect 45836 18572 45888 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 2964 18300 3016 18352
rect 3424 18300 3476 18352
rect 6644 18411 6696 18420
rect 6644 18377 6653 18411
rect 6653 18377 6687 18411
rect 6687 18377 6696 18411
rect 6644 18368 6696 18377
rect 8300 18411 8352 18420
rect 8300 18377 8309 18411
rect 8309 18377 8343 18411
rect 8343 18377 8352 18411
rect 8300 18368 8352 18377
rect 11244 18368 11296 18420
rect 14556 18368 14608 18420
rect 15568 18368 15620 18420
rect 15752 18368 15804 18420
rect 18328 18411 18380 18420
rect 18328 18377 18337 18411
rect 18337 18377 18371 18411
rect 18371 18377 18380 18411
rect 18328 18368 18380 18377
rect 18696 18411 18748 18420
rect 18696 18377 18705 18411
rect 18705 18377 18739 18411
rect 18739 18377 18748 18411
rect 18696 18368 18748 18377
rect 20260 18368 20312 18420
rect 22468 18368 22520 18420
rect 9680 18300 9732 18352
rect 10416 18300 10468 18352
rect 1400 18232 1452 18284
rect 3056 18275 3108 18284
rect 3056 18241 3065 18275
rect 3065 18241 3099 18275
rect 3099 18241 3108 18275
rect 3056 18232 3108 18241
rect 3884 18232 3936 18284
rect 2228 18207 2280 18216
rect 2228 18173 2237 18207
rect 2237 18173 2271 18207
rect 2271 18173 2280 18207
rect 2228 18164 2280 18173
rect 3608 18164 3660 18216
rect 4436 18207 4488 18216
rect 4436 18173 4445 18207
rect 4445 18173 4479 18207
rect 4479 18173 4488 18207
rect 4436 18164 4488 18173
rect 3332 18096 3384 18148
rect 7564 18232 7616 18284
rect 8208 18232 8260 18284
rect 6920 18207 6972 18216
rect 6920 18173 6929 18207
rect 6929 18173 6963 18207
rect 6963 18173 6972 18207
rect 6920 18164 6972 18173
rect 9404 18164 9456 18216
rect 9772 18164 9824 18216
rect 4620 18028 4672 18080
rect 5448 18028 5500 18080
rect 9680 18139 9732 18148
rect 9680 18105 9689 18139
rect 9689 18105 9723 18139
rect 9723 18105 9732 18139
rect 9680 18096 9732 18105
rect 14096 18300 14148 18352
rect 7288 18028 7340 18080
rect 10692 18028 10744 18080
rect 11980 18207 12032 18216
rect 11980 18173 11989 18207
rect 11989 18173 12023 18207
rect 12023 18173 12032 18207
rect 11980 18164 12032 18173
rect 12532 18232 12584 18284
rect 13820 18232 13872 18284
rect 13912 18232 13964 18284
rect 14464 18164 14516 18216
rect 14740 18207 14792 18216
rect 14740 18173 14749 18207
rect 14749 18173 14783 18207
rect 14783 18173 14792 18207
rect 14740 18164 14792 18173
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 15108 18164 15160 18216
rect 15568 18164 15620 18216
rect 15936 18164 15988 18216
rect 16120 18164 16172 18216
rect 15292 18096 15344 18148
rect 16304 18096 16356 18148
rect 16672 18207 16724 18216
rect 16672 18173 16681 18207
rect 16681 18173 16715 18207
rect 16715 18173 16724 18207
rect 16672 18164 16724 18173
rect 19248 18232 19300 18284
rect 21640 18300 21692 18352
rect 24952 18368 25004 18420
rect 29368 18368 29420 18420
rect 22008 18232 22060 18284
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 23020 18275 23072 18284
rect 23020 18241 23029 18275
rect 23029 18241 23063 18275
rect 23063 18241 23072 18275
rect 23020 18232 23072 18241
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 24124 18232 24176 18284
rect 30012 18368 30064 18420
rect 31116 18411 31168 18420
rect 31116 18377 31125 18411
rect 31125 18377 31159 18411
rect 31159 18377 31168 18411
rect 31116 18368 31168 18377
rect 31760 18368 31812 18420
rect 32496 18411 32548 18420
rect 32496 18377 32505 18411
rect 32505 18377 32539 18411
rect 32539 18377 32548 18411
rect 32496 18368 32548 18377
rect 32588 18411 32640 18420
rect 32588 18377 32597 18411
rect 32597 18377 32631 18411
rect 32631 18377 32640 18411
rect 32588 18368 32640 18377
rect 33692 18368 33744 18420
rect 35256 18368 35308 18420
rect 35532 18368 35584 18420
rect 35992 18368 36044 18420
rect 36176 18411 36228 18420
rect 36176 18377 36185 18411
rect 36185 18377 36219 18411
rect 36219 18377 36228 18411
rect 36176 18368 36228 18377
rect 36636 18411 36688 18420
rect 36636 18377 36645 18411
rect 36645 18377 36679 18411
rect 36679 18377 36688 18411
rect 36636 18368 36688 18377
rect 36084 18343 36136 18352
rect 36084 18309 36093 18343
rect 36093 18309 36127 18343
rect 36127 18309 36136 18343
rect 36084 18300 36136 18309
rect 30472 18275 30524 18284
rect 30472 18241 30481 18275
rect 30481 18241 30515 18275
rect 30515 18241 30524 18275
rect 30472 18232 30524 18241
rect 33692 18275 33744 18284
rect 33692 18241 33701 18275
rect 33701 18241 33735 18275
rect 33735 18241 33744 18275
rect 33692 18232 33744 18241
rect 34520 18275 34572 18284
rect 34520 18241 34554 18275
rect 34554 18241 34572 18275
rect 34520 18232 34572 18241
rect 37648 18411 37700 18420
rect 37648 18377 37657 18411
rect 37657 18377 37691 18411
rect 37691 18377 37700 18411
rect 37648 18368 37700 18377
rect 40040 18368 40092 18420
rect 40776 18368 40828 18420
rect 44732 18368 44784 18420
rect 40316 18300 40368 18352
rect 39120 18232 39172 18284
rect 40132 18232 40184 18284
rect 19156 18164 19208 18216
rect 19984 18207 20036 18216
rect 19984 18173 19993 18207
rect 19993 18173 20027 18207
rect 20027 18173 20036 18207
rect 19984 18164 20036 18173
rect 22744 18164 22796 18216
rect 23296 18164 23348 18216
rect 17684 18096 17736 18148
rect 17316 18028 17368 18080
rect 18880 18096 18932 18148
rect 19800 18096 19852 18148
rect 22284 18096 22336 18148
rect 22468 18096 22520 18148
rect 25504 18164 25556 18216
rect 26700 18164 26752 18216
rect 29828 18164 29880 18216
rect 24676 18096 24728 18148
rect 26240 18096 26292 18148
rect 26884 18096 26936 18148
rect 29460 18096 29512 18148
rect 25872 18028 25924 18080
rect 26148 18028 26200 18080
rect 29092 18028 29144 18080
rect 29736 18028 29788 18080
rect 30288 18207 30340 18216
rect 30288 18173 30322 18207
rect 30322 18173 30340 18207
rect 30288 18164 30340 18173
rect 33508 18207 33560 18216
rect 33508 18173 33517 18207
rect 33517 18173 33551 18207
rect 33551 18173 33560 18207
rect 33508 18164 33560 18173
rect 33876 18164 33928 18216
rect 34244 18164 34296 18216
rect 35440 18164 35492 18216
rect 36176 18164 36228 18216
rect 36268 18207 36320 18216
rect 36268 18173 36277 18207
rect 36277 18173 36311 18207
rect 36311 18173 36320 18207
rect 36268 18164 36320 18173
rect 37740 18207 37792 18216
rect 37740 18173 37749 18207
rect 37749 18173 37783 18207
rect 37783 18173 37792 18207
rect 37740 18164 37792 18173
rect 30564 18028 30616 18080
rect 30656 18028 30708 18080
rect 33140 18096 33192 18148
rect 33324 18096 33376 18148
rect 40500 18164 40552 18216
rect 34060 18028 34112 18080
rect 41144 18207 41196 18216
rect 41144 18173 41153 18207
rect 41153 18173 41187 18207
rect 41187 18173 41196 18207
rect 41144 18164 41196 18173
rect 41420 18232 41472 18284
rect 43812 18275 43864 18284
rect 43812 18241 43821 18275
rect 43821 18241 43855 18275
rect 43855 18241 43864 18275
rect 43812 18232 43864 18241
rect 44180 18232 44232 18284
rect 45008 18275 45060 18284
rect 45008 18241 45017 18275
rect 45017 18241 45051 18275
rect 45051 18241 45060 18275
rect 45008 18232 45060 18241
rect 45836 18275 45888 18284
rect 45836 18241 45845 18275
rect 45845 18241 45879 18275
rect 45879 18241 45888 18275
rect 45836 18232 45888 18241
rect 41512 18164 41564 18216
rect 41696 18207 41748 18216
rect 41696 18173 41705 18207
rect 41705 18173 41739 18207
rect 41739 18173 41748 18207
rect 41696 18164 41748 18173
rect 42064 18207 42116 18216
rect 42064 18173 42073 18207
rect 42073 18173 42107 18207
rect 42107 18173 42116 18207
rect 42064 18164 42116 18173
rect 44364 18164 44416 18216
rect 44824 18164 44876 18216
rect 41788 18096 41840 18148
rect 41236 18028 41288 18080
rect 41696 18028 41748 18080
rect 43812 18028 43864 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2964 17867 3016 17876
rect 2964 17833 2973 17867
rect 2973 17833 3007 17867
rect 3007 17833 3016 17867
rect 2964 17824 3016 17833
rect 3884 17867 3936 17876
rect 3884 17833 3893 17867
rect 3893 17833 3927 17867
rect 3927 17833 3936 17867
rect 3884 17824 3936 17833
rect 4712 17824 4764 17876
rect 5816 17824 5868 17876
rect 7564 17867 7616 17876
rect 7564 17833 7573 17867
rect 7573 17833 7607 17867
rect 7607 17833 7616 17867
rect 7564 17824 7616 17833
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 8760 17824 8812 17876
rect 13084 17867 13136 17876
rect 13084 17833 13093 17867
rect 13093 17833 13127 17867
rect 13127 17833 13136 17867
rect 13084 17824 13136 17833
rect 16304 17867 16356 17876
rect 16304 17833 16313 17867
rect 16313 17833 16347 17867
rect 16347 17833 16356 17867
rect 16304 17824 16356 17833
rect 4252 17688 4304 17740
rect 4528 17688 4580 17740
rect 4712 17688 4764 17740
rect 4804 17731 4856 17740
rect 4804 17697 4813 17731
rect 4813 17697 4847 17731
rect 4847 17697 4856 17731
rect 4804 17688 4856 17697
rect 3332 17663 3384 17672
rect 3332 17629 3341 17663
rect 3341 17629 3375 17663
rect 3375 17629 3384 17663
rect 3332 17620 3384 17629
rect 4160 17663 4212 17672
rect 4160 17629 4169 17663
rect 4169 17629 4203 17663
rect 4203 17629 4212 17663
rect 4160 17620 4212 17629
rect 5264 17620 5316 17672
rect 11060 17756 11112 17808
rect 7196 17688 7248 17740
rect 8576 17688 8628 17740
rect 9496 17731 9548 17740
rect 9496 17697 9505 17731
rect 9505 17697 9539 17731
rect 9539 17697 9548 17731
rect 9496 17688 9548 17697
rect 10692 17688 10744 17740
rect 10968 17731 11020 17740
rect 10968 17697 10977 17731
rect 10977 17697 11011 17731
rect 11011 17697 11020 17731
rect 10968 17688 11020 17697
rect 6092 17620 6144 17672
rect 7012 17663 7064 17672
rect 7012 17629 7021 17663
rect 7021 17629 7055 17663
rect 7055 17629 7064 17663
rect 7012 17620 7064 17629
rect 7472 17620 7524 17672
rect 8392 17620 8444 17672
rect 8760 17663 8812 17672
rect 8760 17629 8769 17663
rect 8769 17629 8803 17663
rect 8803 17629 8812 17663
rect 8760 17620 8812 17629
rect 10324 17663 10376 17672
rect 10324 17629 10333 17663
rect 10333 17629 10367 17663
rect 10367 17629 10376 17663
rect 10324 17620 10376 17629
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 11336 17663 11388 17672
rect 11336 17629 11370 17663
rect 11370 17629 11388 17663
rect 11336 17620 11388 17629
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 15844 17756 15896 17808
rect 13636 17731 13688 17740
rect 13636 17697 13645 17731
rect 13645 17697 13679 17731
rect 13679 17697 13688 17731
rect 13636 17688 13688 17697
rect 13820 17688 13872 17740
rect 14464 17688 14516 17740
rect 14648 17688 14700 17740
rect 15108 17688 15160 17740
rect 13912 17620 13964 17672
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 15476 17620 15528 17672
rect 15660 17663 15712 17672
rect 15660 17629 15669 17663
rect 15669 17629 15703 17663
rect 15703 17629 15712 17663
rect 15660 17620 15712 17629
rect 19708 17824 19760 17876
rect 17040 17756 17092 17808
rect 20444 17756 20496 17808
rect 21272 17824 21324 17876
rect 23572 17756 23624 17808
rect 17776 17688 17828 17740
rect 18328 17688 18380 17740
rect 25412 17688 25464 17740
rect 28264 17688 28316 17740
rect 29092 17731 29144 17740
rect 29092 17697 29101 17731
rect 29101 17697 29135 17731
rect 29135 17697 29144 17731
rect 29092 17688 29144 17697
rect 29184 17731 29236 17740
rect 29184 17697 29193 17731
rect 29193 17697 29227 17731
rect 29227 17697 29236 17731
rect 29184 17688 29236 17697
rect 17316 17620 17368 17672
rect 23204 17663 23256 17672
rect 23204 17629 23213 17663
rect 23213 17629 23247 17663
rect 23247 17629 23256 17663
rect 23204 17620 23256 17629
rect 26608 17663 26660 17672
rect 26608 17629 26617 17663
rect 26617 17629 26651 17663
rect 26651 17629 26660 17663
rect 26608 17620 26660 17629
rect 30104 17756 30156 17808
rect 31668 17799 31720 17808
rect 31668 17765 31677 17799
rect 31677 17765 31711 17799
rect 31711 17765 31720 17799
rect 31668 17756 31720 17765
rect 29828 17731 29880 17740
rect 29828 17697 29837 17731
rect 29837 17697 29871 17731
rect 29871 17697 29880 17731
rect 29828 17688 29880 17697
rect 30012 17731 30064 17740
rect 30012 17697 30021 17731
rect 30021 17697 30055 17731
rect 30055 17697 30064 17731
rect 30012 17688 30064 17697
rect 30564 17688 30616 17740
rect 31392 17688 31444 17740
rect 37740 17756 37792 17808
rect 30840 17663 30892 17672
rect 30840 17629 30874 17663
rect 30874 17629 30892 17663
rect 30840 17620 30892 17629
rect 31024 17663 31076 17672
rect 31024 17629 31033 17663
rect 31033 17629 31067 17663
rect 31067 17629 31076 17663
rect 31024 17620 31076 17629
rect 34520 17620 34572 17672
rect 34704 17620 34756 17672
rect 34980 17620 35032 17672
rect 35532 17688 35584 17740
rect 37464 17620 37516 17672
rect 37924 17620 37976 17672
rect 41236 17824 41288 17876
rect 42892 17824 42944 17876
rect 45836 17867 45888 17876
rect 45836 17833 45845 17867
rect 45845 17833 45879 17867
rect 45879 17833 45888 17867
rect 45836 17824 45888 17833
rect 46112 17824 46164 17876
rect 41052 17756 41104 17808
rect 44088 17756 44140 17808
rect 40408 17688 40460 17740
rect 38660 17663 38712 17672
rect 38660 17629 38669 17663
rect 38669 17629 38703 17663
rect 38703 17629 38712 17663
rect 38660 17620 38712 17629
rect 38844 17620 38896 17672
rect 39948 17620 40000 17672
rect 41328 17620 41380 17672
rect 44180 17663 44232 17672
rect 44180 17629 44189 17663
rect 44189 17629 44223 17663
rect 44223 17629 44232 17663
rect 44180 17620 44232 17629
rect 4804 17484 4856 17536
rect 5172 17484 5224 17536
rect 6920 17552 6972 17604
rect 7196 17527 7248 17536
rect 7196 17493 7205 17527
rect 7205 17493 7239 17527
rect 7239 17493 7248 17527
rect 7196 17484 7248 17493
rect 7932 17484 7984 17536
rect 11980 17484 12032 17536
rect 17040 17595 17092 17604
rect 17040 17561 17049 17595
rect 17049 17561 17083 17595
rect 17083 17561 17092 17595
rect 17040 17552 17092 17561
rect 26884 17552 26936 17604
rect 33876 17552 33928 17604
rect 35348 17552 35400 17604
rect 15660 17484 15712 17536
rect 23020 17527 23072 17536
rect 23020 17493 23029 17527
rect 23029 17493 23063 17527
rect 23063 17493 23072 17527
rect 23020 17484 23072 17493
rect 26424 17527 26476 17536
rect 26424 17493 26433 17527
rect 26433 17493 26467 17527
rect 26467 17493 26476 17527
rect 26424 17484 26476 17493
rect 26700 17484 26752 17536
rect 26976 17484 27028 17536
rect 29000 17527 29052 17536
rect 29000 17493 29009 17527
rect 29009 17493 29043 17527
rect 29043 17493 29052 17527
rect 29000 17484 29052 17493
rect 29552 17527 29604 17536
rect 29552 17493 29561 17527
rect 29561 17493 29595 17527
rect 29595 17493 29604 17527
rect 29552 17484 29604 17493
rect 30288 17484 30340 17536
rect 30840 17484 30892 17536
rect 34704 17527 34756 17536
rect 34704 17493 34713 17527
rect 34713 17493 34747 17527
rect 34747 17493 34756 17527
rect 34704 17484 34756 17493
rect 35164 17527 35216 17536
rect 35164 17493 35173 17527
rect 35173 17493 35207 17527
rect 35207 17493 35216 17527
rect 35164 17484 35216 17493
rect 35992 17484 36044 17536
rect 38108 17595 38160 17604
rect 38108 17561 38117 17595
rect 38117 17561 38151 17595
rect 38151 17561 38160 17595
rect 38108 17552 38160 17561
rect 42800 17552 42852 17604
rect 43812 17552 43864 17604
rect 44364 17663 44416 17672
rect 44364 17629 44373 17663
rect 44373 17629 44407 17663
rect 44407 17629 44416 17663
rect 44364 17620 44416 17629
rect 44548 17663 44600 17672
rect 44548 17629 44557 17663
rect 44557 17629 44591 17663
rect 44591 17629 44600 17663
rect 44548 17620 44600 17629
rect 45560 17620 45612 17672
rect 46388 17663 46440 17672
rect 46388 17629 46397 17663
rect 46397 17629 46431 17663
rect 46431 17629 46440 17663
rect 46388 17620 46440 17629
rect 46756 17663 46808 17672
rect 46756 17629 46765 17663
rect 46765 17629 46799 17663
rect 46799 17629 46808 17663
rect 46756 17620 46808 17629
rect 41880 17484 41932 17536
rect 45008 17484 45060 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 2228 17280 2280 17332
rect 3792 17280 3844 17332
rect 6644 17280 6696 17332
rect 7288 17280 7340 17332
rect 8300 17280 8352 17332
rect 14280 17280 14332 17332
rect 14556 17323 14608 17332
rect 14556 17289 14565 17323
rect 14565 17289 14599 17323
rect 14599 17289 14608 17323
rect 14556 17280 14608 17289
rect 15660 17280 15712 17332
rect 21272 17323 21324 17332
rect 6828 17212 6880 17264
rect 21272 17289 21281 17323
rect 21281 17289 21315 17323
rect 21315 17289 21324 17323
rect 21272 17280 21324 17289
rect 20352 17212 20404 17264
rect 940 17144 992 17196
rect 2320 17187 2372 17196
rect 2320 17153 2354 17187
rect 2354 17153 2372 17187
rect 2320 17144 2372 17153
rect 4528 17144 4580 17196
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 7932 17187 7984 17196
rect 7932 17153 7941 17187
rect 7941 17153 7975 17187
rect 7975 17153 7984 17187
rect 7932 17144 7984 17153
rect 14188 17144 14240 17196
rect 14832 17144 14884 17196
rect 19248 17187 19300 17196
rect 19248 17153 19257 17187
rect 19257 17153 19291 17187
rect 19291 17153 19300 17187
rect 19248 17144 19300 17153
rect 22652 17280 22704 17332
rect 23480 17280 23532 17332
rect 24032 17323 24084 17332
rect 24032 17289 24041 17323
rect 24041 17289 24075 17323
rect 24075 17289 24084 17323
rect 24032 17280 24084 17289
rect 26332 17323 26384 17332
rect 26332 17289 26341 17323
rect 26341 17289 26375 17323
rect 26375 17289 26384 17323
rect 26332 17280 26384 17289
rect 26516 17280 26568 17332
rect 29000 17280 29052 17332
rect 30288 17280 30340 17332
rect 34428 17280 34480 17332
rect 38844 17280 38896 17332
rect 39948 17280 40000 17332
rect 40316 17280 40368 17332
rect 41236 17280 41288 17332
rect 41328 17280 41380 17332
rect 42156 17280 42208 17332
rect 42248 17280 42300 17332
rect 42800 17280 42852 17332
rect 44548 17323 44600 17332
rect 44548 17289 44557 17323
rect 44557 17289 44591 17323
rect 44591 17289 44600 17323
rect 44548 17280 44600 17289
rect 23020 17212 23072 17264
rect 24860 17212 24912 17264
rect 26424 17212 26476 17264
rect 29552 17212 29604 17264
rect 29828 17212 29880 17264
rect 32128 17212 32180 17264
rect 38384 17212 38436 17264
rect 22560 17144 22612 17196
rect 4160 17119 4212 17128
rect 4160 17085 4169 17119
rect 4169 17085 4203 17119
rect 4203 17085 4212 17119
rect 4160 17076 4212 17085
rect 4712 17076 4764 17128
rect 5264 17076 5316 17128
rect 5540 17076 5592 17128
rect 6736 17076 6788 17128
rect 7840 17076 7892 17128
rect 16212 17076 16264 17128
rect 18144 17076 18196 17128
rect 18236 17119 18288 17128
rect 18236 17085 18245 17119
rect 18245 17085 18279 17119
rect 18279 17085 18288 17119
rect 18236 17076 18288 17085
rect 18788 17076 18840 17128
rect 19156 17076 19208 17128
rect 19892 17076 19944 17128
rect 4620 17008 4672 17060
rect 2412 16940 2464 16992
rect 12348 17008 12400 17060
rect 17960 17008 18012 17060
rect 18696 17051 18748 17060
rect 18696 17017 18705 17051
rect 18705 17017 18739 17051
rect 18739 17017 18748 17051
rect 18696 17008 18748 17017
rect 5356 16940 5408 16992
rect 6644 16940 6696 16992
rect 7196 16940 7248 16992
rect 7840 16940 7892 16992
rect 11060 16940 11112 16992
rect 13084 16940 13136 16992
rect 16948 16940 17000 16992
rect 20076 16940 20128 16992
rect 20996 16940 21048 16992
rect 21180 16940 21232 16992
rect 21640 16940 21692 16992
rect 25964 16983 26016 16992
rect 25964 16949 25973 16983
rect 25973 16949 26007 16983
rect 26007 16949 26016 16983
rect 25964 16940 26016 16949
rect 26884 17144 26936 17196
rect 31392 17144 31444 17196
rect 26700 17076 26752 17128
rect 26792 17076 26844 17128
rect 28540 17119 28592 17128
rect 28540 17085 28549 17119
rect 28549 17085 28583 17119
rect 28583 17085 28592 17119
rect 28540 17076 28592 17085
rect 29920 17076 29972 17128
rect 31024 17076 31076 17128
rect 33232 17144 33284 17196
rect 34336 17187 34388 17196
rect 34336 17153 34345 17187
rect 34345 17153 34379 17187
rect 34379 17153 34388 17187
rect 34336 17144 34388 17153
rect 34704 17144 34756 17196
rect 36084 17144 36136 17196
rect 29644 17008 29696 17060
rect 30472 17008 30524 17060
rect 33600 17119 33652 17128
rect 33600 17085 33609 17119
rect 33609 17085 33643 17119
rect 33643 17085 33652 17119
rect 33600 17076 33652 17085
rect 34152 17076 34204 17128
rect 35164 17076 35216 17128
rect 34336 17008 34388 17060
rect 31300 16940 31352 16992
rect 32864 16940 32916 16992
rect 34152 16940 34204 16992
rect 34980 16940 35032 16992
rect 35532 16940 35584 16992
rect 38016 16940 38068 16992
rect 38476 16940 38528 16992
rect 38844 17187 38896 17196
rect 38844 17153 38853 17187
rect 38853 17153 38887 17187
rect 38887 17153 38896 17187
rect 38844 17144 38896 17153
rect 42064 17212 42116 17264
rect 40040 17144 40092 17196
rect 39856 17076 39908 17128
rect 38936 17008 38988 17060
rect 41696 17144 41748 17196
rect 41144 17076 41196 17128
rect 41236 17076 41288 17128
rect 43076 17144 43128 17196
rect 44364 17144 44416 17196
rect 40868 17008 40920 17060
rect 43168 17076 43220 17128
rect 43536 17076 43588 17128
rect 44824 17212 44876 17264
rect 44732 17187 44784 17196
rect 44732 17153 44741 17187
rect 44741 17153 44775 17187
rect 44775 17153 44784 17187
rect 44732 17144 44784 17153
rect 42248 17008 42300 17060
rect 43352 17008 43404 17060
rect 44916 17051 44968 17060
rect 44916 17017 44925 17051
rect 44925 17017 44959 17051
rect 44959 17017 44968 17051
rect 44916 17008 44968 17017
rect 40224 16940 40276 16992
rect 42340 16940 42392 16992
rect 44088 16940 44140 16992
rect 45100 16940 45152 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2320 16736 2372 16788
rect 4804 16736 4856 16788
rect 2136 16668 2188 16720
rect 6828 16668 6880 16720
rect 3792 16600 3844 16652
rect 5356 16600 5408 16652
rect 4712 16532 4764 16584
rect 5448 16575 5500 16584
rect 5448 16541 5457 16575
rect 5457 16541 5491 16575
rect 5491 16541 5500 16575
rect 5448 16532 5500 16541
rect 6276 16600 6328 16652
rect 9404 16643 9456 16652
rect 9404 16609 9413 16643
rect 9413 16609 9447 16643
rect 9447 16609 9456 16643
rect 9404 16600 9456 16609
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 12624 16600 12676 16652
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 16948 16668 17000 16720
rect 15936 16600 15988 16652
rect 16212 16600 16264 16652
rect 16672 16600 16724 16652
rect 18236 16736 18288 16788
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 20076 16711 20128 16720
rect 20076 16677 20085 16711
rect 20085 16677 20119 16711
rect 20119 16677 20128 16711
rect 20076 16668 20128 16677
rect 23204 16779 23256 16788
rect 23204 16745 23213 16779
rect 23213 16745 23247 16779
rect 23247 16745 23256 16779
rect 23204 16736 23256 16745
rect 8300 16532 8352 16584
rect 9220 16532 9272 16584
rect 10692 16464 10744 16516
rect 4252 16439 4304 16448
rect 4252 16405 4261 16439
rect 4261 16405 4295 16439
rect 4295 16405 4304 16439
rect 4252 16396 4304 16405
rect 10140 16396 10192 16448
rect 12072 16396 12124 16448
rect 12440 16396 12492 16448
rect 13636 16396 13688 16448
rect 14096 16396 14148 16448
rect 14740 16396 14792 16448
rect 16948 16575 17000 16584
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 16948 16532 17000 16541
rect 20260 16532 20312 16584
rect 17224 16507 17276 16516
rect 17224 16473 17258 16507
rect 17258 16473 17276 16507
rect 17224 16464 17276 16473
rect 20536 16575 20588 16584
rect 20536 16541 20545 16575
rect 20545 16541 20579 16575
rect 20579 16541 20588 16575
rect 20536 16532 20588 16541
rect 23572 16668 23624 16720
rect 24860 16779 24912 16788
rect 24860 16745 24869 16779
rect 24869 16745 24903 16779
rect 24903 16745 24912 16779
rect 24860 16736 24912 16745
rect 26608 16736 26660 16788
rect 32128 16779 32180 16788
rect 32128 16745 32137 16779
rect 32137 16745 32171 16779
rect 32171 16745 32180 16779
rect 32128 16736 32180 16745
rect 34428 16736 34480 16788
rect 39856 16736 39908 16788
rect 30656 16668 30708 16720
rect 23848 16643 23900 16652
rect 23848 16609 23857 16643
rect 23857 16609 23891 16643
rect 23891 16609 23900 16643
rect 23848 16600 23900 16609
rect 26884 16643 26936 16652
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 28448 16600 28500 16652
rect 20996 16532 21048 16584
rect 24032 16532 24084 16584
rect 25964 16532 26016 16584
rect 26516 16532 26568 16584
rect 29092 16532 29144 16584
rect 29644 16532 29696 16584
rect 30288 16532 30340 16584
rect 31576 16532 31628 16584
rect 32864 16575 32916 16584
rect 32864 16541 32873 16575
rect 32873 16541 32907 16575
rect 32907 16541 32916 16575
rect 32864 16532 32916 16541
rect 38016 16643 38068 16652
rect 38016 16609 38025 16643
rect 38025 16609 38059 16643
rect 38059 16609 38068 16643
rect 38016 16600 38068 16609
rect 34336 16532 34388 16584
rect 34612 16532 34664 16584
rect 35532 16532 35584 16584
rect 21272 16464 21324 16516
rect 21824 16464 21876 16516
rect 23940 16464 23992 16516
rect 15292 16439 15344 16448
rect 15292 16405 15301 16439
rect 15301 16405 15335 16439
rect 15335 16405 15344 16439
rect 15292 16396 15344 16405
rect 15844 16396 15896 16448
rect 17960 16396 18012 16448
rect 19156 16396 19208 16448
rect 19340 16396 19392 16448
rect 19800 16396 19852 16448
rect 21180 16396 21232 16448
rect 25136 16464 25188 16516
rect 31116 16464 31168 16516
rect 24308 16396 24360 16448
rect 27068 16396 27120 16448
rect 34060 16464 34112 16516
rect 37280 16575 37332 16584
rect 37280 16541 37289 16575
rect 37289 16541 37323 16575
rect 37323 16541 37332 16575
rect 37280 16532 37332 16541
rect 38292 16575 38344 16584
rect 38292 16541 38301 16575
rect 38301 16541 38335 16575
rect 38335 16541 38344 16575
rect 38292 16532 38344 16541
rect 38476 16575 38528 16584
rect 38476 16541 38485 16575
rect 38485 16541 38519 16575
rect 38519 16541 38528 16575
rect 38476 16532 38528 16541
rect 38844 16575 38896 16584
rect 38844 16541 38853 16575
rect 38853 16541 38887 16575
rect 38887 16541 38896 16575
rect 38844 16532 38896 16541
rect 39948 16532 40000 16584
rect 40684 16668 40736 16720
rect 40868 16668 40920 16720
rect 42064 16736 42116 16788
rect 42708 16736 42760 16788
rect 42800 16736 42852 16788
rect 44732 16779 44784 16788
rect 44732 16745 44741 16779
rect 44741 16745 44775 16779
rect 44775 16745 44784 16779
rect 44732 16736 44784 16745
rect 44824 16736 44876 16788
rect 41052 16600 41104 16652
rect 37924 16464 37976 16516
rect 34244 16396 34296 16448
rect 34428 16396 34480 16448
rect 38936 16439 38988 16448
rect 38936 16405 38945 16439
rect 38945 16405 38979 16439
rect 38979 16405 38988 16439
rect 38936 16396 38988 16405
rect 40040 16396 40092 16448
rect 40316 16507 40368 16516
rect 40316 16473 40325 16507
rect 40325 16473 40359 16507
rect 40359 16473 40368 16507
rect 40316 16464 40368 16473
rect 40776 16532 40828 16584
rect 40960 16575 41012 16584
rect 40960 16541 40969 16575
rect 40969 16541 41003 16575
rect 41003 16541 41012 16575
rect 40960 16532 41012 16541
rect 41236 16575 41288 16584
rect 41236 16541 41245 16575
rect 41245 16541 41279 16575
rect 41279 16541 41288 16575
rect 41236 16532 41288 16541
rect 42616 16643 42668 16652
rect 42616 16609 42625 16643
rect 42625 16609 42659 16643
rect 42659 16609 42668 16643
rect 42616 16600 42668 16609
rect 40776 16396 40828 16448
rect 40960 16396 41012 16448
rect 41328 16396 41380 16448
rect 41604 16396 41656 16448
rect 42156 16575 42208 16584
rect 42156 16541 42165 16575
rect 42165 16541 42199 16575
rect 42199 16541 42208 16575
rect 42156 16532 42208 16541
rect 42340 16575 42392 16584
rect 42340 16541 42349 16575
rect 42349 16541 42383 16575
rect 42383 16541 42392 16575
rect 42340 16532 42392 16541
rect 42524 16575 42576 16584
rect 42524 16541 42533 16575
rect 42533 16541 42567 16575
rect 42567 16541 42576 16575
rect 42524 16532 42576 16541
rect 42708 16532 42760 16584
rect 43352 16643 43404 16652
rect 43352 16609 43361 16643
rect 43361 16609 43395 16643
rect 43395 16609 43404 16643
rect 43352 16600 43404 16609
rect 43076 16532 43128 16584
rect 44088 16668 44140 16720
rect 44916 16668 44968 16720
rect 45376 16600 45428 16652
rect 43812 16575 43864 16584
rect 43812 16541 43821 16575
rect 43821 16541 43855 16575
rect 43855 16541 43864 16575
rect 43812 16532 43864 16541
rect 45008 16575 45060 16584
rect 45008 16541 45017 16575
rect 45017 16541 45051 16575
rect 45051 16541 45060 16575
rect 45008 16532 45060 16541
rect 42708 16396 42760 16448
rect 43260 16439 43312 16448
rect 43260 16405 43269 16439
rect 43269 16405 43303 16439
rect 43303 16405 43312 16439
rect 43260 16396 43312 16405
rect 43536 16507 43588 16516
rect 43536 16473 43545 16507
rect 43545 16473 43579 16507
rect 43579 16473 43588 16507
rect 43536 16464 43588 16473
rect 44364 16464 44416 16516
rect 45744 16507 45796 16516
rect 45744 16473 45753 16507
rect 45753 16473 45787 16507
rect 45787 16473 45796 16507
rect 45744 16464 45796 16473
rect 44732 16396 44784 16448
rect 44824 16396 44876 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 5264 16192 5316 16244
rect 6920 16192 6972 16244
rect 7288 16192 7340 16244
rect 9496 16192 9548 16244
rect 10048 16192 10100 16244
rect 10692 16235 10744 16244
rect 10692 16201 10701 16235
rect 10701 16201 10735 16235
rect 10735 16201 10744 16235
rect 10692 16192 10744 16201
rect 7104 16124 7156 16176
rect 11060 16124 11112 16176
rect 2412 16056 2464 16108
rect 2596 16099 2648 16108
rect 2596 16065 2630 16099
rect 2630 16065 2648 16099
rect 2596 16056 2648 16065
rect 4252 16099 4304 16108
rect 4252 16065 4261 16099
rect 4261 16065 4295 16099
rect 4295 16065 4304 16099
rect 4252 16056 4304 16065
rect 4712 16056 4764 16108
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 3976 15988 4028 16040
rect 6920 15988 6972 16040
rect 5724 15920 5776 15972
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 8760 16031 8812 16040
rect 8760 15997 8769 16031
rect 8769 15997 8803 16031
rect 8803 15997 8812 16031
rect 8760 15988 8812 15997
rect 8944 16031 8996 16040
rect 8944 15997 8953 16031
rect 8953 15997 8987 16031
rect 8987 15997 8996 16031
rect 8944 15988 8996 15997
rect 9956 16099 10008 16108
rect 9956 16065 9965 16099
rect 9965 16065 9999 16099
rect 9999 16065 10008 16099
rect 9956 16056 10008 16065
rect 10692 16056 10744 16108
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 9772 16031 9824 16040
rect 9772 15997 9806 16031
rect 9806 15997 9824 16031
rect 9772 15988 9824 15997
rect 12072 16031 12124 16040
rect 12072 15997 12081 16031
rect 12081 15997 12115 16031
rect 12115 15997 12124 16031
rect 12072 15988 12124 15997
rect 9220 15920 9272 15972
rect 16672 16192 16724 16244
rect 17224 16235 17276 16244
rect 17224 16201 17233 16235
rect 17233 16201 17267 16235
rect 17267 16201 17276 16235
rect 17224 16192 17276 16201
rect 3792 15895 3844 15904
rect 3792 15861 3801 15895
rect 3801 15861 3835 15895
rect 3835 15861 3844 15895
rect 3792 15852 3844 15861
rect 6368 15895 6420 15904
rect 6368 15861 6377 15895
rect 6377 15861 6411 15895
rect 6411 15861 6420 15895
rect 6368 15852 6420 15861
rect 7196 15852 7248 15904
rect 10324 15852 10376 15904
rect 15844 16124 15896 16176
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 14740 16099 14792 16108
rect 14740 16065 14774 16099
rect 14774 16065 14792 16099
rect 14740 16056 14792 16065
rect 15292 16056 15344 16108
rect 14096 16031 14148 16040
rect 14096 15997 14105 16031
rect 14105 15997 14139 16031
rect 14139 15997 14148 16031
rect 14096 15988 14148 15997
rect 17316 16056 17368 16108
rect 17132 15988 17184 16040
rect 20996 16192 21048 16244
rect 21180 16235 21232 16244
rect 21180 16201 21189 16235
rect 21189 16201 21223 16235
rect 21223 16201 21232 16235
rect 21180 16192 21232 16201
rect 21272 16192 21324 16244
rect 21088 16124 21140 16176
rect 18236 16056 18288 16108
rect 19340 16099 19392 16108
rect 19340 16065 19374 16099
rect 19374 16065 19392 16099
rect 19340 16056 19392 16065
rect 20168 16056 20220 16108
rect 21272 16056 21324 16108
rect 21364 16099 21416 16108
rect 21364 16065 21373 16099
rect 21373 16065 21407 16099
rect 21407 16065 21416 16099
rect 21364 16056 21416 16065
rect 21456 16056 21508 16108
rect 21824 16056 21876 16108
rect 22468 16099 22520 16108
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 22468 16056 22520 16065
rect 26700 16192 26752 16244
rect 29184 16192 29236 16244
rect 31116 16235 31168 16244
rect 31116 16201 31125 16235
rect 31125 16201 31159 16235
rect 31159 16201 31168 16235
rect 31116 16192 31168 16201
rect 24216 16124 24268 16176
rect 17776 15988 17828 16040
rect 18328 16031 18380 16040
rect 18328 15997 18337 16031
rect 18337 15997 18371 16031
rect 18371 15997 18380 16031
rect 18328 15988 18380 15997
rect 17960 15920 18012 15972
rect 18788 15920 18840 15972
rect 14648 15852 14700 15904
rect 16304 15895 16356 15904
rect 16304 15861 16313 15895
rect 16313 15861 16347 15895
rect 16347 15861 16356 15895
rect 16304 15852 16356 15861
rect 16672 15852 16724 15904
rect 19984 15852 20036 15904
rect 20536 15988 20588 16040
rect 23664 16099 23716 16108
rect 23664 16065 23673 16099
rect 23673 16065 23707 16099
rect 23707 16065 23716 16099
rect 23664 16056 23716 16065
rect 23940 16099 23992 16108
rect 23940 16065 23949 16099
rect 23949 16065 23983 16099
rect 23983 16065 23992 16099
rect 23940 16056 23992 16065
rect 24860 16099 24912 16108
rect 24860 16065 24869 16099
rect 24869 16065 24903 16099
rect 24903 16065 24912 16099
rect 24860 16056 24912 16065
rect 28908 16124 28960 16176
rect 29092 16124 29144 16176
rect 31944 16124 31996 16176
rect 34060 16235 34112 16244
rect 34060 16201 34069 16235
rect 34069 16201 34103 16235
rect 34103 16201 34112 16235
rect 34060 16192 34112 16201
rect 35348 16192 35400 16244
rect 38292 16192 38344 16244
rect 43812 16192 43864 16244
rect 45376 16235 45428 16244
rect 45376 16201 45385 16235
rect 45385 16201 45419 16235
rect 45419 16201 45428 16235
rect 45376 16192 45428 16201
rect 34612 16167 34664 16176
rect 34612 16133 34646 16167
rect 34646 16133 34664 16167
rect 34612 16124 34664 16133
rect 38936 16124 38988 16176
rect 25136 16056 25188 16108
rect 26516 16099 26568 16108
rect 26516 16065 26525 16099
rect 26525 16065 26559 16099
rect 26559 16065 26568 16099
rect 26516 16056 26568 16065
rect 27068 16099 27120 16108
rect 27068 16065 27077 16099
rect 27077 16065 27111 16099
rect 27111 16065 27120 16099
rect 27068 16056 27120 16065
rect 27712 16056 27764 16108
rect 27896 16099 27948 16108
rect 27896 16065 27905 16099
rect 27905 16065 27939 16099
rect 27939 16065 27948 16099
rect 27896 16056 27948 16065
rect 28264 16099 28316 16108
rect 28264 16065 28273 16099
rect 28273 16065 28307 16099
rect 28307 16065 28316 16099
rect 28264 16056 28316 16065
rect 29000 16099 29052 16108
rect 29000 16065 29009 16099
rect 29009 16065 29043 16099
rect 29043 16065 29052 16099
rect 29000 16056 29052 16065
rect 31300 16099 31352 16108
rect 31300 16065 31309 16099
rect 31309 16065 31343 16099
rect 31343 16065 31352 16099
rect 31300 16056 31352 16065
rect 31576 16056 31628 16108
rect 32404 16099 32456 16108
rect 32404 16065 32438 16099
rect 32438 16065 32456 16099
rect 32404 16056 32456 16065
rect 34244 16099 34296 16108
rect 34244 16065 34253 16099
rect 34253 16065 34287 16099
rect 34287 16065 34296 16099
rect 34244 16056 34296 16065
rect 34336 16099 34388 16108
rect 34336 16065 34345 16099
rect 34345 16065 34379 16099
rect 34379 16065 34388 16099
rect 34336 16056 34388 16065
rect 37556 16099 37608 16108
rect 37556 16065 37565 16099
rect 37565 16065 37599 16099
rect 37599 16065 37608 16099
rect 37556 16056 37608 16065
rect 39396 16056 39448 16108
rect 40224 16056 40276 16108
rect 40776 16099 40828 16108
rect 40776 16065 40785 16099
rect 40785 16065 40819 16099
rect 40819 16065 40828 16099
rect 40776 16056 40828 16065
rect 24032 15988 24084 16040
rect 20812 15852 20864 15904
rect 22008 15852 22060 15904
rect 22560 15852 22612 15904
rect 22652 15895 22704 15904
rect 22652 15861 22661 15895
rect 22661 15861 22695 15895
rect 22695 15861 22704 15895
rect 22652 15852 22704 15861
rect 22836 15895 22888 15904
rect 22836 15861 22845 15895
rect 22845 15861 22879 15895
rect 22879 15861 22888 15895
rect 22836 15852 22888 15861
rect 23296 15895 23348 15904
rect 23296 15861 23305 15895
rect 23305 15861 23339 15895
rect 23339 15861 23348 15895
rect 23296 15852 23348 15861
rect 27712 15920 27764 15972
rect 30104 15920 30156 15972
rect 30288 15920 30340 15972
rect 25320 15852 25372 15904
rect 26056 15852 26108 15904
rect 28172 15852 28224 15904
rect 28448 15895 28500 15904
rect 28448 15861 28457 15895
rect 28457 15861 28491 15895
rect 28491 15861 28500 15895
rect 28448 15852 28500 15861
rect 29644 15852 29696 15904
rect 37280 16031 37332 16040
rect 37280 15997 37289 16031
rect 37289 15997 37323 16031
rect 37323 15997 37332 16031
rect 37280 15988 37332 15997
rect 40316 15988 40368 16040
rect 38844 15920 38896 15972
rect 39028 15920 39080 15972
rect 42156 16056 42208 16108
rect 42708 16099 42760 16108
rect 42708 16065 42717 16099
rect 42717 16065 42751 16099
rect 42751 16065 42760 16099
rect 42708 16056 42760 16065
rect 44732 16056 44784 16108
rect 45836 16056 45888 16108
rect 46480 16099 46532 16108
rect 46480 16065 46489 16099
rect 46489 16065 46523 16099
rect 46523 16065 46532 16099
rect 46480 16056 46532 16065
rect 42524 15920 42576 15972
rect 44824 15988 44876 16040
rect 45100 16031 45152 16040
rect 45100 15997 45109 16031
rect 45109 15997 45143 16031
rect 45143 15997 45152 16031
rect 45100 15988 45152 15997
rect 45468 16031 45520 16040
rect 45468 15997 45477 16031
rect 45477 15997 45511 16031
rect 45511 15997 45520 16031
rect 45468 15988 45520 15997
rect 44916 15920 44968 15972
rect 36084 15852 36136 15904
rect 43720 15852 43772 15904
rect 46664 15895 46716 15904
rect 46664 15861 46673 15895
rect 46673 15861 46707 15895
rect 46707 15861 46716 15895
rect 46664 15852 46716 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2596 15648 2648 15700
rect 8576 15648 8628 15700
rect 8944 15648 8996 15700
rect 7104 15580 7156 15632
rect 3792 15444 3844 15496
rect 4620 15444 4672 15496
rect 5724 15487 5776 15496
rect 5724 15453 5733 15487
rect 5733 15453 5767 15487
rect 5767 15453 5776 15487
rect 5724 15444 5776 15453
rect 5816 15487 5868 15496
rect 5816 15453 5825 15487
rect 5825 15453 5859 15487
rect 5859 15453 5868 15487
rect 5816 15444 5868 15453
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 10140 15648 10192 15700
rect 21456 15648 21508 15700
rect 22468 15648 22520 15700
rect 22560 15648 22612 15700
rect 9496 15512 9548 15564
rect 9680 15512 9732 15564
rect 10508 15512 10560 15564
rect 12072 15512 12124 15564
rect 14648 15580 14700 15632
rect 15844 15580 15896 15632
rect 8760 15444 8812 15496
rect 8944 15487 8996 15496
rect 8944 15453 8953 15487
rect 8953 15453 8987 15487
rect 8987 15453 8996 15487
rect 8944 15444 8996 15453
rect 9956 15487 10008 15496
rect 9956 15453 9990 15487
rect 9990 15453 10008 15487
rect 9956 15444 10008 15453
rect 4160 15351 4212 15360
rect 4160 15317 4169 15351
rect 4169 15317 4203 15351
rect 4203 15317 4212 15351
rect 4160 15308 4212 15317
rect 4712 15308 4764 15360
rect 5264 15308 5316 15360
rect 7196 15376 7248 15428
rect 7748 15351 7800 15360
rect 7748 15317 7757 15351
rect 7757 15317 7791 15351
rect 7791 15317 7800 15351
rect 7748 15308 7800 15317
rect 12532 15376 12584 15428
rect 15292 15376 15344 15428
rect 10232 15308 10284 15360
rect 13176 15308 13228 15360
rect 20352 15623 20404 15632
rect 20352 15589 20361 15623
rect 20361 15589 20395 15623
rect 20395 15589 20404 15623
rect 20352 15580 20404 15589
rect 22008 15580 22060 15632
rect 25136 15580 25188 15632
rect 17776 15512 17828 15564
rect 19340 15512 19392 15564
rect 20076 15512 20128 15564
rect 20904 15555 20956 15564
rect 20904 15521 20913 15555
rect 20913 15521 20947 15555
rect 20947 15521 20956 15555
rect 20904 15512 20956 15521
rect 21272 15512 21324 15564
rect 24124 15512 24176 15564
rect 16212 15351 16264 15360
rect 16212 15317 16221 15351
rect 16221 15317 16255 15351
rect 16255 15317 16264 15351
rect 16212 15308 16264 15317
rect 17132 15308 17184 15360
rect 17224 15351 17276 15360
rect 17224 15317 17233 15351
rect 17233 15317 17267 15351
rect 17267 15317 17276 15351
rect 17224 15308 17276 15317
rect 17316 15308 17368 15360
rect 19524 15444 19576 15496
rect 19708 15487 19760 15496
rect 19708 15453 19717 15487
rect 19717 15453 19751 15487
rect 19751 15453 19760 15487
rect 19708 15444 19760 15453
rect 20720 15487 20772 15496
rect 20720 15453 20754 15487
rect 20754 15453 20772 15487
rect 20720 15444 20772 15453
rect 21916 15444 21968 15496
rect 23480 15444 23532 15496
rect 24860 15444 24912 15496
rect 26792 15444 26844 15496
rect 29368 15487 29420 15496
rect 29368 15453 29377 15487
rect 29377 15453 29411 15487
rect 29411 15453 29420 15487
rect 29368 15444 29420 15453
rect 18328 15376 18380 15428
rect 26332 15419 26384 15428
rect 26332 15385 26366 15419
rect 26366 15385 26384 15419
rect 26332 15376 26384 15385
rect 18236 15308 18288 15360
rect 29092 15376 29144 15428
rect 27344 15308 27396 15360
rect 32404 15691 32456 15700
rect 32404 15657 32413 15691
rect 32413 15657 32447 15691
rect 32447 15657 32456 15691
rect 32404 15648 32456 15657
rect 34244 15648 34296 15700
rect 36268 15648 36320 15700
rect 37004 15648 37056 15700
rect 39856 15648 39908 15700
rect 45744 15648 45796 15700
rect 38108 15580 38160 15632
rect 46480 15580 46532 15632
rect 32036 15512 32088 15564
rect 33692 15512 33744 15564
rect 39212 15512 39264 15564
rect 45560 15555 45612 15564
rect 45560 15521 45569 15555
rect 45569 15521 45603 15555
rect 45603 15521 45612 15555
rect 45560 15512 45612 15521
rect 34428 15444 34480 15496
rect 35992 15444 36044 15496
rect 36544 15444 36596 15496
rect 36912 15487 36964 15496
rect 36912 15453 36921 15487
rect 36921 15453 36955 15487
rect 36955 15453 36964 15487
rect 36912 15444 36964 15453
rect 41236 15444 41288 15496
rect 45192 15444 45244 15496
rect 46388 15487 46440 15496
rect 46388 15453 46397 15487
rect 46397 15453 46431 15487
rect 46431 15453 46440 15487
rect 46388 15444 46440 15453
rect 39764 15376 39816 15428
rect 30932 15351 30984 15360
rect 30932 15317 30941 15351
rect 30941 15317 30975 15351
rect 30975 15317 30984 15351
rect 30932 15308 30984 15317
rect 31944 15351 31996 15360
rect 31944 15317 31953 15351
rect 31953 15317 31987 15351
rect 31987 15317 31996 15351
rect 31944 15308 31996 15317
rect 32496 15308 32548 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 4620 15104 4672 15156
rect 5264 15104 5316 15156
rect 2412 14968 2464 15020
rect 5816 15036 5868 15088
rect 6368 15036 6420 15088
rect 7748 15036 7800 15088
rect 3700 15011 3752 15020
rect 3700 14977 3734 15011
rect 3734 14977 3752 15011
rect 3700 14968 3752 14977
rect 7012 14968 7064 15020
rect 8944 15104 8996 15156
rect 10692 15104 10744 15156
rect 12532 15147 12584 15156
rect 12532 15113 12541 15147
rect 12541 15113 12575 15147
rect 12575 15113 12584 15147
rect 12532 15104 12584 15113
rect 10140 15079 10192 15088
rect 10140 15045 10149 15079
rect 10149 15045 10183 15079
rect 10183 15045 10192 15079
rect 10140 15036 10192 15045
rect 10232 15079 10284 15088
rect 10232 15045 10241 15079
rect 10241 15045 10275 15079
rect 10275 15045 10284 15079
rect 10232 15036 10284 15045
rect 10416 14943 10468 14952
rect 10416 14909 10425 14943
rect 10425 14909 10459 14943
rect 10459 14909 10468 14943
rect 10416 14900 10468 14909
rect 13176 15147 13228 15156
rect 13176 15113 13185 15147
rect 13185 15113 13219 15147
rect 13219 15113 13228 15147
rect 13176 15104 13228 15113
rect 15292 15147 15344 15156
rect 15292 15113 15301 15147
rect 15301 15113 15335 15147
rect 15335 15113 15344 15147
rect 15292 15104 15344 15113
rect 16212 15104 16264 15156
rect 18328 15147 18380 15156
rect 18328 15113 18337 15147
rect 18337 15113 18371 15147
rect 18371 15113 18380 15147
rect 18328 15104 18380 15113
rect 19340 15104 19392 15156
rect 20260 15104 20312 15156
rect 16304 15036 16356 15088
rect 17224 15079 17276 15088
rect 17224 15045 17258 15079
rect 17258 15045 17276 15079
rect 17224 15036 17276 15045
rect 22652 15104 22704 15156
rect 26332 15147 26384 15156
rect 26332 15113 26341 15147
rect 26341 15113 26375 15147
rect 26375 15113 26384 15147
rect 26332 15104 26384 15113
rect 23296 15036 23348 15088
rect 16948 15011 17000 15020
rect 16948 14977 16957 15011
rect 16957 14977 16991 15011
rect 16991 14977 17000 15011
rect 16948 14968 17000 14977
rect 19340 15011 19392 15020
rect 19340 14977 19349 15011
rect 19349 14977 19383 15011
rect 19383 14977 19392 15011
rect 19340 14968 19392 14977
rect 20076 15011 20128 15020
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 20352 15011 20404 15020
rect 20352 14977 20361 15011
rect 20361 14977 20395 15011
rect 20395 14977 20404 15011
rect 20352 14968 20404 14977
rect 20996 14968 21048 15020
rect 26424 14968 26476 15020
rect 29368 15104 29420 15156
rect 30656 15104 30708 15156
rect 30932 15104 30984 15156
rect 45192 15104 45244 15156
rect 46388 15104 46440 15156
rect 28172 15036 28224 15088
rect 29920 15036 29972 15088
rect 31300 15036 31352 15088
rect 27344 15011 27396 15020
rect 27344 14977 27353 15011
rect 27353 14977 27387 15011
rect 27387 14977 27396 15011
rect 27344 14968 27396 14977
rect 28632 14968 28684 15020
rect 33784 15011 33836 15020
rect 33784 14977 33793 15011
rect 33793 14977 33827 15011
rect 33827 14977 33836 15011
rect 33784 14968 33836 14977
rect 35348 14968 35400 15020
rect 37096 14968 37148 15020
rect 38476 14968 38528 15020
rect 40132 15036 40184 15088
rect 13636 14900 13688 14952
rect 15936 14943 15988 14952
rect 15936 14909 15945 14943
rect 15945 14909 15979 14943
rect 15979 14909 15988 14943
rect 15936 14900 15988 14909
rect 19708 14900 19760 14952
rect 20720 14900 20772 14952
rect 21732 14900 21784 14952
rect 26884 14900 26936 14952
rect 27436 14943 27488 14952
rect 27436 14909 27445 14943
rect 27445 14909 27479 14943
rect 27479 14909 27488 14943
rect 27436 14900 27488 14909
rect 28448 14900 28500 14952
rect 29736 14943 29788 14952
rect 29736 14909 29745 14943
rect 29745 14909 29779 14943
rect 29779 14909 29788 14943
rect 29736 14900 29788 14909
rect 18696 14832 18748 14884
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 9588 14764 9640 14816
rect 16212 14764 16264 14816
rect 27804 14832 27856 14884
rect 35900 14900 35952 14952
rect 39304 15011 39356 15020
rect 39304 14977 39313 15011
rect 39313 14977 39347 15011
rect 39347 14977 39356 15011
rect 39304 14968 39356 14977
rect 39396 15011 39448 15020
rect 39396 14977 39405 15011
rect 39405 14977 39439 15011
rect 39439 14977 39448 15011
rect 39396 14968 39448 14977
rect 42156 14968 42208 15020
rect 42524 14968 42576 15020
rect 43260 14968 43312 15020
rect 43720 15011 43772 15020
rect 43720 14977 43729 15011
rect 43729 14977 43763 15011
rect 43763 14977 43772 15011
rect 43720 14968 43772 14977
rect 44272 15036 44324 15088
rect 45192 15011 45244 15020
rect 45192 14977 45201 15011
rect 45201 14977 45235 15011
rect 45235 14977 45244 15011
rect 45192 14968 45244 14977
rect 39212 14832 39264 14884
rect 43628 14875 43680 14884
rect 43628 14841 43637 14875
rect 43637 14841 43671 14875
rect 43671 14841 43680 14875
rect 43628 14832 43680 14841
rect 23388 14764 23440 14816
rect 26516 14764 26568 14816
rect 29092 14764 29144 14816
rect 34152 14764 34204 14816
rect 34336 14764 34388 14816
rect 38660 14807 38712 14816
rect 38660 14773 38669 14807
rect 38669 14773 38703 14807
rect 38703 14773 38712 14807
rect 38660 14764 38712 14773
rect 39672 14807 39724 14816
rect 39672 14773 39681 14807
rect 39681 14773 39715 14807
rect 39715 14773 39724 14807
rect 39672 14764 39724 14773
rect 41144 14807 41196 14816
rect 41144 14773 41153 14807
rect 41153 14773 41187 14807
rect 41187 14773 41196 14807
rect 41144 14764 41196 14773
rect 42984 14764 43036 14816
rect 45468 14807 45520 14816
rect 45468 14773 45477 14807
rect 45477 14773 45511 14807
rect 45511 14773 45520 14807
rect 45468 14764 45520 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3700 14560 3752 14612
rect 6552 14603 6604 14612
rect 6552 14569 6561 14603
rect 6561 14569 6595 14603
rect 6595 14569 6604 14603
rect 6552 14560 6604 14569
rect 10232 14560 10284 14612
rect 6920 14424 6972 14476
rect 18328 14560 18380 14612
rect 19064 14560 19116 14612
rect 20352 14560 20404 14612
rect 24032 14560 24084 14612
rect 26424 14560 26476 14612
rect 19800 14492 19852 14544
rect 20536 14492 20588 14544
rect 27804 14603 27856 14612
rect 27804 14569 27813 14603
rect 27813 14569 27847 14603
rect 27847 14569 27856 14603
rect 27804 14560 27856 14569
rect 28632 14603 28684 14612
rect 28632 14569 28641 14603
rect 28641 14569 28675 14603
rect 28675 14569 28684 14603
rect 28632 14560 28684 14569
rect 28908 14560 28960 14612
rect 30748 14560 30800 14612
rect 33508 14560 33560 14612
rect 37648 14560 37700 14612
rect 38200 14560 38252 14612
rect 39672 14560 39724 14612
rect 40316 14560 40368 14612
rect 41236 14603 41288 14612
rect 41236 14569 41245 14603
rect 41245 14569 41279 14603
rect 41279 14569 41288 14603
rect 41236 14560 41288 14569
rect 22284 14467 22336 14476
rect 22284 14433 22293 14467
rect 22293 14433 22327 14467
rect 22327 14433 22336 14467
rect 22284 14424 22336 14433
rect 25228 14424 25280 14476
rect 26608 14467 26660 14476
rect 26608 14433 26617 14467
rect 26617 14433 26651 14467
rect 26651 14433 26660 14467
rect 26608 14424 26660 14433
rect 26976 14467 27028 14476
rect 26976 14433 27010 14467
rect 27010 14433 27028 14467
rect 26976 14424 27028 14433
rect 27528 14424 27580 14476
rect 29736 14492 29788 14544
rect 42156 14603 42208 14612
rect 42156 14569 42165 14603
rect 42165 14569 42199 14603
rect 42199 14569 42208 14603
rect 42156 14560 42208 14569
rect 45376 14560 45428 14612
rect 29184 14467 29236 14476
rect 29184 14433 29193 14467
rect 29193 14433 29227 14467
rect 29227 14433 29236 14467
rect 29184 14424 29236 14433
rect 30564 14424 30616 14476
rect 30840 14424 30892 14476
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 7196 14356 7248 14408
rect 12164 14356 12216 14408
rect 13636 14356 13688 14408
rect 15384 14356 15436 14408
rect 7748 14288 7800 14340
rect 12440 14331 12492 14340
rect 12440 14297 12449 14331
rect 12449 14297 12483 14331
rect 12483 14297 12492 14331
rect 12440 14288 12492 14297
rect 15936 14288 15988 14340
rect 16120 14331 16172 14340
rect 16120 14297 16129 14331
rect 16129 14297 16163 14331
rect 16163 14297 16172 14331
rect 16120 14288 16172 14297
rect 18604 14356 18656 14408
rect 20076 14356 20128 14408
rect 20444 14288 20496 14340
rect 20812 14288 20864 14340
rect 940 14220 992 14272
rect 19800 14220 19852 14272
rect 21732 14263 21784 14272
rect 21732 14229 21741 14263
rect 21741 14229 21775 14263
rect 21775 14229 21784 14263
rect 21732 14220 21784 14229
rect 22100 14263 22152 14272
rect 22100 14229 22109 14263
rect 22109 14229 22143 14263
rect 22143 14229 22152 14263
rect 22100 14220 22152 14229
rect 22744 14220 22796 14272
rect 23664 14331 23716 14340
rect 23664 14297 23673 14331
rect 23673 14297 23707 14331
rect 23707 14297 23716 14331
rect 23664 14288 23716 14297
rect 25596 14399 25648 14408
rect 25596 14365 25605 14399
rect 25605 14365 25639 14399
rect 25639 14365 25648 14399
rect 25596 14356 25648 14365
rect 25872 14288 25924 14340
rect 24308 14220 24360 14272
rect 24768 14263 24820 14272
rect 24768 14229 24777 14263
rect 24777 14229 24811 14263
rect 24811 14229 24820 14263
rect 24768 14220 24820 14229
rect 24860 14263 24912 14272
rect 24860 14229 24869 14263
rect 24869 14229 24903 14263
rect 24903 14229 24912 14263
rect 24860 14220 24912 14229
rect 25412 14263 25464 14272
rect 25412 14229 25421 14263
rect 25421 14229 25455 14263
rect 25455 14229 25464 14263
rect 25412 14220 25464 14229
rect 26148 14399 26200 14408
rect 26148 14365 26157 14399
rect 26157 14365 26191 14399
rect 26191 14365 26200 14399
rect 26148 14356 26200 14365
rect 26884 14399 26936 14408
rect 26884 14365 26893 14399
rect 26893 14365 26927 14399
rect 26927 14365 26936 14399
rect 26884 14356 26936 14365
rect 27160 14399 27212 14408
rect 27160 14365 27169 14399
rect 27169 14365 27203 14399
rect 27203 14365 27212 14399
rect 27160 14356 27212 14365
rect 29552 14399 29604 14408
rect 29552 14365 29561 14399
rect 29561 14365 29595 14399
rect 29595 14365 29604 14399
rect 29552 14356 29604 14365
rect 31852 14424 31904 14476
rect 32036 14467 32088 14476
rect 32036 14433 32045 14467
rect 32045 14433 32079 14467
rect 32079 14433 32088 14467
rect 32036 14424 32088 14433
rect 32496 14424 32548 14476
rect 34244 14424 34296 14476
rect 37740 14424 37792 14476
rect 38476 14424 38528 14476
rect 40592 14467 40644 14476
rect 40592 14433 40601 14467
rect 40601 14433 40635 14467
rect 40635 14433 40644 14467
rect 40592 14424 40644 14433
rect 30748 14288 30800 14340
rect 35256 14288 35308 14340
rect 26976 14220 27028 14272
rect 27160 14220 27212 14272
rect 28632 14220 28684 14272
rect 31024 14263 31076 14272
rect 31024 14229 31033 14263
rect 31033 14229 31067 14263
rect 31067 14229 31076 14263
rect 31024 14220 31076 14229
rect 31852 14263 31904 14272
rect 31852 14229 31861 14263
rect 31861 14229 31895 14263
rect 31895 14229 31904 14263
rect 31852 14220 31904 14229
rect 34520 14220 34572 14272
rect 35900 14356 35952 14408
rect 38568 14356 38620 14408
rect 39856 14399 39908 14408
rect 39856 14365 39865 14399
rect 39865 14365 39899 14399
rect 39899 14365 39908 14399
rect 39856 14356 39908 14365
rect 40132 14356 40184 14408
rect 40224 14356 40276 14408
rect 40960 14399 41012 14408
rect 40960 14365 40974 14399
rect 40974 14365 41008 14399
rect 41008 14365 41012 14399
rect 40960 14356 41012 14365
rect 36084 14331 36136 14340
rect 36084 14297 36118 14331
rect 36118 14297 36136 14331
rect 36084 14288 36136 14297
rect 37832 14220 37884 14272
rect 38108 14288 38160 14340
rect 43720 14424 43772 14476
rect 45192 14356 45244 14408
rect 38476 14220 38528 14272
rect 40500 14220 40552 14272
rect 40684 14220 40736 14272
rect 43076 14220 43128 14272
rect 44180 14220 44232 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 19708 14016 19760 14068
rect 22100 14016 22152 14068
rect 10232 13991 10284 14000
rect 10232 13957 10241 13991
rect 10241 13957 10275 13991
rect 10275 13957 10284 13991
rect 10232 13948 10284 13957
rect 13360 13948 13412 14000
rect 14648 13948 14700 14000
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 9680 13880 9732 13932
rect 11060 13880 11112 13932
rect 12624 13923 12676 13932
rect 12624 13889 12633 13923
rect 12633 13889 12667 13923
rect 12667 13889 12676 13923
rect 12624 13880 12676 13889
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 19524 13948 19576 14000
rect 19800 13880 19852 13932
rect 20260 13880 20312 13932
rect 20444 13948 20496 14000
rect 23388 14016 23440 14068
rect 24768 14016 24820 14068
rect 31024 14016 31076 14068
rect 12440 13812 12492 13864
rect 19248 13812 19300 13864
rect 25412 13991 25464 14000
rect 25412 13957 25446 13991
rect 25446 13957 25464 13991
rect 25412 13948 25464 13957
rect 27160 13948 27212 14000
rect 26884 13880 26936 13932
rect 25044 13812 25096 13864
rect 26148 13812 26200 13864
rect 7748 13744 7800 13796
rect 8024 13744 8076 13796
rect 12716 13744 12768 13796
rect 22744 13787 22796 13796
rect 22744 13753 22753 13787
rect 22753 13753 22787 13787
rect 22787 13753 22796 13787
rect 22744 13744 22796 13753
rect 26976 13855 27028 13864
rect 26976 13821 26985 13855
rect 26985 13821 27019 13855
rect 27019 13821 27028 13855
rect 26976 13812 27028 13821
rect 27160 13855 27212 13864
rect 27160 13821 27169 13855
rect 27169 13821 27203 13855
rect 27203 13821 27212 13855
rect 27160 13812 27212 13821
rect 28172 13923 28224 13932
rect 28172 13889 28181 13923
rect 28181 13889 28215 13923
rect 28215 13889 28224 13923
rect 28172 13880 28224 13889
rect 29276 13923 29328 13932
rect 29276 13889 29285 13923
rect 29285 13889 29319 13923
rect 29319 13889 29328 13923
rect 29276 13880 29328 13889
rect 30656 13923 30708 13932
rect 30656 13889 30665 13923
rect 30665 13889 30699 13923
rect 30699 13889 30708 13923
rect 30656 13880 30708 13889
rect 30748 13923 30800 13932
rect 30748 13889 30782 13923
rect 30782 13889 30800 13923
rect 30748 13880 30800 13889
rect 32496 14059 32548 14068
rect 32496 14025 32505 14059
rect 32505 14025 32539 14059
rect 32539 14025 32548 14059
rect 32496 14016 32548 14025
rect 35256 14059 35308 14068
rect 35256 14025 35265 14059
rect 35265 14025 35299 14059
rect 35299 14025 35308 14059
rect 35256 14016 35308 14025
rect 37648 14059 37700 14068
rect 37648 14025 37657 14059
rect 37657 14025 37691 14059
rect 37691 14025 37700 14059
rect 37648 14016 37700 14025
rect 37832 14016 37884 14068
rect 40132 14059 40184 14068
rect 40132 14025 40141 14059
rect 40141 14025 40175 14059
rect 40175 14025 40184 14059
rect 40132 14016 40184 14025
rect 40960 14016 41012 14068
rect 42984 14059 43036 14068
rect 42984 14025 42993 14059
rect 42993 14025 43027 14059
rect 43027 14025 43036 14059
rect 42984 14016 43036 14025
rect 40500 13948 40552 14000
rect 27988 13855 28040 13864
rect 27988 13821 28022 13855
rect 28022 13821 28040 13855
rect 27988 13812 28040 13821
rect 28724 13812 28776 13864
rect 27712 13744 27764 13796
rect 29644 13744 29696 13796
rect 30104 13812 30156 13864
rect 30012 13744 30064 13796
rect 30380 13787 30432 13796
rect 30380 13753 30389 13787
rect 30389 13753 30423 13787
rect 30423 13753 30432 13787
rect 30380 13744 30432 13753
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 9312 13719 9364 13728
rect 9312 13685 9321 13719
rect 9321 13685 9355 13719
rect 9355 13685 9364 13719
rect 9312 13676 9364 13685
rect 10324 13719 10376 13728
rect 10324 13685 10333 13719
rect 10333 13685 10367 13719
rect 10367 13685 10376 13719
rect 10324 13676 10376 13685
rect 15016 13676 15068 13728
rect 24584 13676 24636 13728
rect 26516 13719 26568 13728
rect 26516 13685 26525 13719
rect 26525 13685 26559 13719
rect 26559 13685 26568 13719
rect 26516 13676 26568 13685
rect 27068 13676 27120 13728
rect 27988 13676 28040 13728
rect 28908 13719 28960 13728
rect 28908 13685 28917 13719
rect 28917 13685 28951 13719
rect 28951 13685 28960 13719
rect 28908 13676 28960 13685
rect 31116 13812 31168 13864
rect 33232 13880 33284 13932
rect 33324 13880 33376 13932
rect 32680 13855 32732 13864
rect 32680 13821 32689 13855
rect 32689 13821 32723 13855
rect 32723 13821 32732 13855
rect 32680 13812 32732 13821
rect 33508 13812 33560 13864
rect 34612 13923 34664 13932
rect 34612 13889 34621 13923
rect 34621 13889 34655 13923
rect 34655 13889 34664 13923
rect 34612 13880 34664 13889
rect 36268 13880 36320 13932
rect 40684 13880 40736 13932
rect 41144 13923 41196 13932
rect 41144 13889 41153 13923
rect 41153 13889 41187 13923
rect 41187 13889 41196 13923
rect 41144 13880 41196 13889
rect 42248 13880 42300 13932
rect 43076 13923 43128 13932
rect 43076 13889 43085 13923
rect 43085 13889 43119 13923
rect 43119 13889 43128 13923
rect 43076 13880 43128 13889
rect 33968 13812 34020 13864
rect 34152 13812 34204 13864
rect 34428 13855 34480 13864
rect 34428 13821 34462 13855
rect 34462 13821 34480 13855
rect 34428 13812 34480 13821
rect 35716 13855 35768 13864
rect 35716 13821 35725 13855
rect 35725 13821 35759 13855
rect 35759 13821 35768 13855
rect 35716 13812 35768 13821
rect 33876 13744 33928 13796
rect 37004 13744 37056 13796
rect 40960 13855 41012 13864
rect 40960 13821 40969 13855
rect 40969 13821 41003 13855
rect 41003 13821 41012 13855
rect 40960 13812 41012 13821
rect 43168 13812 43220 13864
rect 44180 13923 44232 13932
rect 44180 13889 44189 13923
rect 44189 13889 44223 13923
rect 44223 13889 44232 13923
rect 44180 13880 44232 13889
rect 45192 13880 45244 13932
rect 46848 13812 46900 13864
rect 31944 13676 31996 13728
rect 33416 13676 33468 13728
rect 35348 13676 35400 13728
rect 37096 13719 37148 13728
rect 37096 13685 37105 13719
rect 37105 13685 37139 13719
rect 37139 13685 37148 13719
rect 37096 13676 37148 13685
rect 37280 13719 37332 13728
rect 37280 13685 37289 13719
rect 37289 13685 37323 13719
rect 37323 13685 37332 13719
rect 37280 13676 37332 13685
rect 42800 13719 42852 13728
rect 42800 13685 42809 13719
rect 42809 13685 42843 13719
rect 42843 13685 42852 13719
rect 42800 13676 42852 13685
rect 43260 13676 43312 13728
rect 45376 13676 45428 13728
rect 45468 13719 45520 13728
rect 45468 13685 45477 13719
rect 45477 13685 45511 13719
rect 45511 13685 45520 13719
rect 45468 13676 45520 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 8944 13336 8996 13388
rect 17776 13472 17828 13524
rect 18696 13472 18748 13524
rect 20260 13515 20312 13524
rect 20260 13481 20269 13515
rect 20269 13481 20303 13515
rect 20303 13481 20312 13515
rect 20260 13472 20312 13481
rect 20904 13472 20956 13524
rect 21364 13472 21416 13524
rect 14648 13404 14700 13456
rect 24216 13515 24268 13524
rect 24216 13481 24225 13515
rect 24225 13481 24259 13515
rect 24259 13481 24268 13515
rect 24216 13472 24268 13481
rect 25596 13472 25648 13524
rect 27160 13472 27212 13524
rect 28724 13472 28776 13524
rect 29644 13472 29696 13524
rect 31024 13472 31076 13524
rect 31852 13472 31904 13524
rect 33232 13515 33284 13524
rect 33232 13481 33241 13515
rect 33241 13481 33275 13515
rect 33275 13481 33284 13515
rect 33232 13472 33284 13481
rect 26332 13404 26384 13456
rect 14280 13336 14332 13388
rect 4436 13311 4488 13320
rect 4436 13277 4445 13311
rect 4445 13277 4479 13311
rect 4479 13277 4488 13311
rect 4436 13268 4488 13277
rect 10324 13268 10376 13320
rect 10416 13268 10468 13320
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 14648 13311 14700 13320
rect 14648 13277 14657 13311
rect 14657 13277 14691 13311
rect 14691 13277 14700 13311
rect 14648 13268 14700 13277
rect 15016 13311 15068 13320
rect 15016 13277 15050 13311
rect 15050 13277 15068 13311
rect 15016 13268 15068 13277
rect 16672 13268 16724 13320
rect 20076 13268 20128 13320
rect 21732 13336 21784 13388
rect 20904 13311 20956 13320
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 21180 13311 21232 13320
rect 21180 13277 21189 13311
rect 21189 13277 21223 13311
rect 21223 13277 21232 13311
rect 21180 13268 21232 13277
rect 21916 13268 21968 13320
rect 6920 13200 6972 13252
rect 4252 13175 4304 13184
rect 4252 13141 4261 13175
rect 4261 13141 4295 13175
rect 4295 13141 4304 13175
rect 4252 13132 4304 13141
rect 6552 13132 6604 13184
rect 7840 13175 7892 13184
rect 7840 13141 7849 13175
rect 7849 13141 7883 13175
rect 7883 13141 7892 13175
rect 7840 13132 7892 13141
rect 10692 13175 10744 13184
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 10692 13132 10744 13141
rect 16948 13200 17000 13252
rect 11888 13132 11940 13184
rect 13820 13132 13872 13184
rect 14556 13132 14608 13184
rect 16120 13175 16172 13184
rect 16120 13141 16129 13175
rect 16129 13141 16163 13175
rect 16163 13141 16172 13175
rect 18144 13200 18196 13252
rect 20628 13200 20680 13252
rect 16120 13132 16172 13141
rect 17316 13132 17368 13184
rect 19156 13132 19208 13184
rect 21088 13175 21140 13184
rect 21088 13141 21097 13175
rect 21097 13141 21131 13175
rect 21131 13141 21140 13175
rect 21088 13132 21140 13141
rect 21640 13200 21692 13252
rect 23572 13379 23624 13388
rect 23572 13345 23581 13379
rect 23581 13345 23615 13379
rect 23615 13345 23624 13379
rect 23572 13336 23624 13345
rect 24676 13336 24728 13388
rect 25964 13336 26016 13388
rect 26700 13336 26752 13388
rect 22560 13311 22612 13320
rect 22560 13277 22569 13311
rect 22569 13277 22603 13311
rect 22603 13277 22612 13311
rect 22560 13268 22612 13277
rect 23296 13311 23348 13320
rect 23296 13277 23305 13311
rect 23305 13277 23339 13311
rect 23339 13277 23348 13311
rect 23296 13268 23348 13277
rect 23388 13311 23440 13320
rect 23388 13277 23422 13311
rect 23422 13277 23440 13311
rect 23388 13268 23440 13277
rect 25504 13268 25556 13320
rect 26516 13268 26568 13320
rect 23020 13132 23072 13184
rect 24676 13132 24728 13184
rect 25044 13200 25096 13252
rect 27436 13404 27488 13456
rect 29552 13404 29604 13456
rect 30288 13404 30340 13456
rect 33140 13404 33192 13456
rect 27528 13268 27580 13320
rect 29828 13336 29880 13388
rect 30104 13379 30156 13388
rect 30104 13345 30113 13379
rect 30113 13345 30147 13379
rect 30147 13345 30156 13379
rect 30104 13336 30156 13345
rect 30656 13336 30708 13388
rect 30932 13379 30984 13388
rect 30932 13345 30966 13379
rect 30966 13345 30984 13379
rect 30932 13336 30984 13345
rect 31300 13336 31352 13388
rect 31668 13336 31720 13388
rect 27712 13243 27764 13252
rect 27712 13209 27746 13243
rect 27746 13209 27764 13243
rect 27712 13200 27764 13209
rect 25780 13132 25832 13184
rect 26332 13132 26384 13184
rect 28724 13132 28776 13184
rect 30012 13268 30064 13320
rect 31944 13268 31996 13320
rect 34244 13379 34296 13388
rect 34244 13345 34253 13379
rect 34253 13345 34287 13379
rect 34287 13345 34296 13379
rect 34244 13336 34296 13345
rect 34336 13379 34388 13388
rect 34336 13345 34345 13379
rect 34345 13345 34379 13379
rect 34379 13345 34388 13379
rect 34336 13336 34388 13345
rect 33416 13132 33468 13184
rect 36268 13472 36320 13524
rect 36360 13472 36412 13524
rect 46112 13472 46164 13524
rect 43720 13404 43772 13456
rect 37004 13336 37056 13388
rect 37096 13268 37148 13320
rect 37556 13268 37608 13320
rect 38384 13268 38436 13320
rect 42524 13268 42576 13320
rect 43260 13311 43312 13320
rect 43260 13277 43269 13311
rect 43269 13277 43303 13311
rect 43303 13277 43312 13311
rect 43260 13268 43312 13277
rect 45468 13311 45520 13320
rect 45468 13277 45477 13311
rect 45477 13277 45511 13311
rect 45511 13277 45520 13311
rect 45468 13268 45520 13277
rect 46204 13268 46256 13320
rect 33876 13200 33928 13252
rect 33968 13132 34020 13184
rect 34336 13132 34388 13184
rect 38016 13200 38068 13252
rect 36636 13175 36688 13184
rect 36636 13141 36645 13175
rect 36645 13141 36679 13175
rect 36679 13141 36688 13175
rect 36636 13132 36688 13141
rect 37464 13175 37516 13184
rect 37464 13141 37473 13175
rect 37473 13141 37507 13175
rect 37507 13141 37516 13175
rect 37464 13132 37516 13141
rect 43076 13132 43128 13184
rect 43260 13132 43312 13184
rect 45100 13132 45152 13184
rect 46664 13175 46716 13184
rect 46664 13141 46673 13175
rect 46673 13141 46707 13175
rect 46707 13141 46716 13175
rect 46664 13132 46716 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 4436 12928 4488 12980
rect 7656 12928 7708 12980
rect 9864 12928 9916 12980
rect 4252 12860 4304 12912
rect 1492 12835 1544 12844
rect 1492 12801 1501 12835
rect 1501 12801 1535 12835
rect 1535 12801 1544 12835
rect 1492 12792 1544 12801
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 3700 12767 3752 12776
rect 3700 12733 3709 12767
rect 3709 12733 3743 12767
rect 3743 12733 3752 12767
rect 3700 12724 3752 12733
rect 5632 12767 5684 12776
rect 5632 12733 5641 12767
rect 5641 12733 5675 12767
rect 5675 12733 5684 12767
rect 5632 12724 5684 12733
rect 6276 12860 6328 12912
rect 6460 12860 6512 12912
rect 9312 12860 9364 12912
rect 6736 12792 6788 12844
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 6000 12724 6052 12776
rect 6552 12767 6604 12776
rect 6552 12733 6561 12767
rect 6561 12733 6595 12767
rect 6595 12733 6604 12767
rect 6552 12724 6604 12733
rect 7380 12767 7432 12776
rect 7380 12733 7414 12767
rect 7414 12733 7432 12767
rect 7380 12724 7432 12733
rect 7748 12724 7800 12776
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 10692 12928 10744 12980
rect 10968 12860 11020 12912
rect 11704 12928 11756 12980
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 13820 12928 13872 12937
rect 15292 12928 15344 12980
rect 16120 12971 16172 12980
rect 16120 12937 16129 12971
rect 16129 12937 16163 12971
rect 16163 12937 16172 12971
rect 16120 12928 16172 12937
rect 16948 12928 17000 12980
rect 11612 12792 11664 12844
rect 11888 12792 11940 12844
rect 12716 12835 12768 12844
rect 12716 12801 12725 12835
rect 12725 12801 12759 12835
rect 12759 12801 12768 12835
rect 12716 12792 12768 12801
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 14556 12835 14608 12844
rect 14556 12801 14590 12835
rect 14590 12801 14608 12835
rect 14556 12792 14608 12801
rect 19156 12928 19208 12980
rect 24676 12928 24728 12980
rect 24860 12971 24912 12980
rect 24860 12937 24869 12971
rect 24869 12937 24903 12971
rect 24903 12937 24912 12971
rect 24860 12928 24912 12937
rect 24952 12928 25004 12980
rect 29920 12928 29972 12980
rect 30748 12928 30800 12980
rect 20168 12860 20220 12912
rect 33140 12928 33192 12980
rect 17316 12835 17368 12844
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 18144 12835 18196 12844
rect 18144 12801 18178 12835
rect 18178 12801 18196 12835
rect 18144 12792 18196 12801
rect 18328 12835 18380 12844
rect 18328 12801 18337 12835
rect 18337 12801 18371 12835
rect 18371 12801 18380 12835
rect 18328 12792 18380 12801
rect 19708 12792 19760 12844
rect 20904 12835 20956 12844
rect 20904 12801 20913 12835
rect 20913 12801 20947 12835
rect 20947 12801 20956 12835
rect 20904 12792 20956 12801
rect 6552 12588 6604 12640
rect 7472 12588 7524 12640
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 10324 12631 10376 12640
rect 10324 12597 10333 12631
rect 10333 12597 10367 12631
rect 10367 12597 10376 12631
rect 12624 12724 12676 12776
rect 13912 12767 13964 12776
rect 13912 12733 13921 12767
rect 13921 12733 13955 12767
rect 13955 12733 13964 12767
rect 13912 12724 13964 12733
rect 14004 12767 14056 12776
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 16212 12767 16264 12776
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 16212 12724 16264 12733
rect 16488 12724 16540 12776
rect 16948 12724 17000 12776
rect 17500 12724 17552 12776
rect 17776 12767 17828 12776
rect 17776 12733 17785 12767
rect 17785 12733 17819 12767
rect 17819 12733 17828 12767
rect 17776 12724 17828 12733
rect 17868 12724 17920 12776
rect 18880 12724 18932 12776
rect 19340 12724 19392 12776
rect 10324 12588 10376 12597
rect 12532 12588 12584 12640
rect 15660 12631 15712 12640
rect 15660 12597 15669 12631
rect 15669 12597 15703 12631
rect 15703 12597 15712 12631
rect 15660 12588 15712 12597
rect 21180 12835 21232 12844
rect 21180 12801 21189 12835
rect 21189 12801 21223 12835
rect 21223 12801 21232 12835
rect 21180 12792 21232 12801
rect 22560 12792 22612 12844
rect 23020 12767 23072 12776
rect 23020 12733 23029 12767
rect 23029 12733 23063 12767
rect 23063 12733 23072 12767
rect 23020 12724 23072 12733
rect 23296 12724 23348 12776
rect 23940 12767 23992 12776
rect 23940 12733 23949 12767
rect 23949 12733 23983 12767
rect 23983 12733 23992 12767
rect 23940 12724 23992 12733
rect 24032 12767 24084 12776
rect 24032 12733 24066 12767
rect 24066 12733 24084 12767
rect 24032 12724 24084 12733
rect 24584 12724 24636 12776
rect 25964 12792 26016 12844
rect 27712 12792 27764 12844
rect 28908 12792 28960 12844
rect 29092 12835 29144 12844
rect 29092 12801 29126 12835
rect 29126 12801 29144 12835
rect 29092 12792 29144 12801
rect 31024 12860 31076 12912
rect 32680 12860 32732 12912
rect 30104 12792 30156 12844
rect 30288 12792 30340 12844
rect 30380 12792 30432 12844
rect 33876 12928 33928 12980
rect 34520 12928 34572 12980
rect 36084 12971 36136 12980
rect 36084 12937 36093 12971
rect 36093 12937 36127 12971
rect 36127 12937 36136 12971
rect 36084 12928 36136 12937
rect 39856 12928 39908 12980
rect 43168 12928 43220 12980
rect 20352 12631 20404 12640
rect 20352 12597 20361 12631
rect 20361 12597 20395 12631
rect 20395 12597 20404 12631
rect 20352 12588 20404 12597
rect 23204 12588 23256 12640
rect 23664 12699 23716 12708
rect 23664 12665 23673 12699
rect 23673 12665 23707 12699
rect 23707 12665 23716 12699
rect 23664 12656 23716 12665
rect 27804 12724 27856 12776
rect 28632 12724 28684 12776
rect 29920 12724 29972 12776
rect 24768 12656 24820 12708
rect 24952 12631 25004 12640
rect 24952 12597 24961 12631
rect 24961 12597 24995 12631
rect 24995 12597 25004 12631
rect 24952 12588 25004 12597
rect 27620 12656 27672 12708
rect 29828 12656 29880 12708
rect 33508 12724 33560 12776
rect 34152 12835 34204 12844
rect 34152 12801 34161 12835
rect 34161 12801 34195 12835
rect 34195 12801 34204 12835
rect 34152 12792 34204 12801
rect 34336 12792 34388 12844
rect 37280 12792 37332 12844
rect 39212 12835 39264 12844
rect 39212 12801 39221 12835
rect 39221 12801 39255 12835
rect 39255 12801 39264 12835
rect 39212 12792 39264 12801
rect 33784 12724 33836 12776
rect 33968 12724 34020 12776
rect 31484 12588 31536 12640
rect 33232 12656 33284 12708
rect 39580 12835 39632 12844
rect 39580 12801 39589 12835
rect 39589 12801 39623 12835
rect 39623 12801 39632 12835
rect 39580 12792 39632 12801
rect 39948 12792 40000 12844
rect 45100 12835 45152 12844
rect 45100 12801 45109 12835
rect 45109 12801 45143 12835
rect 45143 12801 45152 12835
rect 45100 12792 45152 12801
rect 39948 12656 40000 12708
rect 40960 12724 41012 12776
rect 41052 12724 41104 12776
rect 42800 12724 42852 12776
rect 43076 12767 43128 12776
rect 43076 12733 43085 12767
rect 43085 12733 43119 12767
rect 43119 12733 43128 12767
rect 43076 12724 43128 12733
rect 43168 12767 43220 12776
rect 43168 12733 43177 12767
rect 43177 12733 43211 12767
rect 43211 12733 43220 12767
rect 43168 12724 43220 12733
rect 44916 12767 44968 12776
rect 44916 12733 44925 12767
rect 44925 12733 44959 12767
rect 44959 12733 44968 12767
rect 44916 12724 44968 12733
rect 41604 12656 41656 12708
rect 36636 12588 36688 12640
rect 40040 12588 40092 12640
rect 43536 12588 43588 12640
rect 44088 12588 44140 12640
rect 44548 12588 44600 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 5264 12384 5316 12436
rect 6920 12384 6972 12436
rect 7104 12384 7156 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 14648 12384 14700 12436
rect 15660 12384 15712 12436
rect 17868 12384 17920 12436
rect 20352 12384 20404 12436
rect 11060 12316 11112 12368
rect 12256 12359 12308 12368
rect 12256 12325 12265 12359
rect 12265 12325 12299 12359
rect 12299 12325 12308 12359
rect 12256 12316 12308 12325
rect 17408 12316 17460 12368
rect 3700 12248 3752 12300
rect 6000 12291 6052 12300
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6000 12248 6052 12257
rect 6460 12291 6512 12300
rect 6460 12257 6469 12291
rect 6469 12257 6503 12291
rect 6503 12257 6512 12291
rect 6460 12248 6512 12257
rect 6552 12248 6604 12300
rect 6920 12248 6972 12300
rect 7380 12248 7432 12300
rect 8024 12248 8076 12300
rect 8484 12248 8536 12300
rect 10416 12248 10468 12300
rect 11612 12291 11664 12300
rect 11612 12257 11621 12291
rect 11621 12257 11655 12291
rect 11655 12257 11664 12291
rect 11612 12248 11664 12257
rect 11888 12248 11940 12300
rect 12532 12291 12584 12300
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 12532 12248 12584 12257
rect 12624 12291 12676 12300
rect 12624 12257 12658 12291
rect 12658 12257 12676 12291
rect 12624 12248 12676 12257
rect 15108 12291 15160 12300
rect 15108 12257 15117 12291
rect 15117 12257 15151 12291
rect 15151 12257 15160 12291
rect 15108 12248 15160 12257
rect 16948 12291 17000 12300
rect 16948 12257 16957 12291
rect 16957 12257 16991 12291
rect 16991 12257 17000 12291
rect 16948 12248 17000 12257
rect 17316 12248 17368 12300
rect 17684 12248 17736 12300
rect 17868 12291 17920 12300
rect 17868 12257 17877 12291
rect 17877 12257 17911 12291
rect 17911 12257 17920 12291
rect 17868 12248 17920 12257
rect 18052 12248 18104 12300
rect 19064 12248 19116 12300
rect 19248 12248 19300 12300
rect 4160 12112 4212 12164
rect 7012 12223 7064 12232
rect 7012 12189 7021 12223
rect 7021 12189 7055 12223
rect 7055 12189 7064 12223
rect 7012 12180 7064 12189
rect 7840 12180 7892 12232
rect 10324 12180 10376 12232
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 15660 12180 15712 12232
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 19524 12223 19576 12232
rect 19524 12189 19533 12223
rect 19533 12189 19567 12223
rect 19567 12189 19576 12223
rect 19524 12180 19576 12189
rect 19892 12223 19944 12232
rect 19892 12189 19901 12223
rect 19901 12189 19935 12223
rect 19935 12189 19944 12223
rect 19892 12180 19944 12189
rect 6736 12044 6788 12096
rect 8208 12087 8260 12096
rect 8208 12053 8217 12087
rect 8217 12053 8251 12087
rect 8251 12053 8260 12087
rect 8208 12044 8260 12053
rect 10968 12044 11020 12096
rect 14464 12044 14516 12096
rect 16212 12044 16264 12096
rect 18696 12044 18748 12096
rect 23388 12316 23440 12368
rect 24032 12316 24084 12368
rect 25780 12427 25832 12436
rect 25780 12393 25789 12427
rect 25789 12393 25823 12427
rect 25823 12393 25832 12427
rect 25780 12384 25832 12393
rect 25964 12384 26016 12436
rect 33692 12384 33744 12436
rect 22928 12248 22980 12300
rect 22468 12180 22520 12232
rect 22744 12180 22796 12232
rect 23296 12180 23348 12232
rect 22008 12112 22060 12164
rect 24492 12180 24544 12232
rect 24676 12223 24728 12232
rect 24676 12189 24710 12223
rect 24710 12189 24728 12223
rect 24676 12180 24728 12189
rect 25504 12180 25556 12232
rect 20720 12044 20772 12096
rect 23112 12087 23164 12096
rect 23112 12053 23121 12087
rect 23121 12053 23155 12087
rect 23155 12053 23164 12087
rect 23112 12044 23164 12053
rect 23480 12087 23532 12096
rect 23480 12053 23489 12087
rect 23489 12053 23523 12087
rect 23523 12053 23532 12087
rect 23480 12044 23532 12053
rect 25044 12112 25096 12164
rect 25872 12155 25924 12164
rect 25872 12121 25881 12155
rect 25881 12121 25915 12155
rect 25915 12121 25924 12155
rect 25872 12112 25924 12121
rect 25504 12044 25556 12096
rect 26700 12044 26752 12096
rect 26792 12044 26844 12096
rect 27252 12112 27304 12164
rect 30472 12316 30524 12368
rect 36452 12359 36504 12368
rect 36452 12325 36461 12359
rect 36461 12325 36495 12359
rect 36495 12325 36504 12359
rect 36452 12316 36504 12325
rect 30288 12248 30340 12300
rect 29920 12180 29972 12232
rect 32772 12180 32824 12232
rect 33600 12112 33652 12164
rect 29276 12044 29328 12096
rect 33692 12044 33744 12096
rect 36544 12180 36596 12232
rect 36728 12180 36780 12232
rect 38752 12384 38804 12436
rect 38844 12384 38896 12436
rect 39212 12384 39264 12436
rect 40040 12427 40092 12436
rect 40040 12393 40049 12427
rect 40049 12393 40083 12427
rect 40083 12393 40092 12427
rect 40040 12384 40092 12393
rect 41604 12427 41656 12436
rect 41604 12393 41613 12427
rect 41613 12393 41647 12427
rect 41647 12393 41656 12427
rect 41604 12384 41656 12393
rect 41696 12384 41748 12436
rect 39488 12316 39540 12368
rect 40868 12316 40920 12368
rect 43076 12384 43128 12436
rect 38016 12248 38068 12300
rect 44088 12316 44140 12368
rect 37464 12044 37516 12096
rect 38844 12180 38896 12232
rect 39120 12112 39172 12164
rect 39764 12180 39816 12232
rect 40408 12180 40460 12232
rect 41696 12180 41748 12232
rect 42248 12223 42300 12232
rect 42248 12189 42257 12223
rect 42257 12189 42291 12223
rect 42291 12189 42300 12223
rect 42248 12180 42300 12189
rect 38844 12087 38896 12096
rect 38844 12053 38853 12087
rect 38853 12053 38887 12087
rect 38887 12053 38896 12087
rect 38844 12044 38896 12053
rect 38936 12044 38988 12096
rect 41052 12112 41104 12164
rect 42708 12180 42760 12232
rect 43352 12248 43404 12300
rect 43628 12180 43680 12232
rect 43812 12223 43864 12232
rect 43812 12189 43821 12223
rect 43821 12189 43855 12223
rect 43855 12189 43864 12223
rect 43812 12180 43864 12189
rect 43996 12180 44048 12232
rect 44180 12223 44232 12232
rect 44180 12189 44189 12223
rect 44189 12189 44223 12223
rect 44223 12189 44232 12223
rect 44180 12180 44232 12189
rect 44548 12223 44600 12232
rect 44548 12189 44557 12223
rect 44557 12189 44591 12223
rect 44591 12189 44600 12223
rect 44548 12180 44600 12189
rect 43168 12112 43220 12164
rect 43260 12112 43312 12164
rect 40224 12087 40276 12096
rect 40224 12053 40233 12087
rect 40233 12053 40267 12087
rect 40267 12053 40276 12087
rect 40224 12044 40276 12053
rect 41420 12087 41472 12096
rect 41420 12053 41429 12087
rect 41429 12053 41463 12087
rect 41463 12053 41472 12087
rect 41420 12044 41472 12053
rect 43536 12044 43588 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 4160 11883 4212 11892
rect 4160 11849 4169 11883
rect 4169 11849 4203 11883
rect 4203 11849 4212 11883
rect 4160 11840 4212 11849
rect 5264 11840 5316 11892
rect 8208 11840 8260 11892
rect 12624 11840 12676 11892
rect 19524 11840 19576 11892
rect 21272 11840 21324 11892
rect 22008 11883 22060 11892
rect 22008 11849 22017 11883
rect 22017 11849 22051 11883
rect 22051 11849 22060 11883
rect 22008 11840 22060 11849
rect 23940 11840 23992 11892
rect 7012 11772 7064 11824
rect 8852 11772 8904 11824
rect 23296 11772 23348 11824
rect 23848 11772 23900 11824
rect 25964 11772 26016 11824
rect 26700 11840 26752 11892
rect 5632 11704 5684 11756
rect 5632 11500 5684 11552
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 8944 11704 8996 11756
rect 9312 11747 9364 11756
rect 9312 11713 9346 11747
rect 9346 11713 9364 11747
rect 9312 11704 9364 11713
rect 10968 11747 11020 11756
rect 10968 11713 10977 11747
rect 10977 11713 11011 11747
rect 11011 11713 11020 11747
rect 10968 11704 11020 11713
rect 14188 11704 14240 11756
rect 23112 11704 23164 11756
rect 7656 11636 7708 11688
rect 26792 11747 26844 11756
rect 26792 11713 26801 11747
rect 26801 11713 26835 11747
rect 26835 11713 26844 11747
rect 26792 11704 26844 11713
rect 24492 11636 24544 11688
rect 27528 11704 27580 11756
rect 29276 11704 29328 11756
rect 31852 11840 31904 11892
rect 30012 11772 30064 11824
rect 31576 11815 31628 11824
rect 31576 11781 31585 11815
rect 31585 11781 31619 11815
rect 31619 11781 31628 11815
rect 31576 11772 31628 11781
rect 34244 11883 34296 11892
rect 34244 11849 34253 11883
rect 34253 11849 34287 11883
rect 34287 11849 34296 11883
rect 34244 11840 34296 11849
rect 38016 11883 38068 11892
rect 38016 11849 38025 11883
rect 38025 11849 38059 11883
rect 38059 11849 38068 11883
rect 38016 11840 38068 11849
rect 34336 11772 34388 11824
rect 29828 11704 29880 11756
rect 30196 11747 30248 11756
rect 30196 11713 30205 11747
rect 30205 11713 30239 11747
rect 30239 11713 30248 11747
rect 30196 11704 30248 11713
rect 30380 11704 30432 11756
rect 31392 11704 31444 11756
rect 32496 11704 32548 11756
rect 34152 11747 34204 11756
rect 34152 11713 34161 11747
rect 34161 11713 34195 11747
rect 34195 11713 34204 11747
rect 34152 11704 34204 11713
rect 37832 11772 37884 11824
rect 30564 11636 30616 11688
rect 33600 11679 33652 11688
rect 33600 11645 33609 11679
rect 33609 11645 33643 11679
rect 33643 11645 33652 11679
rect 33600 11636 33652 11645
rect 33692 11636 33744 11688
rect 38476 11704 38528 11756
rect 41420 11840 41472 11892
rect 41696 11840 41748 11892
rect 38844 11772 38896 11824
rect 43168 11840 43220 11892
rect 39396 11704 39448 11756
rect 6460 11568 6512 11620
rect 8300 11568 8352 11620
rect 10968 11568 11020 11620
rect 7564 11500 7616 11552
rect 10508 11543 10560 11552
rect 10508 11509 10517 11543
rect 10517 11509 10551 11543
rect 10551 11509 10560 11543
rect 10508 11500 10560 11509
rect 18696 11500 18748 11552
rect 19708 11500 19760 11552
rect 23020 11543 23072 11552
rect 23020 11509 23029 11543
rect 23029 11509 23063 11543
rect 23063 11509 23072 11543
rect 23020 11500 23072 11509
rect 23204 11500 23256 11552
rect 25872 11500 25924 11552
rect 35900 11568 35952 11620
rect 27252 11500 27304 11552
rect 27344 11500 27396 11552
rect 28724 11500 28776 11552
rect 31392 11500 31444 11552
rect 32680 11500 32732 11552
rect 34428 11500 34480 11552
rect 38108 11568 38160 11620
rect 38844 11679 38896 11688
rect 38844 11645 38853 11679
rect 38853 11645 38887 11679
rect 38887 11645 38896 11679
rect 38844 11636 38896 11645
rect 43996 11772 44048 11824
rect 40408 11704 40460 11756
rect 42064 11704 42116 11756
rect 43168 11704 43220 11756
rect 43536 11747 43588 11756
rect 43536 11713 43545 11747
rect 43545 11713 43579 11747
rect 43579 11713 43588 11747
rect 43536 11704 43588 11713
rect 43628 11704 43680 11756
rect 42432 11679 42484 11688
rect 42432 11645 42441 11679
rect 42441 11645 42475 11679
rect 42475 11645 42484 11679
rect 42432 11636 42484 11645
rect 42984 11636 43036 11688
rect 43260 11679 43312 11688
rect 43260 11645 43269 11679
rect 43269 11645 43303 11679
rect 43303 11645 43312 11679
rect 43260 11636 43312 11645
rect 43444 11679 43496 11688
rect 43444 11645 43453 11679
rect 43453 11645 43487 11679
rect 43487 11645 43496 11679
rect 43444 11636 43496 11645
rect 43996 11679 44048 11688
rect 43996 11645 44005 11679
rect 44005 11645 44039 11679
rect 44039 11645 44048 11679
rect 43996 11636 44048 11645
rect 44916 11636 44968 11688
rect 38568 11500 38620 11552
rect 40040 11500 40092 11552
rect 42708 11500 42760 11552
rect 43352 11568 43404 11620
rect 43076 11543 43128 11552
rect 43076 11509 43085 11543
rect 43085 11509 43119 11543
rect 43119 11509 43128 11543
rect 43076 11500 43128 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 6736 11339 6788 11348
rect 6736 11305 6745 11339
rect 6745 11305 6779 11339
rect 6779 11305 6788 11339
rect 6736 11296 6788 11305
rect 9312 11296 9364 11348
rect 23204 11296 23256 11348
rect 23940 11296 23992 11348
rect 3700 11160 3752 11212
rect 7564 11160 7616 11212
rect 10968 11203 11020 11212
rect 10968 11169 10977 11203
rect 10977 11169 11011 11203
rect 11011 11169 11020 11203
rect 10968 11160 11020 11169
rect 12440 11160 12492 11212
rect 14464 11203 14516 11212
rect 14464 11169 14473 11203
rect 14473 11169 14507 11203
rect 14507 11169 14516 11203
rect 14464 11160 14516 11169
rect 5632 11135 5684 11144
rect 5632 11101 5666 11135
rect 5666 11101 5684 11135
rect 5632 11092 5684 11101
rect 10508 11092 10560 11144
rect 12808 11092 12860 11144
rect 13544 11092 13596 11144
rect 14740 11160 14792 11212
rect 19708 11228 19760 11280
rect 25136 11271 25188 11280
rect 25136 11237 25145 11271
rect 25145 11237 25179 11271
rect 25179 11237 25188 11271
rect 25136 11228 25188 11237
rect 16488 11160 16540 11212
rect 19340 11160 19392 11212
rect 19800 11203 19852 11212
rect 19800 11169 19809 11203
rect 19809 11169 19843 11203
rect 19843 11169 19852 11203
rect 19800 11160 19852 11169
rect 20168 11160 20220 11212
rect 25044 11160 25096 11212
rect 29276 11296 29328 11348
rect 31576 11296 31628 11348
rect 34336 11296 34388 11348
rect 25872 11271 25924 11280
rect 25872 11237 25881 11271
rect 25881 11237 25915 11271
rect 25915 11237 25924 11271
rect 25872 11228 25924 11237
rect 26332 11271 26384 11280
rect 26332 11237 26341 11271
rect 26341 11237 26375 11271
rect 26375 11237 26384 11271
rect 26332 11228 26384 11237
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 17316 11092 17368 11144
rect 22468 11135 22520 11144
rect 22468 11101 22477 11135
rect 22477 11101 22511 11135
rect 22511 11101 22520 11135
rect 22468 11092 22520 11101
rect 24492 11092 24544 11144
rect 26056 11203 26108 11212
rect 26056 11169 26065 11203
rect 26065 11169 26099 11203
rect 26099 11169 26108 11203
rect 26056 11160 26108 11169
rect 6184 11024 6236 11076
rect 8852 11024 8904 11076
rect 10048 11024 10100 11076
rect 10968 11024 11020 11076
rect 13452 11024 13504 11076
rect 13636 11024 13688 11076
rect 16304 11024 16356 11076
rect 18052 11024 18104 11076
rect 22836 11024 22888 11076
rect 25412 11067 25464 11076
rect 25412 11033 25421 11067
rect 25421 11033 25455 11067
rect 25455 11033 25464 11067
rect 25412 11024 25464 11033
rect 25872 11092 25924 11144
rect 9680 10956 9732 11008
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 15200 10999 15252 11008
rect 15200 10965 15209 10999
rect 15209 10965 15243 10999
rect 15243 10965 15252 10999
rect 15200 10956 15252 10965
rect 15844 10999 15896 11008
rect 15844 10965 15853 10999
rect 15853 10965 15887 10999
rect 15887 10965 15896 10999
rect 15844 10956 15896 10965
rect 17776 10956 17828 11008
rect 20260 10999 20312 11008
rect 20260 10965 20269 10999
rect 20269 10965 20303 10999
rect 20303 10965 20312 10999
rect 20260 10956 20312 10965
rect 25872 10956 25924 11008
rect 29828 11228 29880 11280
rect 30472 11228 30524 11280
rect 30380 11092 30432 11144
rect 31668 11092 31720 11144
rect 27436 11024 27488 11076
rect 31208 11024 31260 11076
rect 32680 11135 32732 11144
rect 32680 11101 32689 11135
rect 32689 11101 32723 11135
rect 32723 11101 32732 11135
rect 32680 11092 32732 11101
rect 35348 11160 35400 11212
rect 36912 11296 36964 11348
rect 38752 11296 38804 11348
rect 39028 11339 39080 11348
rect 39028 11305 39037 11339
rect 39037 11305 39071 11339
rect 39071 11305 39080 11339
rect 39028 11296 39080 11305
rect 42524 11296 42576 11348
rect 43444 11296 43496 11348
rect 38568 11228 38620 11280
rect 39488 11271 39540 11280
rect 34428 11135 34480 11144
rect 34428 11101 34437 11135
rect 34437 11101 34471 11135
rect 34471 11101 34480 11135
rect 34428 11092 34480 11101
rect 35900 11135 35952 11144
rect 35900 11101 35909 11135
rect 35909 11101 35943 11135
rect 35943 11101 35952 11135
rect 35900 11092 35952 11101
rect 37740 11135 37792 11144
rect 37740 11101 37749 11135
rect 37749 11101 37783 11135
rect 37783 11101 37792 11135
rect 37740 11092 37792 11101
rect 37924 11135 37976 11144
rect 37924 11101 37933 11135
rect 37933 11101 37967 11135
rect 37967 11101 37976 11135
rect 37924 11092 37976 11101
rect 38384 11135 38436 11144
rect 38384 11101 38393 11135
rect 38393 11101 38427 11135
rect 38427 11101 38436 11135
rect 38384 11092 38436 11101
rect 39488 11237 39497 11271
rect 39497 11237 39531 11271
rect 39531 11237 39540 11271
rect 39488 11228 39540 11237
rect 43996 11228 44048 11280
rect 38844 11135 38896 11144
rect 38844 11101 38853 11135
rect 38853 11101 38887 11135
rect 38887 11101 38896 11135
rect 38844 11092 38896 11101
rect 39120 11135 39172 11144
rect 39120 11101 39129 11135
rect 39129 11101 39163 11135
rect 39163 11101 39172 11135
rect 39120 11092 39172 11101
rect 33232 11024 33284 11076
rect 26240 10956 26292 11008
rect 34244 10999 34296 11008
rect 34244 10965 34253 10999
rect 34253 10965 34287 10999
rect 34287 10965 34296 10999
rect 34244 10956 34296 10965
rect 39304 11092 39356 11144
rect 40776 11092 40828 11144
rect 43628 11160 43680 11212
rect 42616 11092 42668 11144
rect 42800 11092 42852 11144
rect 43168 11092 43220 11144
rect 43536 11135 43588 11144
rect 43536 11101 43545 11135
rect 43545 11101 43579 11135
rect 43579 11101 43588 11135
rect 43536 11092 43588 11101
rect 35440 10956 35492 11008
rect 38384 10956 38436 11008
rect 39120 10956 39172 11008
rect 39396 10956 39448 11008
rect 39580 10999 39632 11008
rect 39580 10965 39589 10999
rect 39589 10965 39623 10999
rect 39623 10965 39632 10999
rect 39580 10956 39632 10965
rect 43352 11024 43404 11076
rect 43168 10999 43220 11008
rect 43168 10965 43177 10999
rect 43177 10965 43211 10999
rect 43211 10965 43220 10999
rect 43168 10956 43220 10965
rect 43628 10956 43680 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 7748 10752 7800 10804
rect 8668 10752 8720 10804
rect 10784 10752 10836 10804
rect 12624 10752 12676 10804
rect 8668 10659 8720 10668
rect 8668 10625 8702 10659
rect 8702 10625 8720 10659
rect 8668 10616 8720 10625
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 9496 10616 9548 10668
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 14188 10752 14240 10804
rect 14280 10684 14332 10736
rect 15200 10727 15252 10736
rect 15200 10693 15234 10727
rect 15234 10693 15252 10727
rect 15200 10684 15252 10693
rect 15844 10752 15896 10804
rect 18880 10752 18932 10804
rect 20812 10752 20864 10804
rect 22836 10795 22888 10804
rect 22836 10761 22845 10795
rect 22845 10761 22879 10795
rect 22879 10761 22888 10795
rect 22836 10752 22888 10761
rect 30472 10795 30524 10804
rect 30472 10761 30481 10795
rect 30481 10761 30515 10795
rect 30515 10761 30524 10795
rect 30472 10752 30524 10761
rect 31208 10795 31260 10804
rect 31208 10761 31217 10795
rect 31217 10761 31251 10795
rect 31251 10761 31260 10795
rect 31208 10752 31260 10761
rect 34152 10752 34204 10804
rect 37924 10752 37976 10804
rect 38844 10752 38896 10804
rect 39304 10752 39356 10804
rect 40408 10752 40460 10804
rect 41052 10752 41104 10804
rect 42432 10752 42484 10804
rect 15936 10684 15988 10736
rect 25136 10684 25188 10736
rect 34244 10684 34296 10736
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 7564 10548 7616 10600
rect 7656 10591 7708 10600
rect 7656 10557 7665 10591
rect 7665 10557 7699 10591
rect 7699 10557 7708 10591
rect 7656 10548 7708 10557
rect 7840 10591 7892 10600
rect 7840 10557 7849 10591
rect 7849 10557 7883 10591
rect 7883 10557 7892 10591
rect 7840 10548 7892 10557
rect 8300 10591 8352 10600
rect 8300 10557 8309 10591
rect 8309 10557 8343 10591
rect 8343 10557 8352 10591
rect 8300 10548 8352 10557
rect 8576 10591 8628 10600
rect 8576 10557 8585 10591
rect 8585 10557 8619 10591
rect 8619 10557 8628 10591
rect 8576 10548 8628 10557
rect 9036 10548 9088 10600
rect 11244 10548 11296 10600
rect 11612 10548 11664 10600
rect 12256 10548 12308 10600
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 12624 10548 12676 10600
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 12808 10412 12860 10464
rect 13636 10412 13688 10464
rect 14188 10412 14240 10464
rect 15016 10616 15068 10668
rect 17316 10659 17368 10668
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 17776 10659 17828 10668
rect 17776 10625 17785 10659
rect 17785 10625 17819 10659
rect 17819 10625 17828 10659
rect 17776 10616 17828 10625
rect 18052 10659 18104 10668
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 18880 10659 18932 10668
rect 18880 10625 18914 10659
rect 18914 10625 18932 10659
rect 18880 10616 18932 10625
rect 19064 10659 19116 10668
rect 19064 10625 19073 10659
rect 19073 10625 19107 10659
rect 19107 10625 19116 10659
rect 19064 10616 19116 10625
rect 20076 10616 20128 10668
rect 23020 10659 23072 10668
rect 23020 10625 23029 10659
rect 23029 10625 23063 10659
rect 23063 10625 23072 10659
rect 23020 10616 23072 10625
rect 29000 10616 29052 10668
rect 29644 10659 29696 10668
rect 29644 10625 29678 10659
rect 29678 10625 29696 10659
rect 29644 10616 29696 10625
rect 29828 10659 29880 10668
rect 29828 10625 29837 10659
rect 29837 10625 29871 10659
rect 29871 10625 29880 10659
rect 29828 10616 29880 10625
rect 31392 10659 31444 10668
rect 31392 10625 31401 10659
rect 31401 10625 31435 10659
rect 31435 10625 31444 10659
rect 31392 10616 31444 10625
rect 33232 10659 33284 10668
rect 33232 10625 33241 10659
rect 33241 10625 33275 10659
rect 33275 10625 33284 10659
rect 33232 10616 33284 10625
rect 34612 10616 34664 10668
rect 35348 10616 35400 10668
rect 35992 10659 36044 10668
rect 35992 10625 36001 10659
rect 36001 10625 36035 10659
rect 36035 10625 36044 10659
rect 35992 10616 36044 10625
rect 37832 10616 37884 10668
rect 38108 10659 38160 10668
rect 38108 10625 38117 10659
rect 38117 10625 38151 10659
rect 38151 10625 38160 10659
rect 38108 10616 38160 10625
rect 38384 10659 38436 10668
rect 38384 10625 38393 10659
rect 38393 10625 38427 10659
rect 38427 10625 38436 10659
rect 38384 10616 38436 10625
rect 39580 10684 39632 10736
rect 40500 10684 40552 10736
rect 43076 10684 43128 10736
rect 38752 10659 38804 10668
rect 38752 10625 38761 10659
rect 38761 10625 38795 10659
rect 38795 10625 38804 10659
rect 38752 10616 38804 10625
rect 39120 10616 39172 10668
rect 40040 10659 40092 10668
rect 40040 10625 40049 10659
rect 40049 10625 40083 10659
rect 40083 10625 40092 10659
rect 40040 10616 40092 10625
rect 15936 10548 15988 10600
rect 17868 10591 17920 10600
rect 17868 10557 17877 10591
rect 17877 10557 17911 10591
rect 17911 10557 17920 10591
rect 17868 10548 17920 10557
rect 18788 10591 18840 10600
rect 17592 10523 17644 10532
rect 17592 10489 17601 10523
rect 17601 10489 17635 10523
rect 17635 10489 17644 10523
rect 17592 10480 17644 10489
rect 17684 10480 17736 10532
rect 15292 10412 15344 10464
rect 18788 10557 18797 10591
rect 18797 10557 18831 10591
rect 18831 10557 18840 10591
rect 18788 10548 18840 10557
rect 19892 10548 19944 10600
rect 29184 10548 29236 10600
rect 29368 10548 29420 10600
rect 29552 10591 29604 10600
rect 29552 10557 29561 10591
rect 29561 10557 29595 10591
rect 29595 10557 29604 10591
rect 29552 10548 29604 10557
rect 38660 10591 38712 10600
rect 38660 10557 38669 10591
rect 38669 10557 38703 10591
rect 38703 10557 38712 10591
rect 38660 10548 38712 10557
rect 40408 10659 40460 10668
rect 40408 10625 40417 10659
rect 40417 10625 40451 10659
rect 40451 10625 40460 10659
rect 40408 10616 40460 10625
rect 40776 10616 40828 10668
rect 20536 10412 20588 10464
rect 22008 10480 22060 10532
rect 38384 10480 38436 10532
rect 39488 10480 39540 10532
rect 40316 10480 40368 10532
rect 21272 10412 21324 10464
rect 31484 10412 31536 10464
rect 38292 10412 38344 10464
rect 42892 10659 42944 10668
rect 42892 10625 42901 10659
rect 42901 10625 42935 10659
rect 42935 10625 42944 10659
rect 42892 10616 42944 10625
rect 43352 10795 43404 10804
rect 43352 10761 43361 10795
rect 43361 10761 43395 10795
rect 43395 10761 43404 10795
rect 43352 10752 43404 10761
rect 43628 10795 43680 10804
rect 43628 10761 43653 10795
rect 43653 10761 43680 10795
rect 43628 10752 43680 10761
rect 43444 10727 43496 10736
rect 43444 10693 43453 10727
rect 43453 10693 43487 10727
rect 43487 10693 43496 10727
rect 43444 10684 43496 10693
rect 44180 10616 44232 10668
rect 46480 10659 46532 10668
rect 46480 10625 46489 10659
rect 46489 10625 46523 10659
rect 46523 10625 46532 10659
rect 46480 10616 46532 10625
rect 43352 10412 43404 10464
rect 46664 10455 46716 10464
rect 46664 10421 46673 10455
rect 46673 10421 46707 10455
rect 46707 10421 46716 10455
rect 46664 10412 46716 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 6184 10115 6236 10124
rect 6184 10081 6193 10115
rect 6193 10081 6227 10115
rect 6227 10081 6236 10115
rect 6184 10072 6236 10081
rect 7196 10072 7248 10124
rect 8484 10208 8536 10260
rect 9496 10208 9548 10260
rect 10416 10208 10468 10260
rect 9680 10140 9732 10192
rect 6276 10004 6328 10056
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 2228 9979 2280 9988
rect 2228 9945 2237 9979
rect 2237 9945 2271 9979
rect 2271 9945 2280 9979
rect 2228 9936 2280 9945
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 8576 9936 8628 9988
rect 8852 9936 8904 9988
rect 10140 9936 10192 9988
rect 9588 9868 9640 9920
rect 15292 10140 15344 10192
rect 18052 10208 18104 10260
rect 20076 10251 20128 10260
rect 20076 10217 20085 10251
rect 20085 10217 20119 10251
rect 20119 10217 20128 10251
rect 20076 10208 20128 10217
rect 20260 10208 20312 10260
rect 11244 10115 11296 10124
rect 11244 10081 11253 10115
rect 11253 10081 11287 10115
rect 11287 10081 11296 10115
rect 11244 10072 11296 10081
rect 11612 10072 11664 10124
rect 12624 10072 12676 10124
rect 13452 10072 13504 10124
rect 13636 10115 13688 10124
rect 13636 10081 13645 10115
rect 13645 10081 13679 10115
rect 13679 10081 13688 10115
rect 13636 10072 13688 10081
rect 14096 10115 14148 10124
rect 14096 10081 14105 10115
rect 14105 10081 14139 10115
rect 14139 10081 14148 10115
rect 14096 10072 14148 10081
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 12440 10047 12492 10056
rect 12440 10013 12449 10047
rect 12449 10013 12483 10047
rect 12483 10013 12492 10047
rect 12440 10004 12492 10013
rect 13544 10004 13596 10056
rect 14188 10004 14240 10056
rect 16672 10004 16724 10056
rect 17040 10004 17092 10056
rect 17592 10004 17644 10056
rect 19432 10004 19484 10056
rect 20536 10072 20588 10124
rect 20352 10047 20404 10056
rect 20352 10013 20361 10047
rect 20361 10013 20395 10047
rect 20395 10013 20404 10047
rect 20352 10004 20404 10013
rect 20444 10004 20496 10056
rect 21088 10072 21140 10124
rect 20996 10047 21048 10056
rect 20996 10013 21005 10047
rect 21005 10013 21039 10047
rect 21039 10013 21048 10047
rect 20996 10004 21048 10013
rect 21640 10047 21692 10056
rect 21640 10013 21649 10047
rect 21649 10013 21683 10047
rect 21683 10013 21692 10047
rect 21640 10004 21692 10013
rect 26240 10140 26292 10192
rect 22284 10072 22336 10124
rect 22376 10072 22428 10124
rect 23112 10115 23164 10124
rect 23112 10081 23121 10115
rect 23121 10081 23155 10115
rect 23155 10081 23164 10115
rect 23112 10072 23164 10081
rect 22192 10047 22244 10056
rect 22192 10013 22201 10047
rect 22201 10013 22235 10047
rect 22235 10013 22244 10047
rect 22192 10004 22244 10013
rect 20076 9936 20128 9988
rect 11060 9868 11112 9920
rect 12164 9868 12216 9920
rect 16304 9868 16356 9920
rect 20168 9868 20220 9920
rect 21456 9911 21508 9920
rect 21456 9877 21465 9911
rect 21465 9877 21499 9911
rect 21499 9877 21508 9911
rect 21456 9868 21508 9877
rect 21548 9868 21600 9920
rect 22008 9868 22060 9920
rect 22376 9911 22428 9920
rect 22376 9877 22385 9911
rect 22385 9877 22419 9911
rect 22419 9877 22428 9911
rect 22376 9868 22428 9877
rect 23204 10047 23256 10056
rect 23204 10013 23213 10047
rect 23213 10013 23247 10047
rect 23247 10013 23256 10047
rect 23204 10004 23256 10013
rect 27804 10115 27856 10124
rect 27804 10081 27813 10115
rect 27813 10081 27847 10115
rect 27847 10081 27856 10115
rect 27804 10072 27856 10081
rect 29000 10072 29052 10124
rect 29920 10140 29972 10192
rect 30104 10140 30156 10192
rect 31484 10183 31536 10192
rect 31484 10149 31493 10183
rect 31493 10149 31527 10183
rect 31527 10149 31536 10183
rect 31484 10140 31536 10149
rect 29644 10072 29696 10124
rect 30748 10115 30800 10124
rect 30748 10081 30757 10115
rect 30757 10081 30791 10115
rect 30791 10081 30800 10115
rect 30748 10072 30800 10081
rect 31116 10072 31168 10124
rect 32036 10115 32088 10124
rect 32036 10081 32045 10115
rect 32045 10081 32079 10115
rect 32079 10081 32088 10115
rect 32036 10072 32088 10081
rect 27712 10047 27764 10056
rect 27712 10013 27721 10047
rect 27721 10013 27755 10047
rect 27755 10013 27764 10047
rect 27712 10004 27764 10013
rect 29184 10004 29236 10056
rect 29368 10004 29420 10056
rect 30564 10047 30616 10056
rect 30564 10013 30598 10047
rect 30598 10013 30616 10047
rect 30564 10004 30616 10013
rect 29460 9936 29512 9988
rect 29092 9868 29144 9920
rect 29184 9911 29236 9920
rect 29184 9877 29193 9911
rect 29193 9877 29227 9911
rect 29227 9877 29236 9911
rect 29184 9868 29236 9877
rect 29552 9868 29604 9920
rect 37372 10208 37424 10260
rect 40408 10208 40460 10260
rect 37832 10140 37884 10192
rect 43076 10140 43128 10192
rect 39212 10072 39264 10124
rect 35440 10047 35492 10056
rect 35440 10013 35449 10047
rect 35449 10013 35483 10047
rect 35483 10013 35492 10047
rect 35440 10004 35492 10013
rect 39396 10047 39448 10056
rect 39396 10013 39405 10047
rect 39405 10013 39439 10047
rect 39439 10013 39448 10047
rect 39396 10004 39448 10013
rect 39488 10047 39540 10056
rect 39488 10013 39497 10047
rect 39497 10013 39531 10047
rect 39531 10013 39540 10047
rect 39488 10004 39540 10013
rect 40592 10072 40644 10124
rect 40868 10072 40920 10124
rect 30564 9868 30616 9920
rect 33324 9868 33376 9920
rect 38292 9936 38344 9988
rect 41052 10047 41104 10056
rect 41052 10013 41061 10047
rect 41061 10013 41095 10047
rect 41095 10013 41104 10047
rect 41052 10004 41104 10013
rect 42432 10004 42484 10056
rect 43720 10072 43772 10124
rect 42984 10047 43036 10056
rect 42984 10013 42993 10047
rect 42993 10013 43027 10047
rect 43027 10013 43036 10047
rect 42984 10004 43036 10013
rect 44180 10004 44232 10056
rect 42800 9936 42852 9988
rect 37372 9868 37424 9920
rect 39764 9868 39816 9920
rect 43168 9911 43220 9920
rect 43168 9877 43177 9911
rect 43177 9877 43211 9911
rect 43211 9877 43220 9911
rect 43168 9868 43220 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 7748 9707 7800 9716
rect 7748 9673 7757 9707
rect 7757 9673 7791 9707
rect 7791 9673 7800 9707
rect 7748 9664 7800 9673
rect 6368 9596 6420 9648
rect 10048 9639 10100 9648
rect 10048 9605 10057 9639
rect 10057 9605 10091 9639
rect 10091 9605 10100 9639
rect 10048 9596 10100 9605
rect 7840 9528 7892 9580
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 6184 9460 6236 9512
rect 7656 9460 7708 9512
rect 8668 9460 8720 9512
rect 10600 9460 10652 9512
rect 12440 9664 12492 9716
rect 17040 9664 17092 9716
rect 20260 9664 20312 9716
rect 20352 9664 20404 9716
rect 25136 9664 25188 9716
rect 27712 9664 27764 9716
rect 19708 9639 19760 9648
rect 19708 9605 19717 9639
rect 19717 9605 19751 9639
rect 19751 9605 19760 9639
rect 19708 9596 19760 9605
rect 19800 9639 19852 9648
rect 19800 9605 19809 9639
rect 19809 9605 19843 9639
rect 19843 9605 19852 9639
rect 19800 9596 19852 9605
rect 26332 9596 26384 9648
rect 17868 9571 17920 9580
rect 17868 9537 17877 9571
rect 17877 9537 17911 9571
rect 17911 9537 17920 9571
rect 17868 9528 17920 9537
rect 18052 9571 18104 9580
rect 18052 9537 18061 9571
rect 18061 9537 18095 9571
rect 18095 9537 18104 9571
rect 18052 9528 18104 9537
rect 18788 9571 18840 9580
rect 18788 9537 18797 9571
rect 18797 9537 18831 9571
rect 18831 9537 18840 9571
rect 18788 9528 18840 9537
rect 18880 9571 18932 9580
rect 18880 9537 18914 9571
rect 18914 9537 18932 9571
rect 18880 9528 18932 9537
rect 19064 9571 19116 9580
rect 19064 9537 19073 9571
rect 19073 9537 19107 9571
rect 19107 9537 19116 9571
rect 19064 9528 19116 9537
rect 19800 9460 19852 9512
rect 21088 9528 21140 9580
rect 21456 9528 21508 9580
rect 22284 9528 22336 9580
rect 24400 9528 24452 9580
rect 25228 9571 25280 9580
rect 25228 9537 25237 9571
rect 25237 9537 25271 9571
rect 25271 9537 25280 9571
rect 25228 9528 25280 9537
rect 23112 9460 23164 9512
rect 24584 9460 24636 9512
rect 24952 9503 25004 9512
rect 24952 9469 24961 9503
rect 24961 9469 24995 9503
rect 24995 9469 25004 9503
rect 24952 9460 25004 9469
rect 25412 9460 25464 9512
rect 17500 9392 17552 9444
rect 9588 9324 9640 9376
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 16580 9324 16632 9376
rect 17040 9324 17092 9376
rect 20076 9435 20128 9444
rect 20076 9401 20085 9435
rect 20085 9401 20119 9435
rect 20119 9401 20128 9435
rect 20076 9392 20128 9401
rect 21088 9435 21140 9444
rect 21088 9401 21097 9435
rect 21097 9401 21131 9435
rect 21131 9401 21140 9435
rect 21088 9392 21140 9401
rect 24124 9392 24176 9444
rect 19892 9324 19944 9376
rect 22560 9324 22612 9376
rect 26792 9571 26844 9580
rect 26792 9537 26801 9571
rect 26801 9537 26835 9571
rect 26835 9537 26844 9571
rect 26792 9528 26844 9537
rect 27528 9596 27580 9648
rect 29092 9664 29144 9716
rect 35256 9664 35308 9716
rect 36176 9664 36228 9716
rect 39856 9664 39908 9716
rect 46480 9664 46532 9716
rect 29184 9596 29236 9648
rect 29552 9596 29604 9648
rect 28264 9392 28316 9444
rect 29276 9392 29328 9444
rect 27712 9324 27764 9376
rect 28356 9367 28408 9376
rect 28356 9333 28365 9367
rect 28365 9333 28399 9367
rect 28399 9333 28408 9367
rect 28356 9324 28408 9333
rect 29460 9324 29512 9376
rect 31300 9528 31352 9580
rect 31944 9596 31996 9648
rect 35992 9596 36044 9648
rect 36452 9596 36504 9648
rect 40500 9596 40552 9648
rect 41052 9596 41104 9648
rect 38384 9571 38436 9580
rect 38384 9537 38393 9571
rect 38393 9537 38427 9571
rect 38427 9537 38436 9571
rect 38384 9528 38436 9537
rect 38660 9528 38712 9580
rect 40040 9528 40092 9580
rect 32036 9460 32088 9512
rect 32128 9460 32180 9512
rect 32312 9460 32364 9512
rect 35348 9460 35400 9512
rect 35808 9460 35860 9512
rect 39488 9460 39540 9512
rect 40316 9571 40368 9580
rect 40316 9537 40325 9571
rect 40325 9537 40359 9571
rect 40359 9537 40368 9571
rect 40316 9528 40368 9537
rect 40684 9528 40736 9580
rect 41144 9528 41196 9580
rect 43352 9596 43404 9648
rect 40776 9460 40828 9512
rect 34796 9392 34848 9444
rect 37740 9392 37792 9444
rect 41052 9392 41104 9444
rect 42892 9528 42944 9580
rect 43168 9528 43220 9580
rect 43076 9503 43128 9512
rect 43076 9469 43085 9503
rect 43085 9469 43119 9503
rect 43119 9469 43128 9503
rect 43076 9460 43128 9469
rect 43260 9503 43312 9512
rect 43260 9469 43269 9503
rect 43269 9469 43303 9503
rect 43303 9469 43312 9503
rect 43260 9460 43312 9469
rect 42708 9392 42760 9444
rect 38108 9324 38160 9376
rect 38384 9367 38436 9376
rect 38384 9333 38393 9367
rect 38393 9333 38427 9367
rect 38427 9333 38436 9367
rect 38384 9324 38436 9333
rect 41420 9324 41472 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 6184 9120 6236 9172
rect 9772 9120 9824 9172
rect 22376 9120 22428 9172
rect 9680 9052 9732 9104
rect 14556 9052 14608 9104
rect 20904 9052 20956 9104
rect 10140 8984 10192 9036
rect 10416 8984 10468 9036
rect 14188 8984 14240 9036
rect 15016 8984 15068 9036
rect 16488 8984 16540 9036
rect 21824 8984 21876 9036
rect 22192 9027 22244 9036
rect 22192 8993 22201 9027
rect 22201 8993 22235 9027
rect 22235 8993 22244 9027
rect 22192 8984 22244 8993
rect 22468 8984 22520 9036
rect 11060 8916 11112 8968
rect 19616 8916 19668 8968
rect 20352 8916 20404 8968
rect 12624 8848 12676 8900
rect 14004 8848 14056 8900
rect 10968 8780 11020 8832
rect 13820 8780 13872 8832
rect 14832 8780 14884 8832
rect 15568 8823 15620 8832
rect 15568 8789 15577 8823
rect 15577 8789 15611 8823
rect 15611 8789 15620 8823
rect 15568 8780 15620 8789
rect 15660 8823 15712 8832
rect 15660 8789 15669 8823
rect 15669 8789 15703 8823
rect 15703 8789 15712 8823
rect 15660 8780 15712 8789
rect 16120 8780 16172 8832
rect 17132 8848 17184 8900
rect 19340 8848 19392 8900
rect 20628 8848 20680 8900
rect 22008 8959 22060 8968
rect 22008 8925 22017 8959
rect 22017 8925 22051 8959
rect 22051 8925 22060 8959
rect 22008 8916 22060 8925
rect 22284 8959 22336 8968
rect 22284 8925 22293 8959
rect 22293 8925 22327 8959
rect 22327 8925 22336 8959
rect 22284 8916 22336 8925
rect 26792 9120 26844 9172
rect 27528 9120 27580 9172
rect 31944 9120 31996 9172
rect 24860 9052 24912 9104
rect 24952 9052 25004 9104
rect 24400 9027 24452 9036
rect 24400 8993 24409 9027
rect 24409 8993 24443 9027
rect 24443 8993 24452 9027
rect 24400 8984 24452 8993
rect 24584 9027 24636 9036
rect 24584 8993 24593 9027
rect 24593 8993 24627 9027
rect 24627 8993 24636 9027
rect 24584 8984 24636 8993
rect 25044 9027 25096 9036
rect 25044 8993 25053 9027
rect 25053 8993 25087 9027
rect 25087 8993 25096 9027
rect 25044 8984 25096 8993
rect 25964 8984 26016 9036
rect 28264 9052 28316 9104
rect 25412 8959 25464 8968
rect 25412 8925 25446 8959
rect 25446 8925 25464 8959
rect 25412 8916 25464 8925
rect 25596 8959 25648 8968
rect 25596 8925 25605 8959
rect 25605 8925 25639 8959
rect 25639 8925 25648 8959
rect 25596 8916 25648 8925
rect 27252 8984 27304 9036
rect 27528 8984 27580 9036
rect 27804 9027 27856 9036
rect 27804 8993 27813 9027
rect 27813 8993 27847 9027
rect 27847 8993 27856 9027
rect 27804 8984 27856 8993
rect 28356 8916 28408 8968
rect 30840 8984 30892 9036
rect 31024 8916 31076 8968
rect 38384 9120 38436 9172
rect 40776 9120 40828 9172
rect 42800 9120 42852 9172
rect 32220 8916 32272 8968
rect 37372 8984 37424 9036
rect 16580 8780 16632 8832
rect 16948 8780 17000 8832
rect 18880 8780 18932 8832
rect 19064 8780 19116 8832
rect 20444 8780 20496 8832
rect 21732 8823 21784 8832
rect 21732 8789 21741 8823
rect 21741 8789 21775 8823
rect 21775 8789 21784 8823
rect 21732 8780 21784 8789
rect 22468 8780 22520 8832
rect 23572 8780 23624 8832
rect 24032 8823 24084 8832
rect 24032 8789 24041 8823
rect 24041 8789 24075 8823
rect 24075 8789 24084 8823
rect 24032 8780 24084 8789
rect 26240 8823 26292 8832
rect 26240 8789 26249 8823
rect 26249 8789 26283 8823
rect 26283 8789 26292 8823
rect 26240 8780 26292 8789
rect 27528 8780 27580 8832
rect 32404 8891 32456 8900
rect 32404 8857 32438 8891
rect 32438 8857 32456 8891
rect 32404 8848 32456 8857
rect 36452 8959 36504 8968
rect 36452 8925 36461 8959
rect 36461 8925 36495 8959
rect 36495 8925 36504 8959
rect 36452 8916 36504 8925
rect 36544 8959 36596 8968
rect 36544 8925 36558 8959
rect 36558 8925 36592 8959
rect 36592 8925 36596 8959
rect 36544 8916 36596 8925
rect 37372 8848 37424 8900
rect 30748 8823 30800 8832
rect 30748 8789 30757 8823
rect 30757 8789 30791 8823
rect 30791 8789 30800 8823
rect 30748 8780 30800 8789
rect 33048 8780 33100 8832
rect 33600 8780 33652 8832
rect 35808 8780 35860 8832
rect 37740 8959 37792 8968
rect 37740 8925 37749 8959
rect 37749 8925 37783 8959
rect 37783 8925 37792 8959
rect 37740 8916 37792 8925
rect 39672 8959 39724 8968
rect 39672 8925 39681 8959
rect 39681 8925 39715 8959
rect 39715 8925 39724 8959
rect 39672 8916 39724 8925
rect 42708 8959 42760 8968
rect 42708 8925 42717 8959
rect 42717 8925 42751 8959
rect 42751 8925 42760 8959
rect 42708 8916 42760 8925
rect 42892 8959 42944 8968
rect 42892 8925 42901 8959
rect 42901 8925 42935 8959
rect 42935 8925 42944 8959
rect 42892 8916 42944 8925
rect 43260 8916 43312 8968
rect 37924 8848 37976 8900
rect 38476 8780 38528 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 7840 8576 7892 8628
rect 8760 8576 8812 8628
rect 9404 8576 9456 8628
rect 14004 8619 14056 8628
rect 14004 8585 14013 8619
rect 14013 8585 14047 8619
rect 14047 8585 14056 8619
rect 14004 8576 14056 8585
rect 8024 8508 8076 8560
rect 8300 8440 8352 8492
rect 8484 8483 8536 8492
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 11704 8440 11756 8492
rect 12440 8440 12492 8492
rect 13912 8483 13964 8492
rect 13912 8449 13921 8483
rect 13921 8449 13955 8483
rect 13955 8449 13964 8483
rect 13912 8440 13964 8449
rect 12256 8372 12308 8424
rect 14188 8415 14240 8424
rect 14188 8381 14197 8415
rect 14197 8381 14231 8415
rect 14231 8381 14240 8415
rect 14188 8372 14240 8381
rect 15568 8576 15620 8628
rect 18144 8576 18196 8628
rect 20076 8576 20128 8628
rect 20904 8619 20956 8628
rect 20904 8585 20913 8619
rect 20913 8585 20947 8619
rect 20947 8585 20956 8619
rect 20904 8576 20956 8585
rect 22192 8576 22244 8628
rect 24400 8576 24452 8628
rect 25596 8576 25648 8628
rect 25964 8576 26016 8628
rect 31300 8619 31352 8628
rect 31300 8585 31309 8619
rect 31309 8585 31343 8619
rect 31343 8585 31352 8619
rect 31300 8576 31352 8585
rect 32404 8576 32456 8628
rect 34796 8619 34848 8628
rect 34796 8585 34805 8619
rect 34805 8585 34839 8619
rect 34839 8585 34848 8619
rect 34796 8576 34848 8585
rect 37924 8576 37976 8628
rect 39764 8576 39816 8628
rect 39856 8619 39908 8628
rect 39856 8585 39865 8619
rect 39865 8585 39899 8619
rect 39899 8585 39908 8619
rect 39856 8576 39908 8585
rect 21732 8508 21784 8560
rect 14832 8483 14884 8492
rect 14832 8449 14841 8483
rect 14841 8449 14875 8483
rect 14875 8449 14884 8483
rect 14832 8440 14884 8449
rect 16948 8440 17000 8492
rect 18144 8483 18196 8492
rect 18144 8449 18178 8483
rect 18178 8449 18196 8483
rect 18144 8440 18196 8449
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 23112 8483 23164 8492
rect 23112 8449 23121 8483
rect 23121 8449 23155 8483
rect 23155 8449 23164 8483
rect 23112 8440 23164 8449
rect 24032 8508 24084 8560
rect 36084 8508 36136 8560
rect 37556 8508 37608 8560
rect 29552 8440 29604 8492
rect 30656 8483 30708 8492
rect 30656 8449 30665 8483
rect 30665 8449 30699 8483
rect 30699 8449 30708 8483
rect 30656 8440 30708 8449
rect 32496 8483 32548 8492
rect 32496 8449 32505 8483
rect 32505 8449 32539 8483
rect 32539 8449 32548 8483
rect 32496 8440 32548 8449
rect 34152 8483 34204 8492
rect 34152 8449 34161 8483
rect 34161 8449 34195 8483
rect 34195 8449 34204 8483
rect 34152 8440 34204 8449
rect 37648 8483 37700 8492
rect 37648 8449 37657 8483
rect 37657 8449 37691 8483
rect 37691 8449 37700 8483
rect 37648 8440 37700 8449
rect 38016 8440 38068 8492
rect 39672 8508 39724 8560
rect 17224 8372 17276 8424
rect 17684 8372 17736 8424
rect 18052 8415 18104 8424
rect 7288 8304 7340 8356
rect 14280 8304 14332 8356
rect 17500 8304 17552 8356
rect 7748 8279 7800 8288
rect 7748 8245 7757 8279
rect 7757 8245 7791 8279
rect 7791 8245 7800 8279
rect 7748 8236 7800 8245
rect 10508 8279 10560 8288
rect 10508 8245 10517 8279
rect 10517 8245 10551 8279
rect 10551 8245 10560 8279
rect 10508 8236 10560 8245
rect 13820 8236 13872 8288
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 18972 8372 19024 8424
rect 19064 8415 19116 8424
rect 19064 8381 19073 8415
rect 19073 8381 19107 8415
rect 19107 8381 19116 8415
rect 19064 8372 19116 8381
rect 19616 8372 19668 8424
rect 19524 8304 19576 8356
rect 19708 8347 19760 8356
rect 19708 8313 19717 8347
rect 19717 8313 19751 8347
rect 19751 8313 19760 8347
rect 19708 8304 19760 8313
rect 20076 8415 20128 8424
rect 20076 8381 20110 8415
rect 20110 8381 20128 8415
rect 20076 8372 20128 8381
rect 20628 8372 20680 8424
rect 24492 8372 24544 8424
rect 29460 8415 29512 8424
rect 29460 8381 29469 8415
rect 29469 8381 29503 8415
rect 29503 8381 29512 8415
rect 29460 8372 29512 8381
rect 29644 8415 29696 8424
rect 29644 8381 29653 8415
rect 29653 8381 29687 8415
rect 29687 8381 29696 8415
rect 29644 8372 29696 8381
rect 30104 8415 30156 8424
rect 30104 8381 30113 8415
rect 30113 8381 30147 8415
rect 30147 8381 30156 8415
rect 30104 8372 30156 8381
rect 30380 8415 30432 8424
rect 30380 8381 30389 8415
rect 30389 8381 30423 8415
rect 30423 8381 30432 8415
rect 30380 8372 30432 8381
rect 30564 8372 30616 8424
rect 32680 8372 32732 8424
rect 22100 8347 22152 8356
rect 22100 8313 22109 8347
rect 22109 8313 22143 8347
rect 22143 8313 22152 8347
rect 22100 8304 22152 8313
rect 23020 8304 23072 8356
rect 23664 8304 23716 8356
rect 20168 8236 20220 8288
rect 22836 8236 22888 8288
rect 23480 8236 23532 8288
rect 30840 8236 30892 8288
rect 32956 8236 33008 8288
rect 33692 8372 33744 8424
rect 33968 8415 34020 8424
rect 33968 8381 34002 8415
rect 34002 8381 34020 8415
rect 33968 8372 34020 8381
rect 33416 8304 33468 8356
rect 34612 8304 34664 8356
rect 35348 8304 35400 8356
rect 40224 8440 40276 8492
rect 46112 8440 46164 8492
rect 38476 8415 38528 8424
rect 38476 8381 38485 8415
rect 38485 8381 38519 8415
rect 38519 8381 38528 8415
rect 38476 8372 38528 8381
rect 45928 8415 45980 8424
rect 45928 8381 45937 8415
rect 45937 8381 45971 8415
rect 45971 8381 45980 8415
rect 45928 8372 45980 8381
rect 34336 8236 34388 8288
rect 37464 8279 37516 8288
rect 37464 8245 37473 8279
rect 37473 8245 37507 8279
rect 37507 8245 37516 8279
rect 37464 8236 37516 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 8300 8032 8352 8084
rect 11612 8075 11664 8084
rect 11612 8041 11621 8075
rect 11621 8041 11655 8075
rect 11655 8041 11664 8075
rect 11612 8032 11664 8041
rect 11704 8075 11756 8084
rect 11704 8041 11713 8075
rect 11713 8041 11747 8075
rect 11747 8041 11756 8075
rect 11704 8032 11756 8041
rect 13912 8075 13964 8084
rect 13912 8041 13921 8075
rect 13921 8041 13955 8075
rect 13955 8041 13964 8075
rect 13912 8032 13964 8041
rect 8760 8007 8812 8016
rect 8760 7973 8769 8007
rect 8769 7973 8803 8007
rect 8803 7973 8812 8007
rect 8760 7964 8812 7973
rect 8484 7896 8536 7948
rect 9404 7939 9456 7948
rect 9404 7905 9413 7939
rect 9413 7905 9447 7939
rect 9447 7905 9456 7939
rect 9404 7896 9456 7905
rect 9864 7896 9916 7948
rect 9956 7896 10008 7948
rect 10232 7939 10284 7948
rect 10232 7905 10241 7939
rect 10241 7905 10275 7939
rect 10275 7905 10284 7939
rect 10232 7896 10284 7905
rect 12256 7939 12308 7948
rect 12256 7905 12265 7939
rect 12265 7905 12299 7939
rect 12299 7905 12308 7939
rect 12256 7896 12308 7905
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 10508 7871 10560 7880
rect 10508 7837 10542 7871
rect 10542 7837 10560 7871
rect 10508 7828 10560 7837
rect 11612 7828 11664 7880
rect 12440 7828 12492 7880
rect 15660 7896 15712 7948
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 14556 7871 14608 7880
rect 14556 7837 14565 7871
rect 14565 7837 14599 7871
rect 14599 7837 14608 7871
rect 14556 7828 14608 7837
rect 16764 7828 16816 7880
rect 10968 7760 11020 7812
rect 11980 7760 12032 7812
rect 12624 7760 12676 7812
rect 9312 7735 9364 7744
rect 9312 7701 9321 7735
rect 9321 7701 9355 7735
rect 9355 7701 9364 7735
rect 9312 7692 9364 7701
rect 14188 7760 14240 7812
rect 16028 7803 16080 7812
rect 16028 7769 16062 7803
rect 16062 7769 16080 7803
rect 16028 7760 16080 7769
rect 14372 7735 14424 7744
rect 14372 7701 14381 7735
rect 14381 7701 14415 7735
rect 14415 7701 14424 7735
rect 14372 7692 14424 7701
rect 17132 8075 17184 8084
rect 17132 8041 17141 8075
rect 17141 8041 17175 8075
rect 17175 8041 17184 8075
rect 17132 8032 17184 8041
rect 17868 8007 17920 8016
rect 17868 7973 17877 8007
rect 17877 7973 17911 8007
rect 17911 7973 17920 8007
rect 17868 7964 17920 7973
rect 19984 7964 20036 8016
rect 21088 8075 21140 8084
rect 21088 8041 21097 8075
rect 21097 8041 21131 8075
rect 21131 8041 21140 8075
rect 21088 8032 21140 8041
rect 21180 8032 21232 8084
rect 22100 7964 22152 8016
rect 25136 7964 25188 8016
rect 17224 7939 17276 7948
rect 17224 7905 17233 7939
rect 17233 7905 17267 7939
rect 17267 7905 17276 7939
rect 17224 7896 17276 7905
rect 17776 7896 17828 7948
rect 17960 7896 18012 7948
rect 18236 7939 18288 7948
rect 18236 7905 18270 7939
rect 18270 7905 18288 7939
rect 18236 7896 18288 7905
rect 17592 7828 17644 7880
rect 19064 7896 19116 7948
rect 19340 7896 19392 7948
rect 19524 7896 19576 7948
rect 19892 7939 19944 7948
rect 19892 7905 19901 7939
rect 19901 7905 19935 7939
rect 19935 7905 19944 7939
rect 19892 7896 19944 7905
rect 20444 7939 20496 7948
rect 20444 7905 20453 7939
rect 20453 7905 20487 7939
rect 20487 7905 20496 7939
rect 20444 7896 20496 7905
rect 30748 8032 30800 8084
rect 32496 8032 32548 8084
rect 33048 8032 33100 8084
rect 19156 7828 19208 7880
rect 19616 7828 19668 7880
rect 20168 7871 20220 7880
rect 20168 7837 20177 7871
rect 20177 7837 20211 7871
rect 20211 7837 20220 7871
rect 20168 7828 20220 7837
rect 19616 7692 19668 7744
rect 26516 7896 26568 7948
rect 27804 7896 27856 7948
rect 22836 7871 22888 7880
rect 22836 7837 22870 7871
rect 22870 7837 22888 7871
rect 22836 7828 22888 7837
rect 26240 7828 26292 7880
rect 28540 7828 28592 7880
rect 29460 7896 29512 7948
rect 30104 7896 30156 7948
rect 30196 7939 30248 7948
rect 30196 7905 30205 7939
rect 30205 7905 30239 7939
rect 30239 7905 30248 7939
rect 30196 7896 30248 7905
rect 30564 7939 30616 7948
rect 30564 7905 30598 7939
rect 30598 7905 30616 7939
rect 30564 7896 30616 7905
rect 29644 7828 29696 7880
rect 30472 7871 30524 7880
rect 30472 7837 30481 7871
rect 30481 7837 30515 7871
rect 30515 7837 30524 7871
rect 30472 7828 30524 7837
rect 30748 7871 30800 7880
rect 30748 7837 30757 7871
rect 30757 7837 30791 7871
rect 30791 7837 30800 7871
rect 30748 7828 30800 7837
rect 32772 7896 32824 7948
rect 32956 7896 33008 7948
rect 34336 7964 34388 8016
rect 36268 8032 36320 8084
rect 38660 8075 38712 8084
rect 38660 8041 38669 8075
rect 38669 8041 38703 8075
rect 38703 8041 38712 8075
rect 38660 8032 38712 8041
rect 33600 7939 33652 7948
rect 33600 7905 33609 7939
rect 33609 7905 33643 7939
rect 33643 7905 33652 7939
rect 33600 7896 33652 7905
rect 34520 7896 34572 7948
rect 34612 7896 34664 7948
rect 35256 7939 35308 7948
rect 35256 7905 35265 7939
rect 35265 7905 35299 7939
rect 35299 7905 35308 7939
rect 35256 7896 35308 7905
rect 32680 7871 32732 7880
rect 32680 7837 32689 7871
rect 32689 7837 32723 7871
rect 32723 7837 32732 7871
rect 32680 7828 32732 7837
rect 33048 7828 33100 7880
rect 33692 7871 33744 7880
rect 33692 7837 33726 7871
rect 33726 7837 33744 7871
rect 33692 7828 33744 7837
rect 33856 7871 33908 7880
rect 33856 7837 33885 7871
rect 33885 7837 33908 7871
rect 33856 7828 33908 7837
rect 35164 7871 35216 7880
rect 35164 7837 35173 7871
rect 35173 7837 35207 7871
rect 35207 7837 35216 7871
rect 35164 7828 35216 7837
rect 38016 7828 38068 7880
rect 38752 7871 38804 7880
rect 38752 7837 38761 7871
rect 38761 7837 38795 7871
rect 38795 7837 38804 7871
rect 38752 7828 38804 7837
rect 29184 7760 29236 7812
rect 23848 7692 23900 7744
rect 23940 7735 23992 7744
rect 23940 7701 23949 7735
rect 23949 7701 23983 7735
rect 23983 7701 23992 7735
rect 23940 7692 23992 7701
rect 26792 7692 26844 7744
rect 27160 7692 27212 7744
rect 31208 7692 31260 7744
rect 33140 7692 33192 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 7656 7488 7708 7540
rect 9312 7488 9364 7540
rect 9864 7488 9916 7540
rect 10968 7488 11020 7540
rect 11244 7488 11296 7540
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 13820 7531 13872 7540
rect 13820 7497 13829 7531
rect 13829 7497 13863 7531
rect 13863 7497 13872 7531
rect 13820 7488 13872 7497
rect 16028 7488 16080 7540
rect 16580 7488 16632 7540
rect 7748 7463 7800 7472
rect 7748 7429 7782 7463
rect 7782 7429 7800 7463
rect 7748 7420 7800 7429
rect 10232 7395 10284 7404
rect 10232 7361 10266 7395
rect 10266 7361 10284 7395
rect 10232 7352 10284 7361
rect 14372 7420 14424 7472
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 18788 7488 18840 7540
rect 20720 7488 20772 7540
rect 20996 7488 21048 7540
rect 22008 7531 22060 7540
rect 22008 7497 22017 7531
rect 22017 7497 22051 7531
rect 22051 7497 22060 7531
rect 22008 7488 22060 7497
rect 23112 7531 23164 7540
rect 23112 7497 23121 7531
rect 23121 7497 23155 7531
rect 23155 7497 23164 7531
rect 23112 7488 23164 7497
rect 23940 7488 23992 7540
rect 25412 7488 25464 7540
rect 19616 7463 19668 7472
rect 19616 7429 19625 7463
rect 19625 7429 19659 7463
rect 19659 7429 19668 7463
rect 19616 7420 19668 7429
rect 19708 7420 19760 7472
rect 23664 7420 23716 7472
rect 18788 7352 18840 7404
rect 18880 7352 18932 7404
rect 7380 7284 7432 7336
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 10968 7284 11020 7336
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 17316 7284 17368 7336
rect 16764 7216 16816 7268
rect 18972 7216 19024 7268
rect 9956 7148 10008 7200
rect 11520 7191 11572 7200
rect 11520 7157 11529 7191
rect 11529 7157 11563 7191
rect 11563 7157 11572 7191
rect 11520 7148 11572 7157
rect 19064 7148 19116 7200
rect 19524 7395 19576 7404
rect 19524 7361 19533 7395
rect 19533 7361 19567 7395
rect 19567 7361 19576 7395
rect 19524 7352 19576 7361
rect 19892 7352 19944 7404
rect 23388 7352 23440 7404
rect 19432 7284 19484 7336
rect 20168 7284 20220 7336
rect 21180 7284 21232 7336
rect 23480 7284 23532 7336
rect 26516 7420 26568 7472
rect 23848 7352 23900 7404
rect 24676 7352 24728 7404
rect 29184 7531 29236 7540
rect 29184 7497 29193 7531
rect 29193 7497 29227 7531
rect 29227 7497 29236 7531
rect 29184 7488 29236 7497
rect 24216 7284 24268 7336
rect 30196 7420 30248 7472
rect 35164 7488 35216 7540
rect 37464 7488 37516 7540
rect 36268 7463 36320 7472
rect 36268 7429 36277 7463
rect 36277 7429 36311 7463
rect 36311 7429 36320 7463
rect 36268 7420 36320 7429
rect 27160 7395 27212 7404
rect 27160 7361 27169 7395
rect 27169 7361 27203 7395
rect 27203 7361 27212 7395
rect 27160 7352 27212 7361
rect 26240 7216 26292 7268
rect 27068 7284 27120 7336
rect 29552 7352 29604 7404
rect 30012 7352 30064 7404
rect 29276 7327 29328 7336
rect 29276 7293 29285 7327
rect 29285 7293 29319 7327
rect 29319 7293 29328 7327
rect 29276 7284 29328 7293
rect 29828 7284 29880 7336
rect 31944 7395 31996 7404
rect 31944 7361 31953 7395
rect 31953 7361 31987 7395
rect 31987 7361 31996 7395
rect 31944 7352 31996 7361
rect 32220 7352 32272 7404
rect 32680 7352 32732 7404
rect 30472 7216 30524 7268
rect 34428 7395 34480 7404
rect 34428 7361 34437 7395
rect 34437 7361 34471 7395
rect 34471 7361 34480 7395
rect 34428 7352 34480 7361
rect 34520 7352 34572 7404
rect 34060 7327 34112 7336
rect 34060 7293 34069 7327
rect 34069 7293 34103 7327
rect 34103 7293 34112 7327
rect 34060 7284 34112 7293
rect 34244 7327 34296 7336
rect 34244 7293 34253 7327
rect 34253 7293 34287 7327
rect 34287 7293 34296 7327
rect 34244 7284 34296 7293
rect 36544 7327 36596 7336
rect 36544 7293 36553 7327
rect 36553 7293 36587 7327
rect 36587 7293 36596 7327
rect 36544 7284 36596 7293
rect 27252 7148 27304 7200
rect 30840 7148 30892 7200
rect 31208 7148 31260 7200
rect 33232 7148 33284 7200
rect 33508 7191 33560 7200
rect 33508 7157 33517 7191
rect 33517 7157 33551 7191
rect 33551 7157 33560 7191
rect 33508 7148 33560 7157
rect 34336 7148 34388 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 10232 6944 10284 6996
rect 14464 6808 14516 6860
rect 15200 6851 15252 6860
rect 15200 6817 15209 6851
rect 15209 6817 15243 6851
rect 15243 6817 15252 6851
rect 15200 6808 15252 6817
rect 15568 6851 15620 6860
rect 15568 6817 15602 6851
rect 15602 6817 15620 6851
rect 15568 6808 15620 6817
rect 15752 6851 15804 6860
rect 15752 6817 15761 6851
rect 15761 6817 15795 6851
rect 15795 6817 15804 6851
rect 15752 6808 15804 6817
rect 19432 6944 19484 6996
rect 19524 6944 19576 6996
rect 11520 6740 11572 6792
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 14648 6740 14700 6792
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 15660 6604 15712 6656
rect 19064 6783 19116 6792
rect 19064 6749 19073 6783
rect 19073 6749 19107 6783
rect 19107 6749 19116 6783
rect 19064 6740 19116 6749
rect 19156 6740 19208 6792
rect 24676 6851 24728 6860
rect 24676 6817 24685 6851
rect 24685 6817 24719 6851
rect 24719 6817 24728 6851
rect 24676 6808 24728 6817
rect 28540 6987 28592 6996
rect 28540 6953 28549 6987
rect 28549 6953 28583 6987
rect 28583 6953 28592 6987
rect 28540 6944 28592 6953
rect 31944 6944 31996 6996
rect 33048 6944 33100 6996
rect 34612 6944 34664 6996
rect 27068 6740 27120 6792
rect 27252 6740 27304 6792
rect 18972 6672 19024 6724
rect 17316 6647 17368 6656
rect 17316 6613 17325 6647
rect 17325 6613 17359 6647
rect 17359 6613 17368 6647
rect 17316 6604 17368 6613
rect 17684 6647 17736 6656
rect 17684 6613 17693 6647
rect 17693 6613 17727 6647
rect 17727 6613 17736 6647
rect 17684 6604 17736 6613
rect 17868 6604 17920 6656
rect 26516 6672 26568 6724
rect 29828 6876 29880 6928
rect 29736 6851 29788 6860
rect 29736 6817 29745 6851
rect 29745 6817 29779 6851
rect 29779 6817 29788 6851
rect 29736 6808 29788 6817
rect 33140 6876 33192 6928
rect 34060 6876 34112 6928
rect 32588 6851 32640 6860
rect 32588 6817 32597 6851
rect 32597 6817 32631 6851
rect 32631 6817 32640 6851
rect 32588 6808 32640 6817
rect 33232 6808 33284 6860
rect 28908 6740 28960 6792
rect 30840 6783 30892 6792
rect 30840 6749 30849 6783
rect 30849 6749 30883 6783
rect 30883 6749 30892 6783
rect 30840 6740 30892 6749
rect 33508 6740 33560 6792
rect 37464 6876 37516 6928
rect 34336 6783 34388 6792
rect 34336 6749 34345 6783
rect 34345 6749 34379 6783
rect 34379 6749 34388 6783
rect 34336 6740 34388 6749
rect 30748 6672 30800 6724
rect 19156 6604 19208 6656
rect 19892 6604 19944 6656
rect 24860 6604 24912 6656
rect 26148 6604 26200 6656
rect 26424 6604 26476 6656
rect 30288 6604 30340 6656
rect 30656 6647 30708 6656
rect 30656 6613 30665 6647
rect 30665 6613 30699 6647
rect 30699 6613 30708 6647
rect 30656 6604 30708 6613
rect 34520 6604 34572 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 17684 6400 17736 6452
rect 13176 6307 13228 6316
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 14004 6307 14056 6316
rect 14004 6273 14013 6307
rect 14013 6273 14047 6307
rect 14047 6273 14056 6307
rect 14004 6264 14056 6273
rect 14188 6196 14240 6248
rect 12992 6103 13044 6112
rect 12992 6069 13001 6103
rect 13001 6069 13035 6103
rect 13035 6069 13044 6103
rect 12992 6060 13044 6069
rect 14096 6060 14148 6112
rect 14648 6239 14700 6248
rect 14648 6205 14657 6239
rect 14657 6205 14691 6239
rect 14691 6205 14700 6239
rect 14648 6196 14700 6205
rect 15568 6264 15620 6316
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 15384 6239 15436 6248
rect 15384 6205 15393 6239
rect 15393 6205 15427 6239
rect 15427 6205 15436 6239
rect 15384 6196 15436 6205
rect 14556 6128 14608 6180
rect 15016 6128 15068 6180
rect 14924 6060 14976 6112
rect 16764 6307 16816 6316
rect 16764 6273 16773 6307
rect 16773 6273 16807 6307
rect 16807 6273 16816 6307
rect 16764 6264 16816 6273
rect 17040 6307 17092 6316
rect 17040 6273 17074 6307
rect 17074 6273 17092 6307
rect 17040 6264 17092 6273
rect 20352 6332 20404 6384
rect 23664 6443 23716 6452
rect 23664 6409 23673 6443
rect 23673 6409 23707 6443
rect 23707 6409 23716 6443
rect 23664 6400 23716 6409
rect 25596 6443 25648 6452
rect 25596 6409 25605 6443
rect 25605 6409 25639 6443
rect 25639 6409 25648 6443
rect 25596 6400 25648 6409
rect 26424 6400 26476 6452
rect 26516 6443 26568 6452
rect 26516 6409 26525 6443
rect 26525 6409 26559 6443
rect 26559 6409 26568 6443
rect 26516 6400 26568 6409
rect 27068 6400 27120 6452
rect 17408 6060 17460 6112
rect 19248 6060 19300 6112
rect 19340 6060 19392 6112
rect 22192 6264 22244 6316
rect 24216 6307 24268 6316
rect 24216 6273 24225 6307
rect 24225 6273 24259 6307
rect 24259 6273 24268 6307
rect 24216 6264 24268 6273
rect 22100 6196 22152 6248
rect 22468 6239 22520 6248
rect 22468 6205 22477 6239
rect 22477 6205 22511 6239
rect 22511 6205 22520 6239
rect 22468 6196 22520 6205
rect 22560 6196 22612 6248
rect 22836 6239 22888 6248
rect 22836 6205 22870 6239
rect 22870 6205 22888 6239
rect 22836 6196 22888 6205
rect 24492 6307 24544 6316
rect 24492 6273 24526 6307
rect 24526 6273 24544 6307
rect 24492 6264 24544 6273
rect 27344 6332 27396 6384
rect 25964 6264 26016 6316
rect 26148 6307 26200 6316
rect 26148 6273 26157 6307
rect 26157 6273 26191 6307
rect 26191 6273 26200 6307
rect 26148 6264 26200 6273
rect 26700 6307 26752 6316
rect 26700 6273 26709 6307
rect 26709 6273 26743 6307
rect 26743 6273 26752 6307
rect 26700 6264 26752 6273
rect 30196 6400 30248 6452
rect 30656 6332 30708 6384
rect 28908 6307 28960 6316
rect 28908 6273 28917 6307
rect 28917 6273 28951 6307
rect 28951 6273 28960 6307
rect 28908 6264 28960 6273
rect 32128 6332 32180 6384
rect 33048 6332 33100 6384
rect 31484 6307 31536 6316
rect 31484 6273 31493 6307
rect 31493 6273 31527 6307
rect 31527 6273 31536 6307
rect 31484 6264 31536 6273
rect 29000 6196 29052 6248
rect 29184 6239 29236 6248
rect 29184 6205 29193 6239
rect 29193 6205 29227 6239
rect 29227 6205 29236 6239
rect 29184 6196 29236 6205
rect 26700 6128 26752 6180
rect 29828 6128 29880 6180
rect 27344 6060 27396 6112
rect 33876 6128 33928 6180
rect 31300 6103 31352 6112
rect 31300 6069 31309 6103
rect 31309 6069 31343 6103
rect 31343 6069 31352 6103
rect 31300 6060 31352 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 13176 5856 13228 5908
rect 14648 5856 14700 5908
rect 15476 5856 15528 5908
rect 17040 5856 17092 5908
rect 17408 5856 17460 5908
rect 19708 5856 19760 5908
rect 14004 5788 14056 5840
rect 14188 5788 14240 5840
rect 15016 5788 15068 5840
rect 17868 5788 17920 5840
rect 21732 5788 21784 5840
rect 22100 5788 22152 5840
rect 23020 5856 23072 5908
rect 23388 5856 23440 5908
rect 24492 5899 24544 5908
rect 24492 5865 24501 5899
rect 24501 5865 24535 5899
rect 24535 5865 24544 5899
rect 24492 5856 24544 5865
rect 24860 5856 24912 5908
rect 26240 5856 26292 5908
rect 27528 5856 27580 5908
rect 29644 5856 29696 5908
rect 14740 5763 14792 5772
rect 14740 5729 14749 5763
rect 14749 5729 14783 5763
rect 14783 5729 14792 5763
rect 14740 5720 14792 5729
rect 18880 5720 18932 5772
rect 19340 5720 19392 5772
rect 24952 5788 25004 5840
rect 25780 5788 25832 5840
rect 22652 5763 22704 5772
rect 22652 5729 22686 5763
rect 22686 5729 22704 5763
rect 22652 5720 22704 5729
rect 23480 5720 23532 5772
rect 12440 5652 12492 5704
rect 17316 5695 17368 5704
rect 17316 5661 17325 5695
rect 17325 5661 17359 5695
rect 17359 5661 17368 5695
rect 17316 5652 17368 5661
rect 13912 5584 13964 5636
rect 14464 5559 14516 5568
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 14464 5516 14516 5525
rect 22560 5695 22612 5704
rect 22560 5661 22569 5695
rect 22569 5661 22603 5695
rect 22603 5661 22612 5695
rect 22560 5652 22612 5661
rect 22192 5516 22244 5568
rect 22652 5516 22704 5568
rect 25136 5652 25188 5704
rect 28632 5720 28684 5772
rect 29184 5720 29236 5772
rect 24860 5627 24912 5636
rect 24860 5593 24869 5627
rect 24869 5593 24903 5627
rect 24903 5593 24912 5627
rect 24860 5584 24912 5593
rect 25044 5627 25096 5636
rect 25044 5593 25053 5627
rect 25053 5593 25087 5627
rect 25087 5593 25096 5627
rect 25044 5584 25096 5593
rect 25596 5584 25648 5636
rect 29552 5652 29604 5704
rect 29736 5652 29788 5704
rect 31300 5652 31352 5704
rect 35348 5652 35400 5704
rect 44364 5652 44416 5704
rect 31024 5584 31076 5636
rect 24952 5516 25004 5568
rect 25964 5516 26016 5568
rect 35072 5559 35124 5568
rect 35072 5525 35081 5559
rect 35081 5525 35115 5559
rect 35115 5525 35124 5559
rect 35072 5516 35124 5525
rect 46664 5559 46716 5568
rect 46664 5525 46673 5559
rect 46673 5525 46707 5559
rect 46707 5525 46716 5559
rect 46664 5516 46716 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 6092 5244 6144 5296
rect 12992 5244 13044 5296
rect 16856 5312 16908 5364
rect 17500 5312 17552 5364
rect 17868 5312 17920 5364
rect 9864 5176 9916 5228
rect 10692 5176 10744 5228
rect 18788 5244 18840 5296
rect 22100 5312 22152 5364
rect 22836 5312 22888 5364
rect 23480 5312 23532 5364
rect 24768 5312 24820 5364
rect 26148 5312 26200 5364
rect 26792 5355 26844 5364
rect 26792 5321 26801 5355
rect 26801 5321 26835 5355
rect 26835 5321 26844 5355
rect 26792 5312 26844 5321
rect 27528 5312 27580 5364
rect 31484 5312 31536 5364
rect 33324 5312 33376 5364
rect 29828 5244 29880 5296
rect 35072 5287 35124 5296
rect 35072 5253 35106 5287
rect 35106 5253 35124 5287
rect 35072 5244 35124 5253
rect 14096 5219 14148 5228
rect 14096 5185 14105 5219
rect 14105 5185 14139 5219
rect 14139 5185 14148 5219
rect 14096 5176 14148 5185
rect 16764 5176 16816 5228
rect 17224 5176 17276 5228
rect 18696 5176 18748 5228
rect 21640 5219 21692 5228
rect 21640 5185 21649 5219
rect 21649 5185 21683 5219
rect 21683 5185 21692 5219
rect 21640 5176 21692 5185
rect 26148 5219 26200 5228
rect 26148 5185 26157 5219
rect 26157 5185 26191 5219
rect 26191 5185 26200 5219
rect 26148 5176 26200 5185
rect 12440 5151 12492 5160
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 21824 5108 21876 5160
rect 24952 5151 25004 5160
rect 24952 5117 24961 5151
rect 24961 5117 24995 5151
rect 24995 5117 25004 5151
rect 24952 5108 25004 5117
rect 940 4972 992 5024
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 14464 5040 14516 5092
rect 23020 5040 23072 5092
rect 13636 4972 13688 5024
rect 13912 5015 13964 5024
rect 13912 4981 13921 5015
rect 13921 4981 13955 5015
rect 13955 4981 13964 5015
rect 13912 4972 13964 4981
rect 19248 5015 19300 5024
rect 19248 4981 19257 5015
rect 19257 4981 19291 5015
rect 19291 4981 19300 5015
rect 19248 4972 19300 4981
rect 25872 5151 25924 5160
rect 25872 5117 25881 5151
rect 25881 5117 25915 5151
rect 25915 5117 25924 5151
rect 25872 5108 25924 5117
rect 26056 5108 26108 5160
rect 28908 5176 28960 5228
rect 29000 5176 29052 5228
rect 27988 5151 28040 5160
rect 27988 5117 27997 5151
rect 27997 5117 28031 5151
rect 28031 5117 28040 5151
rect 27988 5108 28040 5117
rect 29644 5108 29696 5160
rect 30196 5151 30248 5160
rect 30196 5117 30205 5151
rect 30205 5117 30239 5151
rect 30239 5117 30248 5151
rect 30196 5108 30248 5117
rect 32128 5151 32180 5160
rect 32128 5117 32137 5151
rect 32137 5117 32171 5151
rect 32171 5117 32180 5151
rect 32128 5108 32180 5117
rect 32312 5151 32364 5160
rect 32312 5117 32321 5151
rect 32321 5117 32355 5151
rect 32355 5117 32364 5151
rect 32312 5108 32364 5117
rect 33048 5151 33100 5160
rect 33048 5117 33057 5151
rect 33057 5117 33091 5151
rect 33091 5117 33100 5151
rect 33048 5108 33100 5117
rect 33140 5151 33192 5160
rect 33140 5117 33174 5151
rect 33174 5117 33192 5151
rect 33140 5108 33192 5117
rect 34152 5108 34204 5160
rect 25964 4972 26016 5024
rect 27528 4972 27580 5024
rect 33416 4972 33468 5024
rect 33508 4972 33560 5024
rect 35440 5176 35492 5228
rect 34612 5108 34664 5160
rect 34796 5151 34848 5160
rect 34796 5117 34805 5151
rect 34805 5117 34839 5151
rect 34839 5117 34848 5151
rect 34796 5108 34848 5117
rect 35440 4972 35492 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 10692 4811 10744 4820
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 17224 4811 17276 4820
rect 17224 4777 17233 4811
rect 17233 4777 17267 4811
rect 17267 4777 17276 4811
rect 17224 4768 17276 4777
rect 21640 4768 21692 4820
rect 25780 4768 25832 4820
rect 18236 4632 18288 4684
rect 20352 4632 20404 4684
rect 11520 4564 11572 4616
rect 15016 4564 15068 4616
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 15108 4471 15160 4480
rect 15108 4437 15117 4471
rect 15117 4437 15151 4471
rect 15151 4437 15160 4471
rect 15108 4428 15160 4437
rect 17868 4564 17920 4616
rect 19248 4564 19300 4616
rect 22836 4607 22888 4616
rect 22836 4573 22845 4607
rect 22845 4573 22879 4607
rect 22879 4573 22888 4607
rect 22836 4564 22888 4573
rect 24952 4632 25004 4684
rect 25596 4675 25648 4684
rect 25596 4641 25605 4675
rect 25605 4641 25639 4675
rect 25639 4641 25648 4675
rect 25596 4632 25648 4641
rect 25964 4700 26016 4752
rect 27436 4743 27488 4752
rect 27436 4709 27445 4743
rect 27445 4709 27479 4743
rect 27479 4709 27488 4743
rect 27436 4700 27488 4709
rect 28908 4743 28960 4752
rect 28908 4709 28917 4743
rect 28917 4709 28951 4743
rect 28951 4709 28960 4743
rect 28908 4700 28960 4709
rect 29000 4743 29052 4752
rect 29000 4709 29009 4743
rect 29009 4709 29043 4743
rect 29043 4709 29052 4743
rect 29000 4700 29052 4709
rect 31852 4768 31904 4820
rect 35348 4768 35400 4820
rect 25872 4632 25924 4684
rect 25964 4564 26016 4616
rect 26608 4607 26660 4616
rect 26608 4573 26642 4607
rect 26642 4573 26660 4607
rect 26608 4564 26660 4573
rect 27436 4564 27488 4616
rect 19800 4496 19852 4548
rect 21732 4496 21784 4548
rect 25136 4496 25188 4548
rect 27620 4496 27672 4548
rect 32864 4700 32916 4752
rect 29736 4632 29788 4684
rect 32128 4675 32180 4684
rect 32128 4641 32137 4675
rect 32137 4641 32171 4675
rect 32171 4641 32180 4675
rect 32128 4632 32180 4641
rect 29920 4607 29972 4616
rect 29920 4573 29929 4607
rect 29929 4573 29963 4607
rect 29963 4573 29972 4607
rect 29920 4564 29972 4573
rect 32036 4607 32088 4616
rect 32036 4573 32045 4607
rect 32045 4573 32079 4607
rect 32079 4573 32088 4607
rect 32036 4564 32088 4573
rect 32680 4632 32732 4684
rect 33508 4632 33560 4684
rect 36084 4632 36136 4684
rect 36544 4632 36596 4684
rect 32312 4607 32364 4616
rect 32312 4573 32321 4607
rect 32321 4573 32355 4607
rect 32355 4573 32364 4607
rect 32312 4564 32364 4573
rect 33140 4607 33192 4616
rect 33140 4573 33174 4607
rect 33174 4573 33192 4607
rect 33140 4564 33192 4573
rect 33324 4607 33376 4616
rect 33324 4573 33333 4607
rect 33333 4573 33367 4607
rect 33367 4573 33376 4607
rect 33324 4564 33376 4573
rect 35440 4607 35492 4616
rect 35440 4573 35449 4607
rect 35449 4573 35483 4607
rect 35483 4573 35492 4607
rect 35440 4564 35492 4573
rect 35992 4564 36044 4616
rect 38292 4607 38344 4616
rect 38292 4573 38301 4607
rect 38301 4573 38335 4607
rect 38335 4573 38344 4607
rect 38292 4564 38344 4573
rect 18604 4428 18656 4480
rect 21364 4428 21416 4480
rect 24860 4428 24912 4480
rect 26056 4428 26108 4480
rect 26608 4428 26660 4480
rect 27344 4428 27396 4480
rect 29828 4428 29880 4480
rect 31852 4471 31904 4480
rect 31852 4437 31861 4471
rect 31861 4437 31895 4471
rect 31895 4437 31904 4471
rect 31852 4428 31904 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 17776 4156 17828 4208
rect 19800 4224 19852 4276
rect 22192 4267 22244 4276
rect 22192 4233 22201 4267
rect 22201 4233 22235 4267
rect 22235 4233 22244 4267
rect 22192 4224 22244 4233
rect 22560 4224 22612 4276
rect 25872 4224 25924 4276
rect 25964 4224 26016 4276
rect 27988 4224 28040 4276
rect 36084 4224 36136 4276
rect 14372 4131 14424 4140
rect 14372 4097 14406 4131
rect 14406 4097 14424 4131
rect 14372 4088 14424 4097
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 18604 4131 18656 4140
rect 18604 4097 18613 4131
rect 18613 4097 18647 4131
rect 18647 4097 18656 4131
rect 18604 4088 18656 4097
rect 19248 4156 19300 4208
rect 27344 4156 27396 4208
rect 27436 4156 27488 4208
rect 13636 4020 13688 4072
rect 15844 4020 15896 4072
rect 15108 3952 15160 4004
rect 16672 3952 16724 4004
rect 18236 4020 18288 4072
rect 18328 3952 18380 4004
rect 16948 3884 17000 3936
rect 17316 3884 17368 3936
rect 23480 4088 23532 4140
rect 25780 4088 25832 4140
rect 27528 4131 27580 4140
rect 27528 4097 27537 4131
rect 27537 4097 27571 4131
rect 27571 4097 27580 4131
rect 27528 4088 27580 4097
rect 29000 4156 29052 4208
rect 31852 4156 31904 4208
rect 38292 4156 38344 4208
rect 28632 4131 28684 4140
rect 28632 4097 28641 4131
rect 28641 4097 28675 4131
rect 28675 4097 28684 4131
rect 28632 4088 28684 4097
rect 31024 4131 31076 4140
rect 31024 4097 31033 4131
rect 31033 4097 31067 4131
rect 31067 4097 31076 4131
rect 31024 4088 31076 4097
rect 31944 4088 31996 4140
rect 32220 4088 32272 4140
rect 34796 4088 34848 4140
rect 19340 3884 19392 3936
rect 21088 3927 21140 3936
rect 21088 3893 21097 3927
rect 21097 3893 21131 3927
rect 21131 3893 21140 3927
rect 21088 3884 21140 3893
rect 21180 3884 21232 3936
rect 22468 4063 22520 4072
rect 22468 4029 22477 4063
rect 22477 4029 22511 4063
rect 22511 4029 22520 4063
rect 22468 4020 22520 4029
rect 24032 4020 24084 4072
rect 25044 4063 25096 4072
rect 25044 4029 25053 4063
rect 25053 4029 25087 4063
rect 25087 4029 25096 4063
rect 25044 4020 25096 4029
rect 22744 3884 22796 3936
rect 23756 3927 23808 3936
rect 23756 3893 23765 3927
rect 23765 3893 23799 3927
rect 23799 3893 23808 3927
rect 23756 3884 23808 3893
rect 25136 3884 25188 3936
rect 26056 3884 26108 3936
rect 27620 3952 27672 4004
rect 29920 3952 29972 4004
rect 32772 3952 32824 4004
rect 39212 3995 39264 4004
rect 39212 3961 39221 3995
rect 39221 3961 39255 3995
rect 39255 3961 39264 3995
rect 39212 3952 39264 3961
rect 44548 3952 44600 4004
rect 30748 3884 30800 3936
rect 32128 3884 32180 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 14372 3680 14424 3732
rect 17040 3680 17092 3732
rect 18328 3680 18380 3732
rect 17776 3612 17828 3664
rect 16396 3544 16448 3596
rect 14740 3519 14792 3528
rect 14740 3485 14749 3519
rect 14749 3485 14783 3519
rect 14783 3485 14792 3519
rect 14740 3476 14792 3485
rect 15844 3476 15896 3528
rect 16672 3519 16724 3528
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 16764 3519 16816 3528
rect 16764 3485 16773 3519
rect 16773 3485 16807 3519
rect 16807 3485 16816 3519
rect 16764 3476 16816 3485
rect 17316 3476 17368 3528
rect 14280 3383 14332 3392
rect 14280 3349 14289 3383
rect 14289 3349 14323 3383
rect 14323 3349 14332 3383
rect 14280 3340 14332 3349
rect 15476 3383 15528 3392
rect 15476 3349 15485 3383
rect 15485 3349 15519 3383
rect 15519 3349 15528 3383
rect 15476 3340 15528 3349
rect 16580 3340 16632 3392
rect 18788 3587 18840 3596
rect 18788 3553 18797 3587
rect 18797 3553 18831 3587
rect 18831 3553 18840 3587
rect 18788 3544 18840 3553
rect 18604 3519 18656 3528
rect 18604 3485 18613 3519
rect 18613 3485 18647 3519
rect 18647 3485 18656 3519
rect 18604 3476 18656 3485
rect 18696 3383 18748 3392
rect 18696 3349 18705 3383
rect 18705 3349 18739 3383
rect 18739 3349 18748 3383
rect 18696 3340 18748 3349
rect 19800 3340 19852 3392
rect 21180 3680 21232 3732
rect 22192 3723 22244 3732
rect 22192 3689 22201 3723
rect 22201 3689 22235 3723
rect 22235 3689 22244 3723
rect 22192 3680 22244 3689
rect 23480 3723 23532 3732
rect 23480 3689 23489 3723
rect 23489 3689 23523 3723
rect 23523 3689 23532 3723
rect 23480 3680 23532 3689
rect 25872 3680 25924 3732
rect 22376 3612 22428 3664
rect 20628 3587 20680 3596
rect 20628 3553 20637 3587
rect 20637 3553 20671 3587
rect 20671 3553 20680 3587
rect 20628 3544 20680 3553
rect 22744 3587 22796 3596
rect 22744 3553 22753 3587
rect 22753 3553 22787 3587
rect 22787 3553 22796 3587
rect 22744 3544 22796 3553
rect 22836 3587 22888 3596
rect 22836 3553 22845 3587
rect 22845 3553 22879 3587
rect 22879 3553 22888 3587
rect 22836 3544 22888 3553
rect 24124 3587 24176 3596
rect 24124 3553 24133 3587
rect 24133 3553 24167 3587
rect 24167 3553 24176 3587
rect 27436 3680 27488 3732
rect 24124 3544 24176 3553
rect 20904 3476 20956 3528
rect 21088 3519 21140 3528
rect 21088 3485 21122 3519
rect 21122 3485 21140 3519
rect 21088 3476 21140 3485
rect 21364 3476 21416 3528
rect 21824 3408 21876 3460
rect 22376 3476 22428 3528
rect 24032 3476 24084 3528
rect 24216 3476 24268 3528
rect 29368 3544 29420 3596
rect 30012 3587 30064 3596
rect 30012 3553 30021 3587
rect 30021 3553 30055 3587
rect 30055 3553 30064 3587
rect 30012 3544 30064 3553
rect 30196 3587 30248 3596
rect 30196 3553 30205 3587
rect 30205 3553 30239 3587
rect 30239 3553 30248 3587
rect 30196 3544 30248 3553
rect 31944 3680 31996 3732
rect 32036 3680 32088 3732
rect 32772 3680 32824 3732
rect 31852 3655 31904 3664
rect 31852 3621 31861 3655
rect 31861 3621 31895 3655
rect 31895 3621 31904 3655
rect 31852 3612 31904 3621
rect 33140 3612 33192 3664
rect 34244 3612 34296 3664
rect 31760 3544 31812 3596
rect 32588 3544 32640 3596
rect 33232 3587 33284 3596
rect 33232 3553 33241 3587
rect 33241 3553 33275 3587
rect 33275 3553 33284 3587
rect 33232 3544 33284 3553
rect 33876 3587 33928 3596
rect 33876 3553 33885 3587
rect 33885 3553 33919 3587
rect 33919 3553 33928 3587
rect 33876 3544 33928 3553
rect 35256 3587 35308 3596
rect 35256 3553 35265 3587
rect 35265 3553 35299 3587
rect 35299 3553 35308 3587
rect 35256 3544 35308 3553
rect 22560 3340 22612 3392
rect 22652 3383 22704 3392
rect 22652 3349 22661 3383
rect 22661 3349 22695 3383
rect 22695 3349 22704 3383
rect 22652 3340 22704 3349
rect 23112 3383 23164 3392
rect 23112 3349 23121 3383
rect 23121 3349 23155 3383
rect 23155 3349 23164 3383
rect 23112 3340 23164 3349
rect 24952 3408 25004 3460
rect 26056 3476 26108 3528
rect 27620 3519 27672 3528
rect 27620 3485 27629 3519
rect 27629 3485 27663 3519
rect 27663 3485 27672 3519
rect 27620 3476 27672 3485
rect 29828 3476 29880 3528
rect 30564 3476 30616 3528
rect 30748 3519 30800 3528
rect 30748 3485 30782 3519
rect 30782 3485 30800 3519
rect 30748 3476 30800 3485
rect 24860 3340 24912 3392
rect 25596 3340 25648 3392
rect 29368 3340 29420 3392
rect 31484 3408 31536 3460
rect 33048 3451 33100 3460
rect 33048 3417 33057 3451
rect 33057 3417 33091 3451
rect 33091 3417 33100 3451
rect 33048 3408 33100 3417
rect 31760 3340 31812 3392
rect 31944 3383 31996 3392
rect 31944 3349 31953 3383
rect 31953 3349 31987 3383
rect 31987 3349 31996 3383
rect 31944 3340 31996 3349
rect 32128 3340 32180 3392
rect 33508 3476 33560 3528
rect 34704 3476 34756 3528
rect 34704 3383 34756 3392
rect 34704 3349 34713 3383
rect 34713 3349 34747 3383
rect 34747 3349 34756 3383
rect 34704 3340 34756 3349
rect 35164 3383 35216 3392
rect 35164 3349 35173 3383
rect 35173 3349 35207 3383
rect 35207 3349 35216 3383
rect 35164 3340 35216 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 15476 3136 15528 3188
rect 18696 3136 18748 3188
rect 20904 3179 20956 3188
rect 20904 3145 20913 3179
rect 20913 3145 20947 3179
rect 20947 3145 20956 3179
rect 20904 3136 20956 3145
rect 14280 3068 14332 3120
rect 17132 3068 17184 3120
rect 22468 3136 22520 3188
rect 22652 3136 22704 3188
rect 24860 3179 24912 3188
rect 24860 3145 24869 3179
rect 24869 3145 24903 3179
rect 24903 3145 24912 3179
rect 24860 3136 24912 3145
rect 24952 3179 25004 3188
rect 24952 3145 24961 3179
rect 24961 3145 24995 3179
rect 24995 3145 25004 3179
rect 24952 3136 25004 3145
rect 25780 3179 25832 3188
rect 25780 3145 25789 3179
rect 25789 3145 25823 3179
rect 25823 3145 25832 3179
rect 25780 3136 25832 3145
rect 26332 3136 26384 3188
rect 23112 3068 23164 3120
rect 23756 3111 23808 3120
rect 23756 3077 23790 3111
rect 23790 3077 23808 3111
rect 23756 3068 23808 3077
rect 25596 3068 25648 3120
rect 27620 3068 27672 3120
rect 16764 3000 16816 3052
rect 16948 3043 17000 3052
rect 16948 3009 16982 3043
rect 16982 3009 17000 3043
rect 16948 3000 17000 3009
rect 19340 3000 19392 3052
rect 19800 3043 19852 3052
rect 19800 3009 19834 3043
rect 19834 3009 19852 3043
rect 19800 3000 19852 3009
rect 21824 3043 21876 3052
rect 21824 3009 21833 3043
rect 21833 3009 21867 3043
rect 21867 3009 21876 3043
rect 21824 3000 21876 3009
rect 13636 2932 13688 2984
rect 24216 3000 24268 3052
rect 25136 3043 25188 3052
rect 25136 3009 25145 3043
rect 25145 3009 25179 3043
rect 25179 3009 25188 3043
rect 25136 3000 25188 3009
rect 28632 3000 28684 3052
rect 29184 3043 29236 3052
rect 29184 3009 29218 3043
rect 29218 3009 29236 3043
rect 29184 3000 29236 3009
rect 25044 2932 25096 2984
rect 26332 2975 26384 2984
rect 26332 2941 26341 2975
rect 26341 2941 26375 2975
rect 26375 2941 26384 2975
rect 26332 2932 26384 2941
rect 2228 2907 2280 2916
rect 2228 2873 2237 2907
rect 2237 2873 2271 2907
rect 2271 2873 2280 2907
rect 2228 2864 2280 2873
rect 30012 3136 30064 3188
rect 31024 3179 31076 3188
rect 31024 3145 31033 3179
rect 31033 3145 31067 3179
rect 31067 3145 31076 3179
rect 31024 3136 31076 3145
rect 31852 3136 31904 3188
rect 33324 3136 33376 3188
rect 34612 3136 34664 3188
rect 35164 3136 35216 3188
rect 45560 3136 45612 3188
rect 30564 3068 30616 3120
rect 31484 3111 31536 3120
rect 31484 3077 31493 3111
rect 31493 3077 31527 3111
rect 31527 3077 31536 3111
rect 31484 3068 31536 3077
rect 31944 3068 31996 3120
rect 32036 3000 32088 3052
rect 31760 2932 31812 2984
rect 33416 3000 33468 3052
rect 46572 3043 46624 3052
rect 46572 3009 46581 3043
rect 46581 3009 46615 3043
rect 46615 3009 46624 3043
rect 46572 3000 46624 3009
rect 20 2796 72 2848
rect 18420 2796 18472 2848
rect 22468 2796 22520 2848
rect 22560 2796 22612 2848
rect 28632 2796 28684 2848
rect 31668 2796 31720 2848
rect 33232 2796 33284 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 5908 2592 5960 2644
rect 2688 2524 2740 2576
rect 1952 2388 2004 2440
rect 10784 2524 10836 2576
rect 13268 2524 13320 2576
rect 36452 2592 36504 2644
rect 38752 2592 38804 2644
rect 9404 2499 9456 2508
rect 9404 2465 9413 2499
rect 9413 2465 9447 2499
rect 9447 2465 9456 2499
rect 9404 2456 9456 2465
rect 6460 2388 6512 2440
rect 9036 2388 9088 2440
rect 11336 2388 11388 2440
rect 13544 2388 13596 2440
rect 20720 2456 20772 2508
rect 37648 2524 37700 2576
rect 16120 2388 16172 2440
rect 18696 2388 18748 2440
rect 20996 2431 21048 2440
rect 20996 2397 21005 2431
rect 21005 2397 21039 2431
rect 21039 2397 21048 2431
rect 20996 2388 21048 2397
rect 23204 2388 23256 2440
rect 25136 2388 25188 2440
rect 28632 2388 28684 2440
rect 29368 2431 29420 2440
rect 29368 2397 29377 2431
rect 29377 2397 29411 2431
rect 29411 2397 29420 2431
rect 29368 2388 29420 2397
rect 37188 2456 37240 2508
rect 42708 2499 42760 2508
rect 42708 2465 42717 2499
rect 42717 2465 42751 2499
rect 42751 2465 42760 2499
rect 42708 2456 42760 2465
rect 45468 2456 45520 2508
rect 46204 2499 46256 2508
rect 46204 2465 46213 2499
rect 46213 2465 46247 2499
rect 46247 2465 46256 2499
rect 46204 2456 46256 2465
rect 34704 2388 34756 2440
rect 34888 2431 34940 2440
rect 34888 2397 34897 2431
rect 34897 2397 34931 2431
rect 34931 2397 34940 2431
rect 34888 2388 34940 2397
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 39304 2388 39356 2440
rect 41880 2388 41932 2440
rect 44548 2431 44600 2440
rect 44548 2397 44557 2431
rect 44557 2397 44591 2431
rect 44591 2397 44600 2431
rect 44548 2388 44600 2397
rect 940 2252 992 2304
rect 4528 2252 4580 2304
rect 11612 2252 11664 2304
rect 13636 2252 13688 2304
rect 20628 2320 20680 2372
rect 34612 2320 34664 2372
rect 46388 2320 46440 2372
rect 18696 2252 18748 2304
rect 27712 2252 27764 2304
rect 29184 2295 29236 2304
rect 29184 2261 29193 2295
rect 29193 2261 29227 2295
rect 29227 2261 29236 2295
rect 29184 2252 29236 2261
rect 30380 2295 30432 2304
rect 30380 2261 30389 2295
rect 30389 2261 30423 2295
rect 30423 2261 30432 2295
rect 30380 2252 30432 2261
rect 32220 2252 32272 2304
rect 33416 2295 33468 2304
rect 33416 2261 33425 2295
rect 33425 2261 33459 2295
rect 33459 2261 33468 2295
rect 33416 2252 33468 2261
rect 34796 2252 34848 2304
rect 37372 2252 37424 2304
rect 44456 2252 44508 2304
rect 45652 2295 45704 2304
rect 45652 2261 45661 2295
rect 45661 2261 45695 2295
rect 45695 2261 45704 2295
rect 45652 2252 45704 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 1306 49624 1362 50424
rect 3238 49624 3294 50424
rect 5814 49722 5870 50424
rect 8390 49722 8446 50424
rect 10322 49722 10378 50424
rect 12898 49722 12954 50424
rect 15474 49722 15530 50424
rect 5814 49694 6040 49722
rect 5814 49624 5870 49694
rect 1124 47184 1176 47190
rect 1124 47126 1176 47132
rect 1136 47025 1164 47126
rect 1122 47016 1178 47025
rect 1122 46951 1178 46960
rect 1320 46714 1348 49624
rect 1766 49056 1822 49065
rect 1766 48991 1822 49000
rect 1780 47802 1808 48991
rect 3252 47802 3280 49624
rect 4874 47900 5182 47909
rect 4874 47898 4880 47900
rect 4936 47898 4960 47900
rect 5016 47898 5040 47900
rect 5096 47898 5120 47900
rect 5176 47898 5182 47900
rect 4936 47846 4938 47898
rect 5118 47846 5120 47898
rect 4874 47844 4880 47846
rect 4936 47844 4960 47846
rect 5016 47844 5040 47846
rect 5096 47844 5120 47846
rect 5176 47844 5182 47846
rect 4874 47835 5182 47844
rect 1768 47796 1820 47802
rect 1768 47738 1820 47744
rect 3240 47796 3292 47802
rect 3240 47738 3292 47744
rect 6012 47734 6040 49694
rect 8390 49694 8708 49722
rect 8390 49624 8446 49694
rect 6092 48068 6144 48074
rect 6092 48010 6144 48016
rect 6104 47802 6132 48010
rect 6092 47796 6144 47802
rect 6092 47738 6144 47744
rect 6000 47728 6052 47734
rect 6000 47670 6052 47676
rect 8680 47666 8708 49694
rect 10322 49694 10640 49722
rect 10322 49624 10378 49694
rect 10612 47802 10640 49694
rect 12898 49694 13216 49722
rect 12898 49624 12954 49694
rect 13188 47802 13216 49694
rect 15474 49694 15792 49722
rect 15474 49624 15530 49694
rect 15764 47802 15792 49694
rect 17406 49624 17462 50424
rect 19982 49624 20038 50424
rect 22558 49624 22614 50424
rect 24490 49722 24546 50424
rect 27066 49722 27122 50424
rect 24490 49694 24624 49722
rect 24490 49624 24546 49694
rect 17420 47802 17448 49624
rect 19996 47802 20024 49624
rect 22572 47802 22600 49624
rect 10600 47796 10652 47802
rect 10600 47738 10652 47744
rect 13176 47796 13228 47802
rect 13176 47738 13228 47744
rect 15752 47796 15804 47802
rect 15752 47738 15804 47744
rect 17408 47796 17460 47802
rect 17408 47738 17460 47744
rect 19984 47796 20036 47802
rect 19984 47738 20036 47744
rect 22560 47796 22612 47802
rect 22560 47738 22612 47744
rect 24596 47666 24624 49694
rect 27066 49694 27292 49722
rect 27066 49624 27122 49694
rect 27264 47734 27292 49694
rect 28998 49624 29054 50424
rect 31574 49722 31630 50424
rect 34150 49722 34206 50424
rect 31574 49694 31708 49722
rect 31574 49624 31630 49694
rect 29012 47802 29040 49624
rect 29000 47796 29052 47802
rect 31680 47784 31708 49694
rect 34150 49694 34468 49722
rect 34150 49624 34206 49694
rect 32128 48068 32180 48074
rect 32128 48010 32180 48016
rect 31760 47796 31812 47802
rect 31680 47756 31760 47784
rect 29000 47738 29052 47744
rect 31760 47738 31812 47744
rect 27252 47728 27304 47734
rect 27252 47670 27304 47676
rect 28264 47728 28316 47734
rect 28264 47670 28316 47676
rect 2320 47660 2372 47666
rect 2320 47602 2372 47608
rect 3056 47660 3108 47666
rect 3056 47602 3108 47608
rect 8668 47660 8720 47666
rect 8668 47602 8720 47608
rect 10232 47660 10284 47666
rect 10232 47602 10284 47608
rect 15200 47660 15252 47666
rect 15200 47602 15252 47608
rect 17316 47660 17368 47666
rect 17316 47602 17368 47608
rect 19248 47660 19300 47666
rect 19248 47602 19300 47608
rect 20352 47660 20404 47666
rect 20352 47602 20404 47608
rect 23204 47660 23256 47666
rect 23204 47602 23256 47608
rect 24584 47660 24636 47666
rect 24584 47602 24636 47608
rect 27344 47660 27396 47666
rect 27344 47602 27396 47608
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 1308 46708 1360 46714
rect 1308 46650 1360 46656
rect 1400 44396 1452 44402
rect 1400 44338 1452 44344
rect 938 44296 994 44305
rect 938 44231 940 44240
rect 992 44231 994 44240
rect 940 44202 992 44208
rect 1412 42294 1440 44338
rect 1400 42288 1452 42294
rect 1400 42230 1452 42236
rect 1400 41608 1452 41614
rect 938 41576 994 41585
rect 1400 41550 1452 41556
rect 938 41511 994 41520
rect 952 41478 980 41511
rect 940 41472 992 41478
rect 940 41414 992 41420
rect 940 39840 992 39846
rect 940 39782 992 39788
rect 952 39545 980 39782
rect 938 39536 994 39545
rect 938 39471 994 39480
rect 940 37256 992 37262
rect 940 37198 992 37204
rect 952 36825 980 37198
rect 938 36816 994 36825
rect 938 36751 994 36760
rect 938 32056 994 32065
rect 938 31991 994 32000
rect 952 31890 980 31991
rect 940 31884 992 31890
rect 940 31826 992 31832
rect 940 29640 992 29646
rect 940 29582 992 29588
rect 952 29345 980 29582
rect 938 29336 994 29345
rect 938 29271 994 29280
rect 940 26784 992 26790
rect 940 26726 992 26732
rect 952 26625 980 26726
rect 938 26616 994 26625
rect 938 26551 994 26560
rect 940 24812 992 24818
rect 940 24754 992 24760
rect 952 24585 980 24754
rect 1412 24721 1440 41550
rect 1492 39636 1544 39642
rect 1492 39578 1544 39584
rect 1504 34678 1532 39578
rect 1768 35080 1820 35086
rect 1768 35022 1820 35028
rect 1492 34672 1544 34678
rect 1492 34614 1544 34620
rect 1584 34400 1636 34406
rect 1584 34342 1636 34348
rect 1596 34105 1624 34342
rect 1582 34096 1638 34105
rect 1582 34031 1638 34040
rect 1780 32910 1808 35022
rect 1676 32904 1728 32910
rect 1676 32846 1728 32852
rect 1768 32904 1820 32910
rect 1768 32846 1820 32852
rect 1492 32768 1544 32774
rect 1492 32710 1544 32716
rect 1504 32502 1532 32710
rect 1688 32570 1716 32846
rect 1676 32564 1728 32570
rect 1676 32506 1728 32512
rect 1492 32496 1544 32502
rect 1492 32438 1544 32444
rect 1780 32434 1808 32846
rect 1768 32428 1820 32434
rect 1768 32370 1820 32376
rect 1674 31920 1730 31929
rect 1674 31855 1676 31864
rect 1728 31855 1730 31864
rect 1676 31826 1728 31832
rect 1780 30734 1808 32370
rect 1964 31226 1992 46990
rect 2044 40520 2096 40526
rect 2044 40462 2096 40468
rect 2056 40186 2084 40462
rect 2044 40180 2096 40186
rect 2044 40122 2096 40128
rect 2044 40044 2096 40050
rect 2044 39986 2096 39992
rect 2056 39846 2084 39986
rect 2044 39840 2096 39846
rect 2044 39782 2096 39788
rect 2056 39574 2084 39782
rect 2044 39568 2096 39574
rect 2044 39510 2096 39516
rect 2136 36236 2188 36242
rect 2136 36178 2188 36184
rect 2148 35630 2176 36178
rect 2136 35624 2188 35630
rect 2136 35566 2188 35572
rect 2148 35086 2176 35566
rect 2136 35080 2188 35086
rect 2136 35022 2188 35028
rect 2044 33312 2096 33318
rect 2044 33254 2096 33260
rect 2056 32910 2084 33254
rect 2044 32904 2096 32910
rect 2044 32846 2096 32852
rect 2228 31340 2280 31346
rect 2228 31282 2280 31288
rect 1964 31198 2176 31226
rect 2044 31136 2096 31142
rect 2044 31078 2096 31084
rect 2056 30734 2084 31078
rect 1768 30728 1820 30734
rect 1768 30670 1820 30676
rect 2044 30728 2096 30734
rect 2044 30670 2096 30676
rect 1674 29744 1730 29753
rect 1674 29679 1676 29688
rect 1728 29679 1730 29688
rect 1676 29650 1728 29656
rect 1676 28144 1728 28150
rect 1676 28086 1728 28092
rect 1688 27538 1716 28086
rect 1952 27872 2004 27878
rect 1952 27814 2004 27820
rect 1676 27532 1728 27538
rect 1676 27474 1728 27480
rect 1688 26382 1716 27474
rect 1964 27470 1992 27814
rect 1952 27464 2004 27470
rect 1952 27406 2004 27412
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 1688 25294 1716 26318
rect 2044 26308 2096 26314
rect 2044 26250 2096 26256
rect 2056 26042 2084 26250
rect 2044 26036 2096 26042
rect 2044 25978 2096 25984
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1398 24712 1454 24721
rect 1398 24647 1454 24656
rect 1584 24608 1636 24614
rect 938 24576 994 24585
rect 1584 24550 1636 24556
rect 938 24511 994 24520
rect 940 22024 992 22030
rect 940 21966 992 21972
rect 952 21865 980 21966
rect 938 21856 994 21865
rect 938 21791 994 21800
rect 1306 19816 1362 19825
rect 1306 19751 1362 19760
rect 1320 19514 1348 19751
rect 1308 19508 1360 19514
rect 1308 19450 1360 19456
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 940 17196 992 17202
rect 940 17138 992 17144
rect 952 17105 980 17138
rect 938 17096 994 17105
rect 938 17031 994 17040
rect 1412 14414 1440 18226
rect 1596 17241 1624 24550
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 2056 23118 2084 23462
rect 2148 23322 2176 31198
rect 2240 30394 2268 31282
rect 2228 30388 2280 30394
rect 2228 30330 2280 30336
rect 2332 30274 2360 47602
rect 3068 47258 3096 47602
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 3056 47252 3108 47258
rect 3056 47194 3108 47200
rect 4804 46912 4856 46918
rect 4804 46854 4856 46860
rect 6000 46912 6052 46918
rect 6000 46854 6052 46860
rect 4816 46578 4844 46854
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 6012 46646 6040 46854
rect 6000 46640 6052 46646
rect 6000 46582 6052 46588
rect 4804 46572 4856 46578
rect 4804 46514 4856 46520
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 2688 44464 2740 44470
rect 2688 44406 2740 44412
rect 2596 40384 2648 40390
rect 2596 40326 2648 40332
rect 2608 40186 2636 40326
rect 2596 40180 2648 40186
rect 2596 40122 2648 40128
rect 2700 40066 2728 44406
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4620 43988 4672 43994
rect 4620 43930 4672 43936
rect 4632 43722 4660 43930
rect 3240 43716 3292 43722
rect 3240 43658 3292 43664
rect 4620 43716 4672 43722
rect 4620 43658 4672 43664
rect 2608 40038 2728 40066
rect 2412 37120 2464 37126
rect 2412 37062 2464 37068
rect 2424 30326 2452 37062
rect 2608 35894 2636 40038
rect 2688 39976 2740 39982
rect 2688 39918 2740 39924
rect 2516 35866 2636 35894
rect 2240 30246 2360 30274
rect 2412 30320 2464 30326
rect 2412 30262 2464 30268
rect 2136 23316 2188 23322
rect 2136 23258 2188 23264
rect 1676 23112 1728 23118
rect 1676 23054 1728 23060
rect 2044 23112 2096 23118
rect 2044 23054 2096 23060
rect 1688 22574 1716 23054
rect 2044 22636 2096 22642
rect 2044 22578 2096 22584
rect 1676 22568 1728 22574
rect 1676 22510 1728 22516
rect 1688 20398 1716 22510
rect 2056 22234 2084 22578
rect 2044 22228 2096 22234
rect 2044 22170 2096 22176
rect 2136 20800 2188 20806
rect 2136 20742 2188 20748
rect 2148 20534 2176 20742
rect 2136 20528 2188 20534
rect 2136 20470 2188 20476
rect 1676 20392 1728 20398
rect 2240 20346 2268 30246
rect 2412 30184 2464 30190
rect 2412 30126 2464 30132
rect 2424 29306 2452 30126
rect 2412 29300 2464 29306
rect 2412 29242 2464 29248
rect 2320 28416 2372 28422
rect 2320 28358 2372 28364
rect 2332 28082 2360 28358
rect 2320 28076 2372 28082
rect 2320 28018 2372 28024
rect 2424 26234 2452 29242
rect 2516 26994 2544 35866
rect 2596 30660 2648 30666
rect 2596 30602 2648 30608
rect 2608 30190 2636 30602
rect 2596 30184 2648 30190
rect 2596 30126 2648 30132
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 2424 26206 2544 26234
rect 2516 24750 2544 26206
rect 2412 24744 2464 24750
rect 2412 24686 2464 24692
rect 2504 24744 2556 24750
rect 2504 24686 2556 24692
rect 2424 21894 2452 24686
rect 2412 21888 2464 21894
rect 2412 21830 2464 21836
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 1676 20334 1728 20340
rect 1688 19854 1716 20334
rect 2148 20318 2268 20346
rect 1952 20256 2004 20262
rect 1952 20198 2004 20204
rect 1964 19854 1992 20198
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1952 19848 2004 19854
rect 1952 19790 2004 19796
rect 1688 19378 1716 19790
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1582 17232 1638 17241
rect 1582 17167 1638 17176
rect 2148 16726 2176 20318
rect 2516 19514 2544 20402
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2240 17338 2268 18158
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2332 16794 2360 17138
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2136 16720 2188 16726
rect 2136 16662 2188 16668
rect 2424 16114 2452 16934
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2424 15026 2452 16050
rect 2608 15706 2636 16050
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 1400 14408 1452 14414
rect 938 14376 994 14385
rect 1400 14350 1452 14356
rect 938 14311 994 14320
rect 952 14278 980 14311
rect 940 14272 992 14278
rect 940 14214 992 14220
rect 1492 12844 1544 12850
rect 1492 12786 1544 12792
rect 1504 12345 1532 12786
rect 1676 12776 1728 12782
rect 1674 12744 1676 12753
rect 1728 12744 1730 12753
rect 1674 12679 1730 12688
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 2226 10024 2282 10033
rect 2226 9959 2228 9968
rect 2280 9959 2282 9968
rect 2228 9930 2280 9936
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1596 9625 1624 9862
rect 1582 9616 1638 9625
rect 1582 9551 1638 9560
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6905 1624 7142
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 952 4865 980 4966
rect 938 4856 994 4865
rect 938 4791 994 4800
rect 2226 2952 2282 2961
rect 2226 2887 2228 2896
rect 2280 2887 2282 2896
rect 2228 2858 2280 2864
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 32 800 60 2790
rect 2700 2582 2728 39918
rect 3148 39908 3200 39914
rect 3148 39850 3200 39856
rect 3056 33992 3108 33998
rect 3056 33934 3108 33940
rect 3068 33658 3096 33934
rect 3056 33652 3108 33658
rect 3056 33594 3108 33600
rect 3160 33538 3188 39850
rect 2964 33516 3016 33522
rect 2964 33458 3016 33464
rect 3068 33510 3188 33538
rect 2976 33114 3004 33458
rect 2964 33108 3016 33114
rect 2964 33050 3016 33056
rect 3068 30258 3096 33510
rect 3148 33448 3200 33454
rect 3148 33390 3200 33396
rect 3160 30682 3188 33390
rect 3252 31754 3280 43658
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4632 41414 4660 43658
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 4632 41386 4844 41414
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 3424 40520 3476 40526
rect 3424 40462 3476 40468
rect 3436 37942 3464 40462
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 3516 39092 3568 39098
rect 3516 39034 3568 39040
rect 3424 37936 3476 37942
rect 3424 37878 3476 37884
rect 3332 36032 3384 36038
rect 3332 35974 3384 35980
rect 3344 35698 3372 35974
rect 3332 35692 3384 35698
rect 3332 35634 3384 35640
rect 3424 35216 3476 35222
rect 3424 35158 3476 35164
rect 3436 34678 3464 35158
rect 3424 34672 3476 34678
rect 3424 34614 3476 34620
rect 3252 31726 3372 31754
rect 3160 30654 3280 30682
rect 3148 30592 3200 30598
rect 3148 30534 3200 30540
rect 3160 30394 3188 30534
rect 3148 30388 3200 30394
rect 3148 30330 3200 30336
rect 3056 30252 3108 30258
rect 3056 30194 3108 30200
rect 2964 28416 3016 28422
rect 2964 28358 3016 28364
rect 2976 27674 3004 28358
rect 2964 27668 3016 27674
rect 2964 27610 3016 27616
rect 2872 27124 2924 27130
rect 2872 27066 2924 27072
rect 2780 26580 2832 26586
rect 2780 26522 2832 26528
rect 2792 26042 2820 26522
rect 2884 26042 2912 27066
rect 2976 26858 3004 27610
rect 3068 27538 3096 30194
rect 3252 28626 3280 30654
rect 3240 28620 3292 28626
rect 3240 28562 3292 28568
rect 3148 28076 3200 28082
rect 3148 28018 3200 28024
rect 3160 27674 3188 28018
rect 3148 27668 3200 27674
rect 3148 27610 3200 27616
rect 3056 27532 3108 27538
rect 3056 27474 3108 27480
rect 2964 26852 3016 26858
rect 2964 26794 3016 26800
rect 2780 26036 2832 26042
rect 2780 25978 2832 25984
rect 2872 26036 2924 26042
rect 2872 25978 2924 25984
rect 3238 25256 3294 25265
rect 2780 25220 2832 25226
rect 3344 25242 3372 31726
rect 3294 25214 3372 25242
rect 3238 25191 3294 25200
rect 2780 25162 2832 25168
rect 2792 24954 2820 25162
rect 3252 25158 3280 25191
rect 3240 25152 3292 25158
rect 3240 25094 3292 25100
rect 2780 24948 2832 24954
rect 2780 24890 2832 24896
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 3252 22778 3280 23666
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 2964 22432 3016 22438
rect 2964 22374 3016 22380
rect 2976 22030 3004 22374
rect 3240 22092 3292 22098
rect 3528 22094 3556 39034
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4160 38208 4212 38214
rect 4160 38150 4212 38156
rect 4172 37942 4200 38150
rect 4160 37936 4212 37942
rect 4160 37878 4212 37884
rect 3700 37868 3752 37874
rect 3700 37810 3752 37816
rect 3792 37868 3844 37874
rect 3792 37810 3844 37816
rect 3712 36922 3740 37810
rect 3804 37330 3832 37810
rect 4068 37664 4120 37670
rect 4068 37606 4120 37612
rect 3792 37324 3844 37330
rect 3792 37266 3844 37272
rect 4080 37262 4108 37606
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4068 37256 4120 37262
rect 4068 37198 4120 37204
rect 4712 37188 4764 37194
rect 4712 37130 4764 37136
rect 4436 37120 4488 37126
rect 4436 37062 4488 37068
rect 4448 36922 4476 37062
rect 3700 36916 3752 36922
rect 3700 36858 3752 36864
rect 4436 36916 4488 36922
rect 4488 36876 4660 36904
rect 4436 36858 4488 36864
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 3976 36168 4028 36174
rect 3976 36110 4028 36116
rect 3792 35692 3844 35698
rect 3792 35634 3844 35640
rect 3608 35488 3660 35494
rect 3608 35430 3660 35436
rect 3620 35086 3648 35430
rect 3608 35080 3660 35086
rect 3608 35022 3660 35028
rect 3804 34746 3832 35634
rect 3792 34740 3844 34746
rect 3792 34682 3844 34688
rect 3700 34468 3752 34474
rect 3700 34410 3752 34416
rect 3608 33992 3660 33998
rect 3608 33934 3660 33940
rect 3620 32502 3648 33934
rect 3608 32496 3660 32502
rect 3608 32438 3660 32444
rect 3712 32366 3740 34410
rect 3988 34406 4016 36110
rect 4160 36032 4212 36038
rect 4160 35974 4212 35980
rect 4528 36032 4580 36038
rect 4528 35974 4580 35980
rect 4172 35834 4200 35974
rect 4160 35828 4212 35834
rect 4160 35770 4212 35776
rect 4540 35630 4568 35974
rect 4632 35698 4660 36876
rect 4620 35692 4672 35698
rect 4620 35634 4672 35640
rect 4528 35624 4580 35630
rect 4528 35566 4580 35572
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4528 35284 4580 35290
rect 4528 35226 4580 35232
rect 4540 34762 4568 35226
rect 4632 35154 4660 35634
rect 4724 35562 4752 37130
rect 4712 35556 4764 35562
rect 4712 35498 4764 35504
rect 4620 35148 4672 35154
rect 4620 35090 4672 35096
rect 4724 34950 4752 35498
rect 4712 34944 4764 34950
rect 4712 34886 4764 34892
rect 4540 34734 4752 34762
rect 3976 34400 4028 34406
rect 3976 34342 4028 34348
rect 3884 33856 3936 33862
rect 3884 33798 3936 33804
rect 3896 33522 3924 33798
rect 3988 33522 4016 34342
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4620 33924 4672 33930
rect 4620 33866 4672 33872
rect 3884 33516 3936 33522
rect 3884 33458 3936 33464
rect 3976 33516 4028 33522
rect 3976 33458 4028 33464
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4068 33108 4120 33114
rect 4068 33050 4120 33056
rect 3976 32496 4028 32502
rect 3976 32438 4028 32444
rect 3700 32360 3752 32366
rect 3700 32302 3752 32308
rect 3712 32026 3740 32302
rect 3700 32020 3752 32026
rect 3700 31962 3752 31968
rect 3988 31754 4016 32438
rect 4080 32230 4108 33050
rect 4632 32978 4660 33866
rect 4724 33046 4752 34734
rect 4712 33040 4764 33046
rect 4712 32982 4764 32988
rect 4160 32972 4212 32978
rect 4160 32914 4212 32920
rect 4620 32972 4672 32978
rect 4620 32914 4672 32920
rect 4172 32434 4200 32914
rect 4252 32904 4304 32910
rect 4252 32846 4304 32852
rect 4160 32428 4212 32434
rect 4160 32370 4212 32376
rect 4264 32366 4292 32846
rect 4528 32768 4580 32774
rect 4528 32710 4580 32716
rect 4252 32360 4304 32366
rect 4252 32302 4304 32308
rect 4540 32298 4568 32710
rect 4620 32360 4672 32366
rect 4620 32302 4672 32308
rect 4528 32292 4580 32298
rect 4528 32234 4580 32240
rect 4068 32224 4120 32230
rect 4068 32166 4120 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3988 31726 4108 31754
rect 4080 30818 4108 31726
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4080 30790 4200 30818
rect 4172 30598 4200 30790
rect 4632 30666 4660 32302
rect 4724 31958 4752 32982
rect 4712 31952 4764 31958
rect 4712 31894 4764 31900
rect 4712 31816 4764 31822
rect 4712 31758 4764 31764
rect 4620 30660 4672 30666
rect 4620 30602 4672 30608
rect 3792 30592 3844 30598
rect 3792 30534 3844 30540
rect 4160 30592 4212 30598
rect 4160 30534 4212 30540
rect 3804 30326 3832 30534
rect 4632 30394 4660 30602
rect 4620 30388 4672 30394
rect 4620 30330 4672 30336
rect 3792 30320 3844 30326
rect 3792 30262 3844 30268
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4620 29096 4672 29102
rect 4620 29038 4672 29044
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4436 28552 4488 28558
rect 4436 28494 4488 28500
rect 4528 28552 4580 28558
rect 4528 28494 4580 28500
rect 4068 28416 4120 28422
rect 4068 28358 4120 28364
rect 3976 27872 4028 27878
rect 3976 27814 4028 27820
rect 3608 27532 3660 27538
rect 3608 27474 3660 27480
rect 3240 22034 3292 22040
rect 3436 22066 3556 22094
rect 2964 22024 3016 22030
rect 2964 21966 3016 21972
rect 2964 20800 3016 20806
rect 2964 20742 3016 20748
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 2976 20602 3004 20742
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 2976 19514 3004 19994
rect 3068 19514 3096 20742
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3252 19310 3280 22034
rect 3332 20324 3384 20330
rect 3332 20266 3384 20272
rect 3344 19446 3372 20266
rect 3332 19440 3384 19446
rect 3332 19382 3384 19388
rect 3240 19304 3292 19310
rect 3240 19246 3292 19252
rect 3252 18970 3280 19246
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3436 18358 3464 22066
rect 3516 20256 3568 20262
rect 3516 20198 3568 20204
rect 3528 19854 3556 20198
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 2964 18352 3016 18358
rect 2964 18294 3016 18300
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 2976 17882 3004 18294
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 3068 18193 3096 18226
rect 3620 18222 3648 27474
rect 3988 27470 4016 27814
rect 3976 27464 4028 27470
rect 3976 27406 4028 27412
rect 3988 26874 4016 27406
rect 4080 27334 4108 28358
rect 4448 27860 4476 28494
rect 4540 28150 4568 28494
rect 4528 28144 4580 28150
rect 4528 28086 4580 28092
rect 4632 28082 4660 29038
rect 4620 28076 4672 28082
rect 4620 28018 4672 28024
rect 4448 27832 4660 27860
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27674 4660 27832
rect 4620 27668 4672 27674
rect 4620 27610 4672 27616
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4080 27130 4108 27270
rect 4068 27124 4120 27130
rect 4068 27066 4120 27072
rect 4620 26988 4672 26994
rect 4620 26930 4672 26936
rect 3988 26846 4108 26874
rect 3976 26784 4028 26790
rect 3976 26726 4028 26732
rect 3988 26382 4016 26726
rect 4080 26450 4108 26846
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4528 26580 4580 26586
rect 4528 26522 4580 26528
rect 4068 26444 4120 26450
rect 4068 26386 4120 26392
rect 3976 26376 4028 26382
rect 3976 26318 4028 26324
rect 3884 26240 3936 26246
rect 3884 26182 3936 26188
rect 3896 25294 3924 26182
rect 4080 25906 4108 26386
rect 4252 26376 4304 26382
rect 4252 26318 4304 26324
rect 4068 25900 4120 25906
rect 4068 25842 4120 25848
rect 4264 25838 4292 26318
rect 4540 25945 4568 26522
rect 4632 26450 4660 26930
rect 4724 26625 4752 31758
rect 4816 30818 4844 41386
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 10048 41268 10100 41274
rect 10048 41210 10100 41216
rect 8944 40520 8996 40526
rect 8944 40462 8996 40468
rect 8852 40452 8904 40458
rect 8852 40394 8904 40400
rect 6920 40384 6972 40390
rect 6920 40326 6972 40332
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 6932 39846 6960 40326
rect 8864 40186 8892 40394
rect 8852 40180 8904 40186
rect 8852 40122 8904 40128
rect 6920 39840 6972 39846
rect 6920 39782 6972 39788
rect 6932 39574 6960 39782
rect 6920 39568 6972 39574
rect 6920 39510 6972 39516
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 7656 38956 7708 38962
rect 7656 38898 7708 38904
rect 7380 38752 7432 38758
rect 7380 38694 7432 38700
rect 5356 38548 5408 38554
rect 5356 38490 5408 38496
rect 5264 38344 5316 38350
rect 5264 38286 5316 38292
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 5172 37664 5224 37670
rect 5172 37606 5224 37612
rect 5184 37262 5212 37606
rect 5276 37466 5304 38286
rect 5264 37460 5316 37466
rect 5264 37402 5316 37408
rect 5172 37256 5224 37262
rect 5172 37198 5224 37204
rect 5264 37120 5316 37126
rect 5264 37062 5316 37068
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 5276 36922 5304 37062
rect 5264 36916 5316 36922
rect 5264 36858 5316 36864
rect 5276 36174 5304 36858
rect 5264 36168 5316 36174
rect 5264 36110 5316 36116
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 5276 35894 5304 36110
rect 5368 36038 5396 38490
rect 7392 38350 7420 38694
rect 5632 38344 5684 38350
rect 5632 38286 5684 38292
rect 7380 38344 7432 38350
rect 7380 38286 7432 38292
rect 5644 37806 5672 38286
rect 6000 38276 6052 38282
rect 6000 38218 6052 38224
rect 6012 38010 6040 38218
rect 7012 38208 7064 38214
rect 7012 38150 7064 38156
rect 7024 38010 7052 38150
rect 6000 38004 6052 38010
rect 6000 37946 6052 37952
rect 7012 38004 7064 38010
rect 7012 37946 7064 37952
rect 6460 37936 6512 37942
rect 6460 37878 6512 37884
rect 6276 37868 6328 37874
rect 6276 37810 6328 37816
rect 5632 37800 5684 37806
rect 5632 37742 5684 37748
rect 6288 37262 6316 37810
rect 6472 37398 6500 37878
rect 6460 37392 6512 37398
rect 6460 37334 6512 37340
rect 7024 37262 7052 37946
rect 7196 37324 7248 37330
rect 7196 37266 7248 37272
rect 6276 37256 6328 37262
rect 6276 37198 6328 37204
rect 6644 37256 6696 37262
rect 6644 37198 6696 37204
rect 7012 37256 7064 37262
rect 7012 37198 7064 37204
rect 5448 37188 5500 37194
rect 5448 37130 5500 37136
rect 5460 36718 5488 37130
rect 6656 36922 6684 37198
rect 7104 37188 7156 37194
rect 7104 37130 7156 37136
rect 6644 36916 6696 36922
rect 6644 36858 6696 36864
rect 7116 36854 7144 37130
rect 7104 36848 7156 36854
rect 7104 36790 7156 36796
rect 6920 36780 6972 36786
rect 6920 36722 6972 36728
rect 5448 36712 5500 36718
rect 5448 36654 5500 36660
rect 5356 36032 5408 36038
rect 5356 35974 5408 35980
rect 5276 35866 5396 35894
rect 5264 35828 5316 35834
rect 5264 35770 5316 35776
rect 5276 35698 5304 35770
rect 5264 35692 5316 35698
rect 5264 35634 5316 35640
rect 4988 35624 5040 35630
rect 4988 35566 5040 35572
rect 5172 35624 5224 35630
rect 5172 35566 5224 35572
rect 4896 35488 4948 35494
rect 4896 35430 4948 35436
rect 4908 35154 4936 35430
rect 5000 35290 5028 35566
rect 4988 35284 5040 35290
rect 4988 35226 5040 35232
rect 5184 35154 5212 35566
rect 5276 35154 5304 35634
rect 4896 35148 4948 35154
rect 4896 35090 4948 35096
rect 5172 35148 5224 35154
rect 5172 35090 5224 35096
rect 5264 35148 5316 35154
rect 5264 35090 5316 35096
rect 4908 35034 4936 35090
rect 4908 35006 5304 35034
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 5276 32994 5304 35006
rect 5368 34678 5396 35866
rect 5356 34672 5408 34678
rect 5356 34614 5408 34620
rect 5460 34066 5488 36654
rect 5632 35624 5684 35630
rect 5632 35566 5684 35572
rect 5540 34944 5592 34950
rect 5540 34886 5592 34892
rect 5448 34060 5500 34066
rect 5448 34002 5500 34008
rect 5552 33946 5580 34886
rect 5356 33924 5408 33930
rect 5356 33866 5408 33872
rect 5460 33918 5580 33946
rect 5368 33658 5396 33866
rect 5356 33652 5408 33658
rect 5356 33594 5408 33600
rect 5276 32966 5396 32994
rect 4988 32904 5040 32910
rect 5040 32852 5304 32858
rect 4988 32846 5304 32852
rect 5000 32830 5304 32846
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4988 32564 5040 32570
rect 5276 32552 5304 32830
rect 5368 32774 5396 32966
rect 5356 32768 5408 32774
rect 5356 32710 5408 32716
rect 5040 32524 5304 32552
rect 4988 32506 5040 32512
rect 5000 32434 5028 32506
rect 4988 32428 5040 32434
rect 4988 32370 5040 32376
rect 5264 31952 5316 31958
rect 5264 31894 5316 31900
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4988 31272 5040 31278
rect 4988 31214 5040 31220
rect 5000 30938 5028 31214
rect 5276 30954 5304 31894
rect 5368 31822 5396 32710
rect 5460 32366 5488 33918
rect 5644 32978 5672 35566
rect 6092 35488 6144 35494
rect 6092 35430 6144 35436
rect 6828 35488 6880 35494
rect 6828 35430 6880 35436
rect 6104 35290 6132 35430
rect 6092 35284 6144 35290
rect 6092 35226 6144 35232
rect 6090 35184 6146 35193
rect 6090 35119 6092 35128
rect 6144 35119 6146 35128
rect 6092 35090 6144 35096
rect 6840 35086 6868 35430
rect 6552 35080 6604 35086
rect 6552 35022 6604 35028
rect 6828 35080 6880 35086
rect 6828 35022 6880 35028
rect 6276 34944 6328 34950
rect 6276 34886 6328 34892
rect 6288 34678 6316 34886
rect 6276 34672 6328 34678
rect 6276 34614 6328 34620
rect 6564 34610 6592 35022
rect 6932 34950 6960 36722
rect 7208 36242 7236 37266
rect 7668 37126 7696 38898
rect 8956 38282 8984 40462
rect 10060 40118 10088 41210
rect 10244 41177 10272 47602
rect 11336 47048 11388 47054
rect 11336 46990 11388 46996
rect 11348 41682 11376 46990
rect 13728 44872 13780 44878
rect 13728 44814 13780 44820
rect 13740 43246 13768 44814
rect 15212 43450 15240 47602
rect 17328 47258 17356 47602
rect 18236 47456 18288 47462
rect 18236 47398 18288 47404
rect 17316 47252 17368 47258
rect 17316 47194 17368 47200
rect 17868 47116 17920 47122
rect 17868 47058 17920 47064
rect 17132 46912 17184 46918
rect 17132 46854 17184 46860
rect 17500 46912 17552 46918
rect 17500 46854 17552 46860
rect 17592 46912 17644 46918
rect 17592 46854 17644 46860
rect 16948 46572 17000 46578
rect 16948 46514 17000 46520
rect 15660 46368 15712 46374
rect 15660 46310 15712 46316
rect 15568 45280 15620 45286
rect 15568 45222 15620 45228
rect 15384 44804 15436 44810
rect 15384 44746 15436 44752
rect 15396 44538 15424 44746
rect 15384 44532 15436 44538
rect 15384 44474 15436 44480
rect 15580 44402 15608 45222
rect 15672 44878 15700 46310
rect 16960 46170 16988 46514
rect 16948 46164 17000 46170
rect 16948 46106 17000 46112
rect 17144 45966 17172 46854
rect 17512 46714 17540 46854
rect 17500 46708 17552 46714
rect 17500 46650 17552 46656
rect 17512 45966 17540 46650
rect 17132 45960 17184 45966
rect 17132 45902 17184 45908
rect 17500 45960 17552 45966
rect 17500 45902 17552 45908
rect 17604 45830 17632 46854
rect 17684 46504 17736 46510
rect 17684 46446 17736 46452
rect 17696 45898 17724 46446
rect 17880 46034 17908 47058
rect 18248 47054 18276 47398
rect 19260 47054 19288 47602
rect 19432 47456 19484 47462
rect 19432 47398 19484 47404
rect 18236 47048 18288 47054
rect 18236 46990 18288 46996
rect 18420 47048 18472 47054
rect 18420 46990 18472 46996
rect 19248 47048 19300 47054
rect 19248 46990 19300 46996
rect 17960 46572 18012 46578
rect 17960 46514 18012 46520
rect 17868 46028 17920 46034
rect 17868 45970 17920 45976
rect 17684 45892 17736 45898
rect 17684 45834 17736 45840
rect 15936 45824 15988 45830
rect 15936 45766 15988 45772
rect 17592 45824 17644 45830
rect 17592 45766 17644 45772
rect 15660 44872 15712 44878
rect 15660 44814 15712 44820
rect 15568 44396 15620 44402
rect 15568 44338 15620 44344
rect 15948 43926 15976 45766
rect 16856 45484 16908 45490
rect 16856 45426 16908 45432
rect 16868 45014 16896 45426
rect 17132 45416 17184 45422
rect 17132 45358 17184 45364
rect 17316 45416 17368 45422
rect 17316 45358 17368 45364
rect 17144 45082 17172 45358
rect 17132 45076 17184 45082
rect 17132 45018 17184 45024
rect 16856 45008 16908 45014
rect 16856 44950 16908 44956
rect 16580 44940 16632 44946
rect 16580 44882 16632 44888
rect 16488 44736 16540 44742
rect 16488 44678 16540 44684
rect 16500 44402 16528 44678
rect 16488 44396 16540 44402
rect 16488 44338 16540 44344
rect 15936 43920 15988 43926
rect 15936 43862 15988 43868
rect 15476 43784 15528 43790
rect 15476 43726 15528 43732
rect 15200 43444 15252 43450
rect 15200 43386 15252 43392
rect 15108 43308 15160 43314
rect 15108 43250 15160 43256
rect 13728 43240 13780 43246
rect 13728 43182 13780 43188
rect 13740 42770 13768 43182
rect 13728 42764 13780 42770
rect 13728 42706 13780 42712
rect 13268 42628 13320 42634
rect 13268 42570 13320 42576
rect 13280 42362 13308 42570
rect 13268 42356 13320 42362
rect 13268 42298 13320 42304
rect 12716 42220 12768 42226
rect 12716 42162 12768 42168
rect 13544 42220 13596 42226
rect 13544 42162 13596 42168
rect 11336 41676 11388 41682
rect 11336 41618 11388 41624
rect 11348 41206 11376 41618
rect 11336 41200 11388 41206
rect 10230 41168 10286 41177
rect 11336 41142 11388 41148
rect 10230 41103 10286 41112
rect 12164 41132 12216 41138
rect 10244 40730 10272 41103
rect 12164 41074 12216 41080
rect 10692 40996 10744 41002
rect 10692 40938 10744 40944
rect 10232 40724 10284 40730
rect 10232 40666 10284 40672
rect 10704 40526 10732 40938
rect 10784 40928 10836 40934
rect 10784 40870 10836 40876
rect 11520 40928 11572 40934
rect 11520 40870 11572 40876
rect 10796 40594 10824 40870
rect 10784 40588 10836 40594
rect 10784 40530 10836 40536
rect 10692 40520 10744 40526
rect 10692 40462 10744 40468
rect 10416 40384 10468 40390
rect 10416 40326 10468 40332
rect 10048 40112 10100 40118
rect 10048 40054 10100 40060
rect 10060 39846 10088 40054
rect 10428 40050 10456 40326
rect 11532 40050 11560 40870
rect 12176 40730 12204 41074
rect 12164 40724 12216 40730
rect 12084 40684 12164 40712
rect 11888 40112 11940 40118
rect 11888 40054 11940 40060
rect 10416 40044 10468 40050
rect 10416 39986 10468 39992
rect 10600 40044 10652 40050
rect 10600 39986 10652 39992
rect 11336 40044 11388 40050
rect 11336 39986 11388 39992
rect 11520 40044 11572 40050
rect 11520 39986 11572 39992
rect 10232 39976 10284 39982
rect 10232 39918 10284 39924
rect 10244 39846 10272 39918
rect 9036 39840 9088 39846
rect 9036 39782 9088 39788
rect 10048 39840 10100 39846
rect 10048 39782 10100 39788
rect 10232 39840 10284 39846
rect 10232 39782 10284 39788
rect 9048 39302 9076 39782
rect 9036 39296 9088 39302
rect 9036 39238 9088 39244
rect 8944 38276 8996 38282
rect 8944 38218 8996 38224
rect 8484 38208 8536 38214
rect 8484 38150 8536 38156
rect 8760 38208 8812 38214
rect 8760 38150 8812 38156
rect 8496 37874 8524 38150
rect 8772 37874 8800 38150
rect 8484 37868 8536 37874
rect 8484 37810 8536 37816
rect 8760 37868 8812 37874
rect 8760 37810 8812 37816
rect 7748 37732 7800 37738
rect 7748 37674 7800 37680
rect 7288 37120 7340 37126
rect 7288 37062 7340 37068
rect 7656 37120 7708 37126
rect 7656 37062 7708 37068
rect 7300 36854 7328 37062
rect 7760 36922 7788 37674
rect 8496 37330 8524 37810
rect 8484 37324 8536 37330
rect 8484 37266 8536 37272
rect 8772 37262 8800 37810
rect 8760 37256 8812 37262
rect 8760 37198 8812 37204
rect 7748 36916 7800 36922
rect 7748 36858 7800 36864
rect 7288 36848 7340 36854
rect 7288 36790 7340 36796
rect 8208 36712 8260 36718
rect 8208 36654 8260 36660
rect 7196 36236 7248 36242
rect 7196 36178 7248 36184
rect 7656 36236 7708 36242
rect 7656 36178 7708 36184
rect 7668 35630 7696 36178
rect 7932 35692 7984 35698
rect 7932 35634 7984 35640
rect 7656 35624 7708 35630
rect 7656 35566 7708 35572
rect 6920 34944 6972 34950
rect 6920 34886 6972 34892
rect 6552 34604 6604 34610
rect 6552 34546 6604 34552
rect 6564 33266 6592 34546
rect 6380 33238 6592 33266
rect 5632 32972 5684 32978
rect 5632 32914 5684 32920
rect 5448 32360 5500 32366
rect 5448 32302 5500 32308
rect 5356 31816 5408 31822
rect 5356 31758 5408 31764
rect 5446 31784 5502 31793
rect 5446 31719 5502 31728
rect 5460 31278 5488 31719
rect 5448 31272 5500 31278
rect 5448 31214 5500 31220
rect 4988 30932 5040 30938
rect 5276 30926 5488 30954
rect 4988 30874 5040 30880
rect 5460 30818 5488 30926
rect 4816 30790 5212 30818
rect 5460 30790 5580 30818
rect 4804 30728 4856 30734
rect 4804 30670 4856 30676
rect 4816 30054 4844 30670
rect 5184 30648 5212 30790
rect 5448 30660 5500 30666
rect 5184 30620 5396 30648
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4804 30048 4856 30054
rect 4804 29990 4856 29996
rect 4816 29102 4844 29990
rect 5264 29776 5316 29782
rect 5264 29718 5316 29724
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 5276 27044 5304 29718
rect 5000 27016 5304 27044
rect 4710 26616 4766 26625
rect 4710 26551 4766 26560
rect 4710 26480 4766 26489
rect 4620 26444 4672 26450
rect 4766 26424 4844 26432
rect 4710 26415 4712 26424
rect 4620 26386 4672 26392
rect 4764 26404 4844 26424
rect 4712 26386 4764 26392
rect 4620 26240 4672 26246
rect 4620 26182 4672 26188
rect 4526 25936 4582 25945
rect 4526 25871 4582 25880
rect 4252 25832 4304 25838
rect 4252 25774 4304 25780
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3884 25288 3936 25294
rect 3884 25230 3936 25236
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24290 4660 26182
rect 4712 25764 4764 25770
rect 4712 25706 4764 25712
rect 4448 24262 4660 24290
rect 3700 24132 3752 24138
rect 3700 24074 3752 24080
rect 3712 22710 3740 24074
rect 3790 23624 3846 23633
rect 4448 23610 4476 24262
rect 4528 24200 4580 24206
rect 4528 24142 4580 24148
rect 3790 23559 3846 23568
rect 4080 23582 4476 23610
rect 3804 23254 3832 23559
rect 3792 23248 3844 23254
rect 3792 23190 3844 23196
rect 3804 22778 3832 23190
rect 3792 22772 3844 22778
rect 3792 22714 3844 22720
rect 3700 22704 3752 22710
rect 3700 22646 3752 22652
rect 3712 21894 3740 22646
rect 3792 22568 3844 22574
rect 3792 22510 3844 22516
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 3804 21010 3832 22510
rect 4080 22114 4108 23582
rect 4540 23526 4568 24142
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4528 23520 4580 23526
rect 4528 23462 4580 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23186 4660 24006
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4528 23112 4580 23118
rect 4528 23054 4580 23060
rect 4540 22681 4568 23054
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4526 22672 4582 22681
rect 4526 22607 4582 22616
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4080 22086 4200 22114
rect 4172 21434 4200 22086
rect 4632 22030 4660 22918
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4080 21406 4200 21434
rect 4080 21026 4108 21406
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3792 21004 3844 21010
rect 4080 20998 4200 21026
rect 3792 20946 3844 20952
rect 3608 18216 3660 18222
rect 3054 18184 3110 18193
rect 3608 18158 3660 18164
rect 3054 18119 3110 18128
rect 3332 18148 3384 18154
rect 3332 18090 3384 18096
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 3344 17678 3372 18090
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3804 17338 3832 20946
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 3884 20596 3936 20602
rect 3884 20538 3936 20544
rect 3896 19922 3924 20538
rect 3988 20534 4016 20742
rect 3976 20528 4028 20534
rect 3976 20470 4028 20476
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 3884 19916 3936 19922
rect 3884 19858 3936 19864
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3988 19446 4016 19654
rect 4080 19446 4108 20334
rect 4172 20330 4200 20998
rect 4724 20398 4752 25706
rect 4816 24206 4844 26404
rect 5000 26246 5028 27016
rect 5080 26852 5132 26858
rect 5080 26794 5132 26800
rect 5092 26450 5120 26794
rect 5080 26444 5132 26450
rect 5080 26386 5132 26392
rect 4988 26240 5040 26246
rect 5092 26228 5120 26386
rect 5092 26200 5304 26228
rect 4988 26182 5040 26188
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4894 25936 4950 25945
rect 5276 25922 5304 26200
rect 5092 25906 5304 25922
rect 4894 25871 4896 25880
rect 4948 25871 4950 25880
rect 5080 25900 5304 25906
rect 4896 25842 4948 25848
rect 5132 25894 5304 25900
rect 5368 25922 5396 30620
rect 5448 30602 5500 30608
rect 5460 30394 5488 30602
rect 5448 30388 5500 30394
rect 5448 30330 5500 30336
rect 5552 30274 5580 30790
rect 5460 30246 5580 30274
rect 5460 29594 5488 30246
rect 5460 29566 5580 29594
rect 5448 29504 5500 29510
rect 5448 29446 5500 29452
rect 5460 29238 5488 29446
rect 5448 29232 5500 29238
rect 5448 29174 5500 29180
rect 5552 29050 5580 29566
rect 5460 29022 5580 29050
rect 5460 26024 5488 29022
rect 5644 26586 5672 32914
rect 6380 32366 6408 33238
rect 6564 33114 6592 33238
rect 6552 33108 6604 33114
rect 6552 33050 6604 33056
rect 7668 32978 7696 35566
rect 7944 35222 7972 35634
rect 7932 35216 7984 35222
rect 7932 35158 7984 35164
rect 7944 34762 7972 35158
rect 8220 35154 8248 36654
rect 8944 35692 8996 35698
rect 8944 35634 8996 35640
rect 8300 35488 8352 35494
rect 8300 35430 8352 35436
rect 8208 35148 8260 35154
rect 8208 35090 8260 35096
rect 7944 34734 8064 34762
rect 8036 34678 8064 34734
rect 8024 34672 8076 34678
rect 8024 34614 8076 34620
rect 8220 32978 8248 35090
rect 8312 34610 8340 35430
rect 8956 35290 8984 35634
rect 8944 35284 8996 35290
rect 8944 35226 8996 35232
rect 8668 35148 8720 35154
rect 8668 35090 8720 35096
rect 8392 35012 8444 35018
rect 8392 34954 8444 34960
rect 8404 34746 8432 34954
rect 8392 34740 8444 34746
rect 8392 34682 8444 34688
rect 8300 34604 8352 34610
rect 8300 34546 8352 34552
rect 7104 32972 7156 32978
rect 7104 32914 7156 32920
rect 7656 32972 7708 32978
rect 7656 32914 7708 32920
rect 8208 32972 8260 32978
rect 8208 32914 8260 32920
rect 6736 32768 6788 32774
rect 6736 32710 6788 32716
rect 6920 32768 6972 32774
rect 6920 32710 6972 32716
rect 6748 32502 6776 32710
rect 6736 32496 6788 32502
rect 6736 32438 6788 32444
rect 6368 32360 6420 32366
rect 6420 32308 6776 32314
rect 6368 32302 6776 32308
rect 5724 32292 5776 32298
rect 5724 32234 5776 32240
rect 6380 32286 6776 32302
rect 5736 31754 5764 32234
rect 6276 32020 6328 32026
rect 6276 31962 6328 31968
rect 5736 31726 5856 31754
rect 5632 26580 5684 26586
rect 5632 26522 5684 26528
rect 5724 26512 5776 26518
rect 5724 26454 5776 26460
rect 5460 25996 5672 26024
rect 5368 25894 5580 25922
rect 5080 25842 5132 25848
rect 5356 25832 5408 25838
rect 5408 25792 5488 25820
rect 5356 25774 5408 25780
rect 5172 25696 5224 25702
rect 5172 25638 5224 25644
rect 5184 25498 5212 25638
rect 5172 25492 5224 25498
rect 5172 25434 5224 25440
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5264 24948 5316 24954
rect 5264 24890 5316 24896
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4804 24064 4856 24070
rect 4804 24006 4856 24012
rect 4816 23576 4844 24006
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5276 23848 5304 24890
rect 5184 23820 5304 23848
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 4896 23588 4948 23594
rect 4816 23548 4896 23576
rect 4896 23530 4948 23536
rect 4908 23118 4936 23530
rect 5092 23186 5120 23598
rect 5184 23497 5212 23820
rect 5264 23656 5316 23662
rect 5262 23624 5264 23633
rect 5316 23624 5318 23633
rect 5318 23582 5396 23610
rect 5262 23559 5318 23568
rect 5170 23488 5226 23497
rect 5170 23423 5226 23432
rect 5184 23186 5212 23423
rect 5080 23180 5132 23186
rect 5080 23122 5132 23128
rect 5172 23180 5224 23186
rect 5172 23122 5224 23128
rect 4896 23112 4948 23118
rect 4896 23054 4948 23060
rect 5092 22964 5120 23122
rect 5368 23100 5396 23582
rect 5460 23361 5488 25792
rect 5552 24886 5580 25894
rect 5644 24954 5672 25996
rect 5632 24948 5684 24954
rect 5632 24890 5684 24896
rect 5540 24880 5592 24886
rect 5540 24822 5592 24828
rect 5736 24732 5764 26454
rect 5552 24704 5764 24732
rect 5552 23730 5580 24704
rect 5540 23724 5592 23730
rect 5540 23666 5592 23672
rect 5552 23526 5580 23666
rect 5724 23656 5776 23662
rect 5644 23616 5724 23644
rect 5540 23520 5592 23526
rect 5540 23462 5592 23468
rect 5446 23352 5502 23361
rect 5644 23338 5672 23616
rect 5724 23598 5776 23604
rect 5446 23287 5502 23296
rect 5552 23310 5672 23338
rect 5448 23112 5500 23118
rect 5368 23072 5448 23100
rect 5448 23054 5500 23060
rect 5092 22936 5396 22964
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5368 22778 5396 22936
rect 5446 22944 5502 22953
rect 5446 22879 5502 22888
rect 4804 22772 4856 22778
rect 4804 22714 4856 22720
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 4816 22574 4844 22714
rect 5262 22672 5318 22681
rect 5262 22607 5318 22616
rect 5356 22636 5408 22642
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 4816 22234 4844 22510
rect 5276 22234 5304 22607
rect 5356 22578 5408 22584
rect 5368 22234 5396 22578
rect 4804 22228 4856 22234
rect 4804 22170 4856 22176
rect 5264 22228 5316 22234
rect 5264 22170 5316 22176
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5460 21842 5488 22879
rect 5552 22438 5580 23310
rect 5644 23186 5672 23310
rect 5722 23216 5778 23225
rect 5632 23180 5684 23186
rect 5722 23151 5778 23160
rect 5632 23122 5684 23128
rect 5736 23118 5764 23151
rect 5724 23112 5776 23118
rect 5724 23054 5776 23060
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 5644 22710 5672 22918
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 5632 22704 5684 22710
rect 5632 22646 5684 22652
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 5644 21842 5672 22646
rect 5736 22030 5764 22714
rect 5828 22030 5856 31726
rect 5908 28688 5960 28694
rect 5908 28630 5960 28636
rect 5920 27470 5948 28630
rect 5908 27464 5960 27470
rect 5908 27406 5960 27412
rect 5908 27328 5960 27334
rect 5908 27270 5960 27276
rect 5724 22024 5776 22030
rect 5724 21966 5776 21972
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5816 21888 5868 21894
rect 5460 21814 5580 21842
rect 5644 21814 5764 21842
rect 5816 21830 5868 21836
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 4816 20584 4844 20878
rect 5356 20868 5408 20874
rect 5356 20810 5408 20816
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4816 20556 4936 20584
rect 4436 20392 4488 20398
rect 4712 20392 4764 20398
rect 4488 20340 4660 20346
rect 4436 20334 4660 20340
rect 4764 20340 4844 20346
rect 4712 20334 4844 20340
rect 4160 20324 4212 20330
rect 4448 20318 4660 20334
rect 4724 20318 4844 20334
rect 4160 20266 4212 20272
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4160 19984 4212 19990
rect 4632 19938 4660 20318
rect 4712 20256 4764 20262
rect 4712 20198 4764 20204
rect 4160 19926 4212 19932
rect 3976 19440 4028 19446
rect 3976 19382 4028 19388
rect 4068 19440 4120 19446
rect 4068 19382 4120 19388
rect 4172 19378 4200 19926
rect 4540 19910 4660 19938
rect 4540 19854 4568 19910
rect 4724 19854 4752 20198
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4540 19514 4568 19790
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4816 19378 4844 20318
rect 4908 20262 4936 20556
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4908 19990 4936 20198
rect 5170 20088 5226 20097
rect 5170 20023 5226 20032
rect 5184 19990 5212 20023
rect 4896 19984 4948 19990
rect 4896 19926 4948 19932
rect 5172 19984 5224 19990
rect 5172 19926 5224 19932
rect 5184 19802 5212 19926
rect 5276 19922 5304 20334
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 5184 19774 5304 19802
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 3896 17882 3924 18226
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3804 16658 3832 17274
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3988 16046 4016 18906
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4436 18216 4488 18222
rect 4488 18176 4752 18204
rect 4436 18158 4488 18164
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4528 17740 4580 17746
rect 4632 17728 4660 18022
rect 4724 17882 4752 18176
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 5276 17762 5304 19774
rect 5368 19514 5396 20810
rect 5552 20466 5580 21814
rect 5540 20460 5592 20466
rect 5592 20420 5672 20448
rect 5540 20402 5592 20408
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5460 20058 5488 20334
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5460 19904 5488 19994
rect 5540 19916 5592 19922
rect 5460 19876 5540 19904
rect 5540 19858 5592 19864
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5356 19372 5408 19378
rect 5644 19334 5672 20420
rect 5736 20398 5764 21814
rect 5828 21690 5856 21830
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5356 19314 5408 19320
rect 4580 17700 4660 17728
rect 4712 17740 4764 17746
rect 4528 17682 4580 17688
rect 4712 17682 4764 17688
rect 4804 17740 4856 17746
rect 5000 17734 5304 17762
rect 5000 17728 5028 17734
rect 4856 17700 5028 17728
rect 4804 17682 4856 17688
rect 4160 17672 4212 17678
rect 4264 17649 4292 17682
rect 4160 17614 4212 17620
rect 4250 17640 4306 17649
rect 4172 17134 4200 17614
rect 4250 17575 4306 17584
rect 4540 17202 4568 17682
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 4724 17134 4752 17682
rect 5264 17672 5316 17678
rect 5170 17640 5226 17649
rect 5264 17614 5316 17620
rect 5170 17575 5226 17584
rect 5184 17542 5212 17575
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4620 17060 4672 17066
rect 4620 17002 4672 17008
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4264 16114 4292 16390
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 3804 15502 3832 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15502 4660 17002
rect 4724 16590 4752 17070
rect 4816 16794 4844 17478
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5276 17134 5304 17614
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5276 16250 5304 17070
rect 5368 16998 5396 19314
rect 5460 19306 5672 19334
rect 5460 18170 5488 19306
rect 5460 18142 5580 18170
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5368 16658 5396 16934
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5460 16590 5488 18022
rect 5552 17134 5580 18142
rect 5816 17876 5868 17882
rect 5816 17818 5868 17824
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3712 14618 3740 14962
rect 4172 14906 4200 15302
rect 4632 15162 4660 15438
rect 4724 15366 4752 16050
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 5736 15502 5764 15914
rect 5828 15502 5856 17818
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5276 15162 5304 15302
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5828 15094 5856 15438
rect 5816 15088 5868 15094
rect 5816 15030 5868 15036
rect 4080 14878 4200 14906
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 4080 14414 4108 14878
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4264 12918 4292 13126
rect 4448 12986 4476 13262
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 3712 12306 3740 12718
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3712 11218 3740 12242
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4172 11898 4200 12106
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5276 11898 5304 12378
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5644 11762 5672 12718
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 5644 11150 5672 11494
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5920 2650 5948 27270
rect 6288 26586 6316 31962
rect 6380 31890 6408 32286
rect 6748 32230 6776 32286
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6736 32224 6788 32230
rect 6736 32166 6788 32172
rect 6368 31884 6420 31890
rect 6368 31826 6420 31832
rect 6656 31822 6684 32166
rect 6644 31816 6696 31822
rect 6644 31758 6696 31764
rect 6932 31346 6960 32710
rect 6920 31340 6972 31346
rect 6920 31282 6972 31288
rect 6828 30592 6880 30598
rect 6828 30534 6880 30540
rect 6840 30394 6868 30534
rect 6828 30388 6880 30394
rect 6828 30330 6880 30336
rect 6840 29714 6868 30330
rect 6828 29708 6880 29714
rect 6828 29650 6880 29656
rect 6368 29640 6420 29646
rect 6368 29582 6420 29588
rect 6380 29306 6408 29582
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 6368 29300 6420 29306
rect 6368 29242 6420 29248
rect 6736 29164 6788 29170
rect 6736 29106 6788 29112
rect 6748 28694 6776 29106
rect 6736 28688 6788 28694
rect 6736 28630 6788 28636
rect 6748 28558 6776 28630
rect 6460 28552 6512 28558
rect 6460 28494 6512 28500
rect 6736 28552 6788 28558
rect 6736 28494 6788 28500
rect 6472 27674 6500 28494
rect 6828 28416 6880 28422
rect 6828 28358 6880 28364
rect 6840 28150 6868 28358
rect 6828 28144 6880 28150
rect 6828 28086 6880 28092
rect 6932 28082 6960 29446
rect 7116 28626 7144 32914
rect 7564 32904 7616 32910
rect 7564 32846 7616 32852
rect 7576 32026 7604 32846
rect 7748 32768 7800 32774
rect 7748 32710 7800 32716
rect 7840 32768 7892 32774
rect 7840 32710 7892 32716
rect 8208 32768 8260 32774
rect 8208 32710 8260 32716
rect 8484 32768 8536 32774
rect 8484 32710 8536 32716
rect 7760 32570 7788 32710
rect 7748 32564 7800 32570
rect 7748 32506 7800 32512
rect 7852 32434 7880 32710
rect 7840 32428 7892 32434
rect 7840 32370 7892 32376
rect 8220 32230 8248 32710
rect 8208 32224 8260 32230
rect 8208 32166 8260 32172
rect 8220 32026 8248 32166
rect 7564 32020 7616 32026
rect 7564 31962 7616 31968
rect 8208 32020 8260 32026
rect 8208 31962 8260 31968
rect 8496 31686 8524 32710
rect 8680 31890 8708 35090
rect 8944 32428 8996 32434
rect 8944 32370 8996 32376
rect 8956 32026 8984 32370
rect 8944 32020 8996 32026
rect 8944 31962 8996 31968
rect 8668 31884 8720 31890
rect 8668 31826 8720 31832
rect 8484 31680 8536 31686
rect 8484 31622 8536 31628
rect 7656 31136 7708 31142
rect 7656 31078 7708 31084
rect 7668 30190 7696 31078
rect 8300 30660 8352 30666
rect 8300 30602 8352 30608
rect 8312 30326 8340 30602
rect 8300 30320 8352 30326
rect 8300 30262 8352 30268
rect 7656 30184 7708 30190
rect 7656 30126 7708 30132
rect 7472 29708 7524 29714
rect 7472 29650 7524 29656
rect 7288 29028 7340 29034
rect 7288 28970 7340 28976
rect 7300 28626 7328 28970
rect 7484 28626 7512 29650
rect 7668 29578 7696 30126
rect 8312 29646 8340 30262
rect 8576 30252 8628 30258
rect 8576 30194 8628 30200
rect 8588 29850 8616 30194
rect 8576 29844 8628 29850
rect 8576 29786 8628 29792
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 7656 29572 7708 29578
rect 7656 29514 7708 29520
rect 7668 29170 7696 29514
rect 7656 29164 7708 29170
rect 7656 29106 7708 29112
rect 7840 29164 7892 29170
rect 7840 29106 7892 29112
rect 7852 28762 7880 29106
rect 7840 28756 7892 28762
rect 7840 28698 7892 28704
rect 7104 28620 7156 28626
rect 7104 28562 7156 28568
rect 7288 28620 7340 28626
rect 7288 28562 7340 28568
rect 7472 28620 7524 28626
rect 7472 28562 7524 28568
rect 6920 28076 6972 28082
rect 6920 28018 6972 28024
rect 7380 27872 7432 27878
rect 7380 27814 7432 27820
rect 6460 27668 6512 27674
rect 6460 27610 6512 27616
rect 7012 27464 7064 27470
rect 7012 27406 7064 27412
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6840 26586 6868 26930
rect 6092 26580 6144 26586
rect 6092 26522 6144 26528
rect 6276 26580 6328 26586
rect 6276 26522 6328 26528
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6000 24880 6052 24886
rect 6000 24822 6052 24828
rect 6012 16574 6040 24822
rect 6104 23361 6132 26522
rect 6184 26376 6236 26382
rect 6184 26318 6236 26324
rect 6196 25770 6224 26318
rect 6288 26042 6316 26522
rect 6826 26344 6882 26353
rect 6826 26279 6828 26288
rect 6880 26279 6882 26288
rect 6828 26250 6880 26256
rect 6276 26036 6328 26042
rect 6276 25978 6328 25984
rect 6184 25764 6236 25770
rect 6184 25706 6236 25712
rect 6460 25764 6512 25770
rect 6460 25706 6512 25712
rect 6276 24268 6328 24274
rect 6276 24210 6328 24216
rect 6184 23656 6236 23662
rect 6182 23624 6184 23633
rect 6236 23624 6238 23633
rect 6182 23559 6238 23568
rect 6090 23352 6146 23361
rect 6146 23310 6224 23338
rect 6090 23287 6146 23296
rect 6196 22506 6224 23310
rect 6288 22982 6316 24210
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 6276 22160 6328 22166
rect 6276 22102 6328 22108
rect 6092 22024 6144 22030
rect 6092 21966 6144 21972
rect 6104 19922 6132 21966
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6196 20058 6224 20198
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6288 19990 6316 22102
rect 6472 22094 6500 25706
rect 6828 25696 6880 25702
rect 6828 25638 6880 25644
rect 6840 25294 6868 25638
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6552 25152 6604 25158
rect 6552 25094 6604 25100
rect 6564 24206 6592 25094
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6472 22066 6592 22094
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 6276 19984 6328 19990
rect 6276 19926 6328 19932
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6104 17678 6132 19858
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6288 16658 6316 19926
rect 6380 19854 6408 20742
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6380 19446 6408 19654
rect 6368 19440 6420 19446
rect 6368 19382 6420 19388
rect 6472 19378 6500 19654
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6564 17202 6592 22066
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6932 19922 6960 20538
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6656 19786 6684 19858
rect 6644 19780 6696 19786
rect 6644 19722 6696 19728
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6656 18426 6684 18634
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6932 18222 6960 18702
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6932 17610 6960 18158
rect 7024 17678 7052 27406
rect 7196 27328 7248 27334
rect 7196 27270 7248 27276
rect 7208 26382 7236 27270
rect 7196 26376 7248 26382
rect 7196 26318 7248 26324
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7116 22030 7144 22374
rect 7208 22098 7236 24686
rect 7300 24206 7328 25094
rect 7392 24818 7420 27814
rect 7484 27538 7512 28562
rect 8392 27872 8444 27878
rect 8392 27814 8444 27820
rect 7472 27532 7524 27538
rect 7472 27474 7524 27480
rect 8024 27532 8076 27538
rect 8024 27474 8076 27480
rect 7932 27328 7984 27334
rect 7932 27270 7984 27276
rect 7944 26858 7972 27270
rect 7932 26852 7984 26858
rect 7932 26794 7984 26800
rect 7944 26450 7972 26794
rect 7932 26444 7984 26450
rect 7932 26386 7984 26392
rect 8036 26382 8064 27474
rect 8208 27464 8260 27470
rect 8208 27406 8260 27412
rect 8220 27044 8248 27406
rect 8300 27396 8352 27402
rect 8300 27338 8352 27344
rect 8128 27016 8248 27044
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 7656 25900 7708 25906
rect 7656 25842 7708 25848
rect 7472 25832 7524 25838
rect 7472 25774 7524 25780
rect 7484 25362 7512 25774
rect 7472 25356 7524 25362
rect 7472 25298 7524 25304
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7484 24410 7512 25298
rect 7668 25294 7696 25842
rect 8036 25838 8064 26318
rect 8024 25832 8076 25838
rect 8024 25774 8076 25780
rect 8036 25362 8064 25774
rect 8024 25356 8076 25362
rect 8024 25298 8076 25304
rect 7656 25288 7708 25294
rect 7656 25230 7708 25236
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7288 24200 7340 24206
rect 7288 24142 7340 24148
rect 7380 24064 7432 24070
rect 7380 24006 7432 24012
rect 7196 22092 7248 22098
rect 7196 22034 7248 22040
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7208 21554 7236 22034
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 7208 21010 7236 21490
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 7208 20398 7236 20946
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7196 17740 7248 17746
rect 7196 17682 7248 17688
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6564 16574 6592 17138
rect 6656 16998 6684 17274
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6012 16546 6132 16574
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 6012 12306 6040 12718
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6104 5302 6132 16546
rect 6472 16546 6592 16574
rect 6748 16574 6776 17070
rect 6840 16726 6868 17206
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6932 16574 6960 17546
rect 7208 17542 7236 17682
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17218 7236 17478
rect 7300 17338 7328 18022
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7208 17190 7328 17218
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 6748 16546 6868 16574
rect 6932 16546 7052 16574
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6380 15094 6408 15846
rect 6368 15088 6420 15094
rect 6368 15030 6420 15036
rect 6472 12918 6500 16546
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6564 14618 6592 16050
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 6196 10130 6224 11018
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6196 9518 6224 10066
rect 6288 10062 6316 12854
rect 6564 12782 6592 13126
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6564 12306 6592 12582
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6472 11626 6500 12242
rect 6748 12102 6776 12786
rect 6840 12594 6868 16546
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6932 16046 6960 16186
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6932 14482 6960 15982
rect 7024 15026 7052 16546
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 7116 15638 7144 16118
rect 7208 16046 7236 16934
rect 7300 16250 7328 17190
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 7208 15434 7236 15846
rect 7196 15428 7248 15434
rect 7196 15370 7248 15376
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 7208 14414 7236 15370
rect 7392 15042 7420 24006
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 7840 22500 7892 22506
rect 7840 22442 7892 22448
rect 7472 21548 7524 21554
rect 7472 21490 7524 21496
rect 7484 21146 7512 21490
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7576 17882 7604 18226
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7484 16574 7512 17614
rect 7484 16546 7604 16574
rect 7392 15014 7512 15042
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 13258 6960 13670
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6840 12566 7052 12594
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6932 12306 6960 12378
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 7024 12238 7052 12566
rect 7116 12442 7144 13874
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7392 12306 7420 12718
rect 7484 12646 7512 15014
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11762 6776 12038
rect 7024 11830 7052 12174
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6748 11354 6776 11698
rect 7576 11558 7604 16546
rect 7668 12986 7696 20402
rect 7852 17134 7880 22442
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7944 17202 7972 17478
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7852 16998 7880 17070
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7760 15094 7788 15302
rect 7748 15088 7800 15094
rect 7748 15030 7800 15036
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7760 14346 7788 14758
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 8036 13802 8064 23462
rect 8128 20466 8156 27016
rect 8312 26314 8340 27338
rect 8404 27062 8432 27814
rect 8680 27606 8708 31826
rect 9048 29306 9076 39238
rect 10508 38956 10560 38962
rect 10508 38898 10560 38904
rect 9312 38752 9364 38758
rect 9312 38694 9364 38700
rect 9324 38350 9352 38694
rect 9312 38344 9364 38350
rect 9312 38286 9364 38292
rect 9220 38276 9272 38282
rect 9220 38218 9272 38224
rect 9232 37738 9260 38218
rect 10520 38010 10548 38898
rect 9588 38004 9640 38010
rect 9588 37946 9640 37952
rect 10508 38004 10560 38010
rect 10508 37946 10560 37952
rect 9600 37874 9628 37946
rect 9588 37868 9640 37874
rect 9588 37810 9640 37816
rect 9496 37800 9548 37806
rect 9496 37742 9548 37748
rect 9600 37754 9628 37810
rect 10324 37800 10376 37806
rect 9220 37732 9272 37738
rect 9220 37674 9272 37680
rect 9140 37454 9352 37482
rect 9140 35562 9168 37454
rect 9220 37392 9272 37398
rect 9220 37334 9272 37340
rect 9128 35556 9180 35562
rect 9128 35498 9180 35504
rect 9232 35154 9260 37334
rect 9324 37330 9352 37454
rect 9508 37398 9536 37742
rect 9600 37726 9996 37754
rect 10324 37742 10376 37748
rect 10508 37800 10560 37806
rect 10508 37742 10560 37748
rect 9586 37632 9642 37641
rect 9586 37567 9642 37576
rect 9496 37392 9548 37398
rect 9496 37334 9548 37340
rect 9600 37330 9628 37567
rect 9968 37330 9996 37726
rect 9312 37324 9364 37330
rect 9312 37266 9364 37272
rect 9588 37324 9640 37330
rect 9588 37266 9640 37272
rect 9956 37324 10008 37330
rect 9956 37266 10008 37272
rect 10140 37256 10192 37262
rect 10140 37198 10192 37204
rect 10152 36786 10180 37198
rect 10336 36922 10364 37742
rect 10520 37466 10548 37742
rect 10508 37460 10560 37466
rect 10508 37402 10560 37408
rect 10324 36916 10376 36922
rect 10324 36858 10376 36864
rect 10140 36780 10192 36786
rect 10140 36722 10192 36728
rect 9680 36236 9732 36242
rect 9680 36178 9732 36184
rect 9312 36100 9364 36106
rect 9312 36042 9364 36048
rect 9324 35766 9352 36042
rect 9588 36032 9640 36038
rect 9588 35974 9640 35980
rect 9312 35760 9364 35766
rect 9312 35702 9364 35708
rect 9220 35148 9272 35154
rect 9220 35090 9272 35096
rect 9324 34950 9352 35702
rect 9600 35698 9628 35974
rect 9588 35692 9640 35698
rect 9588 35634 9640 35640
rect 9692 35578 9720 36178
rect 9956 36168 10008 36174
rect 9956 36110 10008 36116
rect 9600 35562 9720 35578
rect 9588 35556 9720 35562
rect 9640 35550 9720 35556
rect 9588 35498 9640 35504
rect 9404 35080 9456 35086
rect 9404 35022 9456 35028
rect 9312 34944 9364 34950
rect 9312 34886 9364 34892
rect 9416 34746 9444 35022
rect 9496 35012 9548 35018
rect 9496 34954 9548 34960
rect 9508 34746 9536 34954
rect 9404 34740 9456 34746
rect 9404 34682 9456 34688
rect 9496 34740 9548 34746
rect 9496 34682 9548 34688
rect 9600 34626 9628 35498
rect 9968 35494 9996 36110
rect 10336 35834 10364 36858
rect 10520 36242 10548 37402
rect 10508 36236 10560 36242
rect 10508 36178 10560 36184
rect 10324 35828 10376 35834
rect 10324 35770 10376 35776
rect 9956 35488 10008 35494
rect 9956 35430 10008 35436
rect 9680 35012 9732 35018
rect 9680 34954 9732 34960
rect 9416 34598 9628 34626
rect 9692 34610 9720 34954
rect 9680 34604 9732 34610
rect 9416 34406 9444 34598
rect 9680 34546 9732 34552
rect 9404 34400 9456 34406
rect 9404 34342 9456 34348
rect 9416 33522 9444 34342
rect 9968 34202 9996 35430
rect 10324 35148 10376 35154
rect 10324 35090 10376 35096
rect 10140 34536 10192 34542
rect 10140 34478 10192 34484
rect 10232 34536 10284 34542
rect 10336 34524 10364 35090
rect 10416 34740 10468 34746
rect 10416 34682 10468 34688
rect 10428 34610 10456 34682
rect 10416 34604 10468 34610
rect 10416 34546 10468 34552
rect 10284 34496 10364 34524
rect 10232 34478 10284 34484
rect 9956 34196 10008 34202
rect 9956 34138 10008 34144
rect 9404 33516 9456 33522
rect 9404 33458 9456 33464
rect 9680 33448 9732 33454
rect 9680 33390 9732 33396
rect 9692 33114 9720 33390
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 9324 32910 9352 33050
rect 9312 32904 9364 32910
rect 9312 32846 9364 32852
rect 9680 32836 9732 32842
rect 9680 32778 9732 32784
rect 9128 32768 9180 32774
rect 9128 32710 9180 32716
rect 9140 32502 9168 32710
rect 9128 32496 9180 32502
rect 9128 32438 9180 32444
rect 9220 32292 9272 32298
rect 9220 32234 9272 32240
rect 9232 31890 9260 32234
rect 9588 31952 9640 31958
rect 9588 31894 9640 31900
rect 9220 31884 9272 31890
rect 9220 31826 9272 31832
rect 9312 30048 9364 30054
rect 9312 29990 9364 29996
rect 9324 29782 9352 29990
rect 9312 29776 9364 29782
rect 9312 29718 9364 29724
rect 9036 29300 9088 29306
rect 9036 29242 9088 29248
rect 9404 29232 9456 29238
rect 9404 29174 9456 29180
rect 9312 29164 9364 29170
rect 9312 29106 9364 29112
rect 9324 28966 9352 29106
rect 9416 28966 9444 29174
rect 9312 28960 9364 28966
rect 9312 28902 9364 28908
rect 9404 28960 9456 28966
rect 9404 28902 9456 28908
rect 9324 28422 9352 28902
rect 9416 28626 9444 28902
rect 9404 28620 9456 28626
rect 9404 28562 9456 28568
rect 9402 28520 9458 28529
rect 9402 28455 9404 28464
rect 9456 28455 9458 28464
rect 9404 28426 9456 28432
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 8668 27600 8720 27606
rect 8668 27542 8720 27548
rect 9128 27532 9180 27538
rect 9128 27474 9180 27480
rect 8392 27056 8444 27062
rect 8392 26998 8444 27004
rect 9140 26926 9168 27474
rect 9324 27402 9352 28358
rect 9312 27396 9364 27402
rect 9312 27338 9364 27344
rect 9128 26920 9180 26926
rect 9128 26862 9180 26868
rect 8576 26512 8628 26518
rect 9600 26489 9628 31894
rect 9692 31482 9720 32778
rect 9864 32768 9916 32774
rect 9864 32710 9916 32716
rect 9876 32434 9904 32710
rect 9864 32428 9916 32434
rect 9864 32370 9916 32376
rect 9772 31884 9824 31890
rect 9876 31872 9904 32370
rect 10152 32298 10180 34478
rect 10520 34202 10548 36178
rect 10324 34196 10376 34202
rect 10324 34138 10376 34144
rect 10508 34196 10560 34202
rect 10508 34138 10560 34144
rect 10232 33380 10284 33386
rect 10232 33322 10284 33328
rect 10140 32292 10192 32298
rect 10140 32234 10192 32240
rect 9956 32224 10008 32230
rect 9956 32166 10008 32172
rect 9968 31890 9996 32166
rect 9824 31844 9904 31872
rect 9772 31826 9824 31832
rect 9876 31482 9904 31844
rect 9956 31884 10008 31890
rect 9956 31826 10008 31832
rect 10140 31680 10192 31686
rect 10140 31622 10192 31628
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 10152 31278 10180 31622
rect 10140 31272 10192 31278
rect 10140 31214 10192 31220
rect 9772 31204 9824 31210
rect 9772 31146 9824 31152
rect 9680 26988 9732 26994
rect 9680 26930 9732 26936
rect 9692 26625 9720 26930
rect 9784 26790 9812 31146
rect 10152 30870 10180 31214
rect 10140 30864 10192 30870
rect 10140 30806 10192 30812
rect 10140 30592 10192 30598
rect 10140 30534 10192 30540
rect 9956 30252 10008 30258
rect 9956 30194 10008 30200
rect 9968 29238 9996 30194
rect 9956 29232 10008 29238
rect 9956 29174 10008 29180
rect 9968 29102 9996 29174
rect 9956 29096 10008 29102
rect 9956 29038 10008 29044
rect 9864 29028 9916 29034
rect 9864 28970 9916 28976
rect 9876 28626 9904 28970
rect 9864 28620 9916 28626
rect 9864 28562 9916 28568
rect 9968 27418 9996 29038
rect 10152 27538 10180 30534
rect 10244 29714 10272 33322
rect 10336 29714 10364 34138
rect 10416 33108 10468 33114
rect 10416 33050 10468 33056
rect 10428 31822 10456 33050
rect 10508 32564 10560 32570
rect 10508 32506 10560 32512
rect 10520 32434 10548 32506
rect 10508 32428 10560 32434
rect 10508 32370 10560 32376
rect 10520 31872 10548 32370
rect 10612 32314 10640 39986
rect 11348 39574 11376 39986
rect 11336 39568 11388 39574
rect 11336 39510 11388 39516
rect 10968 38548 11020 38554
rect 10968 38490 11020 38496
rect 10692 38276 10744 38282
rect 10692 38218 10744 38224
rect 10704 37398 10732 38218
rect 10876 38208 10928 38214
rect 10876 38150 10928 38156
rect 10888 38010 10916 38150
rect 10980 38010 11008 38490
rect 10876 38004 10928 38010
rect 10876 37946 10928 37952
rect 10968 38004 11020 38010
rect 10968 37946 11020 37952
rect 10876 37664 10928 37670
rect 10876 37606 10928 37612
rect 10692 37392 10744 37398
rect 10692 37334 10744 37340
rect 10692 35216 10744 35222
rect 10692 35158 10744 35164
rect 10704 34626 10732 35158
rect 10704 34598 10824 34626
rect 10692 34536 10744 34542
rect 10692 34478 10744 34484
rect 10704 32434 10732 34478
rect 10796 33969 10824 34598
rect 10888 34542 10916 37606
rect 10980 37126 11008 37946
rect 11244 37800 11296 37806
rect 11532 37754 11560 39986
rect 11900 37806 11928 40054
rect 12084 37806 12112 40684
rect 12164 40666 12216 40672
rect 12532 40724 12584 40730
rect 12532 40666 12584 40672
rect 12544 40526 12572 40666
rect 12532 40520 12584 40526
rect 12532 40462 12584 40468
rect 12440 40180 12492 40186
rect 12440 40122 12492 40128
rect 12452 39794 12480 40122
rect 12176 39766 12480 39794
rect 12176 39302 12204 39766
rect 12164 39296 12216 39302
rect 12164 39238 12216 39244
rect 11244 37742 11296 37748
rect 11060 37664 11112 37670
rect 11058 37632 11060 37641
rect 11112 37632 11114 37641
rect 11058 37567 11114 37576
rect 11256 37330 11284 37742
rect 11440 37738 11560 37754
rect 11888 37800 11940 37806
rect 11888 37742 11940 37748
rect 12072 37800 12124 37806
rect 12072 37742 12124 37748
rect 12176 37754 12204 39238
rect 12532 38208 12584 38214
rect 12532 38150 12584 38156
rect 12544 38010 12572 38150
rect 12532 38004 12584 38010
rect 12532 37946 12584 37952
rect 12440 37868 12492 37874
rect 12268 37828 12440 37856
rect 12268 37754 12296 37828
rect 12440 37810 12492 37816
rect 11428 37732 11560 37738
rect 11480 37726 11560 37732
rect 12176 37726 12296 37754
rect 11428 37674 11480 37680
rect 12176 37330 12204 37726
rect 12256 37664 12308 37670
rect 12256 37606 12308 37612
rect 12268 37330 12296 37606
rect 11244 37324 11296 37330
rect 11244 37266 11296 37272
rect 12164 37324 12216 37330
rect 12164 37266 12216 37272
rect 12256 37324 12308 37330
rect 12256 37266 12308 37272
rect 12440 37256 12492 37262
rect 12440 37198 12492 37204
rect 10968 37120 11020 37126
rect 10968 37062 11020 37068
rect 12452 36922 12480 37198
rect 12544 37126 12572 37946
rect 12532 37120 12584 37126
rect 12532 37062 12584 37068
rect 12440 36916 12492 36922
rect 12440 36858 12492 36864
rect 11060 36032 11112 36038
rect 11060 35974 11112 35980
rect 11072 35494 11100 35974
rect 12440 35624 12492 35630
rect 12440 35566 12492 35572
rect 11060 35488 11112 35494
rect 11060 35430 11112 35436
rect 10968 35080 11020 35086
rect 10968 35022 11020 35028
rect 10980 34746 11008 35022
rect 11072 34950 11100 35430
rect 12452 35086 12480 35566
rect 11244 35080 11296 35086
rect 11244 35022 11296 35028
rect 12440 35080 12492 35086
rect 12440 35022 12492 35028
rect 11060 34944 11112 34950
rect 11060 34886 11112 34892
rect 10968 34740 11020 34746
rect 10968 34682 11020 34688
rect 10876 34536 10928 34542
rect 10876 34478 10928 34484
rect 10876 34196 10928 34202
rect 10876 34138 10928 34144
rect 10782 33960 10838 33969
rect 10782 33895 10838 33904
rect 10692 32428 10744 32434
rect 10692 32370 10744 32376
rect 10612 32286 10824 32314
rect 10600 31884 10652 31890
rect 10520 31844 10600 31872
rect 10600 31826 10652 31832
rect 10416 31816 10468 31822
rect 10468 31764 10548 31770
rect 10416 31758 10548 31764
rect 10428 31726 10548 31758
rect 10232 29708 10284 29714
rect 10232 29650 10284 29656
rect 10324 29708 10376 29714
rect 10324 29650 10376 29656
rect 10140 27532 10192 27538
rect 10140 27474 10192 27480
rect 9876 27390 9996 27418
rect 9876 27062 9904 27390
rect 9956 27328 10008 27334
rect 9956 27270 10008 27276
rect 10048 27328 10100 27334
rect 10048 27270 10100 27276
rect 9864 27056 9916 27062
rect 9864 26998 9916 27004
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 9678 26616 9734 26625
rect 9876 26586 9904 26998
rect 9968 26994 9996 27270
rect 10060 27062 10088 27270
rect 10048 27056 10100 27062
rect 10048 26998 10100 27004
rect 9956 26988 10008 26994
rect 9956 26930 10008 26936
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 9678 26551 9734 26560
rect 9864 26580 9916 26586
rect 9864 26522 9916 26528
rect 8576 26454 8628 26460
rect 9586 26480 9642 26489
rect 8300 26308 8352 26314
rect 8300 26250 8352 26256
rect 8588 25906 8616 26454
rect 9586 26415 9642 26424
rect 10060 26382 10088 26726
rect 10048 26376 10100 26382
rect 10048 26318 10100 26324
rect 10428 26314 10456 31726
rect 10508 30184 10560 30190
rect 10508 30126 10560 30132
rect 10520 29646 10548 30126
rect 10692 30116 10744 30122
rect 10692 30058 10744 30064
rect 10704 29714 10732 30058
rect 10692 29708 10744 29714
rect 10692 29650 10744 29656
rect 10508 29640 10560 29646
rect 10508 29582 10560 29588
rect 10600 28416 10652 28422
rect 10600 28358 10652 28364
rect 10612 27538 10640 28358
rect 10600 27532 10652 27538
rect 10600 27474 10652 27480
rect 10796 27418 10824 32286
rect 10888 31793 10916 34138
rect 11256 34134 11284 35022
rect 11796 35012 11848 35018
rect 11796 34954 11848 34960
rect 11520 34944 11572 34950
rect 11520 34886 11572 34892
rect 11532 34542 11560 34886
rect 11808 34746 11836 34954
rect 11796 34740 11848 34746
rect 11796 34682 11848 34688
rect 12452 34542 12480 35022
rect 11520 34536 11572 34542
rect 11520 34478 11572 34484
rect 12440 34536 12492 34542
rect 12440 34478 12492 34484
rect 12624 34536 12676 34542
rect 12624 34478 12676 34484
rect 11244 34128 11296 34134
rect 11244 34070 11296 34076
rect 11428 34060 11480 34066
rect 11428 34002 11480 34008
rect 11152 32224 11204 32230
rect 11152 32166 11204 32172
rect 11336 32224 11388 32230
rect 11336 32166 11388 32172
rect 10874 31784 10930 31793
rect 10874 31719 10930 31728
rect 10888 31278 10916 31719
rect 10876 31272 10928 31278
rect 10876 31214 10928 31220
rect 10968 30796 11020 30802
rect 10968 30738 11020 30744
rect 10980 29102 11008 30738
rect 11060 29164 11112 29170
rect 11060 29106 11112 29112
rect 10968 29096 11020 29102
rect 10968 29038 11020 29044
rect 10980 28694 11008 29038
rect 11072 28762 11100 29106
rect 11060 28756 11112 28762
rect 11060 28698 11112 28704
rect 10968 28688 11020 28694
rect 10968 28630 11020 28636
rect 10876 28620 10928 28626
rect 10876 28562 10928 28568
rect 10888 28234 10916 28562
rect 11060 28416 11112 28422
rect 11058 28384 11060 28393
rect 11112 28384 11114 28393
rect 11058 28319 11114 28328
rect 10888 28206 11008 28234
rect 10980 28014 11008 28206
rect 10968 28008 11020 28014
rect 10968 27950 11020 27956
rect 10980 27674 11008 27950
rect 10968 27668 11020 27674
rect 10968 27610 11020 27616
rect 10796 27390 10916 27418
rect 10784 27328 10836 27334
rect 10784 27270 10836 27276
rect 10796 26994 10824 27270
rect 10784 26988 10836 26994
rect 10784 26930 10836 26936
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 10796 26382 10824 26726
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 10416 26308 10468 26314
rect 10416 26250 10468 26256
rect 10600 26240 10652 26246
rect 10600 26182 10652 26188
rect 9864 25968 9916 25974
rect 9864 25910 9916 25916
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9128 25832 9180 25838
rect 9128 25774 9180 25780
rect 8392 25696 8444 25702
rect 8392 25638 8444 25644
rect 8404 24886 8432 25638
rect 8944 25220 8996 25226
rect 8944 25162 8996 25168
rect 8392 24880 8444 24886
rect 8392 24822 8444 24828
rect 8956 24342 8984 25162
rect 9140 24818 9168 25774
rect 9416 25294 9444 25842
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9784 25362 9812 25774
rect 9876 25362 9904 25910
rect 10612 25906 10640 26182
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 9772 25356 9824 25362
rect 9772 25298 9824 25304
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 9404 25288 9456 25294
rect 9404 25230 9456 25236
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 8944 24336 8996 24342
rect 8944 24278 8996 24284
rect 8300 24064 8352 24070
rect 8300 24006 8352 24012
rect 8208 22568 8260 22574
rect 8208 22510 8260 22516
rect 8220 22234 8248 22510
rect 8208 22228 8260 22234
rect 8208 22170 8260 22176
rect 8312 20534 8340 24006
rect 8760 23520 8812 23526
rect 8760 23462 8812 23468
rect 8772 23118 8800 23462
rect 8956 23118 8984 24278
rect 9312 24132 9364 24138
rect 9312 24074 9364 24080
rect 9128 23724 9180 23730
rect 9128 23666 9180 23672
rect 8760 23112 8812 23118
rect 8760 23054 8812 23060
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 8404 22778 8616 22794
rect 8392 22772 8628 22778
rect 8444 22766 8576 22772
rect 8392 22714 8444 22720
rect 8576 22714 8628 22720
rect 9140 22642 9168 23666
rect 9324 23662 9352 24074
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9232 22778 9260 23598
rect 9220 22772 9272 22778
rect 9220 22714 9272 22720
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 9128 22636 9180 22642
rect 9128 22578 9180 22584
rect 8404 22234 8432 22578
rect 8484 22568 8536 22574
rect 8484 22510 8536 22516
rect 8392 22228 8444 22234
rect 8392 22170 8444 22176
rect 8496 20942 8524 22510
rect 8864 22166 8892 22578
rect 8852 22160 8904 22166
rect 8852 22102 8904 22108
rect 8864 21690 8892 22102
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 8484 20936 8536 20942
rect 8484 20878 8536 20884
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 9220 20324 9272 20330
rect 9220 20266 9272 20272
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8312 19514 8340 20198
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8220 18290 8248 18702
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8312 17338 8340 18362
rect 8404 17678 8432 18566
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 7748 13796 7800 13802
rect 7748 13738 7800 13744
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7668 11694 7696 12922
rect 7760 12782 7788 13738
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7852 12238 7880 13126
rect 8208 12640 8260 12646
rect 8206 12608 8208 12617
rect 8260 12608 8262 12617
rect 8206 12543 8262 12552
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 7576 11218 7604 11494
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7576 10606 7604 11154
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6380 9654 6408 10406
rect 7208 10130 7236 10542
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 7668 9518 7696 10542
rect 7760 9722 7788 10746
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7852 9586 7880 10542
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 6196 9178 6224 9454
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7300 7886 7328 8298
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7342 7420 7822
rect 7668 7546 7696 9454
rect 7852 8634 7880 9522
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 8036 8566 8064 12242
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11898 8248 12038
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8312 11626 8340 16526
rect 8496 12306 8524 19790
rect 8576 18692 8628 18698
rect 8576 18634 8628 18640
rect 8588 17882 8616 18634
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8588 15706 8616 17682
rect 8772 17678 8800 17818
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 9232 16590 9260 20266
rect 9324 20262 9352 23598
rect 9402 23488 9458 23497
rect 9402 23423 9458 23432
rect 9416 23050 9444 23423
rect 9692 23118 9720 24754
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 9404 23044 9456 23050
rect 9404 22986 9456 22992
rect 9416 22710 9444 22986
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 9404 22704 9456 22710
rect 9404 22646 9456 22652
rect 9508 22642 9536 22918
rect 9496 22636 9548 22642
rect 9496 22578 9548 22584
rect 9508 22098 9536 22578
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 9496 22092 9548 22098
rect 9496 22034 9548 22040
rect 9692 22030 9720 22510
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9324 19258 9352 20198
rect 9416 19378 9444 20198
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9324 19230 9536 19258
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9416 16658 9444 18158
rect 9508 17746 9536 19230
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9692 18154 9720 18294
rect 9784 18222 9812 25298
rect 10600 24608 10652 24614
rect 10600 24550 10652 24556
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 10508 22568 10560 22574
rect 10508 22510 10560 22516
rect 10428 22098 10456 22510
rect 10520 22234 10548 22510
rect 10508 22228 10560 22234
rect 10508 22170 10560 22176
rect 10520 22098 10548 22170
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10416 22092 10468 22098
rect 10416 22034 10468 22040
rect 10508 22092 10560 22098
rect 10508 22034 10560 22040
rect 10152 22001 10180 22034
rect 10138 21992 10194 22001
rect 10060 21950 10138 21978
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9876 19718 9904 20402
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8588 15570 8616 15642
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8772 15502 8800 15982
rect 8956 15706 8984 15982
rect 9232 15978 9260 16526
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 9508 15570 9536 16186
rect 9968 16114 9996 20198
rect 10060 16250 10088 21950
rect 10138 21927 10194 21936
rect 10506 21720 10562 21729
rect 10506 21655 10562 21664
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10152 20942 10180 21286
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10428 19990 10456 21354
rect 10520 20346 10548 21655
rect 10612 20942 10640 24550
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 10796 22234 10824 22714
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10692 22024 10744 22030
rect 10690 21992 10692 22001
rect 10744 21992 10746 22001
rect 10690 21927 10746 21936
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10704 21554 10732 21830
rect 10796 21690 10824 22170
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10704 21146 10732 21490
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10520 20318 10640 20346
rect 10508 20256 10560 20262
rect 10508 20198 10560 20204
rect 10416 19984 10468 19990
rect 10520 19961 10548 20198
rect 10416 19926 10468 19932
rect 10506 19952 10562 19961
rect 10324 18896 10376 18902
rect 10324 18838 10376 18844
rect 10336 18766 10364 18838
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10336 17678 10364 18702
rect 10428 18358 10456 19926
rect 10506 19887 10562 19896
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10520 19514 10548 19654
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10416 18352 10468 18358
rect 10416 18294 10468 18300
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 9956 16108 10008 16114
rect 10008 16068 10088 16096
rect 9956 16050 10008 16056
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9692 15570 9720 15982
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8956 15162 8984 15438
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 9508 14634 9536 15506
rect 9784 15450 9812 15982
rect 9956 15496 10008 15502
rect 9600 15444 9956 15450
rect 9600 15438 10008 15444
rect 9600 15422 9996 15438
rect 9600 14822 9628 15422
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9508 14606 9628 14634
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 8944 13388 8996 13394
rect 8944 13330 8996 13336
rect 8956 12850 8984 13330
rect 9324 12918 9352 13670
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8312 10606 8340 11562
rect 8864 11082 8892 11766
rect 8956 11762 8984 12786
rect 8944 11756 8996 11762
rect 9312 11756 9364 11762
rect 8996 11716 9076 11744
rect 8944 11698 8996 11704
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8680 10674 8708 10746
rect 8864 10674 8892 11018
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 8496 8498 8524 10202
rect 8588 9994 8616 10542
rect 8576 9988 8628 9994
rect 8576 9930 8628 9936
rect 8680 9518 8708 10610
rect 9048 10606 9076 11716
rect 9312 11698 9364 11704
rect 9324 11354 9352 11698
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 9508 10266 9536 10610
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 8864 9586 8892 9930
rect 9600 9926 9628 14606
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9692 12442 9720 13874
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 10198 9720 10950
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 9600 9382 9628 9862
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9692 9110 9720 9998
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9784 9178 9812 9318
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7760 7478 7788 8230
rect 8312 8090 8340 8434
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8496 7954 8524 8434
rect 8772 8022 8800 8570
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 9416 7954 9444 8570
rect 9876 7954 9904 12922
rect 10060 11082 10088 16068
rect 10152 15706 10180 16390
rect 10324 15904 10376 15910
rect 10244 15852 10324 15858
rect 10244 15846 10376 15852
rect 10244 15830 10364 15846
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10152 15094 10180 15642
rect 10244 15366 10272 15830
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10244 15094 10272 15302
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10428 14958 10456 18294
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10520 15450 10548 15506
rect 10612 15450 10640 20318
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10704 18086 10732 18702
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10704 17746 10732 18022
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 10704 16250 10732 16458
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10520 15422 10640 15450
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10244 14006 10272 14554
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10244 13410 10272 13942
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10152 13382 10272 13410
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10152 10962 10180 13382
rect 10336 13326 10364 13670
rect 10324 13320 10376 13326
rect 10060 10934 10180 10962
rect 10244 13280 10324 13308
rect 10060 9654 10088 10934
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10152 9382 10180 9930
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10152 9042 10180 9318
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10244 7954 10272 13280
rect 10324 13262 10376 13268
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12986 10456 13262
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10336 12238 10364 12582
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10428 10266 10456 12242
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10520 11150 10548 11494
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10428 9042 10456 10202
rect 10612 9518 10640 15422
rect 10704 15162 10732 16050
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12986 10732 13126
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10810 10824 10950
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7546 9352 7686
rect 9876 7546 9904 7890
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 9968 7342 9996 7890
rect 10520 7886 10548 8230
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9968 7206 9996 7278
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9968 6914 9996 7142
rect 10244 7002 10272 7346
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10888 6914 10916 27390
rect 10968 26852 11020 26858
rect 10968 26794 11020 26800
rect 10980 25702 11008 26794
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 10980 23730 11008 25638
rect 10968 23724 11020 23730
rect 10968 23666 11020 23672
rect 11164 23361 11192 32166
rect 11348 31890 11376 32166
rect 11336 31884 11388 31890
rect 11336 31826 11388 31832
rect 11336 28960 11388 28966
rect 11336 28902 11388 28908
rect 11348 28626 11376 28902
rect 11336 28620 11388 28626
rect 11336 28562 11388 28568
rect 11348 27946 11376 28562
rect 11336 27940 11388 27946
rect 11336 27882 11388 27888
rect 11348 27402 11376 27882
rect 11336 27396 11388 27402
rect 11336 27338 11388 27344
rect 11150 23352 11206 23361
rect 11150 23287 11206 23296
rect 11164 22778 11192 23287
rect 11152 22772 11204 22778
rect 11152 22714 11204 22720
rect 11440 22094 11468 34002
rect 11532 31754 11560 34478
rect 12164 33312 12216 33318
rect 12164 33254 12216 33260
rect 12176 32910 12204 33254
rect 12164 32904 12216 32910
rect 12164 32846 12216 32852
rect 11796 32836 11848 32842
rect 11796 32778 11848 32784
rect 11612 32428 11664 32434
rect 11612 32370 11664 32376
rect 11520 31748 11572 31754
rect 11520 31690 11572 31696
rect 11532 31482 11560 31690
rect 11624 31686 11652 32370
rect 11808 32366 11836 32778
rect 12072 32564 12124 32570
rect 12072 32506 12124 32512
rect 12084 32434 12112 32506
rect 12072 32428 12124 32434
rect 12072 32370 12124 32376
rect 11796 32360 11848 32366
rect 11796 32302 11848 32308
rect 11796 32224 11848 32230
rect 11796 32166 11848 32172
rect 11808 31754 11836 32166
rect 11716 31726 11836 31754
rect 11612 31680 11664 31686
rect 11612 31622 11664 31628
rect 11520 31476 11572 31482
rect 11520 31418 11572 31424
rect 11532 24750 11560 31418
rect 11612 30048 11664 30054
rect 11612 29990 11664 29996
rect 11624 29646 11652 29990
rect 11612 29640 11664 29646
rect 11612 29582 11664 29588
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11532 23866 11560 24686
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11348 22066 11468 22094
rect 11348 21978 11376 22066
rect 11716 21978 11744 31726
rect 12164 31204 12216 31210
rect 12164 31146 12216 31152
rect 11980 30252 12032 30258
rect 11980 30194 12032 30200
rect 11992 28218 12020 30194
rect 11980 28212 12032 28218
rect 11980 28154 12032 28160
rect 11980 27532 12032 27538
rect 11980 27474 12032 27480
rect 11796 27328 11848 27334
rect 11796 27270 11848 27276
rect 11808 27130 11836 27270
rect 11992 27130 12020 27474
rect 11796 27124 11848 27130
rect 11796 27066 11848 27072
rect 11980 27124 12032 27130
rect 11980 27066 12032 27072
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11808 25838 11836 26862
rect 11796 25832 11848 25838
rect 11796 25774 11848 25780
rect 12176 25294 12204 31146
rect 12256 26988 12308 26994
rect 12256 26930 12308 26936
rect 12268 26858 12296 26930
rect 12348 26920 12400 26926
rect 12348 26862 12400 26868
rect 12256 26852 12308 26858
rect 12256 26794 12308 26800
rect 12360 26450 12388 26862
rect 12348 26444 12400 26450
rect 12348 26386 12400 26392
rect 12256 26240 12308 26246
rect 12254 26208 12256 26217
rect 12308 26208 12310 26217
rect 12254 26143 12310 26152
rect 12164 25288 12216 25294
rect 12164 25230 12216 25236
rect 12072 25152 12124 25158
rect 12072 25094 12124 25100
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11900 22642 11928 22986
rect 11888 22636 11940 22642
rect 11888 22578 11940 22584
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11794 21992 11850 22001
rect 11348 21950 11468 21978
rect 11716 21950 11794 21978
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 11348 21690 11376 21830
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11440 21010 11468 21950
rect 11900 21962 11928 22578
rect 11992 22098 12020 22578
rect 11980 22092 12032 22098
rect 11980 22034 12032 22040
rect 11794 21927 11850 21936
rect 11888 21956 11940 21962
rect 11808 21894 11836 21927
rect 11888 21898 11940 21904
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 11900 21078 11928 21898
rect 11888 21072 11940 21078
rect 11888 21014 11940 21020
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11900 20942 11928 21014
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 10980 17746 11008 20810
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 11164 18902 11192 20402
rect 11900 20398 11928 20878
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11428 19372 11480 19378
rect 11624 19360 11652 19790
rect 11992 19786 12020 22034
rect 12084 20602 12112 25094
rect 12452 24818 12480 34478
rect 12636 32842 12664 34478
rect 12624 32836 12676 32842
rect 12624 32778 12676 32784
rect 12636 32570 12664 32778
rect 12624 32564 12676 32570
rect 12624 32506 12676 32512
rect 12532 32224 12584 32230
rect 12532 32166 12584 32172
rect 12544 32026 12572 32166
rect 12532 32020 12584 32026
rect 12532 31962 12584 31968
rect 12532 31884 12584 31890
rect 12532 31826 12584 31832
rect 12544 31249 12572 31826
rect 12530 31240 12586 31249
rect 12530 31175 12586 31184
rect 12728 30122 12756 42162
rect 13556 41818 13584 42162
rect 13740 42158 13768 42706
rect 15120 42634 15148 43250
rect 15212 42770 15240 43386
rect 15488 42906 15516 43726
rect 16592 43654 16620 44882
rect 16868 44878 16896 44950
rect 17328 44946 17356 45358
rect 17316 44940 17368 44946
rect 17316 44882 17368 44888
rect 16856 44872 16908 44878
rect 16856 44814 16908 44820
rect 17040 44192 17092 44198
rect 17040 44134 17092 44140
rect 16764 43784 16816 43790
rect 16764 43726 16816 43732
rect 16948 43784 17000 43790
rect 17052 43772 17080 44134
rect 17000 43744 17080 43772
rect 16948 43726 17000 43732
rect 16028 43648 16080 43654
rect 16028 43590 16080 43596
rect 16580 43648 16632 43654
rect 16580 43590 16632 43596
rect 15476 42900 15528 42906
rect 15476 42842 15528 42848
rect 15200 42764 15252 42770
rect 15200 42706 15252 42712
rect 15108 42628 15160 42634
rect 15108 42570 15160 42576
rect 15844 42560 15896 42566
rect 15844 42502 15896 42508
rect 15856 42362 15884 42502
rect 15844 42356 15896 42362
rect 15844 42298 15896 42304
rect 13728 42152 13780 42158
rect 13728 42094 13780 42100
rect 13544 41812 13596 41818
rect 13544 41754 13596 41760
rect 12900 41608 12952 41614
rect 12900 41550 12952 41556
rect 12808 32020 12860 32026
rect 12808 31962 12860 31968
rect 12820 31822 12848 31962
rect 12808 31816 12860 31822
rect 12808 31758 12860 31764
rect 12716 30116 12768 30122
rect 12716 30058 12768 30064
rect 12624 29504 12676 29510
rect 12624 29446 12676 29452
rect 12636 28626 12664 29446
rect 12716 28960 12768 28966
rect 12716 28902 12768 28908
rect 12624 28620 12676 28626
rect 12624 28562 12676 28568
rect 12636 28082 12664 28562
rect 12728 28218 12756 28902
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12636 27606 12664 28018
rect 12716 27872 12768 27878
rect 12716 27814 12768 27820
rect 12624 27600 12676 27606
rect 12624 27542 12676 27548
rect 12532 27328 12584 27334
rect 12532 27270 12584 27276
rect 12544 27062 12572 27270
rect 12728 27062 12756 27814
rect 12532 27056 12584 27062
rect 12716 27056 12768 27062
rect 12584 27016 12664 27044
rect 12532 26998 12584 27004
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12544 26042 12572 26318
rect 12532 26036 12584 26042
rect 12532 25978 12584 25984
rect 12636 25838 12664 27016
rect 12716 26998 12768 27004
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12728 26217 12756 26318
rect 12714 26208 12770 26217
rect 12820 26194 12848 31758
rect 12912 30938 12940 41550
rect 15856 41414 15884 42298
rect 15764 41386 15884 41414
rect 13636 41132 13688 41138
rect 13636 41074 13688 41080
rect 14464 41132 14516 41138
rect 14464 41074 14516 41080
rect 13268 41064 13320 41070
rect 13268 41006 13320 41012
rect 13176 40520 13228 40526
rect 13176 40462 13228 40468
rect 13188 40186 13216 40462
rect 13176 40180 13228 40186
rect 13176 40122 13228 40128
rect 13084 39636 13136 39642
rect 13084 39578 13136 39584
rect 13096 39506 13124 39578
rect 13084 39500 13136 39506
rect 13084 39442 13136 39448
rect 13176 39432 13228 39438
rect 13176 39374 13228 39380
rect 13084 37800 13136 37806
rect 13004 37760 13084 37788
rect 13004 36786 13032 37760
rect 13084 37742 13136 37748
rect 13084 37324 13136 37330
rect 13084 37266 13136 37272
rect 12992 36780 13044 36786
rect 12992 36722 13044 36728
rect 13096 35834 13124 37266
rect 13084 35828 13136 35834
rect 13084 35770 13136 35776
rect 13084 35488 13136 35494
rect 13084 35430 13136 35436
rect 13096 35154 13124 35430
rect 13084 35148 13136 35154
rect 13084 35090 13136 35096
rect 13188 33844 13216 39374
rect 13096 33816 13216 33844
rect 12992 33516 13044 33522
rect 12992 33458 13044 33464
rect 13004 33114 13032 33458
rect 13096 33454 13124 33816
rect 13176 33584 13228 33590
rect 13176 33526 13228 33532
rect 13084 33448 13136 33454
rect 13084 33390 13136 33396
rect 12992 33108 13044 33114
rect 12992 33050 13044 33056
rect 13188 31890 13216 33526
rect 13280 31890 13308 41006
rect 13544 40384 13596 40390
rect 13544 40326 13596 40332
rect 13556 40186 13584 40326
rect 13544 40180 13596 40186
rect 13544 40122 13596 40128
rect 13648 39982 13676 41074
rect 14004 41064 14056 41070
rect 14004 41006 14056 41012
rect 14016 40730 14044 41006
rect 14004 40724 14056 40730
rect 14004 40666 14056 40672
rect 14016 40594 14044 40666
rect 14004 40588 14056 40594
rect 14004 40530 14056 40536
rect 13636 39976 13688 39982
rect 13636 39918 13688 39924
rect 13648 39302 13676 39918
rect 14016 39438 14044 40530
rect 14476 40186 14504 41074
rect 15384 40928 15436 40934
rect 15384 40870 15436 40876
rect 15108 40520 15160 40526
rect 15108 40462 15160 40468
rect 14464 40180 14516 40186
rect 14464 40122 14516 40128
rect 15016 39908 15068 39914
rect 15016 39850 15068 39856
rect 14004 39432 14056 39438
rect 14004 39374 14056 39380
rect 13636 39296 13688 39302
rect 13636 39238 13688 39244
rect 14016 38418 14044 39374
rect 14740 39364 14792 39370
rect 14740 39306 14792 39312
rect 14752 38758 14780 39306
rect 14096 38752 14148 38758
rect 14096 38694 14148 38700
rect 14740 38752 14792 38758
rect 14740 38694 14792 38700
rect 14004 38412 14056 38418
rect 14004 38354 14056 38360
rect 13360 38344 13412 38350
rect 13360 38286 13412 38292
rect 13636 38344 13688 38350
rect 13636 38286 13688 38292
rect 13912 38344 13964 38350
rect 13912 38286 13964 38292
rect 13372 37466 13400 38286
rect 13648 38010 13676 38286
rect 13820 38208 13872 38214
rect 13820 38150 13872 38156
rect 13636 38004 13688 38010
rect 13636 37946 13688 37952
rect 13832 37874 13860 38150
rect 13820 37868 13872 37874
rect 13820 37810 13872 37816
rect 13924 37466 13952 38286
rect 14016 37942 14044 38354
rect 14004 37936 14056 37942
rect 14004 37878 14056 37884
rect 13360 37460 13412 37466
rect 13360 37402 13412 37408
rect 13912 37460 13964 37466
rect 13912 37402 13964 37408
rect 14108 37126 14136 38694
rect 14740 37800 14792 37806
rect 14740 37742 14792 37748
rect 14752 37126 14780 37742
rect 14924 37664 14976 37670
rect 14924 37606 14976 37612
rect 14832 37460 14884 37466
rect 14832 37402 14884 37408
rect 14096 37120 14148 37126
rect 14096 37062 14148 37068
rect 14280 37120 14332 37126
rect 14280 37062 14332 37068
rect 14740 37120 14792 37126
rect 14740 37062 14792 37068
rect 13728 36168 13780 36174
rect 13728 36110 13780 36116
rect 13740 35290 13768 36110
rect 14108 36106 14136 37062
rect 14096 36100 14148 36106
rect 14096 36042 14148 36048
rect 14292 36038 14320 37062
rect 14464 36848 14516 36854
rect 14462 36816 14464 36825
rect 14516 36816 14518 36825
rect 14462 36751 14518 36760
rect 14280 36032 14332 36038
rect 14280 35974 14332 35980
rect 13820 35760 13872 35766
rect 13820 35702 13872 35708
rect 13728 35284 13780 35290
rect 13728 35226 13780 35232
rect 13636 35080 13688 35086
rect 13636 35022 13688 35028
rect 13360 34604 13412 34610
rect 13360 34546 13412 34552
rect 13372 34202 13400 34546
rect 13360 34196 13412 34202
rect 13360 34138 13412 34144
rect 13360 32564 13412 32570
rect 13360 32506 13412 32512
rect 13176 31884 13228 31890
rect 13176 31826 13228 31832
rect 13268 31884 13320 31890
rect 13268 31826 13320 31832
rect 12900 30932 12952 30938
rect 12900 30874 12952 30880
rect 13176 30048 13228 30054
rect 13176 29990 13228 29996
rect 13084 29164 13136 29170
rect 13084 29106 13136 29112
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 12912 28150 12940 28494
rect 12900 28144 12952 28150
rect 12900 28086 12952 28092
rect 12900 27396 12952 27402
rect 12900 27338 12952 27344
rect 12912 27130 12940 27338
rect 12900 27124 12952 27130
rect 12900 27066 12952 27072
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 12912 26314 12940 26862
rect 12992 26580 13044 26586
rect 12992 26522 13044 26528
rect 12900 26308 12952 26314
rect 12900 26250 12952 26256
rect 12820 26166 12940 26194
rect 12714 26143 12770 26152
rect 12624 25832 12676 25838
rect 12624 25774 12676 25780
rect 12728 25650 12756 26143
rect 12728 25622 12848 25650
rect 12714 25528 12770 25537
rect 12714 25463 12770 25472
rect 12728 25430 12756 25463
rect 12716 25424 12768 25430
rect 12716 25366 12768 25372
rect 12820 25362 12848 25622
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12452 23730 12480 24754
rect 12164 23724 12216 23730
rect 12164 23666 12216 23672
rect 12440 23724 12492 23730
rect 12440 23666 12492 23672
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11980 19780 12032 19786
rect 11980 19722 12032 19728
rect 11716 19514 11744 19722
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11480 19332 11652 19360
rect 11428 19314 11480 19320
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11244 18828 11296 18834
rect 11244 18770 11296 18776
rect 11256 18426 11284 18770
rect 11520 18760 11572 18766
rect 11348 18708 11520 18714
rect 11348 18702 11572 18708
rect 11348 18686 11560 18702
rect 11348 18630 11376 18686
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11058 17912 11114 17921
rect 11058 17847 11114 17856
rect 11072 17814 11100 17847
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 11256 17678 11284 18362
rect 11348 17678 11376 18566
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11520 17672 11572 17678
rect 11624 17660 11652 19332
rect 11704 19236 11756 19242
rect 11704 19178 11756 19184
rect 11716 18834 11744 19178
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11572 17632 11652 17660
rect 11520 17614 11572 17620
rect 11992 17542 12020 18158
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 16182 11100 16934
rect 12084 16454 12112 20538
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 12070 16144 12126 16153
rect 12070 16079 12126 16088
rect 12084 16046 12112 16079
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12084 15570 12112 15982
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12176 14414 12204 23666
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10980 12102 11008 12854
rect 11072 12374 11100 13874
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11716 12986 11744 13262
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11900 12850 11928 13126
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 11624 12306 11652 12786
rect 11900 12306 11928 12786
rect 12268 12374 12296 20946
rect 12544 20942 12572 22578
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12636 20398 12664 25230
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 12820 22642 12848 24074
rect 12912 23866 12940 26166
rect 13004 25838 13032 26522
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 13096 25498 13124 29106
rect 13188 29034 13216 29990
rect 13280 29345 13308 31826
rect 13372 31822 13400 32506
rect 13648 32026 13676 35022
rect 13832 34950 13860 35702
rect 14740 35624 14792 35630
rect 14740 35566 14792 35572
rect 14372 35488 14424 35494
rect 14372 35430 14424 35436
rect 14384 35086 14412 35430
rect 14752 35154 14780 35566
rect 14740 35148 14792 35154
rect 14740 35090 14792 35096
rect 14372 35080 14424 35086
rect 14094 35048 14150 35057
rect 14372 35022 14424 35028
rect 14094 34983 14096 34992
rect 14148 34983 14150 34992
rect 14096 34954 14148 34960
rect 13820 34944 13872 34950
rect 13820 34886 13872 34892
rect 13832 33658 13860 34886
rect 14188 34740 14240 34746
rect 14188 34682 14240 34688
rect 14096 34536 14148 34542
rect 14016 34484 14096 34490
rect 14016 34478 14148 34484
rect 14016 34462 14136 34478
rect 13820 33652 13872 33658
rect 13820 33594 13872 33600
rect 13912 32972 13964 32978
rect 13912 32914 13964 32920
rect 13924 32774 13952 32914
rect 13912 32768 13964 32774
rect 13912 32710 13964 32716
rect 14016 32502 14044 34462
rect 14200 32978 14228 34682
rect 14556 34400 14608 34406
rect 14556 34342 14608 34348
rect 14568 33998 14596 34342
rect 14556 33992 14608 33998
rect 14556 33934 14608 33940
rect 14844 33318 14872 37402
rect 14936 37262 14964 37606
rect 14924 37256 14976 37262
rect 14924 37198 14976 37204
rect 15028 35442 15056 39850
rect 15120 38962 15148 40462
rect 15396 40390 15424 40870
rect 15476 40452 15528 40458
rect 15476 40394 15528 40400
rect 15200 40384 15252 40390
rect 15200 40326 15252 40332
rect 15384 40384 15436 40390
rect 15384 40326 15436 40332
rect 15212 40118 15240 40326
rect 15200 40112 15252 40118
rect 15200 40054 15252 40060
rect 15108 38956 15160 38962
rect 15108 38898 15160 38904
rect 15292 37188 15344 37194
rect 15292 37130 15344 37136
rect 15200 36236 15252 36242
rect 15200 36178 15252 36184
rect 15212 35630 15240 36178
rect 15304 35714 15332 37130
rect 15396 36802 15424 40326
rect 15488 39914 15516 40394
rect 15476 39908 15528 39914
rect 15476 39850 15528 39856
rect 15488 39302 15516 39850
rect 15476 39296 15528 39302
rect 15476 39238 15528 39244
rect 15476 38208 15528 38214
rect 15476 38150 15528 38156
rect 15488 38010 15516 38150
rect 15476 38004 15528 38010
rect 15476 37946 15528 37952
rect 15488 36938 15516 37946
rect 15660 37256 15712 37262
rect 15660 37198 15712 37204
rect 15488 36910 15608 36938
rect 15396 36774 15516 36802
rect 15488 36174 15516 36774
rect 15476 36168 15528 36174
rect 15476 36110 15528 36116
rect 15488 35834 15516 36110
rect 15580 35834 15608 36910
rect 15672 36650 15700 37198
rect 15660 36644 15712 36650
rect 15660 36586 15712 36592
rect 15476 35828 15528 35834
rect 15476 35770 15528 35776
rect 15568 35828 15620 35834
rect 15568 35770 15620 35776
rect 15304 35686 15516 35714
rect 15580 35698 15608 35770
rect 15672 35698 15700 36586
rect 15200 35624 15252 35630
rect 15200 35566 15252 35572
rect 15292 35556 15344 35562
rect 15292 35498 15344 35504
rect 15304 35465 15332 35498
rect 15290 35456 15346 35465
rect 15028 35414 15148 35442
rect 15016 34604 15068 34610
rect 15016 34546 15068 34552
rect 15028 33862 15056 34546
rect 15120 34542 15148 35414
rect 15290 35391 15346 35400
rect 15108 34536 15160 34542
rect 15108 34478 15160 34484
rect 15120 33930 15148 34478
rect 15304 34066 15332 35391
rect 15292 34060 15344 34066
rect 15292 34002 15344 34008
rect 15108 33924 15160 33930
rect 15108 33866 15160 33872
rect 15016 33856 15068 33862
rect 15016 33798 15068 33804
rect 15028 33590 15056 33798
rect 15016 33584 15068 33590
rect 15016 33526 15068 33532
rect 14832 33312 14884 33318
rect 14832 33254 14884 33260
rect 14280 33108 14332 33114
rect 14280 33050 14332 33056
rect 14188 32972 14240 32978
rect 14188 32914 14240 32920
rect 14096 32904 14148 32910
rect 14096 32846 14148 32852
rect 14004 32496 14056 32502
rect 13924 32456 14004 32484
rect 13820 32428 13872 32434
rect 13820 32370 13872 32376
rect 13636 32020 13688 32026
rect 13636 31962 13688 31968
rect 13360 31816 13412 31822
rect 13360 31758 13412 31764
rect 13832 31482 13860 32370
rect 13924 32026 13952 32456
rect 14004 32438 14056 32444
rect 14108 32366 14136 32846
rect 14200 32366 14228 32914
rect 14292 32842 14320 33050
rect 14648 33040 14700 33046
rect 14648 32982 14700 32988
rect 14280 32836 14332 32842
rect 14280 32778 14332 32784
rect 14660 32366 14688 32982
rect 14832 32972 14884 32978
rect 14832 32914 14884 32920
rect 14096 32360 14148 32366
rect 14096 32302 14148 32308
rect 14188 32360 14240 32366
rect 14188 32302 14240 32308
rect 14648 32360 14700 32366
rect 14648 32302 14700 32308
rect 14108 32212 14136 32302
rect 14280 32224 14332 32230
rect 14108 32184 14228 32212
rect 14200 32026 14228 32184
rect 14280 32166 14332 32172
rect 13912 32020 13964 32026
rect 13912 31962 13964 31968
rect 14188 32020 14240 32026
rect 14188 31962 14240 31968
rect 14004 31952 14056 31958
rect 14004 31894 14056 31900
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 13360 30932 13412 30938
rect 13360 30874 13412 30880
rect 13372 30666 13400 30874
rect 13636 30796 13688 30802
rect 13636 30738 13688 30744
rect 13360 30660 13412 30666
rect 13360 30602 13412 30608
rect 13544 30592 13596 30598
rect 13544 30534 13596 30540
rect 13556 30433 13584 30534
rect 13542 30424 13598 30433
rect 13542 30359 13598 30368
rect 13648 30054 13676 30738
rect 13728 30184 13780 30190
rect 13728 30126 13780 30132
rect 13636 30048 13688 30054
rect 13636 29990 13688 29996
rect 13266 29336 13322 29345
rect 13266 29271 13322 29280
rect 13176 29028 13228 29034
rect 13176 28970 13228 28976
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 13096 24342 13124 25434
rect 13084 24336 13136 24342
rect 13084 24278 13136 24284
rect 13188 24274 13216 28970
rect 13636 28552 13688 28558
rect 13636 28494 13688 28500
rect 13452 28416 13504 28422
rect 13452 28358 13504 28364
rect 13268 27464 13320 27470
rect 13268 27406 13320 27412
rect 13280 27334 13308 27406
rect 13268 27328 13320 27334
rect 13268 27270 13320 27276
rect 13280 26246 13308 27270
rect 13464 27130 13492 28358
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 13464 26994 13492 27066
rect 13648 26994 13676 28494
rect 13452 26988 13504 26994
rect 13372 26948 13452 26976
rect 13268 26240 13320 26246
rect 13268 26182 13320 26188
rect 13268 25968 13320 25974
rect 13268 25910 13320 25916
rect 13280 24954 13308 25910
rect 13372 25684 13400 26948
rect 13636 26988 13688 26994
rect 13452 26930 13504 26936
rect 13556 26948 13636 26976
rect 13556 26382 13584 26948
rect 13636 26930 13688 26936
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13544 26376 13596 26382
rect 13544 26318 13596 26324
rect 13556 26058 13584 26318
rect 13648 26314 13676 26726
rect 13636 26308 13688 26314
rect 13636 26250 13688 26256
rect 13464 26030 13584 26058
rect 13464 25974 13492 26030
rect 13452 25968 13504 25974
rect 13452 25910 13504 25916
rect 13544 25696 13596 25702
rect 13372 25656 13544 25684
rect 13544 25638 13596 25644
rect 13268 24948 13320 24954
rect 13268 24890 13320 24896
rect 13636 24336 13688 24342
rect 13636 24278 13688 24284
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13648 24138 13676 24278
rect 13636 24132 13688 24138
rect 13636 24074 13688 24080
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12900 23656 12952 23662
rect 12900 23598 12952 23604
rect 12912 22778 12940 23598
rect 13004 23322 13032 23666
rect 13176 23520 13228 23526
rect 13176 23462 13228 23468
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 13188 23225 13216 23462
rect 13174 23216 13230 23225
rect 13174 23151 13230 23160
rect 12900 22772 12952 22778
rect 12900 22714 12952 22720
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 13004 22094 13032 22714
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 13188 22234 13216 22578
rect 13176 22228 13228 22234
rect 13176 22170 13228 22176
rect 12912 22066 13032 22094
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12544 20058 12572 20334
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12544 18290 12572 18702
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12348 17060 12400 17066
rect 12348 17002 12400 17008
rect 12360 16658 12388 17002
rect 12636 16658 12664 20334
rect 12912 19786 12940 22066
rect 12992 20868 13044 20874
rect 12992 20810 13044 20816
rect 13004 20602 13032 20810
rect 12992 20596 13044 20602
rect 12992 20538 13044 20544
rect 12900 19780 12952 19786
rect 12900 19722 12952 19728
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12820 18766 12848 19110
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 14346 12480 16390
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12544 15162 12572 15370
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12452 13870 12480 14282
rect 12636 13938 12664 16594
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12256 12368 12308 12374
rect 12256 12310 12308 12316
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10980 11762 11008 12038
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10980 11218 11008 11562
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10980 8838 11008 11018
rect 12268 10606 12296 12310
rect 12452 11218 12480 13806
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12728 12850 12756 13738
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12544 12306 12572 12582
rect 12636 12306 12664 12718
rect 12912 12434 12940 19722
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 13096 17882 13124 19314
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13096 16658 13124 16934
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13188 15162 13216 15302
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 12820 12406 12940 12434
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12636 11898 12664 12242
rect 12820 12238 12848 12406
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12820 11778 12848 12174
rect 12728 11750 12848 11778
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12636 10606 12664 10746
rect 12728 10674 12756 11750
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 12256 10600 12308 10606
rect 12440 10600 12492 10606
rect 12256 10542 12308 10548
rect 12360 10548 12440 10554
rect 12360 10542 12492 10548
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 11256 10130 11284 10542
rect 11624 10130 11652 10542
rect 12360 10526 12480 10542
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 8974 11100 9862
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10980 7818 11008 8774
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 11256 7546 11284 10066
rect 11624 8090 11652 10066
rect 12164 10056 12216 10062
rect 12360 10044 12388 10526
rect 12636 10130 12664 10542
rect 12820 10470 12848 11086
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12216 10016 12388 10044
rect 12440 10056 12492 10062
rect 12164 9998 12216 10004
rect 12440 9998 12492 10004
rect 12176 9926 12204 9998
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12452 9722 12480 9998
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 11716 8090 11744 8434
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11624 7886 11652 8026
rect 12268 7954 12296 8366
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 12452 7886 12480 8434
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11992 7546 12020 7754
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 10980 7342 11008 7482
rect 12452 7342 12480 7822
rect 12636 7818 12664 8842
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 9876 6886 9996 6914
rect 10796 6886 10916 6914
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 9876 5234 9904 6886
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10704 4826 10732 5170
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 9402 2680 9458 2689
rect 5908 2644 5960 2650
rect 9402 2615 9458 2624
rect 5908 2586 5960 2592
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 9416 2514 9444 2615
rect 10796 2582 10824 6886
rect 11532 6798 11560 7142
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 12452 5710 12480 7278
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12452 5166 12480 5646
rect 13004 5302 13032 6054
rect 13188 5914 13216 6258
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 11348 2446 11376 4966
rect 11532 4622 11560 4966
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 13280 2582 13308 24006
rect 13372 23730 13400 24006
rect 13648 23730 13676 24074
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13372 23050 13400 23666
rect 13360 23044 13412 23050
rect 13360 22986 13412 22992
rect 13372 14006 13400 22986
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13648 20466 13676 21830
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13648 17746 13676 20402
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13648 16454 13676 17682
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13648 14958 13676 16390
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 13372 9761 13400 13942
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13464 10130 13492 11018
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13556 10062 13584 11086
rect 13648 11082 13676 14350
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13648 10130 13676 10406
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13358 9752 13414 9761
rect 13358 9687 13414 9696
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4078 13676 4966
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13648 2990 13676 4014
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13740 2774 13768 30126
rect 14016 30122 14044 31894
rect 14292 31822 14320 32166
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 14004 30116 14056 30122
rect 14004 30058 14056 30064
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14108 28762 14136 29106
rect 14096 28756 14148 28762
rect 14096 28698 14148 28704
rect 14004 28688 14056 28694
rect 14004 28630 14056 28636
rect 14278 28656 14334 28665
rect 13820 28484 13872 28490
rect 13820 28426 13872 28432
rect 13832 28150 13860 28426
rect 14016 28422 14044 28630
rect 14278 28591 14334 28600
rect 14292 28558 14320 28591
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13912 28144 13964 28150
rect 13912 28086 13964 28092
rect 13820 27668 13872 27674
rect 13820 27610 13872 27616
rect 13832 26926 13860 27610
rect 13924 27606 13952 28086
rect 14016 28082 14044 28358
rect 14292 28218 14320 28494
rect 14464 28416 14516 28422
rect 14464 28358 14516 28364
rect 14280 28212 14332 28218
rect 14280 28154 14332 28160
rect 14372 28144 14424 28150
rect 14372 28086 14424 28092
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 13912 27600 13964 27606
rect 13912 27542 13964 27548
rect 13820 26920 13872 26926
rect 13820 26862 13872 26868
rect 13818 26616 13874 26625
rect 13818 26551 13874 26560
rect 13832 26518 13860 26551
rect 13820 26512 13872 26518
rect 13820 26454 13872 26460
rect 13832 19922 13860 26454
rect 13924 26246 13952 27542
rect 14280 27532 14332 27538
rect 14280 27474 14332 27480
rect 14292 26790 14320 27474
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 13912 26240 13964 26246
rect 13912 26182 13964 26188
rect 14292 25906 14320 26726
rect 14384 25906 14412 28086
rect 14476 28082 14504 28358
rect 14464 28076 14516 28082
rect 14464 28018 14516 28024
rect 14476 26994 14504 28018
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 14568 27305 14596 27950
rect 14660 27538 14780 27554
rect 14648 27532 14780 27538
rect 14700 27526 14780 27532
rect 14648 27474 14700 27480
rect 14648 27396 14700 27402
rect 14648 27338 14700 27344
rect 14554 27296 14610 27305
rect 14554 27231 14610 27240
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 14568 26586 14596 27066
rect 14556 26580 14608 26586
rect 14556 26522 14608 26528
rect 14660 26382 14688 27338
rect 14752 27130 14780 27526
rect 14740 27124 14792 27130
rect 14740 27066 14792 27072
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14752 26382 14780 26930
rect 14648 26376 14700 26382
rect 14648 26318 14700 26324
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14280 25900 14332 25906
rect 14280 25842 14332 25848
rect 14372 25900 14424 25906
rect 14372 25842 14424 25848
rect 14096 25832 14148 25838
rect 14096 25774 14148 25780
rect 14108 25294 14136 25774
rect 14188 25696 14240 25702
rect 14188 25638 14240 25644
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 14096 24676 14148 24682
rect 14096 24618 14148 24624
rect 14108 24206 14136 24618
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 13912 22500 13964 22506
rect 13912 22442 13964 22448
rect 13924 22030 13952 22442
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13924 20602 13952 21082
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18290 13952 18566
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13832 17746 13860 18226
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13924 17678 13952 18226
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12986 13860 13126
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 14016 12782 14044 19858
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 18358 14136 18566
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 14094 17776 14150 17785
rect 14094 17711 14150 17720
rect 14108 17678 14136 17711
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14200 17202 14228 25638
rect 14384 25498 14412 25842
rect 14372 25492 14424 25498
rect 14372 25434 14424 25440
rect 14372 24404 14424 24410
rect 14372 24346 14424 24352
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14292 17338 14320 18702
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14108 16046 14136 16390
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14384 15994 14412 24346
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14568 22982 14596 24006
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14568 21554 14596 22918
rect 14660 22030 14688 26318
rect 14752 25974 14780 26318
rect 14844 26042 14872 32914
rect 15200 32904 15252 32910
rect 15200 32846 15252 32852
rect 15384 32904 15436 32910
rect 15384 32846 15436 32852
rect 15108 32768 15160 32774
rect 15108 32710 15160 32716
rect 14924 32564 14976 32570
rect 14924 32506 14976 32512
rect 14936 32434 14964 32506
rect 15120 32434 15148 32710
rect 15212 32570 15240 32846
rect 15200 32564 15252 32570
rect 15200 32506 15252 32512
rect 14924 32428 14976 32434
rect 14924 32370 14976 32376
rect 15108 32428 15160 32434
rect 15108 32370 15160 32376
rect 15120 31754 15148 32370
rect 15396 32337 15424 32846
rect 15382 32328 15438 32337
rect 15382 32263 15438 32272
rect 15292 31952 15344 31958
rect 15292 31894 15344 31900
rect 15028 31726 15148 31754
rect 15028 28218 15056 31726
rect 15304 31482 15332 31894
rect 15292 31476 15344 31482
rect 15292 31418 15344 31424
rect 15488 31278 15516 35686
rect 15568 35692 15620 35698
rect 15568 35634 15620 35640
rect 15660 35692 15712 35698
rect 15660 35634 15712 35640
rect 15764 31754 15792 41386
rect 15936 38956 15988 38962
rect 15936 38898 15988 38904
rect 15948 38554 15976 38898
rect 15936 38548 15988 38554
rect 15936 38490 15988 38496
rect 15936 37324 15988 37330
rect 15936 37266 15988 37272
rect 15844 36712 15896 36718
rect 15844 36654 15896 36660
rect 15856 36242 15884 36654
rect 15948 36394 15976 37266
rect 16040 36530 16068 43590
rect 16776 43450 16804 43726
rect 16764 43444 16816 43450
rect 16764 43386 16816 43392
rect 17052 43382 17080 43744
rect 17040 43376 17092 43382
rect 17040 43318 17092 43324
rect 17328 43314 17356 44882
rect 17696 44180 17724 45834
rect 17880 45490 17908 45970
rect 17868 45484 17920 45490
rect 17868 45426 17920 45432
rect 17972 45354 18000 46514
rect 18052 46096 18104 46102
rect 18052 46038 18104 46044
rect 18064 45490 18092 46038
rect 18052 45484 18104 45490
rect 18052 45426 18104 45432
rect 17960 45348 18012 45354
rect 17960 45290 18012 45296
rect 17776 44192 17828 44198
rect 17696 44152 17776 44180
rect 17776 44134 17828 44140
rect 17788 43908 17816 44134
rect 17960 43920 18012 43926
rect 17788 43880 17960 43908
rect 17960 43862 18012 43868
rect 16580 43308 16632 43314
rect 16580 43250 16632 43256
rect 17316 43308 17368 43314
rect 17316 43250 17368 43256
rect 16592 42906 16620 43250
rect 17328 42906 17356 43250
rect 18052 43104 18104 43110
rect 18052 43046 18104 43052
rect 16580 42900 16632 42906
rect 16580 42842 16632 42848
rect 17316 42900 17368 42906
rect 17316 42842 17368 42848
rect 16212 42764 16264 42770
rect 16212 42706 16264 42712
rect 16224 37913 16252 42706
rect 18064 42702 18092 43046
rect 18052 42696 18104 42702
rect 18052 42638 18104 42644
rect 17592 42628 17644 42634
rect 17592 42570 17644 42576
rect 17040 41676 17092 41682
rect 17040 41618 17092 41624
rect 16948 41132 17000 41138
rect 16948 41074 17000 41080
rect 16580 40928 16632 40934
rect 16580 40870 16632 40876
rect 16592 40526 16620 40870
rect 16672 40724 16724 40730
rect 16672 40666 16724 40672
rect 16580 40520 16632 40526
rect 16580 40462 16632 40468
rect 16396 39024 16448 39030
rect 16396 38966 16448 38972
rect 16408 38554 16436 38966
rect 16684 38842 16712 40666
rect 16960 40186 16988 41074
rect 17052 41070 17080 41618
rect 17316 41608 17368 41614
rect 17316 41550 17368 41556
rect 17328 41414 17356 41550
rect 17328 41386 17448 41414
rect 17420 41206 17448 41386
rect 17408 41200 17460 41206
rect 17408 41142 17460 41148
rect 17040 41064 17092 41070
rect 17040 41006 17092 41012
rect 17052 40458 17080 41006
rect 17040 40452 17092 40458
rect 17040 40394 17092 40400
rect 16948 40180 17000 40186
rect 16948 40122 17000 40128
rect 17316 39500 17368 39506
rect 17316 39442 17368 39448
rect 16764 39296 16816 39302
rect 16764 39238 16816 39244
rect 17132 39296 17184 39302
rect 17132 39238 17184 39244
rect 16592 38814 16712 38842
rect 16396 38548 16448 38554
rect 16396 38490 16448 38496
rect 16210 37904 16266 37913
rect 16210 37839 16266 37848
rect 16224 37466 16252 37839
rect 16212 37460 16264 37466
rect 16212 37402 16264 37408
rect 16488 36916 16540 36922
rect 16488 36858 16540 36864
rect 16500 36786 16528 36858
rect 16488 36780 16540 36786
rect 16488 36722 16540 36728
rect 16488 36644 16540 36650
rect 16488 36586 16540 36592
rect 16040 36502 16252 36530
rect 15948 36366 16160 36394
rect 15844 36236 15896 36242
rect 15844 36178 15896 36184
rect 15844 35624 15896 35630
rect 15844 35566 15896 35572
rect 15752 31748 15804 31754
rect 15752 31690 15804 31696
rect 15476 31272 15528 31278
rect 15476 31214 15528 31220
rect 15764 30666 15792 31690
rect 15752 30660 15804 30666
rect 15752 30602 15804 30608
rect 15384 30048 15436 30054
rect 15384 29990 15436 29996
rect 15660 30048 15712 30054
rect 15660 29990 15712 29996
rect 15108 29708 15160 29714
rect 15108 29650 15160 29656
rect 15120 29578 15148 29650
rect 15396 29646 15424 29990
rect 15672 29646 15700 29990
rect 15384 29640 15436 29646
rect 15384 29582 15436 29588
rect 15660 29640 15712 29646
rect 15660 29582 15712 29588
rect 15108 29572 15160 29578
rect 15108 29514 15160 29520
rect 15120 29102 15148 29514
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15212 29238 15240 29446
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 15200 29232 15252 29238
rect 15200 29174 15252 29180
rect 15108 29096 15160 29102
rect 15488 29073 15516 29242
rect 15108 29038 15160 29044
rect 15474 29064 15530 29073
rect 15474 28999 15530 29008
rect 15108 28960 15160 28966
rect 15108 28902 15160 28908
rect 15120 28490 15148 28902
rect 15108 28484 15160 28490
rect 15108 28426 15160 28432
rect 15016 28212 15068 28218
rect 15016 28154 15068 28160
rect 15120 27538 15148 28426
rect 15384 28416 15436 28422
rect 15384 28358 15436 28364
rect 15200 28008 15252 28014
rect 15200 27950 15252 27956
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 15212 27470 15240 27950
rect 15200 27464 15252 27470
rect 15200 27406 15252 27412
rect 14922 27296 14978 27305
rect 14922 27231 14978 27240
rect 14832 26036 14884 26042
rect 14832 25978 14884 25984
rect 14740 25968 14792 25974
rect 14740 25910 14792 25916
rect 14936 23338 14964 27231
rect 15396 27062 15424 28358
rect 15856 28098 15884 35566
rect 16028 34944 16080 34950
rect 16028 34886 16080 34892
rect 16040 34678 16068 34886
rect 16028 34672 16080 34678
rect 16028 34614 16080 34620
rect 15936 32836 15988 32842
rect 15936 32778 15988 32784
rect 15948 31822 15976 32778
rect 16028 32224 16080 32230
rect 16028 32166 16080 32172
rect 16040 31822 16068 32166
rect 15936 31816 15988 31822
rect 15936 31758 15988 31764
rect 16028 31816 16080 31822
rect 16028 31758 16080 31764
rect 15948 31482 15976 31758
rect 16028 31680 16080 31686
rect 16028 31622 16080 31628
rect 15936 31476 15988 31482
rect 15936 31418 15988 31424
rect 16040 30734 16068 31622
rect 16028 30728 16080 30734
rect 16028 30670 16080 30676
rect 16040 30326 16068 30670
rect 16132 30326 16160 36366
rect 16224 31754 16252 36502
rect 16500 36258 16528 36586
rect 16592 36394 16620 38814
rect 16672 38752 16724 38758
rect 16672 38694 16724 38700
rect 16684 38350 16712 38694
rect 16776 38350 16804 39238
rect 16856 38888 16908 38894
rect 16856 38830 16908 38836
rect 16672 38344 16724 38350
rect 16672 38286 16724 38292
rect 16764 38344 16816 38350
rect 16764 38286 16816 38292
rect 16868 38214 16896 38830
rect 16948 38412 17000 38418
rect 16948 38354 17000 38360
rect 17040 38412 17092 38418
rect 17040 38354 17092 38360
rect 16856 38208 16908 38214
rect 16856 38150 16908 38156
rect 16868 36922 16896 38150
rect 16856 36916 16908 36922
rect 16856 36858 16908 36864
rect 16764 36848 16816 36854
rect 16762 36816 16764 36825
rect 16816 36816 16818 36825
rect 16762 36751 16818 36760
rect 16764 36576 16816 36582
rect 16764 36518 16816 36524
rect 16592 36366 16712 36394
rect 16500 36242 16620 36258
rect 16500 36236 16632 36242
rect 16500 36230 16580 36236
rect 16580 36178 16632 36184
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 16500 35834 16528 36110
rect 16488 35828 16540 35834
rect 16488 35770 16540 35776
rect 16304 34604 16356 34610
rect 16304 34546 16356 34552
rect 16316 34202 16344 34546
rect 16684 34490 16712 36366
rect 16776 35698 16804 36518
rect 16764 35692 16816 35698
rect 16764 35634 16816 35640
rect 16684 34462 16804 34490
rect 16672 34400 16724 34406
rect 16672 34342 16724 34348
rect 16304 34196 16356 34202
rect 16304 34138 16356 34144
rect 16684 33998 16712 34342
rect 16776 34066 16804 34462
rect 16764 34060 16816 34066
rect 16764 34002 16816 34008
rect 16672 33992 16724 33998
rect 16672 33934 16724 33940
rect 16960 33946 16988 38354
rect 17052 37874 17080 38354
rect 17040 37868 17092 37874
rect 17040 37810 17092 37816
rect 16580 33448 16632 33454
rect 16580 33390 16632 33396
rect 16304 33312 16356 33318
rect 16304 33254 16356 33260
rect 16316 32212 16344 33254
rect 16396 32428 16448 32434
rect 16396 32370 16448 32376
rect 16408 32337 16436 32370
rect 16394 32328 16450 32337
rect 16394 32263 16450 32272
rect 16396 32224 16448 32230
rect 16316 32184 16396 32212
rect 16396 32166 16448 32172
rect 16408 31890 16436 32166
rect 16396 31884 16448 31890
rect 16396 31826 16448 31832
rect 16224 31726 16436 31754
rect 16408 30410 16436 31726
rect 16488 30728 16540 30734
rect 16488 30670 16540 30676
rect 16224 30382 16436 30410
rect 16028 30320 16080 30326
rect 16028 30262 16080 30268
rect 16120 30320 16172 30326
rect 16120 30262 16172 30268
rect 15936 30252 15988 30258
rect 15936 30194 15988 30200
rect 15948 29492 15976 30194
rect 16120 30184 16172 30190
rect 16224 30138 16252 30382
rect 16304 30252 16356 30258
rect 16304 30194 16356 30200
rect 16172 30132 16252 30138
rect 16120 30126 16252 30132
rect 16132 30110 16252 30126
rect 16316 30002 16344 30194
rect 16408 30190 16436 30382
rect 16500 30326 16528 30670
rect 16488 30320 16540 30326
rect 16488 30262 16540 30268
rect 16396 30184 16448 30190
rect 16396 30126 16448 30132
rect 16224 29974 16344 30002
rect 16120 29504 16172 29510
rect 15948 29464 16120 29492
rect 15948 29306 15976 29464
rect 16120 29446 16172 29452
rect 15936 29300 15988 29306
rect 15936 29242 15988 29248
rect 15580 28070 15884 28098
rect 15476 28008 15528 28014
rect 15474 27976 15476 27985
rect 15528 27976 15530 27985
rect 15474 27911 15530 27920
rect 15384 27056 15436 27062
rect 15384 26998 15436 27004
rect 15200 26920 15252 26926
rect 15200 26862 15252 26868
rect 15108 26580 15160 26586
rect 15108 26522 15160 26528
rect 15120 26489 15148 26522
rect 15212 26518 15240 26862
rect 15200 26512 15252 26518
rect 15106 26480 15162 26489
rect 15200 26454 15252 26460
rect 15476 26512 15528 26518
rect 15476 26454 15528 26460
rect 15106 26415 15162 26424
rect 15488 25906 15516 26454
rect 15476 25900 15528 25906
rect 15476 25842 15528 25848
rect 15580 24154 15608 28070
rect 16224 28014 16252 29974
rect 16304 28144 16356 28150
rect 16304 28086 16356 28092
rect 15844 28008 15896 28014
rect 15844 27950 15896 27956
rect 16028 28008 16080 28014
rect 16028 27950 16080 27956
rect 16212 28008 16264 28014
rect 16212 27950 16264 27956
rect 15856 27334 15884 27950
rect 15844 27328 15896 27334
rect 15844 27270 15896 27276
rect 15750 27024 15806 27033
rect 15750 26959 15806 26968
rect 15764 26450 15792 26959
rect 16040 26790 16068 27950
rect 16316 27674 16344 28086
rect 16396 28076 16448 28082
rect 16396 28018 16448 28024
rect 16488 28076 16540 28082
rect 16488 28018 16540 28024
rect 16304 27668 16356 27674
rect 16304 27610 16356 27616
rect 16028 26784 16080 26790
rect 16028 26726 16080 26732
rect 15752 26444 15804 26450
rect 15752 26386 15804 26392
rect 16040 26314 16068 26726
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 16028 26308 16080 26314
rect 16028 26250 16080 26256
rect 15752 26036 15804 26042
rect 15752 25978 15804 25984
rect 15304 24126 15608 24154
rect 15016 24064 15068 24070
rect 15016 24006 15068 24012
rect 15028 23730 15056 24006
rect 15016 23724 15068 23730
rect 15016 23666 15068 23672
rect 15108 23520 15160 23526
rect 15108 23462 15160 23468
rect 14844 23310 14964 23338
rect 14740 23180 14792 23186
rect 14740 23122 14792 23128
rect 14752 22658 14780 23122
rect 14844 23066 14872 23310
rect 14844 23038 15056 23066
rect 15120 23050 15148 23462
rect 14752 22630 14964 22658
rect 14936 22574 14964 22630
rect 14832 22568 14884 22574
rect 14832 22510 14884 22516
rect 14924 22568 14976 22574
rect 14924 22510 14976 22516
rect 14844 22166 14872 22510
rect 14832 22160 14884 22166
rect 14832 22102 14884 22108
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14556 21548 14608 21554
rect 14556 21490 14608 21496
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14476 18222 14504 18770
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14476 16153 14504 17682
rect 14568 17338 14596 18362
rect 14660 17746 14688 21966
rect 14936 21894 14964 22510
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 14740 20868 14792 20874
rect 14740 20810 14792 20816
rect 14752 20602 14780 20810
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14844 18834 14872 19178
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14752 18222 14780 18702
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 15028 17218 15056 23038
rect 15108 23044 15160 23050
rect 15108 22986 15160 22992
rect 15304 22778 15332 24126
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15488 23730 15516 24006
rect 15384 23724 15436 23730
rect 15384 23666 15436 23672
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15396 23322 15424 23666
rect 15384 23316 15436 23322
rect 15384 23258 15436 23264
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 15488 22094 15516 23666
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15580 22778 15608 23054
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15672 22234 15700 23054
rect 15660 22228 15712 22234
rect 15660 22170 15712 22176
rect 15488 22066 15608 22094
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15212 19938 15240 20742
rect 15120 19910 15240 19938
rect 15120 19258 15148 19910
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 15212 19446 15240 19722
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 15120 19230 15240 19258
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 15120 18222 15148 18770
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14936 17190 15056 17218
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14462 16144 14518 16153
rect 14752 16114 14780 16390
rect 14462 16079 14464 16088
rect 14516 16079 14518 16088
rect 14740 16108 14792 16114
rect 14464 16050 14516 16056
rect 14740 16050 14792 16056
rect 14384 15966 14780 15994
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14660 15638 14688 15846
rect 14648 15632 14700 15638
rect 14648 15574 14700 15580
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14660 13462 14688 13942
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14292 12850 14320 13330
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14568 12850 14596 13126
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 13924 12434 13952 12718
rect 13924 12406 14228 12434
rect 14200 11762 14228 12406
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14200 10810 14228 11698
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14292 10742 14320 12786
rect 14660 12442 14688 13262
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11218 14504 12038
rect 14752 11218 14780 15966
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14280 10736 14332 10742
rect 14108 10684 14280 10690
rect 14108 10678 14332 10684
rect 14108 10662 14320 10678
rect 14108 10130 14136 10662
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14200 10062 14228 10406
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14556 9104 14608 9110
rect 14844 9058 14872 17138
rect 14556 9046 14608 9052
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13832 8294 13860 8774
rect 14016 8634 14044 8842
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 7546 13860 8230
rect 13924 8090 13952 8434
rect 14200 8430 14228 8978
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 14292 7886 14320 8298
rect 14568 7886 14596 9046
rect 14752 9030 14872 9058
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14016 5846 14044 6258
rect 14200 6254 14228 7754
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14384 7478 14412 7686
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13912 5636 13964 5642
rect 13912 5578 13964 5584
rect 13924 5030 13952 5578
rect 14108 5234 14136 6054
rect 14200 5846 14228 6190
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14476 5574 14504 6802
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14568 6186 14596 6734
rect 14660 6254 14688 6734
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14660 5914 14688 6190
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14752 5778 14780 9030
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14844 8498 14872 8774
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14936 6118 14964 17190
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13326 15056 13670
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 15120 12306 15148 17682
rect 15212 12434 15240 19230
rect 15304 18154 15332 20878
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15292 18148 15344 18154
rect 15292 18090 15344 18096
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15304 16114 15332 16390
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15304 15162 15332 15370
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15396 14414 15424 19654
rect 15580 19310 15608 22066
rect 15764 21486 15792 25978
rect 16132 24970 16160 26386
rect 16212 26376 16264 26382
rect 16212 26318 16264 26324
rect 16224 25430 16252 26318
rect 16316 25974 16344 27610
rect 16408 27402 16436 28018
rect 16500 27878 16528 28018
rect 16488 27872 16540 27878
rect 16488 27814 16540 27820
rect 16396 27396 16448 27402
rect 16396 27338 16448 27344
rect 16408 26994 16436 27338
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 16304 25968 16356 25974
rect 16304 25910 16356 25916
rect 16212 25424 16264 25430
rect 16212 25366 16264 25372
rect 16316 25294 16344 25910
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 16132 24942 16436 24970
rect 16028 24744 16080 24750
rect 16028 24686 16080 24692
rect 16040 24274 16068 24686
rect 16028 24268 16080 24274
rect 16028 24210 16080 24216
rect 15936 24200 15988 24206
rect 15936 24142 15988 24148
rect 15948 23866 15976 24142
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 16212 22568 16264 22574
rect 16212 22510 16264 22516
rect 16224 22438 16252 22510
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 15752 21480 15804 21486
rect 15750 21448 15752 21457
rect 15804 21448 15806 21457
rect 15750 21383 15806 21392
rect 15764 20806 15792 21383
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15856 20806 15884 21286
rect 16132 20806 16160 21490
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 15856 20602 15884 20742
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15948 19990 15976 20402
rect 16224 20398 16252 22374
rect 16212 20392 16264 20398
rect 16212 20334 16264 20340
rect 15936 19984 15988 19990
rect 15936 19926 15988 19932
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15580 18222 15608 18362
rect 15672 18272 15700 19790
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15764 18426 15792 19314
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15752 18284 15804 18290
rect 15672 18244 15752 18272
rect 15752 18226 15804 18232
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15856 17814 15884 19314
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 16040 18766 16068 19110
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 16028 18760 16080 18766
rect 16080 18708 16160 18714
rect 16028 18702 16160 18708
rect 15948 18222 15976 18702
rect 16040 18686 16160 18702
rect 16132 18222 16160 18686
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 16118 18048 16174 18057
rect 16118 17983 16174 17992
rect 15844 17808 15896 17814
rect 15844 17750 15896 17756
rect 15476 17672 15528 17678
rect 15474 17640 15476 17649
rect 15660 17672 15712 17678
rect 15528 17640 15530 17649
rect 15660 17614 15712 17620
rect 15474 17575 15530 17584
rect 15672 17542 15700 17614
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 17338 15700 17478
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15856 16182 15884 16390
rect 15844 16176 15896 16182
rect 15844 16118 15896 16124
rect 15856 15638 15884 16118
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15948 14958 15976 16594
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 16132 14346 16160 17983
rect 16224 17134 16252 20334
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16316 17882 16344 18090
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16224 16658 16252 17070
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16212 15360 16264 15366
rect 16212 15302 16264 15308
rect 16224 15162 16252 15302
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16224 14822 16252 15098
rect 16316 15094 16344 15846
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 16120 14340 16172 14346
rect 16120 14282 16172 14288
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15304 12986 15332 13874
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15672 12442 15700 12582
rect 15660 12436 15712 12442
rect 15212 12406 15332 12434
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15120 10690 15148 12242
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15212 10742 15240 10950
rect 15028 10674 15148 10690
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15016 10668 15148 10674
rect 15068 10662 15148 10668
rect 15016 10610 15068 10616
rect 15028 9042 15056 10610
rect 15304 10588 15332 12406
rect 15948 12434 15976 14282
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16132 12986 16160 13126
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 15660 12378 15712 12384
rect 15764 12406 15976 12434
rect 15672 12238 15700 12378
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15212 10560 15332 10588
rect 15212 9081 15240 10560
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15304 10198 15332 10406
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15198 9072 15254 9081
rect 15016 9036 15068 9042
rect 15198 9007 15254 9016
rect 15016 8978 15068 8984
rect 15212 6866 15240 9007
rect 15764 8945 15792 12406
rect 16224 12102 16252 12718
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15856 10810 15884 10950
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15948 10742 15976 11086
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15948 10606 15976 10678
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 16316 9926 16344 11018
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 15750 8936 15806 8945
rect 15750 8871 15806 8880
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15580 8634 15608 8774
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15672 7954 15700 8774
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15764 6866 15792 8871
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16028 7812 16080 7818
rect 16028 7754 16080 7760
rect 16040 7546 16068 7754
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16132 7410 16160 8774
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15384 6248 15436 6254
rect 15488 6236 15516 6734
rect 15580 6322 15608 6802
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15672 6322 15700 6598
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15436 6208 15516 6236
rect 15384 6190 15436 6196
rect 15016 6180 15068 6186
rect 15016 6122 15068 6128
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 15028 6066 15056 6122
rect 15028 6038 15148 6066
rect 15016 5840 15068 5846
rect 15016 5782 15068 5788
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14476 5098 14504 5510
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 15028 4622 15056 5782
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 15120 4486 15148 6038
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14384 3738 14412 4082
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14752 3534 14780 4422
rect 15120 4010 15148 4422
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 15488 3398 15516 5850
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15856 4078 15884 4558
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15856 3534 15884 4014
rect 16408 3602 16436 24942
rect 16500 22642 16528 27814
rect 16592 27674 16620 33390
rect 16684 31754 16712 33934
rect 16960 33918 17080 33946
rect 16948 33856 17000 33862
rect 16948 33798 17000 33804
rect 16960 33017 16988 33798
rect 16946 33008 17002 33017
rect 17052 32978 17080 33918
rect 16946 32943 16948 32952
rect 17000 32943 17002 32952
rect 17040 32972 17092 32978
rect 16948 32914 17000 32920
rect 17040 32914 17092 32920
rect 16684 31726 16804 31754
rect 16776 29714 16804 31726
rect 17040 30252 17092 30258
rect 17040 30194 17092 30200
rect 17052 30054 17080 30194
rect 17040 30048 17092 30054
rect 17040 29990 17092 29996
rect 17052 29850 17080 29990
rect 17040 29844 17092 29850
rect 17040 29786 17092 29792
rect 16764 29708 16816 29714
rect 16764 29650 16816 29656
rect 16764 29028 16816 29034
rect 16764 28970 16816 28976
rect 16580 27668 16632 27674
rect 16580 27610 16632 27616
rect 16672 27328 16724 27334
rect 16672 27270 16724 27276
rect 16580 27056 16632 27062
rect 16684 27044 16712 27270
rect 16776 27130 16804 28970
rect 17040 27600 17092 27606
rect 17040 27542 17092 27548
rect 17052 27470 17080 27542
rect 16948 27464 17000 27470
rect 16948 27406 17000 27412
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 16764 27124 16816 27130
rect 16764 27066 16816 27072
rect 16960 27062 16988 27406
rect 16632 27016 16712 27044
rect 16948 27056 17000 27062
rect 16580 26998 16632 27004
rect 16948 26998 17000 27004
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16500 12782 16528 22578
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16500 11218 16528 12718
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16500 9042 16528 11154
rect 16592 9382 16620 26998
rect 16764 26920 16816 26926
rect 16948 26920 17000 26926
rect 16764 26862 16816 26868
rect 16868 26880 16948 26908
rect 16776 26450 16804 26862
rect 16764 26444 16816 26450
rect 16764 26386 16816 26392
rect 16776 25362 16804 26386
rect 16868 26314 16896 26880
rect 16948 26862 17000 26868
rect 17052 26518 17080 27406
rect 17040 26512 17092 26518
rect 17040 26454 17092 26460
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16776 18902 16804 21966
rect 16764 18896 16816 18902
rect 16764 18838 16816 18844
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 16684 18222 16712 18770
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16684 16658 16712 18158
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16684 15910 16712 16186
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16684 10062 16712 13262
rect 16868 12434 16896 26250
rect 17052 26246 17080 26318
rect 17040 26240 17092 26246
rect 17040 26182 17092 26188
rect 17052 25294 17080 26182
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 17052 22642 17080 22918
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 17144 22094 17172 39238
rect 17328 38894 17356 39442
rect 17316 38888 17368 38894
rect 17316 38830 17368 38836
rect 17224 38752 17276 38758
rect 17224 38694 17276 38700
rect 17236 37806 17264 38694
rect 17224 37800 17276 37806
rect 17224 37742 17276 37748
rect 17236 37330 17264 37742
rect 17224 37324 17276 37330
rect 17224 37266 17276 37272
rect 17420 35766 17448 41142
rect 17500 39364 17552 39370
rect 17500 39306 17552 39312
rect 17512 38826 17540 39306
rect 17500 38820 17552 38826
rect 17500 38762 17552 38768
rect 17500 37800 17552 37806
rect 17500 37742 17552 37748
rect 17408 35760 17460 35766
rect 17408 35702 17460 35708
rect 17316 35216 17368 35222
rect 17316 35158 17368 35164
rect 17328 34746 17356 35158
rect 17316 34740 17368 34746
rect 17316 34682 17368 34688
rect 17224 32768 17276 32774
rect 17224 32710 17276 32716
rect 17236 32434 17264 32710
rect 17224 32428 17276 32434
rect 17224 32370 17276 32376
rect 17512 31872 17540 37742
rect 17328 31844 17540 31872
rect 17224 29708 17276 29714
rect 17224 29650 17276 29656
rect 17236 29170 17264 29650
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17328 29102 17356 31844
rect 17604 31754 17632 42570
rect 18064 42362 18092 42638
rect 18052 42356 18104 42362
rect 18052 42298 18104 42304
rect 18052 41472 18104 41478
rect 18248 41460 18276 46990
rect 18328 43648 18380 43654
rect 18328 43590 18380 43596
rect 18340 43314 18368 43590
rect 18328 43308 18380 43314
rect 18328 43250 18380 43256
rect 18104 41432 18276 41460
rect 18052 41414 18104 41420
rect 17684 40384 17736 40390
rect 17684 40326 17736 40332
rect 17776 40384 17828 40390
rect 17776 40326 17828 40332
rect 17696 40186 17724 40326
rect 17684 40180 17736 40186
rect 17684 40122 17736 40128
rect 17696 38486 17724 40122
rect 17788 39982 17816 40326
rect 17776 39976 17828 39982
rect 17776 39918 17828 39924
rect 17776 39840 17828 39846
rect 17776 39782 17828 39788
rect 17788 39030 17816 39782
rect 17776 39024 17828 39030
rect 17776 38966 17828 38972
rect 17960 38888 18012 38894
rect 17960 38830 18012 38836
rect 17684 38480 17736 38486
rect 17684 38422 17736 38428
rect 17776 38412 17828 38418
rect 17776 38354 17828 38360
rect 17868 38412 17920 38418
rect 17868 38354 17920 38360
rect 17682 38040 17738 38049
rect 17682 37975 17738 37984
rect 17696 37806 17724 37975
rect 17788 37856 17816 38354
rect 17880 38321 17908 38354
rect 17866 38312 17922 38321
rect 17866 38247 17922 38256
rect 17972 37874 18000 38830
rect 17868 37868 17920 37874
rect 17788 37828 17868 37856
rect 17868 37810 17920 37816
rect 17960 37868 18012 37874
rect 17960 37810 18012 37816
rect 17684 37800 17736 37806
rect 17684 37742 17736 37748
rect 17776 37324 17828 37330
rect 17776 37266 17828 37272
rect 17684 35080 17736 35086
rect 17684 35022 17736 35028
rect 17696 34610 17724 35022
rect 17684 34604 17736 34610
rect 17684 34546 17736 34552
rect 17788 31754 17816 37266
rect 17960 36780 18012 36786
rect 17960 36722 18012 36728
rect 17972 35834 18000 36722
rect 17960 35828 18012 35834
rect 17960 35770 18012 35776
rect 18064 35698 18092 41414
rect 18432 41206 18460 46990
rect 19444 46374 19472 47398
rect 20260 47116 20312 47122
rect 20180 47076 20260 47104
rect 20180 46510 20208 47076
rect 20260 47058 20312 47064
rect 20364 46986 20392 47602
rect 21364 47048 21416 47054
rect 21364 46990 21416 46996
rect 20352 46980 20404 46986
rect 20352 46922 20404 46928
rect 20260 46708 20312 46714
rect 20260 46650 20312 46656
rect 20168 46504 20220 46510
rect 20168 46446 20220 46452
rect 19432 46368 19484 46374
rect 19432 46310 19484 46316
rect 19444 46034 19472 46310
rect 19432 46028 19484 46034
rect 19432 45970 19484 45976
rect 19984 45824 20036 45830
rect 19984 45766 20036 45772
rect 20168 45824 20220 45830
rect 20168 45766 20220 45772
rect 19996 45490 20024 45766
rect 20180 45490 20208 45766
rect 19984 45484 20036 45490
rect 19984 45426 20036 45432
rect 20168 45484 20220 45490
rect 20168 45426 20220 45432
rect 20180 44402 20208 45426
rect 19708 44396 19760 44402
rect 19708 44338 19760 44344
rect 20168 44396 20220 44402
rect 20168 44338 20220 44344
rect 19720 43994 19748 44338
rect 19984 44192 20036 44198
rect 19984 44134 20036 44140
rect 19708 43988 19760 43994
rect 19708 43930 19760 43936
rect 19156 43920 19208 43926
rect 19156 43862 19208 43868
rect 19064 43784 19116 43790
rect 19062 43752 19064 43761
rect 19116 43752 19118 43761
rect 19062 43687 19118 43696
rect 19076 43654 19104 43687
rect 19064 43648 19116 43654
rect 19064 43590 19116 43596
rect 19064 42560 19116 42566
rect 19064 42502 19116 42508
rect 19076 42362 19104 42502
rect 19064 42356 19116 42362
rect 19064 42298 19116 42304
rect 19064 42016 19116 42022
rect 19064 41958 19116 41964
rect 19076 41614 19104 41958
rect 19168 41682 19196 43862
rect 19708 43376 19760 43382
rect 19708 43318 19760 43324
rect 19616 43308 19668 43314
rect 19616 43250 19668 43256
rect 19628 42702 19656 43250
rect 19720 42770 19748 43318
rect 19708 42764 19760 42770
rect 19708 42706 19760 42712
rect 19892 42764 19944 42770
rect 19892 42706 19944 42712
rect 19616 42696 19668 42702
rect 19616 42638 19668 42644
rect 19248 42560 19300 42566
rect 19248 42502 19300 42508
rect 19708 42560 19760 42566
rect 19708 42502 19760 42508
rect 19260 42226 19288 42502
rect 19248 42220 19300 42226
rect 19248 42162 19300 42168
rect 19524 42016 19576 42022
rect 19524 41958 19576 41964
rect 19156 41676 19208 41682
rect 19156 41618 19208 41624
rect 19536 41614 19564 41958
rect 19064 41608 19116 41614
rect 19064 41550 19116 41556
rect 19524 41608 19576 41614
rect 19524 41550 19576 41556
rect 18880 41472 18932 41478
rect 18880 41414 18932 41420
rect 18892 41206 18920 41414
rect 18420 41200 18472 41206
rect 18420 41142 18472 41148
rect 18880 41200 18932 41206
rect 18880 41142 18932 41148
rect 18604 41132 18656 41138
rect 18604 41074 18656 41080
rect 18236 40928 18288 40934
rect 18236 40870 18288 40876
rect 18248 40594 18276 40870
rect 18236 40588 18288 40594
rect 18236 40530 18288 40536
rect 18248 38978 18276 40530
rect 18616 40390 18644 41074
rect 18696 40588 18748 40594
rect 18696 40530 18748 40536
rect 18604 40384 18656 40390
rect 18604 40326 18656 40332
rect 18156 38950 18276 38978
rect 18156 38214 18184 38950
rect 18236 38888 18288 38894
rect 18236 38830 18288 38836
rect 18248 38418 18276 38830
rect 18236 38412 18288 38418
rect 18236 38354 18288 38360
rect 18420 38344 18472 38350
rect 18420 38286 18472 38292
rect 18144 38208 18196 38214
rect 18144 38150 18196 38156
rect 18156 38010 18184 38150
rect 18432 38010 18460 38286
rect 18144 38004 18196 38010
rect 18144 37946 18196 37952
rect 18420 38004 18472 38010
rect 18420 37946 18472 37952
rect 18328 37800 18380 37806
rect 18380 37760 18460 37788
rect 18328 37742 18380 37748
rect 18236 36168 18288 36174
rect 18236 36110 18288 36116
rect 18052 35692 18104 35698
rect 18052 35634 18104 35640
rect 17868 32972 17920 32978
rect 17868 32914 17920 32920
rect 17972 32932 18184 32960
rect 17880 32881 17908 32914
rect 17866 32872 17922 32881
rect 17866 32807 17922 32816
rect 17972 32774 18000 32932
rect 18052 32836 18104 32842
rect 18052 32778 18104 32784
rect 17960 32768 18012 32774
rect 17960 32710 18012 32716
rect 18064 32570 18092 32778
rect 18156 32570 18184 32932
rect 17960 32564 18012 32570
rect 17960 32506 18012 32512
rect 18052 32564 18104 32570
rect 18052 32506 18104 32512
rect 18144 32564 18196 32570
rect 18144 32506 18196 32512
rect 17512 31726 17632 31754
rect 17696 31726 17816 31754
rect 17408 29640 17460 29646
rect 17408 29582 17460 29588
rect 17420 29306 17448 29582
rect 17408 29300 17460 29306
rect 17408 29242 17460 29248
rect 17512 29238 17540 31726
rect 17696 30190 17724 31726
rect 17972 31482 18000 32506
rect 18142 32328 18198 32337
rect 18142 32263 18198 32272
rect 18156 32230 18184 32263
rect 18144 32224 18196 32230
rect 18144 32166 18196 32172
rect 18248 31793 18276 36110
rect 18328 35012 18380 35018
rect 18328 34954 18380 34960
rect 18340 34202 18368 34954
rect 18328 34196 18380 34202
rect 18328 34138 18380 34144
rect 18328 33924 18380 33930
rect 18328 33866 18380 33872
rect 18234 31784 18290 31793
rect 18064 31742 18234 31770
rect 17960 31476 18012 31482
rect 17960 31418 18012 31424
rect 17958 30968 18014 30977
rect 17958 30903 17960 30912
rect 18012 30903 18014 30912
rect 17960 30874 18012 30880
rect 17684 30184 17736 30190
rect 17684 30126 17736 30132
rect 17960 30184 18012 30190
rect 17960 30126 18012 30132
rect 17500 29232 17552 29238
rect 17500 29174 17552 29180
rect 17316 29096 17368 29102
rect 17316 29038 17368 29044
rect 17696 29034 17724 30126
rect 17972 29832 18000 30126
rect 17788 29804 18000 29832
rect 17788 29714 17816 29804
rect 17776 29708 17828 29714
rect 17776 29650 17828 29656
rect 17960 29708 18012 29714
rect 17960 29650 18012 29656
rect 17972 29102 18000 29650
rect 17960 29096 18012 29102
rect 17960 29038 18012 29044
rect 17684 29028 17736 29034
rect 17684 28970 17736 28976
rect 17592 28008 17644 28014
rect 17592 27950 17644 27956
rect 17604 27674 17632 27950
rect 17696 27674 17724 28970
rect 18064 27878 18092 31742
rect 18234 31719 18290 31728
rect 18340 30394 18368 33866
rect 18432 31754 18460 37760
rect 18708 37754 18736 40530
rect 19064 40452 19116 40458
rect 19064 40394 19116 40400
rect 19076 38350 19104 40394
rect 19720 39438 19748 42502
rect 19904 42158 19932 42706
rect 19892 42152 19944 42158
rect 19892 42094 19944 42100
rect 19904 41818 19932 42094
rect 19892 41812 19944 41818
rect 19892 41754 19944 41760
rect 19708 39432 19760 39438
rect 19708 39374 19760 39380
rect 19524 38956 19576 38962
rect 19524 38898 19576 38904
rect 19340 38752 19392 38758
rect 19340 38694 19392 38700
rect 19064 38344 19116 38350
rect 19064 38286 19116 38292
rect 18972 38276 19024 38282
rect 18972 38218 19024 38224
rect 18984 38049 19012 38218
rect 18970 38040 19026 38049
rect 18970 37975 19026 37984
rect 19076 37874 19104 38286
rect 19352 37942 19380 38694
rect 19432 38208 19484 38214
rect 19432 38150 19484 38156
rect 19340 37936 19392 37942
rect 19340 37878 19392 37884
rect 19064 37868 19116 37874
rect 19064 37810 19116 37816
rect 18708 37726 18920 37754
rect 18604 37664 18656 37670
rect 18604 37606 18656 37612
rect 18696 37664 18748 37670
rect 18696 37606 18748 37612
rect 18512 36304 18564 36310
rect 18512 36246 18564 36252
rect 18524 35714 18552 36246
rect 18616 36106 18644 37606
rect 18708 36310 18736 37606
rect 18696 36304 18748 36310
rect 18696 36246 18748 36252
rect 18604 36100 18656 36106
rect 18604 36042 18656 36048
rect 18788 36032 18840 36038
rect 18788 35974 18840 35980
rect 18524 35686 18736 35714
rect 18512 35624 18564 35630
rect 18512 35566 18564 35572
rect 18524 35086 18552 35566
rect 18512 35080 18564 35086
rect 18512 35022 18564 35028
rect 18524 34678 18552 35022
rect 18512 34672 18564 34678
rect 18512 34614 18564 34620
rect 18708 34626 18736 35686
rect 18800 35290 18828 35974
rect 18788 35284 18840 35290
rect 18788 35226 18840 35232
rect 18524 34490 18552 34614
rect 18708 34598 18828 34626
rect 18696 34536 18748 34542
rect 18524 34462 18644 34490
rect 18696 34478 18748 34484
rect 18512 34400 18564 34406
rect 18512 34342 18564 34348
rect 18524 33998 18552 34342
rect 18512 33992 18564 33998
rect 18512 33934 18564 33940
rect 18616 33590 18644 34462
rect 18604 33584 18656 33590
rect 18604 33526 18656 33532
rect 18708 33436 18736 34478
rect 18524 33408 18736 33436
rect 18524 33017 18552 33408
rect 18604 33312 18656 33318
rect 18604 33254 18656 33260
rect 18510 33008 18566 33017
rect 18510 32943 18566 32952
rect 18524 32774 18552 32943
rect 18616 32910 18644 33254
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 18512 32768 18564 32774
rect 18800 32722 18828 34598
rect 18892 32978 18920 37726
rect 19248 37392 19300 37398
rect 19248 37334 19300 37340
rect 19156 36712 19208 36718
rect 19156 36654 19208 36660
rect 19168 35873 19196 36654
rect 19260 36106 19288 37334
rect 19444 36650 19472 38150
rect 19536 37126 19564 38898
rect 19800 38004 19852 38010
rect 19800 37946 19852 37952
rect 19812 37466 19840 37946
rect 19800 37460 19852 37466
rect 19800 37402 19852 37408
rect 19524 37120 19576 37126
rect 19524 37062 19576 37068
rect 19432 36644 19484 36650
rect 19432 36586 19484 36592
rect 19708 36576 19760 36582
rect 19708 36518 19760 36524
rect 19432 36372 19484 36378
rect 19432 36314 19484 36320
rect 19524 36372 19576 36378
rect 19524 36314 19576 36320
rect 19340 36168 19392 36174
rect 19340 36110 19392 36116
rect 19248 36100 19300 36106
rect 19248 36042 19300 36048
rect 19154 35864 19210 35873
rect 19210 35822 19288 35850
rect 19154 35799 19210 35808
rect 19156 35624 19208 35630
rect 19154 35592 19156 35601
rect 19208 35592 19210 35601
rect 19154 35527 19210 35536
rect 19064 34944 19116 34950
rect 19064 34886 19116 34892
rect 19076 34678 19104 34886
rect 19064 34672 19116 34678
rect 19064 34614 19116 34620
rect 18972 33312 19024 33318
rect 18972 33254 19024 33260
rect 18880 32972 18932 32978
rect 18880 32914 18932 32920
rect 18512 32710 18564 32716
rect 18708 32694 18828 32722
rect 18512 32428 18564 32434
rect 18512 32370 18564 32376
rect 18524 32026 18552 32370
rect 18708 32065 18736 32694
rect 18892 32609 18920 32914
rect 18878 32600 18934 32609
rect 18788 32564 18840 32570
rect 18878 32535 18934 32544
rect 18788 32506 18840 32512
rect 18694 32056 18750 32065
rect 18512 32020 18564 32026
rect 18694 31991 18750 32000
rect 18512 31962 18564 31968
rect 18432 31726 18644 31754
rect 18328 30388 18380 30394
rect 18328 30330 18380 30336
rect 18512 30184 18564 30190
rect 18512 30126 18564 30132
rect 18524 30054 18552 30126
rect 18144 30048 18196 30054
rect 18144 29990 18196 29996
rect 18420 30048 18472 30054
rect 18420 29990 18472 29996
rect 18512 30048 18564 30054
rect 18512 29990 18564 29996
rect 18156 29714 18184 29990
rect 18144 29708 18196 29714
rect 18144 29650 18196 29656
rect 18328 29640 18380 29646
rect 18328 29582 18380 29588
rect 18340 29510 18368 29582
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 18326 29336 18382 29345
rect 18326 29271 18382 29280
rect 18144 29028 18196 29034
rect 18144 28970 18196 28976
rect 18052 27872 18104 27878
rect 18052 27814 18104 27820
rect 17592 27668 17644 27674
rect 17592 27610 17644 27616
rect 17684 27668 17736 27674
rect 17684 27610 17736 27616
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17236 26246 17264 26930
rect 17420 26450 17448 26930
rect 17408 26444 17460 26450
rect 17408 26386 17460 26392
rect 17224 26240 17276 26246
rect 17224 26182 17276 26188
rect 17316 25764 17368 25770
rect 17316 25706 17368 25712
rect 17328 25537 17356 25706
rect 17314 25528 17370 25537
rect 17314 25463 17370 25472
rect 17316 25424 17368 25430
rect 17316 25366 17368 25372
rect 17328 25294 17356 25366
rect 17420 25294 17448 26386
rect 17592 26308 17644 26314
rect 17592 26250 17644 26256
rect 17604 25974 17632 26250
rect 17592 25968 17644 25974
rect 17592 25910 17644 25916
rect 17500 25696 17552 25702
rect 17500 25638 17552 25644
rect 18052 25696 18104 25702
rect 18052 25638 18104 25644
rect 17512 25430 17540 25638
rect 17500 25424 17552 25430
rect 17500 25366 17552 25372
rect 18064 25294 18092 25638
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 18052 25288 18104 25294
rect 18052 25230 18104 25236
rect 17776 25152 17828 25158
rect 17776 25094 17828 25100
rect 17788 24750 17816 25094
rect 18064 24954 18092 25230
rect 18052 24948 18104 24954
rect 18052 24890 18104 24896
rect 17776 24744 17828 24750
rect 17696 24704 17776 24732
rect 17592 24404 17644 24410
rect 17420 24364 17592 24392
rect 17420 24070 17448 24364
rect 17592 24346 17644 24352
rect 17498 24304 17554 24313
rect 17498 24239 17554 24248
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17420 23866 17448 24006
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 17236 22574 17264 23598
rect 17408 23248 17460 23254
rect 17408 23190 17460 23196
rect 17420 23050 17448 23190
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17512 22794 17540 24239
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17604 23798 17632 24006
rect 17592 23792 17644 23798
rect 17592 23734 17644 23740
rect 17696 23118 17724 24704
rect 17776 24686 17828 24692
rect 18050 23216 18106 23225
rect 18050 23151 18106 23160
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17684 23112 17736 23118
rect 17684 23054 17736 23060
rect 17420 22766 17540 22794
rect 17604 22778 17632 23054
rect 17592 22772 17644 22778
rect 17224 22568 17276 22574
rect 17224 22510 17276 22516
rect 16960 22066 17172 22094
rect 17420 22094 17448 22766
rect 17592 22714 17644 22720
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 17512 22234 17540 22646
rect 17500 22228 17552 22234
rect 17500 22170 17552 22176
rect 17696 22166 17724 23054
rect 18064 23050 18092 23151
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 17684 22160 17736 22166
rect 17684 22102 17736 22108
rect 17420 22066 17632 22094
rect 16960 17218 16988 22066
rect 17316 21956 17368 21962
rect 17316 21898 17368 21904
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 17224 21480 17276 21486
rect 17224 21422 17276 21428
rect 17144 20942 17172 21422
rect 17236 21010 17264 21422
rect 17224 21004 17276 21010
rect 17224 20946 17276 20952
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17052 20058 17080 20402
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17144 19961 17172 20878
rect 17130 19952 17186 19961
rect 17130 19887 17186 19896
rect 17328 19854 17356 21898
rect 17604 21010 17632 22066
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17316 18896 17368 18902
rect 17316 18838 17368 18844
rect 17328 18698 17356 18838
rect 17316 18692 17368 18698
rect 17316 18634 17368 18640
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17038 17912 17094 17921
rect 17038 17847 17094 17856
rect 17052 17814 17080 17847
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 17328 17678 17356 18022
rect 17316 17672 17368 17678
rect 17038 17640 17094 17649
rect 17316 17614 17368 17620
rect 17038 17575 17040 17584
rect 17092 17575 17094 17584
rect 17040 17546 17092 17552
rect 16960 17190 17080 17218
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16726 16988 16934
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16960 15026 16988 16526
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16960 12986 16988 13194
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16776 12406 16896 12434
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16592 7546 16620 8774
rect 16776 7970 16804 12406
rect 16960 12306 16988 12718
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 17052 10146 17080 17190
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17236 16250 17264 16458
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17144 15366 17172 15982
rect 17328 15366 17356 16050
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17236 15094 17264 15302
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17328 12850 17356 13126
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17328 12306 17356 12786
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 10674 17356 11086
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 16684 7942 16804 7970
rect 16868 10118 17080 10146
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16684 4162 16712 7942
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16776 7274 16804 7822
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16776 6322 16804 7210
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16868 5370 16896 10118
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17052 9722 17080 9998
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16960 8498 16988 8774
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 17052 7970 17080 9318
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 17144 8090 17172 8842
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17052 7942 17172 7970
rect 17236 7954 17264 8366
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17052 5914 17080 6258
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16592 4134 16712 4162
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 16592 3398 16620 4134
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16684 3534 16712 3946
rect 16776 3534 16804 5170
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 14292 3126 14320 3334
rect 15488 3194 15516 3334
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 16776 3058 16804 3470
rect 16960 3058 16988 3878
rect 17052 3738 17080 4082
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 17144 3126 17172 7942
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17328 7342 17356 10610
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17328 5710 17356 6598
rect 17420 6202 17448 12310
rect 17512 9450 17540 12718
rect 17604 12434 17632 20946
rect 17696 20466 17724 22102
rect 18156 21894 18184 28970
rect 18340 28506 18368 29271
rect 18432 28558 18460 29990
rect 18512 29504 18564 29510
rect 18512 29446 18564 29452
rect 18524 29170 18552 29446
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 18616 29102 18644 31726
rect 18800 30394 18828 32506
rect 18880 32224 18932 32230
rect 18880 32166 18932 32172
rect 18892 31260 18920 32166
rect 18984 31754 19012 33254
rect 19076 32434 19104 34614
rect 19156 32768 19208 32774
rect 19156 32710 19208 32716
rect 19168 32434 19196 32710
rect 19064 32428 19116 32434
rect 19064 32370 19116 32376
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 19076 31890 19104 32370
rect 19168 31958 19196 32370
rect 19260 32230 19288 35822
rect 19248 32224 19300 32230
rect 19248 32166 19300 32172
rect 19246 32056 19302 32065
rect 19246 31991 19302 32000
rect 19156 31952 19208 31958
rect 19156 31894 19208 31900
rect 19064 31884 19116 31890
rect 19064 31826 19116 31832
rect 18984 31726 19104 31754
rect 18892 31232 19012 31260
rect 18696 30388 18748 30394
rect 18696 30330 18748 30336
rect 18788 30388 18840 30394
rect 18788 30330 18840 30336
rect 18604 29096 18656 29102
rect 18604 29038 18656 29044
rect 18616 28994 18644 29038
rect 18524 28966 18644 28994
rect 18708 28966 18736 30330
rect 18984 30190 19012 31232
rect 18880 30184 18932 30190
rect 18880 30126 18932 30132
rect 18972 30184 19024 30190
rect 18972 30126 19024 30132
rect 18788 30048 18840 30054
rect 18788 29990 18840 29996
rect 18800 29102 18828 29990
rect 18892 29510 18920 30126
rect 18880 29504 18932 29510
rect 18880 29446 18932 29452
rect 18788 29096 18840 29102
rect 18788 29038 18840 29044
rect 18248 28478 18368 28506
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 18248 27062 18276 28478
rect 18524 27554 18552 28966
rect 18696 28960 18748 28966
rect 18696 28902 18748 28908
rect 18708 27606 18736 28902
rect 18880 27872 18932 27878
rect 18880 27814 18932 27820
rect 18340 27526 18552 27554
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 18236 27056 18288 27062
rect 18236 26998 18288 27004
rect 18248 26897 18276 26998
rect 18234 26888 18290 26897
rect 18234 26823 18290 26832
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 18248 24886 18276 25230
rect 18236 24880 18288 24886
rect 18236 24822 18288 24828
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 17972 21434 18000 21830
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 17880 21418 18000 21434
rect 17868 21412 18000 21418
rect 17920 21406 18000 21412
rect 17868 21354 17920 21360
rect 18064 21146 18092 21490
rect 18156 21350 18184 21490
rect 18248 21434 18276 24822
rect 18340 21962 18368 27526
rect 18420 27464 18472 27470
rect 18420 27406 18472 27412
rect 18696 27464 18748 27470
rect 18696 27406 18748 27412
rect 18432 27130 18460 27406
rect 18420 27124 18472 27130
rect 18420 27066 18472 27072
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18340 21593 18368 21898
rect 18326 21584 18382 21593
rect 18326 21519 18328 21528
rect 18380 21519 18382 21528
rect 18328 21490 18380 21496
rect 18248 21406 18368 21434
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 17960 20936 18012 20942
rect 18064 20924 18092 21082
rect 18156 20942 18184 21286
rect 18012 20896 18092 20924
rect 18144 20936 18196 20942
rect 17960 20878 18012 20884
rect 18144 20878 18196 20884
rect 18340 20856 18368 21406
rect 18248 20828 18368 20856
rect 17684 20460 17736 20466
rect 17684 20402 17736 20408
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17684 19508 17736 19514
rect 17684 19450 17736 19456
rect 17696 18834 17724 19450
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17696 18154 17724 18634
rect 17684 18148 17736 18154
rect 17684 18090 17736 18096
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17788 16046 17816 17682
rect 17972 17066 18000 19654
rect 18248 19378 18276 20828
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18248 17785 18276 19314
rect 18340 18426 18368 19858
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18234 17776 18290 17785
rect 18340 17746 18368 18362
rect 18234 17711 18290 17720
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17788 15570 17816 15982
rect 17972 15978 18000 16390
rect 18156 15994 18184 17070
rect 18248 16794 18276 17070
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18248 16114 18276 16730
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18328 16040 18380 16046
rect 18156 15988 18328 15994
rect 18156 15982 18380 15988
rect 17960 15972 18012 15978
rect 18156 15966 18368 15982
rect 17960 15914 18012 15920
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 18248 15366 18276 15966
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 18340 15162 18368 15370
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17788 12782 17816 13466
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18156 12850 18184 13194
rect 18340 12850 18368 14554
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17880 12442 17908 12718
rect 17868 12436 17920 12442
rect 17604 12406 17724 12434
rect 17696 12306 17724 12406
rect 18156 12434 18184 12786
rect 17868 12378 17920 12384
rect 18064 12406 18184 12434
rect 17880 12306 17908 12378
rect 18064 12306 18092 12406
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17696 10538 17724 12242
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17788 10674 17816 10950
rect 18064 10674 18092 11018
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17592 10532 17644 10538
rect 17592 10474 17644 10480
rect 17684 10532 17736 10538
rect 17684 10474 17736 10480
rect 17604 10062 17632 10474
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17880 9586 17908 10542
rect 18064 10266 18092 10610
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18064 9586 18092 10202
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 17500 9444 17552 9450
rect 17500 9386 17552 9392
rect 17512 8362 17540 9386
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18156 8498 18184 8570
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17592 7880 17644 7886
rect 17696 7834 17724 8366
rect 17866 8256 17922 8265
rect 17866 8191 17922 8200
rect 17880 8022 17908 8191
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17960 7948 18012 7954
rect 18064 7936 18092 8366
rect 18012 7908 18092 7936
rect 18156 7936 18184 8434
rect 18236 7948 18288 7954
rect 18156 7908 18236 7936
rect 17960 7890 18012 7896
rect 18236 7890 18288 7896
rect 17644 7828 17724 7834
rect 17592 7822 17724 7828
rect 17604 7806 17724 7822
rect 17696 6662 17724 7806
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17696 6458 17724 6598
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17420 6174 17540 6202
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17420 5914 17448 6054
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17512 5370 17540 6174
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17236 4826 17264 5170
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17788 4214 17816 7890
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17880 5846 17908 6598
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17880 4622 17908 5306
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17776 4208 17828 4214
rect 17776 4150 17828 4156
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17328 3534 17356 3878
rect 17788 3670 17816 4150
rect 18248 4078 18276 4626
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18328 4004 18380 4010
rect 18328 3946 18380 3952
rect 18340 3738 18368 3946
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 18432 2854 18460 27066
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 18616 26382 18644 26930
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 18708 25498 18736 27406
rect 18786 27160 18842 27169
rect 18786 27095 18842 27104
rect 18800 27062 18828 27095
rect 18788 27056 18840 27062
rect 18788 26998 18840 27004
rect 18696 25492 18748 25498
rect 18696 25434 18748 25440
rect 18604 24948 18656 24954
rect 18604 24890 18656 24896
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18524 20602 18552 20742
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 18524 19854 18552 20538
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18616 14414 18644 24890
rect 18708 22098 18736 25434
rect 18892 24732 18920 27814
rect 18984 27606 19012 30126
rect 19076 30054 19104 31726
rect 19260 30240 19288 31991
rect 19352 30682 19380 36110
rect 19444 35698 19472 36314
rect 19536 36174 19564 36314
rect 19616 36236 19668 36242
rect 19616 36178 19668 36184
rect 19524 36168 19576 36174
rect 19524 36110 19576 36116
rect 19522 36000 19578 36009
rect 19522 35935 19578 35944
rect 19432 35692 19484 35698
rect 19432 35634 19484 35640
rect 19536 35494 19564 35935
rect 19524 35488 19576 35494
rect 19524 35430 19576 35436
rect 19628 35222 19656 36178
rect 19720 35698 19748 36518
rect 19708 35692 19760 35698
rect 19708 35634 19760 35640
rect 19812 35578 19840 37402
rect 19892 36168 19944 36174
rect 19892 36110 19944 36116
rect 19904 35698 19932 36110
rect 19892 35692 19944 35698
rect 19892 35634 19944 35640
rect 19720 35550 19840 35578
rect 19616 35216 19668 35222
rect 19616 35158 19668 35164
rect 19720 35068 19748 35550
rect 19800 35488 19852 35494
rect 19800 35430 19852 35436
rect 19812 35290 19840 35430
rect 19800 35284 19852 35290
rect 19800 35226 19852 35232
rect 19996 35154 20024 44134
rect 20168 43376 20220 43382
rect 20168 43318 20220 43324
rect 20180 39302 20208 43318
rect 20168 39296 20220 39302
rect 20168 39238 20220 39244
rect 20168 38888 20220 38894
rect 20168 38830 20220 38836
rect 20180 38554 20208 38830
rect 20168 38548 20220 38554
rect 20168 38490 20220 38496
rect 20180 38010 20208 38490
rect 20168 38004 20220 38010
rect 20168 37946 20220 37952
rect 20180 37194 20208 37946
rect 20168 37188 20220 37194
rect 20168 37130 20220 37136
rect 20272 36174 20300 46650
rect 20364 45966 20392 46922
rect 20904 46912 20956 46918
rect 20904 46854 20956 46860
rect 20536 46708 20588 46714
rect 20536 46650 20588 46656
rect 20352 45960 20404 45966
rect 20352 45902 20404 45908
rect 20548 45830 20576 46650
rect 20916 46646 20944 46854
rect 20904 46640 20956 46646
rect 20904 46582 20956 46588
rect 21376 46170 21404 46990
rect 22376 46980 22428 46986
rect 22376 46922 22428 46928
rect 22388 46714 22416 46922
rect 23216 46918 23244 47602
rect 24860 47592 24912 47598
rect 24860 47534 24912 47540
rect 23480 47048 23532 47054
rect 23480 46990 23532 46996
rect 24400 47048 24452 47054
rect 24400 46990 24452 46996
rect 22928 46912 22980 46918
rect 22928 46854 22980 46860
rect 23204 46912 23256 46918
rect 23256 46860 23336 46866
rect 23204 46854 23336 46860
rect 22376 46708 22428 46714
rect 22376 46650 22428 46656
rect 22744 46572 22796 46578
rect 22744 46514 22796 46520
rect 22652 46504 22704 46510
rect 22652 46446 22704 46452
rect 22664 46170 22692 46446
rect 21180 46164 21232 46170
rect 21180 46106 21232 46112
rect 21364 46164 21416 46170
rect 21364 46106 21416 46112
rect 22652 46164 22704 46170
rect 22652 46106 22704 46112
rect 20904 45960 20956 45966
rect 20904 45902 20956 45908
rect 20536 45824 20588 45830
rect 20536 45766 20588 45772
rect 20916 45626 20944 45902
rect 20904 45620 20956 45626
rect 20904 45562 20956 45568
rect 20628 45076 20680 45082
rect 20628 45018 20680 45024
rect 20640 44878 20668 45018
rect 20916 45014 20944 45562
rect 21192 45082 21220 46106
rect 22756 46102 22784 46514
rect 22940 46374 22968 46854
rect 23216 46838 23336 46854
rect 23308 46594 23336 46838
rect 23020 46572 23072 46578
rect 23020 46514 23072 46520
rect 23112 46572 23164 46578
rect 23112 46514 23164 46520
rect 23216 46566 23336 46594
rect 23492 46578 23520 46990
rect 23480 46572 23532 46578
rect 22928 46368 22980 46374
rect 22928 46310 22980 46316
rect 23032 46186 23060 46514
rect 22848 46158 23060 46186
rect 22744 46096 22796 46102
rect 22744 46038 22796 46044
rect 22756 45966 22784 46038
rect 22744 45960 22796 45966
rect 22744 45902 22796 45908
rect 22376 45824 22428 45830
rect 22376 45766 22428 45772
rect 22388 45558 22416 45766
rect 22376 45552 22428 45558
rect 22376 45494 22428 45500
rect 21364 45280 21416 45286
rect 21364 45222 21416 45228
rect 21180 45076 21232 45082
rect 21180 45018 21232 45024
rect 20720 45008 20772 45014
rect 20720 44950 20772 44956
rect 20904 45008 20956 45014
rect 20904 44950 20956 44956
rect 21272 45008 21324 45014
rect 21272 44950 21324 44956
rect 20628 44872 20680 44878
rect 20628 44814 20680 44820
rect 20536 44804 20588 44810
rect 20536 44746 20588 44752
rect 20352 44736 20404 44742
rect 20352 44678 20404 44684
rect 20364 44538 20392 44678
rect 20352 44532 20404 44538
rect 20548 44520 20576 44746
rect 20548 44492 20668 44520
rect 20352 44474 20404 44480
rect 20536 44192 20588 44198
rect 20536 44134 20588 44140
rect 20548 43790 20576 44134
rect 20536 43784 20588 43790
rect 20536 43726 20588 43732
rect 20640 43654 20668 44492
rect 20732 44402 20760 44950
rect 21180 44872 21232 44878
rect 21180 44814 21232 44820
rect 21088 44804 21140 44810
rect 21088 44746 21140 44752
rect 21100 44402 21128 44746
rect 20720 44396 20772 44402
rect 20720 44338 20772 44344
rect 21088 44396 21140 44402
rect 21088 44338 21140 44344
rect 20628 43648 20680 43654
rect 20628 43590 20680 43596
rect 20352 43308 20404 43314
rect 20352 43250 20404 43256
rect 20364 42090 20392 43250
rect 21100 43178 21128 44338
rect 21192 43722 21220 44814
rect 21284 43994 21312 44950
rect 21376 44878 21404 45222
rect 22756 45082 22784 45902
rect 22848 45558 22876 46158
rect 23124 46102 23152 46514
rect 23112 46096 23164 46102
rect 23112 46038 23164 46044
rect 23216 45966 23244 46566
rect 23480 46514 23532 46520
rect 23296 46504 23348 46510
rect 23296 46446 23348 46452
rect 23308 46102 23336 46446
rect 23296 46096 23348 46102
rect 23296 46038 23348 46044
rect 23308 45966 23336 46038
rect 23492 46016 23520 46514
rect 23572 46028 23624 46034
rect 23492 45988 23572 46016
rect 23112 45960 23164 45966
rect 23112 45902 23164 45908
rect 23204 45960 23256 45966
rect 23204 45902 23256 45908
rect 23296 45960 23348 45966
rect 23296 45902 23348 45908
rect 22928 45824 22980 45830
rect 22928 45766 22980 45772
rect 22836 45552 22888 45558
rect 22836 45494 22888 45500
rect 22940 45098 22968 45766
rect 22744 45076 22796 45082
rect 22744 45018 22796 45024
rect 22848 45070 22968 45098
rect 22652 44940 22704 44946
rect 22652 44882 22704 44888
rect 21364 44872 21416 44878
rect 21364 44814 21416 44820
rect 21548 44872 21600 44878
rect 21548 44814 21600 44820
rect 22192 44872 22244 44878
rect 22192 44814 22244 44820
rect 22284 44872 22336 44878
rect 22284 44814 22336 44820
rect 22560 44872 22612 44878
rect 22560 44814 22612 44820
rect 21560 44538 21588 44814
rect 21824 44736 21876 44742
rect 21824 44678 21876 44684
rect 21548 44532 21600 44538
rect 21548 44474 21600 44480
rect 21836 44470 21864 44678
rect 21824 44464 21876 44470
rect 21824 44406 21876 44412
rect 22204 44402 22232 44814
rect 22296 44538 22324 44814
rect 22284 44532 22336 44538
rect 22284 44474 22336 44480
rect 22192 44396 22244 44402
rect 22192 44338 22244 44344
rect 22100 44260 22152 44266
rect 22100 44202 22152 44208
rect 21272 43988 21324 43994
rect 21272 43930 21324 43936
rect 21180 43716 21232 43722
rect 21180 43658 21232 43664
rect 21284 43314 21312 43930
rect 21364 43920 21416 43926
rect 21364 43862 21416 43868
rect 21376 43314 21404 43862
rect 22112 43790 22140 44202
rect 22204 43790 22232 44338
rect 22284 44260 22336 44266
rect 22284 44202 22336 44208
rect 22100 43784 22152 43790
rect 22100 43726 22152 43732
rect 22192 43784 22244 43790
rect 22192 43726 22244 43732
rect 21732 43716 21784 43722
rect 21732 43658 21784 43664
rect 21744 43450 21772 43658
rect 21824 43648 21876 43654
rect 21824 43590 21876 43596
rect 21732 43444 21784 43450
rect 21732 43386 21784 43392
rect 21272 43308 21324 43314
rect 21272 43250 21324 43256
rect 21364 43308 21416 43314
rect 21364 43250 21416 43256
rect 21456 43308 21508 43314
rect 21456 43250 21508 43256
rect 21088 43172 21140 43178
rect 21088 43114 21140 43120
rect 20444 42628 20496 42634
rect 20444 42570 20496 42576
rect 20456 42090 20484 42570
rect 21468 42362 21496 43250
rect 21836 43110 21864 43590
rect 22112 43450 22140 43726
rect 22192 43648 22244 43654
rect 22192 43590 22244 43596
rect 22100 43444 22152 43450
rect 22100 43386 22152 43392
rect 21916 43376 21968 43382
rect 21916 43318 21968 43324
rect 21928 43246 21956 43318
rect 22204 43246 22232 43590
rect 22296 43314 22324 44202
rect 22572 43722 22600 44814
rect 22664 44266 22692 44882
rect 22756 44470 22784 45018
rect 22744 44464 22796 44470
rect 22744 44406 22796 44412
rect 22848 44402 22876 45070
rect 23124 44878 23152 45902
rect 23216 44946 23244 45902
rect 23296 45552 23348 45558
rect 23296 45494 23348 45500
rect 23308 44946 23336 45494
rect 23204 44940 23256 44946
rect 23204 44882 23256 44888
rect 23296 44940 23348 44946
rect 23296 44882 23348 44888
rect 23112 44872 23164 44878
rect 23112 44814 23164 44820
rect 23020 44464 23072 44470
rect 23020 44406 23072 44412
rect 22836 44396 22888 44402
rect 22836 44338 22888 44344
rect 22652 44260 22704 44266
rect 22652 44202 22704 44208
rect 22664 43926 22692 44202
rect 22848 43926 22876 44338
rect 23032 43994 23060 44406
rect 23124 43994 23152 44814
rect 23308 44198 23336 44882
rect 23296 44192 23348 44198
rect 23296 44134 23348 44140
rect 23388 44192 23440 44198
rect 23388 44134 23440 44140
rect 23020 43988 23072 43994
rect 23020 43930 23072 43936
rect 23112 43988 23164 43994
rect 23112 43930 23164 43936
rect 22652 43920 22704 43926
rect 22652 43862 22704 43868
rect 22836 43920 22888 43926
rect 22836 43862 22888 43868
rect 22744 43784 22796 43790
rect 22744 43726 22796 43732
rect 22560 43716 22612 43722
rect 22560 43658 22612 43664
rect 22652 43648 22704 43654
rect 22652 43590 22704 43596
rect 22284 43308 22336 43314
rect 22284 43250 22336 43256
rect 22560 43308 22612 43314
rect 22560 43250 22612 43256
rect 21916 43240 21968 43246
rect 21916 43182 21968 43188
rect 22192 43240 22244 43246
rect 22192 43182 22244 43188
rect 21824 43104 21876 43110
rect 21824 43046 21876 43052
rect 22572 42906 22600 43250
rect 22560 42900 22612 42906
rect 22560 42842 22612 42848
rect 22664 42838 22692 43590
rect 22756 43246 22784 43726
rect 22744 43240 22796 43246
rect 22744 43182 22796 43188
rect 22652 42832 22704 42838
rect 22652 42774 22704 42780
rect 23400 42702 23428 44134
rect 23492 43790 23520 45988
rect 23572 45970 23624 45976
rect 24412 45966 24440 46990
rect 24400 45960 24452 45966
rect 24400 45902 24452 45908
rect 24308 43920 24360 43926
rect 24228 43880 24308 43908
rect 24228 43790 24256 43880
rect 24308 43862 24360 43868
rect 23480 43784 23532 43790
rect 23480 43726 23532 43732
rect 24216 43784 24268 43790
rect 24216 43726 24268 43732
rect 23388 42696 23440 42702
rect 23388 42638 23440 42644
rect 21456 42356 21508 42362
rect 21456 42298 21508 42304
rect 20352 42084 20404 42090
rect 20352 42026 20404 42032
rect 20444 42084 20496 42090
rect 20444 42026 20496 42032
rect 21640 42016 21692 42022
rect 21640 41958 21692 41964
rect 21272 41744 21324 41750
rect 21272 41686 21324 41692
rect 20904 41608 20956 41614
rect 20904 41550 20956 41556
rect 20720 41472 20772 41478
rect 20720 41414 20772 41420
rect 20732 41206 20760 41414
rect 20720 41200 20772 41206
rect 20720 41142 20772 41148
rect 20916 40730 20944 41550
rect 20996 40928 21048 40934
rect 20996 40870 21048 40876
rect 20904 40724 20956 40730
rect 20904 40666 20956 40672
rect 20444 40588 20496 40594
rect 20444 40530 20496 40536
rect 20456 40050 20484 40530
rect 20628 40384 20680 40390
rect 20628 40326 20680 40332
rect 20640 40089 20668 40326
rect 20626 40080 20682 40089
rect 20444 40044 20496 40050
rect 20626 40015 20682 40024
rect 20444 39986 20496 39992
rect 20628 38956 20680 38962
rect 20628 38898 20680 38904
rect 20640 38554 20668 38898
rect 20904 38752 20956 38758
rect 20904 38694 20956 38700
rect 20628 38548 20680 38554
rect 20628 38490 20680 38496
rect 20916 38350 20944 38694
rect 20904 38344 20956 38350
rect 20904 38286 20956 38292
rect 20444 37664 20496 37670
rect 20444 37606 20496 37612
rect 20456 37262 20484 37606
rect 20444 37256 20496 37262
rect 20444 37198 20496 37204
rect 20352 36712 20404 36718
rect 20352 36654 20404 36660
rect 20260 36168 20312 36174
rect 20260 36110 20312 36116
rect 20076 35692 20128 35698
rect 20076 35634 20128 35640
rect 20168 35692 20220 35698
rect 20168 35634 20220 35640
rect 19984 35148 20036 35154
rect 19984 35090 20036 35096
rect 19628 35040 19748 35068
rect 19628 32178 19656 35040
rect 19996 35018 20024 35090
rect 19984 35012 20036 35018
rect 19984 34954 20036 34960
rect 20088 34066 20116 35634
rect 20180 35193 20208 35634
rect 20166 35184 20222 35193
rect 20166 35119 20222 35128
rect 19708 34060 19760 34066
rect 19708 34002 19760 34008
rect 20076 34060 20128 34066
rect 20076 34002 20128 34008
rect 19720 32756 19748 34002
rect 20272 32978 20300 36110
rect 20364 35222 20392 36654
rect 20444 36304 20496 36310
rect 20444 36246 20496 36252
rect 20456 35562 20484 36246
rect 20628 36168 20680 36174
rect 20628 36110 20680 36116
rect 20640 35630 20668 36110
rect 20628 35624 20680 35630
rect 20628 35566 20680 35572
rect 20444 35556 20496 35562
rect 20444 35498 20496 35504
rect 20812 35556 20864 35562
rect 20812 35498 20864 35504
rect 20352 35216 20404 35222
rect 20352 35158 20404 35164
rect 20442 35184 20498 35193
rect 20364 34610 20392 35158
rect 20824 35154 20852 35498
rect 20904 35488 20956 35494
rect 20904 35430 20956 35436
rect 20442 35119 20444 35128
rect 20496 35119 20498 35128
rect 20812 35148 20864 35154
rect 20444 35090 20496 35096
rect 20812 35090 20864 35096
rect 20916 35086 20944 35430
rect 20904 35080 20956 35086
rect 20904 35022 20956 35028
rect 20536 34944 20588 34950
rect 20536 34886 20588 34892
rect 20352 34604 20404 34610
rect 20352 34546 20404 34552
rect 20352 33924 20404 33930
rect 20352 33866 20404 33872
rect 20260 32972 20312 32978
rect 20260 32914 20312 32920
rect 19800 32904 19852 32910
rect 19798 32872 19800 32881
rect 19852 32872 19854 32881
rect 19798 32807 19854 32816
rect 19720 32728 19840 32756
rect 19706 32464 19762 32473
rect 19706 32399 19762 32408
rect 19720 32298 19748 32399
rect 19708 32292 19760 32298
rect 19708 32234 19760 32240
rect 19628 32150 19748 32178
rect 19524 31884 19576 31890
rect 19524 31826 19576 31832
rect 19352 30654 19472 30682
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 19352 30394 19380 30534
rect 19340 30388 19392 30394
rect 19340 30330 19392 30336
rect 19168 30212 19288 30240
rect 19064 30048 19116 30054
rect 19064 29990 19116 29996
rect 19168 29492 19196 30212
rect 19340 30184 19392 30190
rect 19444 30172 19472 30654
rect 19536 30172 19564 31826
rect 19392 30161 19472 30172
rect 19392 30152 19486 30161
rect 19392 30144 19430 30152
rect 19340 30126 19392 30132
rect 19248 30116 19300 30122
rect 19430 30087 19486 30096
rect 19527 30144 19564 30172
rect 19248 30058 19300 30064
rect 19076 29464 19196 29492
rect 18972 27600 19024 27606
rect 18972 27542 19024 27548
rect 19076 27130 19104 29464
rect 19260 29306 19288 30058
rect 19340 30048 19392 30054
rect 19338 30016 19340 30025
rect 19527 30036 19555 30144
rect 19392 30016 19394 30025
rect 19527 30008 19564 30036
rect 19338 29951 19394 29960
rect 19338 29880 19394 29889
rect 19338 29815 19394 29824
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 19260 28762 19288 29106
rect 19248 28756 19300 28762
rect 19248 28698 19300 28704
rect 19352 28626 19380 29815
rect 19340 28620 19392 28626
rect 19340 28562 19392 28568
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 19444 28150 19472 28562
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 19536 27946 19564 30008
rect 19720 30002 19748 32150
rect 19628 29974 19748 30002
rect 19524 27940 19576 27946
rect 19524 27882 19576 27888
rect 19340 27872 19392 27878
rect 19340 27814 19392 27820
rect 19154 27296 19210 27305
rect 19154 27231 19210 27240
rect 19064 27124 19116 27130
rect 19064 27066 19116 27072
rect 18972 24744 19024 24750
rect 18892 24704 18972 24732
rect 18972 24686 19024 24692
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 18786 24168 18842 24177
rect 18786 24103 18842 24112
rect 18800 23866 18828 24103
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 18786 23352 18842 23361
rect 18786 23287 18788 23296
rect 18840 23287 18842 23296
rect 18788 23258 18840 23264
rect 18892 22574 18920 24210
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 18880 22568 18932 22574
rect 18880 22510 18932 22516
rect 18800 22234 18828 22510
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 18696 22092 18748 22098
rect 18696 22034 18748 22040
rect 18800 22030 18828 22170
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18708 21078 18736 21830
rect 18892 21434 18920 22510
rect 18800 21406 18920 21434
rect 18696 21072 18748 21078
rect 18696 21014 18748 21020
rect 18800 19922 18828 21406
rect 18984 21010 19012 24686
rect 19076 24313 19104 27066
rect 19168 27033 19196 27231
rect 19154 27024 19210 27033
rect 19154 26959 19210 26968
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19062 24304 19118 24313
rect 19062 24239 19118 24248
rect 19168 24206 19196 24550
rect 19156 24200 19208 24206
rect 19156 24142 19208 24148
rect 19248 23588 19300 23594
rect 19248 23530 19300 23536
rect 19156 22092 19208 22098
rect 19156 22034 19208 22040
rect 19062 21584 19118 21593
rect 19062 21519 19064 21528
rect 19116 21519 19118 21528
rect 19064 21490 19116 21496
rect 18972 21004 19024 21010
rect 18972 20946 19024 20952
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18696 18692 18748 18698
rect 18696 18634 18748 18640
rect 18708 18426 18736 18634
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18880 18148 18932 18154
rect 18880 18090 18932 18096
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18696 17060 18748 17066
rect 18696 17002 18748 17008
rect 18708 14890 18736 17002
rect 18800 15978 18828 17070
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18708 13530 18736 14826
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18892 12782 18920 18090
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18984 12322 19012 20946
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19076 19786 19104 20334
rect 19064 19780 19116 19786
rect 19064 19722 19116 19728
rect 19064 19236 19116 19242
rect 19064 19178 19116 19184
rect 19076 18902 19104 19178
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 19076 17218 19104 18702
rect 19168 18222 19196 22034
rect 19260 21622 19288 23530
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19260 20330 19288 20742
rect 19248 20324 19300 20330
rect 19248 20266 19300 20272
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19260 18290 19288 18566
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 19076 17202 19288 17218
rect 19076 17196 19300 17202
rect 19076 17190 19248 17196
rect 19076 14618 19104 17190
rect 19248 17138 19300 17144
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19168 16454 19196 17070
rect 19352 16454 19380 27814
rect 19536 26296 19564 27882
rect 19628 27878 19656 29974
rect 19708 29844 19760 29850
rect 19708 29786 19760 29792
rect 19616 27872 19668 27878
rect 19616 27814 19668 27820
rect 19720 26790 19748 29786
rect 19812 28694 19840 32728
rect 19892 32360 19944 32366
rect 19892 32302 19944 32308
rect 19984 32360 20036 32366
rect 19984 32302 20036 32308
rect 20168 32360 20220 32366
rect 20168 32302 20220 32308
rect 19904 31872 19932 32302
rect 19996 32026 20024 32302
rect 20180 32201 20208 32302
rect 20364 32230 20392 33866
rect 20352 32224 20404 32230
rect 20166 32192 20222 32201
rect 20352 32166 20404 32172
rect 20166 32127 20222 32136
rect 19984 32020 20036 32026
rect 19984 31962 20036 31968
rect 20260 32020 20312 32026
rect 20260 31962 20312 31968
rect 20352 32020 20404 32026
rect 20352 31962 20404 31968
rect 20272 31890 20300 31962
rect 20168 31884 20220 31890
rect 19904 31844 20168 31872
rect 20168 31826 20220 31832
rect 20260 31884 20312 31890
rect 20260 31826 20312 31832
rect 20166 31648 20222 31657
rect 20166 31583 20222 31592
rect 20180 31346 20208 31583
rect 20258 31512 20314 31521
rect 20258 31447 20314 31456
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 19984 30320 20036 30326
rect 19984 30262 20036 30268
rect 19892 30184 19944 30190
rect 19892 30126 19944 30132
rect 19904 30025 19932 30126
rect 19890 30016 19946 30025
rect 19890 29951 19946 29960
rect 19892 29708 19944 29714
rect 19892 29650 19944 29656
rect 19800 28688 19852 28694
rect 19800 28630 19852 28636
rect 19812 27606 19840 28630
rect 19904 27878 19932 29650
rect 19996 29238 20024 30262
rect 19984 29232 20036 29238
rect 19984 29174 20036 29180
rect 20272 28762 20300 31447
rect 20364 30394 20392 31962
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 20456 31521 20484 31758
rect 20442 31512 20498 31521
rect 20442 31447 20498 31456
rect 20444 31408 20496 31414
rect 20442 31376 20444 31385
rect 20496 31376 20498 31385
rect 20442 31311 20498 31320
rect 20548 30394 20576 34886
rect 21008 33930 21036 40870
rect 21180 38412 21232 38418
rect 21180 38354 21232 38360
rect 21192 37806 21220 38354
rect 21180 37800 21232 37806
rect 21180 37742 21232 37748
rect 21088 35624 21140 35630
rect 21088 35566 21140 35572
rect 20996 33924 21048 33930
rect 20996 33866 21048 33872
rect 20996 33584 21048 33590
rect 20996 33526 21048 33532
rect 21008 32978 21036 33526
rect 20996 32972 21048 32978
rect 20996 32914 21048 32920
rect 20720 32768 20772 32774
rect 20720 32710 20772 32716
rect 20812 32768 20864 32774
rect 20812 32710 20864 32716
rect 20732 32366 20760 32710
rect 20824 32570 20852 32710
rect 20812 32564 20864 32570
rect 20812 32506 20864 32512
rect 20904 32428 20956 32434
rect 20904 32370 20956 32376
rect 20720 32360 20772 32366
rect 20916 32337 20944 32370
rect 20720 32302 20772 32308
rect 20902 32328 20958 32337
rect 20812 32292 20864 32298
rect 20902 32263 20958 32272
rect 20812 32234 20864 32240
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20352 30388 20404 30394
rect 20352 30330 20404 30336
rect 20536 30388 20588 30394
rect 20536 30330 20588 30336
rect 20534 30152 20590 30161
rect 20534 30087 20590 30096
rect 20444 29708 20496 29714
rect 20444 29650 20496 29656
rect 20260 28756 20312 28762
rect 20260 28698 20312 28704
rect 20168 28484 20220 28490
rect 20168 28426 20220 28432
rect 19982 28112 20038 28121
rect 20180 28082 20208 28426
rect 20352 28416 20404 28422
rect 20352 28358 20404 28364
rect 19982 28047 20038 28056
rect 20168 28076 20220 28082
rect 19996 28014 20024 28047
rect 20168 28018 20220 28024
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19892 27872 19944 27878
rect 19890 27840 19892 27849
rect 19944 27840 19946 27849
rect 19890 27775 19946 27784
rect 19800 27600 19852 27606
rect 19800 27542 19852 27548
rect 20364 27402 20392 28358
rect 20352 27396 20404 27402
rect 20352 27338 20404 27344
rect 20168 27328 20220 27334
rect 20168 27270 20220 27276
rect 19708 26784 19760 26790
rect 19708 26726 19760 26732
rect 19616 26308 19668 26314
rect 19536 26268 19616 26296
rect 19616 26250 19668 26256
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19444 24410 19472 24754
rect 19524 24744 19576 24750
rect 19524 24686 19576 24692
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19536 24206 19564 24686
rect 19616 24676 19668 24682
rect 19616 24618 19668 24624
rect 19628 24410 19656 24618
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 19720 24290 19748 26726
rect 19984 26308 20036 26314
rect 19984 26250 20036 26256
rect 19800 25696 19852 25702
rect 19800 25638 19852 25644
rect 19628 24262 19748 24290
rect 19812 24970 19840 25638
rect 19812 24954 19932 24970
rect 19812 24948 19944 24954
rect 19812 24942 19892 24948
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19536 23866 19564 24142
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 19156 16448 19208 16454
rect 19156 16390 19208 16396
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19168 16096 19196 16390
rect 19340 16108 19392 16114
rect 19168 16068 19340 16096
rect 19340 16050 19392 16056
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19352 15162 19380 15506
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19352 15026 19380 15098
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 19076 12434 19104 14554
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 19168 12986 19196 13126
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19076 12406 19196 12434
rect 18984 12306 19104 12322
rect 18984 12300 19116 12306
rect 18984 12294 19064 12300
rect 19064 12242 19116 12248
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18708 11558 18736 12038
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18708 5234 18736 11494
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18892 10674 18920 10746
rect 19076 10674 19104 12242
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18800 9586 18828 10542
rect 18892 9586 18920 10610
rect 19168 9602 19196 12406
rect 19260 12306 19288 13806
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19352 11218 19380 12718
rect 19444 12238 19472 23734
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 19536 17218 19564 23462
rect 19628 21865 19656 24262
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19720 24041 19748 24074
rect 19706 24032 19762 24041
rect 19706 23967 19762 23976
rect 19812 23798 19840 24942
rect 19892 24890 19944 24896
rect 19996 24834 20024 26250
rect 19904 24806 20024 24834
rect 19800 23792 19852 23798
rect 19706 23760 19762 23769
rect 19800 23734 19852 23740
rect 19706 23695 19762 23704
rect 19720 23594 19748 23695
rect 19708 23588 19760 23594
rect 19708 23530 19760 23536
rect 19800 23588 19852 23594
rect 19800 23530 19852 23536
rect 19708 22568 19760 22574
rect 19708 22510 19760 22516
rect 19720 22030 19748 22510
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19614 21856 19670 21865
rect 19614 21791 19670 21800
rect 19628 20777 19656 21791
rect 19614 20768 19670 20777
rect 19614 20703 19670 20712
rect 19812 18834 19840 23530
rect 19904 23338 19932 24806
rect 20180 24732 20208 27270
rect 20352 26512 20404 26518
rect 20350 26480 20352 26489
rect 20404 26480 20406 26489
rect 20350 26415 20406 26424
rect 20456 26330 20484 29650
rect 20548 26450 20576 30087
rect 20732 29850 20760 31282
rect 20824 31142 20852 32234
rect 20904 32224 20956 32230
rect 20904 32166 20956 32172
rect 20812 31136 20864 31142
rect 20812 31078 20864 31084
rect 20916 30716 20944 32166
rect 21008 31754 21036 32914
rect 21100 31958 21128 35566
rect 21180 34060 21232 34066
rect 21180 34002 21232 34008
rect 21088 31952 21140 31958
rect 21088 31894 21140 31900
rect 21192 31822 21220 34002
rect 21284 33998 21312 41686
rect 21652 41002 21680 41958
rect 21824 41608 21876 41614
rect 21824 41550 21876 41556
rect 24308 41608 24360 41614
rect 24308 41550 24360 41556
rect 21732 41064 21784 41070
rect 21732 41006 21784 41012
rect 21640 40996 21692 41002
rect 21640 40938 21692 40944
rect 21652 40526 21680 40938
rect 21640 40520 21692 40526
rect 21640 40462 21692 40468
rect 21744 38962 21772 41006
rect 21836 40730 21864 41550
rect 23940 41540 23992 41546
rect 23940 41482 23992 41488
rect 22100 41472 22152 41478
rect 22100 41414 22152 41420
rect 22112 41206 22140 41414
rect 23952 41274 23980 41482
rect 23940 41268 23992 41274
rect 23940 41210 23992 41216
rect 22100 41200 22152 41206
rect 22100 41142 22152 41148
rect 24216 41200 24268 41206
rect 24216 41142 24268 41148
rect 24032 41132 24084 41138
rect 24032 41074 24084 41080
rect 22008 40928 22060 40934
rect 22008 40870 22060 40876
rect 21824 40724 21876 40730
rect 21824 40666 21876 40672
rect 22020 40526 22048 40870
rect 22560 40724 22612 40730
rect 22560 40666 22612 40672
rect 22468 40588 22520 40594
rect 22468 40530 22520 40536
rect 22008 40520 22060 40526
rect 22480 40497 22508 40530
rect 22008 40462 22060 40468
rect 22466 40488 22522 40497
rect 21732 38956 21784 38962
rect 21732 38898 21784 38904
rect 21456 38548 21508 38554
rect 21456 38490 21508 38496
rect 21468 37942 21496 38490
rect 21916 38208 21968 38214
rect 21916 38150 21968 38156
rect 21456 37936 21508 37942
rect 21456 37878 21508 37884
rect 21928 37806 21956 38150
rect 22020 37942 22048 40462
rect 22572 40458 22600 40666
rect 22466 40423 22522 40432
rect 22560 40452 22612 40458
rect 22560 40394 22612 40400
rect 23020 40452 23072 40458
rect 23020 40394 23072 40400
rect 22284 40384 22336 40390
rect 22284 40326 22336 40332
rect 22296 40118 22324 40326
rect 23032 40186 23060 40394
rect 23572 40384 23624 40390
rect 23572 40326 23624 40332
rect 23020 40180 23072 40186
rect 23020 40122 23072 40128
rect 22284 40112 22336 40118
rect 22284 40054 22336 40060
rect 23204 40044 23256 40050
rect 23204 39986 23256 39992
rect 23216 39642 23244 39986
rect 23204 39636 23256 39642
rect 23204 39578 23256 39584
rect 23584 39438 23612 40326
rect 24044 40186 24072 41074
rect 24228 41002 24256 41142
rect 24320 41070 24348 41550
rect 24492 41472 24544 41478
rect 24492 41414 24544 41420
rect 24400 41132 24452 41138
rect 24400 41074 24452 41080
rect 24308 41064 24360 41070
rect 24308 41006 24360 41012
rect 24216 40996 24268 41002
rect 24216 40938 24268 40944
rect 24320 40594 24348 41006
rect 24308 40588 24360 40594
rect 24308 40530 24360 40536
rect 24032 40180 24084 40186
rect 24032 40122 24084 40128
rect 23572 39432 23624 39438
rect 23572 39374 23624 39380
rect 22100 38956 22152 38962
rect 22100 38898 22152 38904
rect 22008 37936 22060 37942
rect 22008 37878 22060 37884
rect 21916 37800 21968 37806
rect 21916 37742 21968 37748
rect 22112 37738 22140 38898
rect 23204 38752 23256 38758
rect 23204 38694 23256 38700
rect 22928 38480 22980 38486
rect 22928 38422 22980 38428
rect 22744 38412 22796 38418
rect 22744 38354 22796 38360
rect 22192 38344 22244 38350
rect 22192 38286 22244 38292
rect 22376 38344 22428 38350
rect 22376 38286 22428 38292
rect 22466 38312 22522 38321
rect 22100 37732 22152 37738
rect 22100 37674 22152 37680
rect 21456 37324 21508 37330
rect 21456 37266 21508 37272
rect 21468 35630 21496 37266
rect 22204 37262 22232 38286
rect 22388 37670 22416 38286
rect 22466 38247 22522 38256
rect 22480 37738 22508 38247
rect 22756 37874 22784 38354
rect 22744 37868 22796 37874
rect 22744 37810 22796 37816
rect 22836 37800 22888 37806
rect 22836 37742 22888 37748
rect 22468 37732 22520 37738
rect 22468 37674 22520 37680
rect 22376 37664 22428 37670
rect 22376 37606 22428 37612
rect 22480 37262 22508 37674
rect 22848 37330 22876 37742
rect 22836 37324 22888 37330
rect 22836 37266 22888 37272
rect 22192 37256 22244 37262
rect 22192 37198 22244 37204
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 22008 36712 22060 36718
rect 22008 36654 22060 36660
rect 22020 36174 22048 36654
rect 22100 36304 22152 36310
rect 22100 36246 22152 36252
rect 22008 36168 22060 36174
rect 22008 36110 22060 36116
rect 22020 35834 22048 36110
rect 22008 35828 22060 35834
rect 22008 35770 22060 35776
rect 22112 35766 22140 36246
rect 22560 36236 22612 36242
rect 22560 36178 22612 36184
rect 22284 36032 22336 36038
rect 22284 35974 22336 35980
rect 22296 35834 22324 35974
rect 22284 35828 22336 35834
rect 22284 35770 22336 35776
rect 22100 35760 22152 35766
rect 22100 35702 22152 35708
rect 21916 35692 21968 35698
rect 21916 35634 21968 35640
rect 21456 35624 21508 35630
rect 21456 35566 21508 35572
rect 21732 35624 21784 35630
rect 21732 35566 21784 35572
rect 21272 33992 21324 33998
rect 21272 33934 21324 33940
rect 21546 33960 21602 33969
rect 21180 31816 21232 31822
rect 21180 31758 21232 31764
rect 21284 31754 21312 33934
rect 21546 33895 21548 33904
rect 21600 33895 21602 33904
rect 21548 33866 21600 33872
rect 21640 32836 21692 32842
rect 21640 32778 21692 32784
rect 21546 32600 21602 32609
rect 21456 32564 21508 32570
rect 21546 32535 21548 32544
rect 21456 32506 21508 32512
rect 21600 32535 21602 32544
rect 21548 32506 21600 32512
rect 21468 32298 21496 32506
rect 21456 32292 21508 32298
rect 21456 32234 21508 32240
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 21376 32026 21404 32166
rect 21652 32042 21680 32778
rect 21364 32020 21416 32026
rect 21364 31962 21416 31968
rect 21560 32014 21680 32042
rect 21744 32026 21772 35566
rect 21928 35329 21956 35634
rect 22192 35488 22244 35494
rect 22192 35430 22244 35436
rect 21914 35320 21970 35329
rect 21914 35255 21970 35264
rect 21928 35222 21956 35255
rect 21916 35216 21968 35222
rect 21916 35158 21968 35164
rect 21916 33992 21968 33998
rect 21916 33934 21968 33940
rect 21928 33658 21956 33934
rect 21916 33652 21968 33658
rect 21916 33594 21968 33600
rect 21732 32020 21784 32026
rect 21456 31952 21508 31958
rect 21456 31894 21508 31900
rect 21008 31726 21128 31754
rect 21284 31726 21404 31754
rect 20996 31680 21048 31686
rect 20996 31622 21048 31628
rect 21008 30870 21036 31622
rect 21100 31226 21128 31726
rect 21180 31680 21232 31686
rect 21178 31648 21180 31657
rect 21232 31648 21234 31657
rect 21178 31583 21234 31592
rect 21100 31210 21312 31226
rect 21100 31204 21324 31210
rect 21100 31198 21272 31204
rect 21272 31146 21324 31152
rect 21088 31136 21140 31142
rect 21088 31078 21140 31084
rect 21100 30938 21128 31078
rect 21088 30932 21140 30938
rect 21088 30874 21140 30880
rect 20996 30864 21048 30870
rect 20996 30806 21048 30812
rect 20916 30688 21036 30716
rect 20812 30592 20864 30598
rect 20812 30534 20864 30540
rect 20720 29844 20772 29850
rect 20720 29786 20772 29792
rect 20824 29170 20852 30534
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 20916 29646 20944 30194
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 20904 29504 20956 29510
rect 20904 29446 20956 29452
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 20812 28756 20864 28762
rect 20812 28698 20864 28704
rect 20720 28484 20772 28490
rect 20720 28426 20772 28432
rect 20732 28257 20760 28426
rect 20718 28248 20774 28257
rect 20718 28183 20774 28192
rect 20628 28008 20680 28014
rect 20628 27950 20680 27956
rect 20536 26444 20588 26450
rect 20536 26386 20588 26392
rect 19996 24704 20208 24732
rect 20364 26302 20484 26330
rect 19996 23730 20024 24704
rect 20260 24676 20312 24682
rect 20260 24618 20312 24624
rect 20166 24304 20222 24313
rect 20166 24239 20168 24248
rect 20220 24239 20222 24248
rect 20168 24210 20220 24216
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19996 23526 20024 23666
rect 20180 23526 20208 24006
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 19904 23310 20024 23338
rect 19892 22976 19944 22982
rect 19892 22918 19944 22924
rect 19904 22574 19932 22918
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19904 22098 19932 22510
rect 19996 22148 20024 23310
rect 20272 22574 20300 24618
rect 20260 22568 20312 22574
rect 20260 22510 20312 22516
rect 20272 22438 20300 22510
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 20168 22160 20220 22166
rect 19996 22120 20168 22148
rect 20168 22102 20220 22108
rect 19892 22092 19944 22098
rect 19892 22034 19944 22040
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 19904 19922 19932 21490
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19720 17882 19748 18566
rect 19812 18154 19840 18770
rect 19800 18148 19852 18154
rect 19800 18090 19852 18096
rect 19708 17876 19760 17882
rect 19708 17818 19760 17824
rect 19536 17190 19656 17218
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19536 14006 19564 15438
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19076 9586 19196 9602
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 19064 9580 19196 9586
rect 19116 9574 19196 9580
rect 19064 9522 19116 9528
rect 19076 8838 19104 9522
rect 19352 9024 19380 11154
rect 19444 10062 19472 12174
rect 19536 11898 19564 12174
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19352 8996 19472 9024
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18800 7410 18828 7482
rect 18892 7410 18920 8774
rect 19076 8514 19104 8774
rect 18984 8486 19104 8514
rect 18984 8430 19012 8486
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19076 7954 19104 8366
rect 19352 8106 19380 8842
rect 19168 8078 19380 8106
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 19168 7886 19196 8078
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18892 5778 18920 7346
rect 18984 7274 19196 7290
rect 18972 7268 19196 7274
rect 19024 7262 19196 7268
rect 18972 7210 19024 7216
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 19076 6798 19104 7142
rect 19168 6798 19196 7262
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 18984 6610 19012 6666
rect 19156 6656 19208 6662
rect 18984 6604 19156 6610
rect 18984 6598 19208 6604
rect 18984 6582 19196 6598
rect 19352 6118 19380 7890
rect 19444 7342 19472 8996
rect 19628 8974 19656 17190
rect 19904 17134 19932 19858
rect 19996 19718 20024 20402
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 20088 19514 20116 19790
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19996 18222 20024 19246
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19800 16448 19852 16454
rect 19800 16390 19852 16396
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19720 14958 19748 15438
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19720 14074 19748 14894
rect 19812 14550 19840 16390
rect 19800 14544 19852 14550
rect 19800 14486 19852 14492
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19812 13938 19840 14214
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19720 11558 19748 12786
rect 19904 12238 19932 17070
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20088 16726 20116 16934
rect 20076 16720 20128 16726
rect 20076 16662 20128 16668
rect 20180 16114 20208 22102
rect 20364 22094 20392 26302
rect 20548 24834 20576 26386
rect 20640 26382 20668 27950
rect 20824 27878 20852 28698
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 20824 26790 20852 27814
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20812 26512 20864 26518
rect 20810 26480 20812 26489
rect 20864 26480 20866 26489
rect 20810 26415 20866 26424
rect 20628 26376 20680 26382
rect 20628 26318 20680 26324
rect 20718 26208 20774 26217
rect 20718 26143 20774 26152
rect 20732 25974 20760 26143
rect 20720 25968 20772 25974
rect 20720 25910 20772 25916
rect 20812 25968 20864 25974
rect 20812 25910 20864 25916
rect 20824 25362 20852 25910
rect 20812 25356 20864 25362
rect 20812 25298 20864 25304
rect 20548 24806 20668 24834
rect 20444 24744 20496 24750
rect 20444 24686 20496 24692
rect 20536 24744 20588 24750
rect 20536 24686 20588 24692
rect 20456 24206 20484 24686
rect 20548 24274 20576 24686
rect 20536 24268 20588 24274
rect 20536 24210 20588 24216
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20456 23662 20484 24142
rect 20640 23769 20668 24806
rect 20720 24608 20772 24614
rect 20720 24550 20772 24556
rect 20732 24274 20760 24550
rect 20720 24268 20772 24274
rect 20720 24210 20772 24216
rect 20916 23798 20944 29446
rect 21008 28150 21036 30688
rect 21088 30592 21140 30598
rect 21088 30534 21140 30540
rect 21100 30054 21128 30534
rect 21376 30410 21404 31726
rect 21468 31668 21496 31894
rect 21560 31822 21588 32014
rect 21732 31962 21784 31968
rect 21928 31906 21956 33594
rect 22204 33522 22232 35430
rect 22192 33516 22244 33522
rect 22192 33458 22244 33464
rect 22204 32586 22232 33458
rect 22572 32978 22600 36178
rect 22744 35080 22796 35086
rect 22744 35022 22796 35028
rect 22652 34400 22704 34406
rect 22652 34342 22704 34348
rect 22376 32972 22428 32978
rect 22376 32914 22428 32920
rect 22560 32972 22612 32978
rect 22560 32914 22612 32920
rect 22112 32558 22232 32586
rect 22112 32314 22140 32558
rect 22192 32428 22244 32434
rect 22192 32370 22244 32376
rect 22020 32286 22140 32314
rect 22020 32026 22048 32286
rect 22100 32224 22152 32230
rect 22100 32166 22152 32172
rect 22008 32020 22060 32026
rect 22008 31962 22060 31968
rect 21928 31878 22048 31906
rect 21548 31816 21600 31822
rect 21548 31758 21600 31764
rect 21640 31816 21692 31822
rect 21640 31758 21692 31764
rect 21732 31816 21784 31822
rect 21732 31758 21784 31764
rect 21652 31668 21680 31758
rect 21468 31640 21680 31668
rect 21468 30598 21496 31640
rect 21548 31476 21600 31482
rect 21548 31418 21600 31424
rect 21456 30592 21508 30598
rect 21456 30534 21508 30540
rect 21376 30382 21496 30410
rect 21364 30252 21416 30258
rect 21364 30194 21416 30200
rect 21088 30048 21140 30054
rect 21088 29990 21140 29996
rect 21180 30048 21232 30054
rect 21180 29990 21232 29996
rect 21100 29714 21128 29990
rect 21192 29850 21220 29990
rect 21180 29844 21232 29850
rect 21180 29786 21232 29792
rect 21088 29708 21140 29714
rect 21088 29650 21140 29656
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 20996 28144 21048 28150
rect 20996 28086 21048 28092
rect 21192 27010 21220 29582
rect 21272 28552 21324 28558
rect 21272 28494 21324 28500
rect 21284 27130 21312 28494
rect 21272 27124 21324 27130
rect 21272 27066 21324 27072
rect 21008 26982 21220 27010
rect 21376 26994 21404 30194
rect 21468 29714 21496 30382
rect 21456 29708 21508 29714
rect 21456 29650 21508 29656
rect 21456 29572 21508 29578
rect 21456 29514 21508 29520
rect 21468 29034 21496 29514
rect 21456 29028 21508 29034
rect 21456 28970 21508 28976
rect 21560 28506 21588 31418
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 21652 30938 21680 31282
rect 21744 31278 21772 31758
rect 21824 31680 21876 31686
rect 21824 31622 21876 31628
rect 21732 31272 21784 31278
rect 21732 31214 21784 31220
rect 21640 30932 21692 30938
rect 21640 30874 21692 30880
rect 21652 30258 21680 30874
rect 21732 30660 21784 30666
rect 21732 30602 21784 30608
rect 21744 30326 21772 30602
rect 21732 30320 21784 30326
rect 21732 30262 21784 30268
rect 21640 30252 21692 30258
rect 21640 30194 21692 30200
rect 21468 28478 21588 28506
rect 21468 27146 21496 28478
rect 21548 28416 21600 28422
rect 21548 28358 21600 28364
rect 21560 27470 21588 28358
rect 21548 27464 21600 27470
rect 21548 27406 21600 27412
rect 21468 27118 21588 27146
rect 21008 26926 21036 26982
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 21088 26920 21140 26926
rect 21088 26862 21140 26868
rect 20996 26784 21048 26790
rect 20996 26726 21048 26732
rect 20812 23792 20864 23798
rect 20626 23760 20682 23769
rect 20626 23695 20682 23704
rect 20810 23760 20812 23769
rect 20904 23792 20956 23798
rect 20864 23760 20866 23769
rect 20904 23734 20956 23740
rect 20810 23695 20866 23704
rect 20444 23656 20496 23662
rect 20444 23598 20496 23604
rect 20628 23588 20680 23594
rect 20628 23530 20680 23536
rect 20640 23361 20668 23530
rect 20626 23352 20682 23361
rect 20626 23287 20682 23296
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20732 22574 20760 22714
rect 20628 22568 20680 22574
rect 20628 22510 20680 22516
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20904 22568 20956 22574
rect 20904 22510 20956 22516
rect 20640 22098 20668 22510
rect 20732 22098 20760 22510
rect 20364 22066 20484 22094
rect 20260 20528 20312 20534
rect 20260 20470 20312 20476
rect 20272 18766 20300 20470
rect 20456 20466 20484 22066
rect 20628 22092 20680 22098
rect 20628 22034 20680 22040
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 21146 20852 21286
rect 20916 21146 20944 22510
rect 21008 22094 21036 26726
rect 21100 23730 21128 26862
rect 21192 26382 21220 26982
rect 21364 26988 21416 26994
rect 21364 26930 21416 26936
rect 21456 26988 21508 26994
rect 21456 26930 21508 26936
rect 21180 26376 21232 26382
rect 21468 26353 21496 26930
rect 21180 26318 21232 26324
rect 21454 26344 21510 26353
rect 21454 26279 21510 26288
rect 21560 25514 21588 27118
rect 21652 26976 21680 30194
rect 21836 28994 21864 31622
rect 22020 31464 22048 31878
rect 22112 31822 22140 32166
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 22020 31436 22140 31464
rect 22112 30818 22140 31436
rect 22204 31210 22232 32370
rect 22282 32192 22338 32201
rect 22282 32127 22338 32136
rect 22296 31482 22324 32127
rect 22388 31822 22416 32914
rect 22468 32836 22520 32842
rect 22468 32778 22520 32784
rect 22480 32230 22508 32778
rect 22468 32224 22520 32230
rect 22468 32166 22520 32172
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22376 31680 22428 31686
rect 22376 31622 22428 31628
rect 22388 31482 22416 31622
rect 22480 31482 22508 32166
rect 22664 31754 22692 34342
rect 22756 33862 22784 35022
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22756 32502 22784 33798
rect 22940 32994 22968 38422
rect 23216 38350 23244 38694
rect 23204 38344 23256 38350
rect 23204 38286 23256 38292
rect 23020 38208 23072 38214
rect 23020 38150 23072 38156
rect 23112 38208 23164 38214
rect 23112 38150 23164 38156
rect 23032 36310 23060 38150
rect 23124 38010 23152 38150
rect 23112 38004 23164 38010
rect 23112 37946 23164 37952
rect 23204 37800 23256 37806
rect 23204 37742 23256 37748
rect 23216 37466 23244 37742
rect 23584 37738 23612 39374
rect 23664 39296 23716 39302
rect 23664 39238 23716 39244
rect 23676 38894 23704 39238
rect 23664 38888 23716 38894
rect 23664 38830 23716 38836
rect 23676 38418 23704 38830
rect 24124 38752 24176 38758
rect 24124 38694 24176 38700
rect 23664 38412 23716 38418
rect 23664 38354 23716 38360
rect 23848 38412 23900 38418
rect 23848 38354 23900 38360
rect 23572 37732 23624 37738
rect 23572 37674 23624 37680
rect 23664 37664 23716 37670
rect 23664 37606 23716 37612
rect 23204 37460 23256 37466
rect 23204 37402 23256 37408
rect 23020 36304 23072 36310
rect 23020 36246 23072 36252
rect 23216 36242 23244 37402
rect 23676 36310 23704 37606
rect 23756 37120 23808 37126
rect 23756 37062 23808 37068
rect 23768 36786 23796 37062
rect 23756 36780 23808 36786
rect 23756 36722 23808 36728
rect 23664 36304 23716 36310
rect 23664 36246 23716 36252
rect 23204 36236 23256 36242
rect 23204 36178 23256 36184
rect 23388 36100 23440 36106
rect 23388 36042 23440 36048
rect 23296 35080 23348 35086
rect 23296 35022 23348 35028
rect 23020 34944 23072 34950
rect 23018 34912 23020 34921
rect 23072 34912 23074 34921
rect 23018 34847 23074 34856
rect 23308 34746 23336 35022
rect 23296 34740 23348 34746
rect 23296 34682 23348 34688
rect 23400 34626 23428 36042
rect 23480 36032 23532 36038
rect 23480 35974 23532 35980
rect 23492 35290 23520 35974
rect 23768 35766 23796 36722
rect 23860 35873 23888 38354
rect 24136 38350 24164 38694
rect 24320 38418 24348 40530
rect 24412 40186 24440 41074
rect 24400 40180 24452 40186
rect 24400 40122 24452 40128
rect 24504 40118 24532 41414
rect 24492 40112 24544 40118
rect 24492 40054 24544 40060
rect 24676 40112 24728 40118
rect 24676 40054 24728 40060
rect 24308 38412 24360 38418
rect 24308 38354 24360 38360
rect 24124 38344 24176 38350
rect 24124 38286 24176 38292
rect 24504 37874 24532 40054
rect 24492 37868 24544 37874
rect 24492 37810 24544 37816
rect 24504 37330 24532 37810
rect 24584 37800 24636 37806
rect 24584 37742 24636 37748
rect 24596 37330 24624 37742
rect 24492 37324 24544 37330
rect 24492 37266 24544 37272
rect 24584 37324 24636 37330
rect 24584 37266 24636 37272
rect 24124 37256 24176 37262
rect 24124 37198 24176 37204
rect 23846 35864 23902 35873
rect 23846 35799 23902 35808
rect 23756 35760 23808 35766
rect 23756 35702 23808 35708
rect 23860 35630 23888 35799
rect 23848 35624 23900 35630
rect 23848 35566 23900 35572
rect 23480 35284 23532 35290
rect 23480 35226 23532 35232
rect 23308 34610 23428 34626
rect 23296 34604 23428 34610
rect 23348 34598 23428 34604
rect 23296 34546 23348 34552
rect 23112 33516 23164 33522
rect 23112 33458 23164 33464
rect 23124 33114 23152 33458
rect 23112 33108 23164 33114
rect 23112 33050 23164 33056
rect 22940 32966 23060 32994
rect 22928 32836 22980 32842
rect 22848 32796 22928 32824
rect 22744 32496 22796 32502
rect 22744 32438 22796 32444
rect 22572 31726 22692 31754
rect 22284 31476 22336 31482
rect 22284 31418 22336 31424
rect 22376 31476 22428 31482
rect 22376 31418 22428 31424
rect 22468 31476 22520 31482
rect 22468 31418 22520 31424
rect 22376 31272 22428 31278
rect 22376 31214 22428 31220
rect 22192 31204 22244 31210
rect 22192 31146 22244 31152
rect 22020 30790 22140 30818
rect 21916 30728 21968 30734
rect 21916 30670 21968 30676
rect 21928 30394 21956 30670
rect 21916 30388 21968 30394
rect 21916 30330 21968 30336
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 21928 29646 21956 30194
rect 21916 29640 21968 29646
rect 21916 29582 21968 29588
rect 21836 28966 21956 28994
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21732 28416 21784 28422
rect 21732 28358 21784 28364
rect 21744 28218 21772 28358
rect 21836 28218 21864 28494
rect 21732 28212 21784 28218
rect 21732 28154 21784 28160
rect 21824 28212 21876 28218
rect 21824 28154 21876 28160
rect 21732 26988 21784 26994
rect 21652 26948 21732 26976
rect 21732 26930 21784 26936
rect 21468 25486 21588 25514
rect 21270 25392 21326 25401
rect 21192 25336 21270 25344
rect 21192 25316 21272 25336
rect 21088 23724 21140 23730
rect 21088 23666 21140 23672
rect 21088 22094 21140 22098
rect 21008 22092 21140 22094
rect 21008 22066 21088 22092
rect 21088 22034 21140 22040
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20904 21140 20956 21146
rect 20904 21082 20956 21088
rect 21100 21026 21128 22034
rect 20824 20998 21128 21026
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20628 20800 20680 20806
rect 20534 20768 20590 20777
rect 20628 20742 20680 20748
rect 20534 20703 20590 20712
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20352 18964 20404 18970
rect 20352 18906 20404 18912
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 20364 18698 20392 18906
rect 20456 18766 20484 20402
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 20272 16590 20300 18362
rect 20456 17814 20484 18566
rect 20444 17808 20496 17814
rect 20444 17750 20496 17756
rect 20548 17626 20576 20703
rect 20456 17598 20576 17626
rect 20352 17264 20404 17270
rect 20352 17206 20404 17212
rect 20364 16794 20392 17206
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20350 16552 20406 16561
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20180 15994 20208 16050
rect 19996 15966 20208 15994
rect 19996 15910 20024 15966
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20088 15026 20116 15506
rect 20272 15162 20300 16526
rect 20350 16487 20406 16496
rect 20364 15638 20392 16487
rect 20456 15858 20484 17598
rect 20640 16674 20668 20742
rect 20732 20262 20760 20878
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20732 19718 20760 19790
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20548 16646 20668 16674
rect 20548 16590 20576 16646
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20548 16046 20576 16526
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20456 15830 20668 15858
rect 20352 15632 20404 15638
rect 20352 15574 20404 15580
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20088 13326 20116 14350
rect 20272 14056 20300 15098
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20364 14618 20392 14962
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20548 14385 20576 14486
rect 20534 14376 20590 14385
rect 20444 14340 20496 14346
rect 20534 14311 20590 14320
rect 20444 14282 20496 14288
rect 20180 14028 20300 14056
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20180 12918 20208 14028
rect 20456 14006 20484 14282
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20272 13530 20300 13874
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20548 13138 20576 14311
rect 20640 13258 20668 15830
rect 20732 15722 20760 19654
rect 20824 15910 20852 20998
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21008 19786 21036 20878
rect 21192 19922 21220 25316
rect 21324 25327 21326 25336
rect 21272 25298 21324 25304
rect 21272 24880 21324 24886
rect 21272 24822 21324 24828
rect 21284 24041 21312 24822
rect 21468 24750 21496 25486
rect 21548 25424 21600 25430
rect 21548 25366 21600 25372
rect 21456 24744 21508 24750
rect 21376 24704 21456 24732
rect 21270 24032 21326 24041
rect 21270 23967 21326 23976
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 21284 23633 21312 23666
rect 21270 23624 21326 23633
rect 21270 23559 21326 23568
rect 21272 22568 21324 22574
rect 21376 22522 21404 24704
rect 21456 24686 21508 24692
rect 21560 24410 21588 25366
rect 21548 24404 21600 24410
rect 21548 24346 21600 24352
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21456 23792 21508 23798
rect 21454 23760 21456 23769
rect 21508 23760 21510 23769
rect 21652 23730 21680 24074
rect 21454 23695 21510 23704
rect 21640 23724 21692 23730
rect 21640 23666 21692 23672
rect 21456 23656 21508 23662
rect 21456 23598 21508 23604
rect 21324 22516 21404 22522
rect 21272 22510 21404 22516
rect 21284 22494 21404 22510
rect 21272 22092 21324 22098
rect 21468 22094 21496 23598
rect 21548 23248 21600 23254
rect 21548 23190 21600 23196
rect 21560 22778 21588 23190
rect 21652 23186 21680 23666
rect 21640 23180 21692 23186
rect 21640 23122 21692 23128
rect 21548 22772 21600 22778
rect 21548 22714 21600 22720
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21272 22034 21324 22040
rect 21376 22066 21496 22094
rect 21284 20534 21312 22034
rect 21272 20528 21324 20534
rect 21272 20470 21324 20476
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 21178 19816 21234 19825
rect 20996 19780 21048 19786
rect 21178 19751 21234 19760
rect 20996 19722 21048 19728
rect 21192 19718 21220 19751
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 20994 19000 21050 19009
rect 20994 18935 21050 18944
rect 21008 18834 21036 18935
rect 21192 18902 21220 19110
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 21180 18896 21232 18902
rect 21180 18838 21232 18844
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 21008 16590 21036 16934
rect 20996 16584 21048 16590
rect 20902 16552 20958 16561
rect 20996 16526 21048 16532
rect 20902 16487 20958 16496
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20732 15694 20852 15722
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20732 14958 20760 15438
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20824 14346 20852 15694
rect 20916 15570 20944 16487
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 21008 15026 21036 16186
rect 21100 16182 21128 18838
rect 21192 16998 21220 18838
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 21284 17338 21312 17818
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 16250 21220 16390
rect 21284 16250 21312 16458
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21088 16176 21140 16182
rect 21088 16118 21140 16124
rect 21376 16114 21404 22066
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21468 20466 21496 21490
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21468 19174 21496 20402
rect 21456 19168 21508 19174
rect 21456 19110 21508 19116
rect 21560 18850 21588 22510
rect 21744 22012 21772 26930
rect 21928 24698 21956 28966
rect 22020 26042 22048 30790
rect 22284 29504 22336 29510
rect 22284 29446 22336 29452
rect 22192 28688 22244 28694
rect 22192 28630 22244 28636
rect 22204 28540 22232 28630
rect 22112 28512 22232 28540
rect 22112 27878 22140 28512
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 22100 27872 22152 27878
rect 22100 27814 22152 27820
rect 22204 27554 22232 28086
rect 22112 27526 22232 27554
rect 22112 27470 22140 27526
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 22204 26994 22232 27270
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 22008 26036 22060 26042
rect 22008 25978 22060 25984
rect 22020 25838 22048 25978
rect 22008 25832 22060 25838
rect 22008 25774 22060 25780
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 22112 24750 22140 25230
rect 21836 24670 21956 24698
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 21836 22166 21864 24670
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21928 24342 21956 24550
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 21916 23656 21968 23662
rect 21916 23598 21968 23604
rect 21824 22160 21876 22166
rect 21824 22102 21876 22108
rect 21652 21984 21772 22012
rect 21652 21554 21680 21984
rect 21640 21548 21692 21554
rect 21640 21490 21692 21496
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21560 18822 21772 18850
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21652 18358 21680 18702
rect 21640 18352 21692 18358
rect 21640 18294 21692 18300
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21284 15570 21312 16050
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 21376 13530 21404 16050
rect 21468 15706 21496 16050
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 20916 13326 20944 13466
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 20548 13110 20668 13138
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19720 9654 19748 11222
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19812 9654 19840 11154
rect 19904 10606 19932 12174
rect 20180 11218 20208 12854
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20364 12442 20392 12582
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19892 10600 19944 10606
rect 19892 10542 19944 10548
rect 20088 10266 20116 10610
rect 20272 10266 20300 10950
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20180 10118 20484 10146
rect 20548 10130 20576 10406
rect 20076 9988 20128 9994
rect 20076 9930 20128 9936
rect 20088 9897 20116 9930
rect 20180 9926 20208 10118
rect 20456 10062 20484 10118
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20168 9920 20220 9926
rect 20074 9888 20130 9897
rect 20168 9862 20220 9868
rect 20074 9823 20130 9832
rect 20364 9722 20392 9998
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 20352 9716 20404 9722
rect 20352 9658 20404 9664
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19800 9648 19852 9654
rect 19800 9590 19852 9596
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19706 8392 19762 8401
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19536 7954 19564 8298
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19536 7410 19564 7890
rect 19628 7886 19656 8366
rect 19706 8327 19708 8336
rect 19760 8327 19762 8336
rect 19708 8298 19760 8304
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19628 7478 19656 7686
rect 19616 7472 19668 7478
rect 19616 7414 19668 7420
rect 19708 7472 19760 7478
rect 19708 7414 19760 7420
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19444 7002 19472 7278
rect 19536 7002 19564 7346
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19260 5930 19288 6054
rect 19260 5902 19380 5930
rect 19720 5914 19748 7414
rect 19352 5778 19380 5902
rect 19708 5908 19760 5914
rect 19708 5850 19760 5856
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 18788 5296 18840 5302
rect 18788 5238 18840 5244
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 18616 4146 18644 4422
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18602 3632 18658 3641
rect 18800 3602 18828 5238
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19260 4622 19288 4966
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19260 4214 19288 4558
rect 19248 4208 19300 4214
rect 19248 4150 19300 4156
rect 19352 3942 19380 5714
rect 19812 4554 19840 9454
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19904 7954 19932 9318
rect 20088 8634 20116 9386
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20076 8424 20128 8430
rect 19996 8384 20076 8412
rect 19996 8022 20024 8384
rect 20076 8366 20128 8372
rect 20168 8288 20220 8294
rect 20168 8230 20220 8236
rect 19984 8016 20036 8022
rect 19984 7958 20036 7964
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 20180 7886 20208 8230
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20272 7698 20300 9658
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20180 7670 20300 7698
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19904 6662 19932 7346
rect 20180 7342 20208 7670
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 20364 6390 20392 8910
rect 20640 8906 20668 13110
rect 20916 12850 20944 13262
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 21100 12617 21128 13126
rect 21192 12850 21220 13262
rect 21652 13258 21680 16934
rect 21744 14958 21772 18822
rect 21836 16522 21864 21490
rect 21928 18834 21956 23598
rect 22008 23180 22060 23186
rect 22008 23122 22060 23128
rect 22020 22982 22048 23122
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 22008 22500 22060 22506
rect 22008 22442 22060 22448
rect 22020 22166 22048 22442
rect 22008 22160 22060 22166
rect 22008 22102 22060 22108
rect 22112 21486 22140 24686
rect 22296 24585 22324 29446
rect 22388 28626 22416 31214
rect 22480 30802 22508 31418
rect 22468 30796 22520 30802
rect 22468 30738 22520 30744
rect 22468 30184 22520 30190
rect 22468 30126 22520 30132
rect 22480 29646 22508 30126
rect 22468 29640 22520 29646
rect 22468 29582 22520 29588
rect 22572 29510 22600 31726
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22560 29504 22612 29510
rect 22560 29446 22612 29452
rect 22376 28620 22428 28626
rect 22376 28562 22428 28568
rect 22388 26926 22416 28562
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22468 28008 22520 28014
rect 22468 27950 22520 27956
rect 22480 27674 22508 27950
rect 22468 27668 22520 27674
rect 22468 27610 22520 27616
rect 22468 27328 22520 27334
rect 22468 27270 22520 27276
rect 22480 27062 22508 27270
rect 22468 27056 22520 27062
rect 22468 26998 22520 27004
rect 22376 26920 22428 26926
rect 22376 26862 22428 26868
rect 22480 26858 22508 26998
rect 22468 26852 22520 26858
rect 22468 26794 22520 26800
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22282 24576 22338 24585
rect 22282 24511 22338 24520
rect 22296 24018 22324 24511
rect 22388 24410 22416 24754
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22376 24404 22428 24410
rect 22376 24346 22428 24352
rect 22376 24200 22428 24206
rect 22480 24188 22508 24550
rect 22428 24160 22508 24188
rect 22376 24142 22428 24148
rect 22296 23990 22416 24018
rect 22100 21480 22152 21486
rect 22192 21480 22244 21486
rect 22100 21422 22152 21428
rect 22190 21448 22192 21457
rect 22244 21448 22246 21457
rect 22190 21383 22246 21392
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22296 20942 22324 21286
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 21836 16114 21864 16458
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21928 15502 21956 18770
rect 22112 18290 22140 19110
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22020 18193 22048 18226
rect 22006 18184 22062 18193
rect 22006 18119 22062 18128
rect 22284 18148 22336 18154
rect 22284 18090 22336 18096
rect 22008 15904 22060 15910
rect 22008 15846 22060 15852
rect 22020 15638 22048 15846
rect 22008 15632 22060 15638
rect 22008 15574 22060 15580
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 21732 14952 21784 14958
rect 21784 14900 21864 14906
rect 21732 14894 21864 14900
rect 21744 14878 21864 14894
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21744 13394 21772 14214
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 21640 13252 21692 13258
rect 21640 13194 21692 13200
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21086 12608 21142 12617
rect 21086 12543 21142 12552
rect 20718 12200 20774 12209
rect 20718 12135 20774 12144
rect 20732 12102 20760 12135
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20456 7954 20484 8774
rect 20640 8430 20668 8842
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20732 7546 20760 12038
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 20810 11248 20866 11257
rect 20810 11183 20866 11192
rect 20824 10810 20852 11183
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20352 6384 20404 6390
rect 20352 6326 20404 6332
rect 20364 4690 20392 6326
rect 20352 4684 20404 4690
rect 20352 4626 20404 4632
rect 19800 4548 19852 4554
rect 19800 4490 19852 4496
rect 19812 4282 19840 4490
rect 19800 4276 19852 4282
rect 19800 4218 19852 4224
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 18602 3567 18658 3576
rect 18788 3596 18840 3602
rect 18616 3534 18644 3567
rect 18788 3538 18840 3544
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 18708 3194 18736 3334
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 13648 2746 13768 2774
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 940 2304 992 2310
rect 940 2246 992 2252
rect 952 2145 980 2246
rect 938 2136 994 2145
rect 938 2071 994 2080
rect 1964 800 1992 2382
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4540 800 4568 2246
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 6472 800 6500 2382
rect 9048 800 9076 2382
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 800 11652 2246
rect 13556 800 13584 2382
rect 13648 2310 13676 2746
rect 18708 2446 18736 3130
rect 19352 3058 19380 3878
rect 20626 3632 20682 3641
rect 20626 3567 20628 3576
rect 20680 3567 20682 3576
rect 20628 3538 20680 3544
rect 19800 3392 19852 3398
rect 19800 3334 19852 3340
rect 19812 3058 19840 3334
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 20824 2774 20852 10746
rect 21284 10470 21312 11834
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21652 10169 21680 13194
rect 21638 10160 21694 10169
rect 21088 10124 21140 10130
rect 21638 10095 21694 10104
rect 21088 10066 21140 10072
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 20904 9104 20956 9110
rect 20904 9046 20956 9052
rect 20916 8634 20944 9046
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 21008 7546 21036 9998
rect 21100 9586 21128 10066
rect 21652 10062 21680 10095
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21456 9920 21508 9926
rect 21548 9920 21600 9926
rect 21456 9862 21508 9868
rect 21546 9888 21548 9897
rect 21600 9888 21602 9897
rect 21178 9752 21234 9761
rect 21178 9687 21234 9696
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 21100 8090 21128 9386
rect 21192 8090 21220 9687
rect 21468 9586 21496 9862
rect 21546 9823 21602 9832
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 21836 9042 21864 14878
rect 21928 13326 21956 15438
rect 22296 14482 22324 18090
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 22112 14074 22140 14214
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 22008 12164 22060 12170
rect 22008 12106 22060 12112
rect 22020 11898 22048 12106
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 22020 9926 22048 10474
rect 22190 10160 22246 10169
rect 22388 10130 22416 23990
rect 22572 23066 22600 28494
rect 22480 23038 22600 23066
rect 22480 22574 22508 23038
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22572 22710 22600 22918
rect 22560 22704 22612 22710
rect 22560 22646 22612 22652
rect 22468 22568 22520 22574
rect 22468 22510 22520 22516
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22480 21962 22508 22374
rect 22468 21956 22520 21962
rect 22468 21898 22520 21904
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22468 21412 22520 21418
rect 22468 21354 22520 21360
rect 22480 21146 22508 21354
rect 22572 21350 22600 21490
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22468 21140 22520 21146
rect 22468 21082 22520 21088
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22468 18692 22520 18698
rect 22468 18634 22520 18640
rect 22480 18426 22508 18634
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22466 18184 22522 18193
rect 22466 18119 22468 18128
rect 22520 18119 22522 18128
rect 22468 18090 22520 18096
rect 22572 17202 22600 18702
rect 22664 17338 22692 29582
rect 22756 28994 22784 32438
rect 22848 31958 22876 32796
rect 22928 32778 22980 32784
rect 23032 32722 23060 32966
rect 23112 32972 23164 32978
rect 23112 32914 23164 32920
rect 22940 32694 23060 32722
rect 22836 31952 22888 31958
rect 22836 31894 22888 31900
rect 22848 30802 22876 31894
rect 22940 31142 22968 32694
rect 22928 31136 22980 31142
rect 22928 31078 22980 31084
rect 22836 30796 22888 30802
rect 22836 30738 22888 30744
rect 22756 28966 23060 28994
rect 22928 28484 22980 28490
rect 22928 28426 22980 28432
rect 22744 28076 22796 28082
rect 22744 28018 22796 28024
rect 22756 27334 22784 28018
rect 22940 28014 22968 28426
rect 22928 28008 22980 28014
rect 22928 27950 22980 27956
rect 22836 27940 22888 27946
rect 22836 27882 22888 27888
rect 22848 27470 22876 27882
rect 22836 27464 22888 27470
rect 22836 27406 22888 27412
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22940 26926 22968 27950
rect 22928 26920 22980 26926
rect 22928 26862 22980 26868
rect 22928 26308 22980 26314
rect 22928 26250 22980 26256
rect 22836 25832 22888 25838
rect 22836 25774 22888 25780
rect 22848 24342 22876 25774
rect 22836 24336 22888 24342
rect 22836 24278 22888 24284
rect 22744 23112 22796 23118
rect 22744 23054 22796 23060
rect 22756 22778 22784 23054
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 22940 22574 22968 26250
rect 23032 25906 23060 28966
rect 23124 28082 23152 32914
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 23216 31793 23244 31962
rect 23202 31784 23258 31793
rect 23202 31719 23258 31728
rect 23308 28558 23336 34546
rect 23664 34536 23716 34542
rect 23664 34478 23716 34484
rect 23572 34468 23624 34474
rect 23572 34410 23624 34416
rect 23584 34066 23612 34410
rect 23572 34060 23624 34066
rect 23572 34002 23624 34008
rect 23676 33658 23704 34478
rect 23664 33652 23716 33658
rect 23664 33594 23716 33600
rect 23480 33584 23532 33590
rect 23480 33526 23532 33532
rect 23492 29646 23520 33526
rect 23572 31272 23624 31278
rect 23572 31214 23624 31220
rect 23756 31272 23808 31278
rect 23756 31214 23808 31220
rect 23584 30258 23612 31214
rect 23664 31204 23716 31210
rect 23664 31146 23716 31152
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23112 28076 23164 28082
rect 23112 28018 23164 28024
rect 23388 28008 23440 28014
rect 23388 27950 23440 27956
rect 23204 27668 23256 27674
rect 23204 27610 23256 27616
rect 23110 27432 23166 27441
rect 23216 27402 23244 27610
rect 23400 27538 23428 27950
rect 23388 27532 23440 27538
rect 23388 27474 23440 27480
rect 23110 27367 23112 27376
rect 23164 27367 23166 27376
rect 23204 27396 23256 27402
rect 23112 27338 23164 27344
rect 23204 27338 23256 27344
rect 23296 26988 23348 26994
rect 23400 26976 23428 27474
rect 23348 26948 23428 26976
rect 23296 26930 23348 26936
rect 23572 26852 23624 26858
rect 23572 26794 23624 26800
rect 23480 26444 23532 26450
rect 23480 26386 23532 26392
rect 23112 26036 23164 26042
rect 23112 25978 23164 25984
rect 23020 25900 23072 25906
rect 23020 25842 23072 25848
rect 23124 25294 23152 25978
rect 23492 25922 23520 26386
rect 23400 25906 23520 25922
rect 23296 25900 23348 25906
rect 23296 25842 23348 25848
rect 23388 25900 23520 25906
rect 23440 25894 23520 25900
rect 23388 25842 23440 25848
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23110 24712 23166 24721
rect 23110 24647 23166 24656
rect 23124 24614 23152 24647
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 23124 23866 23152 24346
rect 23204 24200 23256 24206
rect 23202 24168 23204 24177
rect 23256 24168 23258 24177
rect 23202 24103 23258 24112
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23216 23866 23244 24006
rect 23112 23860 23164 23866
rect 23112 23802 23164 23808
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 23202 23352 23258 23361
rect 23202 23287 23258 23296
rect 23216 23186 23244 23287
rect 23204 23180 23256 23186
rect 23204 23122 23256 23128
rect 22744 22568 22796 22574
rect 22744 22510 22796 22516
rect 22928 22568 22980 22574
rect 22928 22510 22980 22516
rect 22756 21418 22784 22510
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 22744 21412 22796 21418
rect 22744 21354 22796 21360
rect 22848 19922 22876 21966
rect 22928 21548 22980 21554
rect 22928 21490 22980 21496
rect 22940 21146 22968 21490
rect 22928 21140 22980 21146
rect 22928 21082 22980 21088
rect 23308 20806 23336 25842
rect 23388 25696 23440 25702
rect 23388 25638 23440 25644
rect 23400 25294 23428 25638
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23400 23118 23428 24210
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 23400 20482 23428 23054
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23492 22234 23520 22578
rect 23480 22228 23532 22234
rect 23480 22170 23532 22176
rect 23584 21962 23612 26794
rect 23676 22574 23704 31146
rect 23768 30938 23796 31214
rect 23860 31142 23888 35566
rect 24136 35494 24164 37198
rect 24688 35714 24716 40054
rect 24768 39976 24820 39982
rect 24768 39918 24820 39924
rect 24780 39302 24808 39918
rect 24768 39296 24820 39302
rect 24768 39238 24820 39244
rect 24228 35686 24716 35714
rect 24228 35630 24256 35686
rect 24216 35624 24268 35630
rect 24216 35566 24268 35572
rect 24032 35488 24084 35494
rect 24032 35430 24084 35436
rect 24124 35488 24176 35494
rect 24124 35430 24176 35436
rect 24044 35086 24072 35430
rect 24412 35154 24440 35686
rect 24676 35624 24728 35630
rect 24676 35566 24728 35572
rect 24688 35442 24716 35566
rect 24688 35414 24808 35442
rect 24400 35148 24452 35154
rect 24400 35090 24452 35096
rect 24780 35086 24808 35414
rect 24032 35080 24084 35086
rect 24032 35022 24084 35028
rect 24216 35080 24268 35086
rect 24216 35022 24268 35028
rect 24768 35080 24820 35086
rect 24768 35022 24820 35028
rect 23940 34944 23992 34950
rect 23940 34886 23992 34892
rect 23952 34610 23980 34886
rect 23940 34604 23992 34610
rect 23940 34546 23992 34552
rect 24124 34196 24176 34202
rect 24124 34138 24176 34144
rect 23848 31136 23900 31142
rect 23848 31078 23900 31084
rect 23756 30932 23808 30938
rect 23756 30874 23808 30880
rect 23768 30190 23796 30874
rect 23756 30184 23808 30190
rect 23756 30126 23808 30132
rect 23848 30116 23900 30122
rect 23848 30058 23900 30064
rect 23860 27946 23888 30058
rect 24136 29889 24164 34138
rect 24228 32473 24256 35022
rect 24780 34542 24808 35022
rect 24768 34536 24820 34542
rect 24768 34478 24820 34484
rect 24584 33448 24636 33454
rect 24584 33390 24636 33396
rect 24400 33312 24452 33318
rect 24400 33254 24452 33260
rect 24412 32774 24440 33254
rect 24596 32910 24624 33390
rect 24584 32904 24636 32910
rect 24584 32846 24636 32852
rect 24768 32836 24820 32842
rect 24768 32778 24820 32784
rect 24400 32768 24452 32774
rect 24400 32710 24452 32716
rect 24584 32768 24636 32774
rect 24584 32710 24636 32716
rect 24676 32768 24728 32774
rect 24676 32710 24728 32716
rect 24214 32464 24270 32473
rect 24214 32399 24270 32408
rect 24228 31278 24256 32399
rect 24216 31272 24268 31278
rect 24216 31214 24268 31220
rect 24412 31260 24440 32710
rect 24596 32570 24624 32710
rect 24584 32564 24636 32570
rect 24584 32506 24636 32512
rect 24688 32450 24716 32710
rect 24780 32570 24808 32778
rect 24768 32564 24820 32570
rect 24768 32506 24820 32512
rect 24688 32422 24808 32450
rect 24676 32360 24728 32366
rect 24676 32302 24728 32308
rect 24584 31680 24636 31686
rect 24584 31622 24636 31628
rect 24596 31278 24624 31622
rect 24492 31272 24544 31278
rect 24412 31232 24492 31260
rect 24412 30258 24440 31232
rect 24492 31214 24544 31220
rect 24584 31272 24636 31278
rect 24584 31214 24636 31220
rect 24492 30932 24544 30938
rect 24492 30874 24544 30880
rect 24400 30252 24452 30258
rect 24400 30194 24452 30200
rect 24216 30184 24268 30190
rect 24216 30126 24268 30132
rect 24122 29880 24178 29889
rect 24122 29815 24178 29824
rect 24228 29510 24256 30126
rect 24216 29504 24268 29510
rect 24216 29446 24268 29452
rect 24400 28688 24452 28694
rect 24400 28630 24452 28636
rect 24412 28014 24440 28630
rect 23940 28008 23992 28014
rect 23940 27950 23992 27956
rect 24308 28008 24360 28014
rect 24308 27950 24360 27956
rect 24400 28008 24452 28014
rect 24400 27950 24452 27956
rect 23848 27940 23900 27946
rect 23848 27882 23900 27888
rect 23848 26920 23900 26926
rect 23952 26908 23980 27950
rect 24032 27668 24084 27674
rect 24032 27610 24084 27616
rect 24044 27470 24072 27610
rect 24032 27464 24084 27470
rect 24216 27464 24268 27470
rect 24032 27406 24084 27412
rect 24214 27432 24216 27441
rect 24268 27432 24270 27441
rect 24214 27367 24270 27376
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 23900 26880 23980 26908
rect 23848 26862 23900 26868
rect 24044 26790 24072 26930
rect 24124 26920 24176 26926
rect 24124 26862 24176 26868
rect 24032 26784 24084 26790
rect 24032 26726 24084 26732
rect 24136 26466 24164 26862
rect 24320 26790 24348 27950
rect 24308 26784 24360 26790
rect 24308 26726 24360 26732
rect 23860 26438 24164 26466
rect 23756 26240 23808 26246
rect 23756 26182 23808 26188
rect 23768 25838 23796 26182
rect 23756 25832 23808 25838
rect 23756 25774 23808 25780
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23768 23118 23796 24142
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23860 21690 23888 26438
rect 23940 26376 23992 26382
rect 23940 26318 23992 26324
rect 23952 24206 23980 26318
rect 24124 25424 24176 25430
rect 24122 25392 24124 25401
rect 24176 25392 24178 25401
rect 24122 25327 24178 25336
rect 23940 24200 23992 24206
rect 23940 24142 23992 24148
rect 24032 24132 24084 24138
rect 24032 24074 24084 24080
rect 23940 24064 23992 24070
rect 23940 24006 23992 24012
rect 23952 23730 23980 24006
rect 24044 23798 24072 24074
rect 24032 23792 24084 23798
rect 24032 23734 24084 23740
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 23940 22772 23992 22778
rect 23940 22714 23992 22720
rect 23952 22098 23980 22714
rect 24032 22500 24084 22506
rect 24032 22442 24084 22448
rect 23940 22092 23992 22098
rect 23940 22034 23992 22040
rect 24044 21962 24072 22442
rect 23940 21956 23992 21962
rect 23940 21898 23992 21904
rect 24032 21956 24084 21962
rect 24032 21898 24084 21904
rect 23848 21684 23900 21690
rect 23848 21626 23900 21632
rect 23860 21146 23888 21626
rect 23952 21418 23980 21898
rect 23940 21412 23992 21418
rect 23940 21354 23992 21360
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 23952 21078 23980 21354
rect 23940 21072 23992 21078
rect 23940 21014 23992 21020
rect 23216 20454 23428 20482
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 23032 19310 23060 19654
rect 22928 19304 22980 19310
rect 22928 19246 22980 19252
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22756 18222 22784 18702
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22480 15706 22508 16050
rect 22834 16008 22890 16017
rect 22834 15943 22890 15952
rect 22848 15910 22876 15943
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22836 15904 22888 15910
rect 22836 15846 22888 15852
rect 22572 15706 22600 15846
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22664 15162 22692 15846
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22756 13802 22784 14214
rect 22744 13796 22796 13802
rect 22744 13738 22796 13744
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22572 12850 22600 13262
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22756 12238 22784 13738
rect 22940 12306 22968 19246
rect 23032 18290 23060 19246
rect 23216 19242 23244 20454
rect 23294 20360 23350 20369
rect 23294 20295 23296 20304
rect 23348 20295 23350 20304
rect 23296 20266 23348 20272
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23400 19854 23428 20198
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23492 19530 23520 19790
rect 24136 19666 24164 25327
rect 24504 24886 24532 30874
rect 24596 30258 24624 31214
rect 24688 30802 24716 32302
rect 24780 31226 24808 32422
rect 24872 31328 24900 47534
rect 27160 47524 27212 47530
rect 27160 47466 27212 47472
rect 25688 47252 25740 47258
rect 25688 47194 25740 47200
rect 25700 46578 25728 47194
rect 26700 47048 26752 47054
rect 26700 46990 26752 46996
rect 27068 47048 27120 47054
rect 27068 46990 27120 46996
rect 26148 46980 26200 46986
rect 26148 46922 26200 46928
rect 25320 46572 25372 46578
rect 25320 46514 25372 46520
rect 25688 46572 25740 46578
rect 25688 46514 25740 46520
rect 25332 46170 25360 46514
rect 25872 46368 25924 46374
rect 25872 46310 25924 46316
rect 25320 46164 25372 46170
rect 25320 46106 25372 46112
rect 25596 45960 25648 45966
rect 25596 45902 25648 45908
rect 25780 45960 25832 45966
rect 25780 45902 25832 45908
rect 25608 44878 25636 45902
rect 25792 45082 25820 45902
rect 25780 45076 25832 45082
rect 25780 45018 25832 45024
rect 25596 44872 25648 44878
rect 25780 44872 25832 44878
rect 25596 44814 25648 44820
rect 25686 44840 25742 44849
rect 25320 44804 25372 44810
rect 25320 44746 25372 44752
rect 25332 44470 25360 44746
rect 25320 44464 25372 44470
rect 25320 44406 25372 44412
rect 25410 44432 25466 44441
rect 25410 44367 25412 44376
rect 25464 44367 25466 44376
rect 25412 44338 25464 44344
rect 25504 43716 25556 43722
rect 25504 43658 25556 43664
rect 25516 43450 25544 43658
rect 25504 43444 25556 43450
rect 25504 43386 25556 43392
rect 25608 43314 25636 44814
rect 25780 44814 25832 44820
rect 25686 44775 25742 44784
rect 25700 44742 25728 44775
rect 25688 44736 25740 44742
rect 25688 44678 25740 44684
rect 25700 44402 25728 44678
rect 25688 44396 25740 44402
rect 25688 44338 25740 44344
rect 25596 43308 25648 43314
rect 25596 43250 25648 43256
rect 24952 40180 25004 40186
rect 24952 40122 25004 40128
rect 24964 37806 24992 40122
rect 25700 39574 25728 44338
rect 25792 43994 25820 44814
rect 25780 43988 25832 43994
rect 25780 43930 25832 43936
rect 25884 42634 25912 46310
rect 26160 46170 26188 46922
rect 26332 46368 26384 46374
rect 26332 46310 26384 46316
rect 26148 46164 26200 46170
rect 26148 46106 26200 46112
rect 26344 45966 26372 46310
rect 25964 45960 26016 45966
rect 25964 45902 26016 45908
rect 26332 45960 26384 45966
rect 26332 45902 26384 45908
rect 25976 45626 26004 45902
rect 25964 45620 26016 45626
rect 25964 45562 26016 45568
rect 26712 44946 26740 46990
rect 27080 46918 27108 46990
rect 27068 46912 27120 46918
rect 27068 46854 27120 46860
rect 27080 46578 27108 46854
rect 27068 46572 27120 46578
rect 27068 46514 27120 46520
rect 26884 46436 26936 46442
rect 26884 46378 26936 46384
rect 26700 44940 26752 44946
rect 26700 44882 26752 44888
rect 26608 44872 26660 44878
rect 26608 44814 26660 44820
rect 26792 44872 26844 44878
rect 26792 44814 26844 44820
rect 26424 44804 26476 44810
rect 26424 44746 26476 44752
rect 26054 44432 26110 44441
rect 26436 44402 26464 44746
rect 26054 44367 26110 44376
rect 26424 44396 26476 44402
rect 25964 44192 26016 44198
rect 25964 44134 26016 44140
rect 25976 43314 26004 44134
rect 26068 43314 26096 44367
rect 26424 44338 26476 44344
rect 26516 44328 26568 44334
rect 26516 44270 26568 44276
rect 26424 44260 26476 44266
rect 26424 44202 26476 44208
rect 26436 43790 26464 44202
rect 26424 43784 26476 43790
rect 26424 43726 26476 43732
rect 26240 43716 26292 43722
rect 26240 43658 26292 43664
rect 26252 43450 26280 43658
rect 26240 43444 26292 43450
rect 26240 43386 26292 43392
rect 26528 43314 26556 44270
rect 26620 43450 26648 44814
rect 26804 44305 26832 44814
rect 26790 44296 26846 44305
rect 26790 44231 26846 44240
rect 26700 43648 26752 43654
rect 26700 43590 26752 43596
rect 26792 43648 26844 43654
rect 26792 43590 26844 43596
rect 26608 43444 26660 43450
rect 26608 43386 26660 43392
rect 26712 43314 26740 43590
rect 26804 43382 26832 43590
rect 26896 43382 26924 46378
rect 26976 44396 27028 44402
rect 26976 44338 27028 44344
rect 26988 43790 27016 44338
rect 26976 43784 27028 43790
rect 26976 43726 27028 43732
rect 27080 43636 27108 46514
rect 27172 45966 27200 47466
rect 27356 47258 27384 47602
rect 27436 47524 27488 47530
rect 27436 47466 27488 47472
rect 27344 47252 27396 47258
rect 27344 47194 27396 47200
rect 27356 46714 27384 47194
rect 27448 47025 27476 47466
rect 28276 47122 28304 47670
rect 31392 47456 31444 47462
rect 31392 47398 31444 47404
rect 31484 47456 31536 47462
rect 31484 47398 31536 47404
rect 29184 47252 29236 47258
rect 29184 47194 29236 47200
rect 30104 47252 30156 47258
rect 30104 47194 30156 47200
rect 28264 47116 28316 47122
rect 28264 47058 28316 47064
rect 27896 47048 27948 47054
rect 27434 47016 27490 47025
rect 27896 46990 27948 46996
rect 27434 46951 27490 46960
rect 27344 46708 27396 46714
rect 27344 46650 27396 46656
rect 27252 46572 27304 46578
rect 27252 46514 27304 46520
rect 27264 46170 27292 46514
rect 27344 46368 27396 46374
rect 27620 46368 27672 46374
rect 27344 46310 27396 46316
rect 27540 46328 27620 46356
rect 27252 46164 27304 46170
rect 27252 46106 27304 46112
rect 27160 45960 27212 45966
rect 27160 45902 27212 45908
rect 27160 43784 27212 43790
rect 27158 43752 27160 43761
rect 27212 43752 27214 43761
rect 27158 43687 27214 43696
rect 26988 43608 27108 43636
rect 26792 43376 26844 43382
rect 26792 43318 26844 43324
rect 26884 43376 26936 43382
rect 26884 43318 26936 43324
rect 25964 43308 26016 43314
rect 25964 43250 26016 43256
rect 26056 43308 26108 43314
rect 26056 43250 26108 43256
rect 26516 43308 26568 43314
rect 26516 43250 26568 43256
rect 26700 43308 26752 43314
rect 26700 43250 26752 43256
rect 25872 42628 25924 42634
rect 25872 42570 25924 42576
rect 26068 41274 26096 43250
rect 26988 42770 27016 43608
rect 27250 43344 27306 43353
rect 27250 43279 27252 43288
rect 27304 43279 27306 43288
rect 27252 43250 27304 43256
rect 27356 43217 27384 46310
rect 27540 45966 27568 46328
rect 27620 46310 27672 46316
rect 27712 46164 27764 46170
rect 27712 46106 27764 46112
rect 27528 45960 27580 45966
rect 27528 45902 27580 45908
rect 27620 45960 27672 45966
rect 27724 45914 27752 46106
rect 27672 45908 27752 45914
rect 27620 45902 27752 45908
rect 27632 45886 27752 45902
rect 27632 45830 27660 45886
rect 27620 45824 27672 45830
rect 27620 45766 27672 45772
rect 27712 45076 27764 45082
rect 27712 45018 27764 45024
rect 27724 44742 27752 45018
rect 27804 44872 27856 44878
rect 27804 44814 27856 44820
rect 27712 44736 27764 44742
rect 27712 44678 27764 44684
rect 27724 44577 27752 44678
rect 27710 44568 27766 44577
rect 27710 44503 27766 44512
rect 27724 43722 27752 44503
rect 27816 44402 27844 44814
rect 27804 44396 27856 44402
rect 27804 44338 27856 44344
rect 27712 43716 27764 43722
rect 27712 43658 27764 43664
rect 27620 43648 27672 43654
rect 27620 43590 27672 43596
rect 27342 43208 27398 43217
rect 27342 43143 27398 43152
rect 27068 43104 27120 43110
rect 27068 43046 27120 43052
rect 27080 42945 27108 43046
rect 27066 42936 27122 42945
rect 27066 42871 27122 42880
rect 26976 42764 27028 42770
rect 26976 42706 27028 42712
rect 26884 42084 26936 42090
rect 26884 42026 26936 42032
rect 26896 41614 26924 42026
rect 26884 41608 26936 41614
rect 26884 41550 26936 41556
rect 27356 41546 27384 43143
rect 27632 42702 27660 43590
rect 27620 42696 27672 42702
rect 27620 42638 27672 42644
rect 27344 41540 27396 41546
rect 27344 41482 27396 41488
rect 26056 41268 26108 41274
rect 26056 41210 26108 41216
rect 27804 41064 27856 41070
rect 27908 41052 27936 46990
rect 28356 46980 28408 46986
rect 28356 46922 28408 46928
rect 28368 46374 28396 46922
rect 28540 46640 28592 46646
rect 28540 46582 28592 46588
rect 28356 46368 28408 46374
rect 28356 46310 28408 46316
rect 28172 46164 28224 46170
rect 28172 46106 28224 46112
rect 27988 45960 28040 45966
rect 27988 45902 28040 45908
rect 28000 45626 28028 45902
rect 27988 45620 28040 45626
rect 27988 45562 28040 45568
rect 27988 45076 28040 45082
rect 27988 45018 28040 45024
rect 28000 44810 28028 45018
rect 27988 44804 28040 44810
rect 27988 44746 28040 44752
rect 28000 44198 28028 44746
rect 27988 44192 28040 44198
rect 27988 44134 28040 44140
rect 28080 44192 28132 44198
rect 28080 44134 28132 44140
rect 27988 43852 28040 43858
rect 27988 43794 28040 43800
rect 28000 43654 28028 43794
rect 28092 43790 28120 44134
rect 28184 43858 28212 46106
rect 28264 46028 28316 46034
rect 28264 45970 28316 45976
rect 28276 45286 28304 45970
rect 28356 45892 28408 45898
rect 28356 45834 28408 45840
rect 28264 45280 28316 45286
rect 28264 45222 28316 45228
rect 28276 44810 28304 45222
rect 28264 44804 28316 44810
rect 28264 44746 28316 44752
rect 28276 43858 28304 44746
rect 28172 43852 28224 43858
rect 28172 43794 28224 43800
rect 28264 43852 28316 43858
rect 28264 43794 28316 43800
rect 28080 43784 28132 43790
rect 28080 43726 28132 43732
rect 27988 43648 28040 43654
rect 27988 43590 28040 43596
rect 28184 43382 28212 43794
rect 28368 43790 28396 45834
rect 28446 44976 28502 44985
rect 28446 44911 28448 44920
rect 28500 44911 28502 44920
rect 28448 44882 28500 44888
rect 28356 43784 28408 43790
rect 28354 43752 28356 43761
rect 28408 43752 28410 43761
rect 28354 43687 28410 43696
rect 28172 43376 28224 43382
rect 28172 43318 28224 43324
rect 28552 43110 28580 46582
rect 29196 46510 29224 47194
rect 29828 47184 29880 47190
rect 29828 47126 29880 47132
rect 29276 46912 29328 46918
rect 29276 46854 29328 46860
rect 29288 46714 29316 46854
rect 29276 46708 29328 46714
rect 29276 46650 29328 46656
rect 29288 46510 29316 46650
rect 29840 46578 29868 47126
rect 30116 47054 30144 47194
rect 31404 47122 31432 47398
rect 31392 47116 31444 47122
rect 31392 47058 31444 47064
rect 31496 47054 31524 47398
rect 31944 47184 31996 47190
rect 31944 47126 31996 47132
rect 30104 47048 30156 47054
rect 30104 46990 30156 46996
rect 30288 47048 30340 47054
rect 30288 46990 30340 46996
rect 31484 47048 31536 47054
rect 31484 46990 31536 46996
rect 30012 46980 30064 46986
rect 30012 46922 30064 46928
rect 29828 46572 29880 46578
rect 29828 46514 29880 46520
rect 29184 46504 29236 46510
rect 29184 46446 29236 46452
rect 29276 46504 29328 46510
rect 29276 46446 29328 46452
rect 29460 46504 29512 46510
rect 29460 46446 29512 46452
rect 28632 46368 28684 46374
rect 28632 46310 28684 46316
rect 28644 45626 28672 46310
rect 29196 45966 29224 46446
rect 29288 46034 29316 46446
rect 29472 46102 29500 46446
rect 30024 46442 30052 46922
rect 30300 46714 30328 46990
rect 30288 46708 30340 46714
rect 30288 46650 30340 46656
rect 31956 46578 31984 47126
rect 32140 46594 32168 48010
rect 34440 47802 34468 49694
rect 36082 49624 36138 50424
rect 38658 49624 38714 50424
rect 41234 49722 41290 50424
rect 43166 49722 43222 50424
rect 45742 49722 45798 50424
rect 41234 49694 41368 49722
rect 41234 49624 41290 49694
rect 35594 47900 35902 47909
rect 35594 47898 35600 47900
rect 35656 47898 35680 47900
rect 35736 47898 35760 47900
rect 35816 47898 35840 47900
rect 35896 47898 35902 47900
rect 35656 47846 35658 47898
rect 35838 47846 35840 47898
rect 35594 47844 35600 47846
rect 35656 47844 35680 47846
rect 35736 47844 35760 47846
rect 35816 47844 35840 47846
rect 35896 47844 35902 47846
rect 35594 47835 35902 47844
rect 36096 47802 36124 49624
rect 34428 47796 34480 47802
rect 34428 47738 34480 47744
rect 36084 47796 36136 47802
rect 36084 47738 36136 47744
rect 38384 47728 38436 47734
rect 38384 47670 38436 47676
rect 32220 47660 32272 47666
rect 32220 47602 32272 47608
rect 34336 47660 34388 47666
rect 34336 47602 34388 47608
rect 36912 47660 36964 47666
rect 36912 47602 36964 47608
rect 32232 47258 32260 47602
rect 32404 47592 32456 47598
rect 32404 47534 32456 47540
rect 32220 47252 32272 47258
rect 32220 47194 32272 47200
rect 32220 47048 32272 47054
rect 32220 46990 32272 46996
rect 32232 46714 32260 46990
rect 32220 46708 32272 46714
rect 32220 46650 32272 46656
rect 30288 46572 30340 46578
rect 30288 46514 30340 46520
rect 31944 46572 31996 46578
rect 32140 46566 32260 46594
rect 31944 46514 31996 46520
rect 29552 46436 29604 46442
rect 29552 46378 29604 46384
rect 30012 46436 30064 46442
rect 30012 46378 30064 46384
rect 29460 46096 29512 46102
rect 29460 46038 29512 46044
rect 29276 46028 29328 46034
rect 29276 45970 29328 45976
rect 29184 45960 29236 45966
rect 29184 45902 29236 45908
rect 29472 45642 29500 46038
rect 29564 45830 29592 46378
rect 29644 46368 29696 46374
rect 29644 46310 29696 46316
rect 29552 45824 29604 45830
rect 29552 45766 29604 45772
rect 28632 45620 28684 45626
rect 28632 45562 28684 45568
rect 28816 45620 28868 45626
rect 28816 45562 28868 45568
rect 29196 45614 29500 45642
rect 28724 45484 28776 45490
rect 28644 45444 28724 45472
rect 28644 45014 28672 45444
rect 28724 45426 28776 45432
rect 28632 45008 28684 45014
rect 28630 44976 28632 44985
rect 28684 44976 28686 44985
rect 28630 44911 28686 44920
rect 28828 44878 28856 45562
rect 28908 45484 28960 45490
rect 28908 45426 28960 45432
rect 28920 45370 28948 45426
rect 28920 45342 29040 45370
rect 28908 45076 28960 45082
rect 28908 45018 28960 45024
rect 28632 44872 28684 44878
rect 28630 44840 28632 44849
rect 28816 44872 28868 44878
rect 28684 44840 28686 44849
rect 28686 44798 28764 44826
rect 28816 44814 28868 44820
rect 28630 44775 28686 44784
rect 28632 44736 28684 44742
rect 28630 44704 28632 44713
rect 28684 44704 28686 44713
rect 28630 44639 28686 44648
rect 28630 44568 28686 44577
rect 28630 44503 28686 44512
rect 28644 43790 28672 44503
rect 28736 44266 28764 44798
rect 28920 44334 28948 45018
rect 29012 45014 29040 45342
rect 29092 45348 29144 45354
rect 29092 45290 29144 45296
rect 29000 45008 29052 45014
rect 29000 44950 29052 44956
rect 29012 44402 29040 44950
rect 29104 44742 29132 45290
rect 29196 45286 29224 45614
rect 29276 45484 29328 45490
rect 29276 45426 29328 45432
rect 29184 45280 29236 45286
rect 29184 45222 29236 45228
rect 29196 44878 29224 45222
rect 29184 44872 29236 44878
rect 29184 44814 29236 44820
rect 29288 44742 29316 45426
rect 29368 45416 29420 45422
rect 29368 45358 29420 45364
rect 29460 45416 29512 45422
rect 29460 45358 29512 45364
rect 29380 45082 29408 45358
rect 29472 45286 29500 45358
rect 29460 45280 29512 45286
rect 29460 45222 29512 45228
rect 29368 45076 29420 45082
rect 29368 45018 29420 45024
rect 29368 44872 29420 44878
rect 29368 44814 29420 44820
rect 29092 44736 29144 44742
rect 29092 44678 29144 44684
rect 29276 44736 29328 44742
rect 29276 44678 29328 44684
rect 29104 44402 29132 44678
rect 29288 44538 29316 44678
rect 29276 44532 29328 44538
rect 29276 44474 29328 44480
rect 29380 44470 29408 44814
rect 29460 44804 29512 44810
rect 29460 44746 29512 44752
rect 29472 44538 29500 44746
rect 29460 44532 29512 44538
rect 29460 44474 29512 44480
rect 29368 44464 29420 44470
rect 29368 44406 29420 44412
rect 29000 44396 29052 44402
rect 29000 44338 29052 44344
rect 29092 44396 29144 44402
rect 29092 44338 29144 44344
rect 28908 44328 28960 44334
rect 28908 44270 28960 44276
rect 28724 44260 28776 44266
rect 28724 44202 28776 44208
rect 29104 44198 29132 44338
rect 29092 44192 29144 44198
rect 29092 44134 29144 44140
rect 28632 43784 28684 43790
rect 29092 43784 29144 43790
rect 28632 43726 28684 43732
rect 28998 43752 29054 43761
rect 29092 43726 29144 43732
rect 29184 43784 29236 43790
rect 29184 43726 29236 43732
rect 28998 43687 29054 43696
rect 29012 43654 29040 43687
rect 29104 43654 29132 43726
rect 29000 43648 29052 43654
rect 29000 43590 29052 43596
rect 29092 43648 29144 43654
rect 29092 43590 29144 43596
rect 28540 43104 28592 43110
rect 28540 43046 28592 43052
rect 29196 42838 29224 43726
rect 29564 43382 29592 45766
rect 29656 45558 29684 46310
rect 30300 46170 30328 46514
rect 30840 46368 30892 46374
rect 30840 46310 30892 46316
rect 30288 46164 30340 46170
rect 30288 46106 30340 46112
rect 30852 45966 30880 46310
rect 30472 45960 30524 45966
rect 30472 45902 30524 45908
rect 30564 45960 30616 45966
rect 30564 45902 30616 45908
rect 30840 45960 30892 45966
rect 30840 45902 30892 45908
rect 30380 45824 30432 45830
rect 30380 45766 30432 45772
rect 29644 45552 29696 45558
rect 29644 45494 29696 45500
rect 30392 45422 30420 45766
rect 30380 45416 30432 45422
rect 30484 45404 30512 45902
rect 30576 45626 30604 45902
rect 30656 45824 30708 45830
rect 30656 45766 30708 45772
rect 30564 45620 30616 45626
rect 30564 45562 30616 45568
rect 30564 45416 30616 45422
rect 30484 45376 30564 45404
rect 30380 45358 30432 45364
rect 30564 45358 30616 45364
rect 29736 45348 29788 45354
rect 29736 45290 29788 45296
rect 29748 44334 29776 45290
rect 30576 45286 30604 45358
rect 30564 45280 30616 45286
rect 30564 45222 30616 45228
rect 30472 45076 30524 45082
rect 30472 45018 30524 45024
rect 29828 45008 29880 45014
rect 29828 44950 29880 44956
rect 29840 44554 29868 44950
rect 30484 44878 30512 45018
rect 30576 44878 30604 45222
rect 30472 44872 30524 44878
rect 30472 44814 30524 44820
rect 30564 44872 30616 44878
rect 30564 44814 30616 44820
rect 30104 44804 30156 44810
rect 30104 44746 30156 44752
rect 29920 44736 29972 44742
rect 29972 44696 30052 44724
rect 29920 44678 29972 44684
rect 29840 44526 29960 44554
rect 29932 44334 29960 44526
rect 29736 44328 29788 44334
rect 29736 44270 29788 44276
rect 29920 44328 29972 44334
rect 29920 44270 29972 44276
rect 29828 44192 29880 44198
rect 29828 44134 29880 44140
rect 29840 43858 29868 44134
rect 29932 43858 29960 44270
rect 30024 43858 30052 44696
rect 30116 44470 30144 44746
rect 30668 44713 30696 45766
rect 30654 44704 30710 44713
rect 30654 44639 30710 44648
rect 30104 44464 30156 44470
rect 30104 44406 30156 44412
rect 29828 43852 29880 43858
rect 29828 43794 29880 43800
rect 29920 43852 29972 43858
rect 29920 43794 29972 43800
rect 30012 43852 30064 43858
rect 30012 43794 30064 43800
rect 29734 43480 29790 43489
rect 29734 43415 29790 43424
rect 29552 43376 29604 43382
rect 29552 43318 29604 43324
rect 29748 43314 29776 43415
rect 30116 43314 30144 44406
rect 30288 44396 30340 44402
rect 30288 44338 30340 44344
rect 30196 43920 30248 43926
rect 30196 43862 30248 43868
rect 29736 43308 29788 43314
rect 29736 43250 29788 43256
rect 29920 43308 29972 43314
rect 29920 43250 29972 43256
rect 30104 43308 30156 43314
rect 30104 43250 30156 43256
rect 29552 43240 29604 43246
rect 29472 43200 29552 43228
rect 29184 42832 29236 42838
rect 29184 42774 29236 42780
rect 29472 42702 29500 43200
rect 29552 43182 29604 43188
rect 29460 42696 29512 42702
rect 29460 42638 29512 42644
rect 28816 42628 28868 42634
rect 28816 42570 28868 42576
rect 27988 41540 28040 41546
rect 27988 41482 28040 41488
rect 27856 41024 27936 41052
rect 27804 41006 27856 41012
rect 25872 40928 25924 40934
rect 25872 40870 25924 40876
rect 25884 40186 25912 40870
rect 27252 40520 27304 40526
rect 27436 40520 27488 40526
rect 27304 40480 27436 40508
rect 27252 40462 27304 40468
rect 27436 40462 27488 40468
rect 27526 40488 27582 40497
rect 26240 40452 26292 40458
rect 26240 40394 26292 40400
rect 26252 40186 26280 40394
rect 27068 40384 27120 40390
rect 27068 40326 27120 40332
rect 27080 40186 27108 40326
rect 25872 40180 25924 40186
rect 25872 40122 25924 40128
rect 26240 40180 26292 40186
rect 26240 40122 26292 40128
rect 26884 40180 26936 40186
rect 27068 40180 27120 40186
rect 26936 40140 27068 40168
rect 26884 40122 26936 40128
rect 27068 40122 27120 40128
rect 27448 40118 27476 40462
rect 27526 40423 27582 40432
rect 27436 40112 27488 40118
rect 27436 40054 27488 40060
rect 27540 39982 27568 40423
rect 26240 39976 26292 39982
rect 26240 39918 26292 39924
rect 27436 39976 27488 39982
rect 27436 39918 27488 39924
rect 27528 39976 27580 39982
rect 27528 39918 27580 39924
rect 26252 39574 26280 39918
rect 25688 39568 25740 39574
rect 25688 39510 25740 39516
rect 26240 39568 26292 39574
rect 26240 39510 26292 39516
rect 27448 39506 27476 39918
rect 26792 39500 26844 39506
rect 26792 39442 26844 39448
rect 27436 39500 27488 39506
rect 27436 39442 27488 39448
rect 25320 38956 25372 38962
rect 25320 38898 25372 38904
rect 25780 38956 25832 38962
rect 25780 38898 25832 38904
rect 25332 37874 25360 38898
rect 25792 38554 25820 38898
rect 25780 38548 25832 38554
rect 25780 38490 25832 38496
rect 26608 38276 26660 38282
rect 26608 38218 26660 38224
rect 26620 38010 26648 38218
rect 26608 38004 26660 38010
rect 26608 37946 26660 37952
rect 26148 37936 26200 37942
rect 25976 37896 26148 37924
rect 25320 37868 25372 37874
rect 25320 37810 25372 37816
rect 24952 37800 25004 37806
rect 24952 37742 25004 37748
rect 25044 37732 25096 37738
rect 25044 37674 25096 37680
rect 25056 37466 25084 37674
rect 25044 37460 25096 37466
rect 25044 37402 25096 37408
rect 25056 35986 25084 37402
rect 25332 37330 25360 37810
rect 25976 37806 26004 37896
rect 26148 37878 26200 37884
rect 26700 37868 26752 37874
rect 26700 37810 26752 37816
rect 25412 37800 25464 37806
rect 25412 37742 25464 37748
rect 25964 37800 26016 37806
rect 25964 37742 26016 37748
rect 26148 37800 26200 37806
rect 26148 37742 26200 37748
rect 25424 37330 25452 37742
rect 25136 37324 25188 37330
rect 25136 37266 25188 37272
rect 25320 37324 25372 37330
rect 25320 37266 25372 37272
rect 25412 37324 25464 37330
rect 25412 37266 25464 37272
rect 24964 35958 25084 35986
rect 24964 31754 24992 35958
rect 25044 35828 25096 35834
rect 25044 35770 25096 35776
rect 25056 35698 25084 35770
rect 25044 35692 25096 35698
rect 25044 35634 25096 35640
rect 25044 35148 25096 35154
rect 25148 35136 25176 37266
rect 25596 37256 25648 37262
rect 25596 37198 25648 37204
rect 25504 36236 25556 36242
rect 25504 36178 25556 36184
rect 25320 35828 25372 35834
rect 25320 35770 25372 35776
rect 25228 35624 25280 35630
rect 25228 35566 25280 35572
rect 25240 35329 25268 35566
rect 25226 35320 25282 35329
rect 25226 35255 25282 35264
rect 25096 35108 25176 35136
rect 25044 35090 25096 35096
rect 25332 35086 25360 35770
rect 25516 35630 25544 36178
rect 25504 35624 25556 35630
rect 25504 35566 25556 35572
rect 25410 35320 25466 35329
rect 25410 35255 25466 35264
rect 25424 35086 25452 35255
rect 25608 35086 25636 37198
rect 25688 36236 25740 36242
rect 25688 36178 25740 36184
rect 25320 35080 25372 35086
rect 25320 35022 25372 35028
rect 25412 35080 25464 35086
rect 25412 35022 25464 35028
rect 25596 35080 25648 35086
rect 25596 35022 25648 35028
rect 25412 32768 25464 32774
rect 25412 32710 25464 32716
rect 25424 32570 25452 32710
rect 25412 32564 25464 32570
rect 25412 32506 25464 32512
rect 25608 32201 25636 35022
rect 25700 34610 25728 36178
rect 25872 34944 25924 34950
rect 25792 34904 25872 34932
rect 25688 34604 25740 34610
rect 25688 34546 25740 34552
rect 25792 34542 25820 34904
rect 25872 34886 25924 34892
rect 25780 34536 25832 34542
rect 25780 34478 25832 34484
rect 25792 33114 25820 34478
rect 25780 33108 25832 33114
rect 25780 33050 25832 33056
rect 25594 32192 25650 32201
rect 25594 32127 25650 32136
rect 24964 31726 25268 31754
rect 24872 31300 25084 31328
rect 24780 31198 24900 31226
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24676 30796 24728 30802
rect 24676 30738 24728 30744
rect 24780 30784 24808 31078
rect 24872 30938 24900 31198
rect 24860 30932 24912 30938
rect 24860 30874 24912 30880
rect 24952 30796 25004 30802
rect 24780 30756 24952 30784
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 24676 30184 24728 30190
rect 24676 30126 24728 30132
rect 24688 28694 24716 30126
rect 24676 28688 24728 28694
rect 24676 28630 24728 28636
rect 24780 27402 24808 30756
rect 24952 30738 25004 30744
rect 24952 30388 25004 30394
rect 25056 30376 25084 31300
rect 25136 30388 25188 30394
rect 25056 30348 25136 30376
rect 24952 30330 25004 30336
rect 25136 30330 25188 30336
rect 24964 29578 24992 30330
rect 25240 30274 25268 31726
rect 25608 31278 25636 32127
rect 25792 31278 25820 33050
rect 25596 31272 25648 31278
rect 25596 31214 25648 31220
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 25148 30246 25268 30274
rect 25320 30252 25372 30258
rect 24952 29572 25004 29578
rect 24952 29514 25004 29520
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 24872 27441 24900 28494
rect 24858 27432 24914 27441
rect 24768 27396 24820 27402
rect 24858 27367 24914 27376
rect 24768 27338 24820 27344
rect 25044 26988 25096 26994
rect 25044 26930 25096 26936
rect 24768 26784 24820 26790
rect 24768 26726 24820 26732
rect 24780 26518 24808 26726
rect 24768 26512 24820 26518
rect 24768 26454 24820 26460
rect 24492 24880 24544 24886
rect 24492 24822 24544 24828
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24688 24206 24716 24550
rect 24308 24200 24360 24206
rect 24308 24142 24360 24148
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24320 22438 24348 24142
rect 24492 23248 24544 23254
rect 24492 23190 24544 23196
rect 25056 23202 25084 26930
rect 25148 26625 25176 30246
rect 25320 30194 25372 30200
rect 25332 29782 25360 30194
rect 25412 30184 25464 30190
rect 25412 30126 25464 30132
rect 25424 29850 25452 30126
rect 25504 30048 25556 30054
rect 25504 29990 25556 29996
rect 25688 30048 25740 30054
rect 25688 29990 25740 29996
rect 25412 29844 25464 29850
rect 25412 29786 25464 29792
rect 25516 29782 25544 29990
rect 25700 29850 25728 29990
rect 25688 29844 25740 29850
rect 25688 29786 25740 29792
rect 25320 29776 25372 29782
rect 25320 29718 25372 29724
rect 25504 29776 25556 29782
rect 25504 29718 25556 29724
rect 25228 29572 25280 29578
rect 25228 29514 25280 29520
rect 25240 28014 25268 29514
rect 25228 28008 25280 28014
rect 25228 27950 25280 27956
rect 25240 26908 25268 27950
rect 25332 27062 25360 29718
rect 25596 27872 25648 27878
rect 25596 27814 25648 27820
rect 25320 27056 25372 27062
rect 25320 26998 25372 27004
rect 25608 26926 25636 27814
rect 25596 26920 25648 26926
rect 25240 26880 25360 26908
rect 25228 26784 25280 26790
rect 25228 26726 25280 26732
rect 25134 26616 25190 26625
rect 25240 26586 25268 26726
rect 25134 26551 25190 26560
rect 25228 26580 25280 26586
rect 25228 26522 25280 26528
rect 25228 25152 25280 25158
rect 25228 25094 25280 25100
rect 25240 24954 25268 25094
rect 25228 24948 25280 24954
rect 25228 24890 25280 24896
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25240 23866 25268 24754
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25228 23588 25280 23594
rect 25228 23530 25280 23536
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24308 22432 24360 22438
rect 24308 22374 24360 22380
rect 24320 22030 24348 22374
rect 24308 22024 24360 22030
rect 24308 21966 24360 21972
rect 24412 21622 24440 22578
rect 24504 22166 24532 23190
rect 24676 23180 24728 23186
rect 25056 23174 25176 23202
rect 24676 23122 24728 23128
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24492 22160 24544 22166
rect 24492 22102 24544 22108
rect 24492 21888 24544 21894
rect 24492 21830 24544 21836
rect 24400 21616 24452 21622
rect 24400 21558 24452 21564
rect 24504 21554 24532 21830
rect 24596 21690 24624 22578
rect 24688 22098 24716 23122
rect 24952 22976 25004 22982
rect 24952 22918 25004 22924
rect 24780 22234 24900 22250
rect 24780 22228 24912 22234
rect 24780 22222 24860 22228
rect 24780 22098 24808 22222
rect 24860 22170 24912 22176
rect 24676 22092 24728 22098
rect 24676 22034 24728 22040
rect 24768 22092 24820 22098
rect 24964 22094 24992 22918
rect 24768 22034 24820 22040
rect 24872 22066 24992 22094
rect 25148 22080 25176 23174
rect 25240 22137 25268 23530
rect 24768 21956 24820 21962
rect 24768 21898 24820 21904
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24584 21684 24636 21690
rect 24584 21626 24636 21632
rect 24308 21548 24360 21554
rect 24308 21490 24360 21496
rect 24492 21548 24544 21554
rect 24688 21536 24716 21830
rect 24780 21690 24808 21898
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24768 21548 24820 21554
rect 24688 21508 24768 21536
rect 24492 21490 24544 21496
rect 24768 21490 24820 21496
rect 24320 20942 24348 21490
rect 24872 20942 24900 22066
rect 25056 22052 25176 22080
rect 25226 22128 25282 22137
rect 25226 22063 25282 22072
rect 24952 21888 25004 21894
rect 24952 21830 25004 21836
rect 24964 21486 24992 21830
rect 25056 21486 25084 22052
rect 24952 21480 25004 21486
rect 24952 21422 25004 21428
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 24308 20936 24360 20942
rect 24308 20878 24360 20884
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24320 20330 24348 20878
rect 24768 20868 24820 20874
rect 24768 20810 24820 20816
rect 24400 20460 24452 20466
rect 24400 20402 24452 20408
rect 24308 20324 24360 20330
rect 24308 20266 24360 20272
rect 23768 19638 24164 19666
rect 23308 19502 23612 19530
rect 23308 19446 23336 19502
rect 23296 19440 23348 19446
rect 23296 19382 23348 19388
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23204 19236 23256 19242
rect 23204 19178 23256 19184
rect 23020 18284 23072 18290
rect 23020 18226 23072 18232
rect 23308 18222 23336 19246
rect 23492 18630 23520 19314
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23584 17814 23612 19502
rect 23664 19236 23716 19242
rect 23664 19178 23716 19184
rect 23676 18834 23704 19178
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23020 17536 23072 17542
rect 23020 17478 23072 17484
rect 23032 17270 23060 17478
rect 23020 17264 23072 17270
rect 23020 17206 23072 17212
rect 23216 16794 23244 17614
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23492 16096 23520 17274
rect 23584 16726 23612 17750
rect 23572 16720 23624 16726
rect 23572 16662 23624 16668
rect 23664 16108 23716 16114
rect 23492 16068 23664 16096
rect 23664 16050 23716 16056
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23308 15094 23336 15846
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23296 15088 23348 15094
rect 23296 15030 23348 15036
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23400 14074 23428 14758
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23020 13184 23072 13190
rect 23020 13126 23072 13132
rect 23032 12782 23060 13126
rect 23308 12782 23336 13262
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 23296 12776 23348 12782
rect 23296 12718 23348 12724
rect 23204 12640 23256 12646
rect 23204 12582 23256 12588
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22480 11150 22508 12174
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23124 11762 23152 12038
rect 23112 11756 23164 11762
rect 23112 11698 23164 11704
rect 23216 11558 23244 12582
rect 23400 12374 23428 13262
rect 23388 12368 23440 12374
rect 23388 12310 23440 12316
rect 23296 12232 23348 12238
rect 23296 12174 23348 12180
rect 23308 11830 23336 12174
rect 23400 12084 23428 12310
rect 23492 12186 23520 15438
rect 23664 14340 23716 14346
rect 23664 14282 23716 14288
rect 23570 13696 23626 13705
rect 23570 13631 23626 13640
rect 23584 13394 23612 13631
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23676 12889 23704 14282
rect 23662 12880 23718 12889
rect 23662 12815 23718 12824
rect 23676 12714 23704 12815
rect 23664 12708 23716 12714
rect 23664 12650 23716 12656
rect 23676 12594 23704 12650
rect 23584 12566 23704 12594
rect 23584 12434 23612 12566
rect 23584 12406 23704 12434
rect 23492 12158 23612 12186
rect 23480 12096 23532 12102
rect 23400 12056 23480 12084
rect 23480 12038 23532 12044
rect 23296 11824 23348 11830
rect 23296 11766 23348 11772
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 22848 10810 22876 11018
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 23032 10674 23060 11494
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 22190 10095 22246 10104
rect 22284 10124 22336 10130
rect 22204 10062 22232 10095
rect 22284 10066 22336 10072
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 22192 10056 22244 10062
rect 22192 9998 22244 10004
rect 22296 10010 22324 10066
rect 22296 9982 22508 10010
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 21744 8566 21772 8774
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21836 8498 21864 8978
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 21192 7342 21220 8026
rect 22020 7546 22048 8910
rect 22204 8634 22232 8978
rect 22296 8974 22324 9522
rect 22388 9178 22416 9862
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22480 9042 22508 9982
rect 23124 9518 23152 10066
rect 23216 10062 23244 11290
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23112 9512 23164 9518
rect 23112 9454 23164 9460
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22468 9036 22520 9042
rect 22468 8978 22520 8984
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22468 8832 22520 8838
rect 22572 8820 22600 9318
rect 23584 8838 23612 12158
rect 22520 8792 22600 8820
rect 23572 8832 23624 8838
rect 22468 8774 22520 8780
rect 23572 8774 23624 8780
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 23020 8356 23072 8362
rect 23020 8298 23072 8304
rect 22112 8022 22140 8298
rect 22836 8288 22888 8294
rect 22836 8230 22888 8236
rect 22466 8120 22522 8129
rect 22466 8055 22522 8064
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 21180 7336 21232 7342
rect 21180 7278 21232 7284
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22112 5846 22140 6190
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 22100 5840 22152 5846
rect 22100 5782 22152 5788
rect 20902 5672 20958 5681
rect 20902 5607 20958 5616
rect 20916 3534 20944 5607
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 21652 4826 21680 5170
rect 21640 4820 21692 4826
rect 21640 4762 21692 4768
rect 21744 4554 21772 5782
rect 22112 5370 22140 5782
rect 22204 5574 22232 6258
rect 22480 6254 22508 8055
rect 22848 7886 22876 8230
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 22560 6248 22612 6254
rect 22836 6248 22888 6254
rect 22560 6190 22612 6196
rect 22664 6208 22836 6236
rect 22572 5710 22600 6190
rect 22664 5778 22692 6208
rect 22836 6190 22888 6196
rect 23032 5914 23060 8298
rect 23124 7546 23152 8434
rect 23676 8362 23704 12406
rect 23768 10033 23796 19638
rect 24124 19508 24176 19514
rect 24124 19450 24176 19456
rect 24136 19310 24164 19450
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 23940 18284 23992 18290
rect 24044 18272 24072 19246
rect 24136 18970 24164 19246
rect 24216 19168 24268 19174
rect 24216 19110 24268 19116
rect 24228 18970 24256 19110
rect 24124 18964 24176 18970
rect 24124 18906 24176 18912
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24136 18290 24164 18906
rect 24320 18834 24348 20266
rect 24412 20058 24440 20402
rect 24676 20256 24728 20262
rect 24676 20198 24728 20204
rect 24400 20052 24452 20058
rect 24400 19994 24452 20000
rect 24688 19922 24716 20198
rect 24780 20058 24808 20810
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24688 19310 24716 19722
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 24308 18828 24360 18834
rect 24308 18770 24360 18776
rect 23992 18244 24072 18272
rect 23940 18226 23992 18232
rect 24044 17338 24072 18244
rect 24124 18284 24176 18290
rect 24124 18226 24176 18232
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 23860 11830 23888 16594
rect 24044 16590 24072 17274
rect 24032 16584 24084 16590
rect 24032 16526 24084 16532
rect 23940 16516 23992 16522
rect 23940 16458 23992 16464
rect 23952 16114 23980 16458
rect 24320 16454 24348 18770
rect 24688 18154 24716 19246
rect 24676 18148 24728 18154
rect 24676 18090 24728 18096
rect 24780 18034 24808 19790
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24872 18834 24900 19110
rect 24860 18828 24912 18834
rect 24860 18770 24912 18776
rect 24952 18692 25004 18698
rect 24952 18634 25004 18640
rect 24964 18426 24992 18634
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 24688 18006 24808 18034
rect 24308 16448 24360 16454
rect 24308 16390 24360 16396
rect 24216 16176 24268 16182
rect 24216 16118 24268 16124
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 24044 14618 24072 15982
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 23952 11898 23980 12718
rect 24044 12374 24072 12718
rect 24032 12368 24084 12374
rect 24032 12310 24084 12316
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 23848 11824 23900 11830
rect 23848 11766 23900 11772
rect 23952 11354 23980 11834
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 23754 10024 23810 10033
rect 23754 9959 23810 9968
rect 24136 9450 24164 15506
rect 24228 13530 24256 16118
rect 24320 14278 24348 16390
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24596 12782 24624 13670
rect 24688 13394 24716 18006
rect 24860 17264 24912 17270
rect 24860 17206 24912 17212
rect 24872 16794 24900 17206
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24860 16108 24912 16114
rect 25056 16096 25084 21422
rect 25136 16516 25188 16522
rect 25136 16458 25188 16464
rect 25148 16114 25176 16458
rect 24912 16068 25084 16096
rect 25136 16108 25188 16114
rect 24860 16050 24912 16056
rect 25136 16050 25188 16056
rect 24872 15502 24900 16050
rect 25136 15632 25188 15638
rect 25136 15574 25188 15580
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24780 14074 24808 14214
rect 24768 14068 24820 14074
rect 24768 14010 24820 14016
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 24688 12986 24716 13126
rect 24872 12986 24900 14214
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 25056 13258 25084 13806
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 24964 12889 24992 12922
rect 24950 12880 25006 12889
rect 24950 12815 25006 12824
rect 24584 12776 24636 12782
rect 24584 12718 24636 12724
rect 24596 12434 24624 12718
rect 24768 12708 24820 12714
rect 24768 12650 24820 12656
rect 24780 12434 24808 12650
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 24596 12406 24808 12434
rect 24492 12232 24544 12238
rect 24492 12174 24544 12180
rect 24504 11694 24532 12174
rect 24492 11688 24544 11694
rect 24492 11630 24544 11636
rect 24504 11150 24532 11630
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 24124 9444 24176 9450
rect 24124 9386 24176 9392
rect 24412 9042 24440 9522
rect 24400 9036 24452 9042
rect 24400 8978 24452 8984
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 24044 8566 24072 8774
rect 24412 8634 24440 8978
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24032 8560 24084 8566
rect 24032 8502 24084 8508
rect 24504 8430 24532 11086
rect 24596 9602 24624 12406
rect 24964 12322 24992 12582
rect 25148 12434 25176 15574
rect 25240 14482 25268 22063
rect 25332 15910 25360 26880
rect 25596 26862 25648 26868
rect 25688 25900 25740 25906
rect 25688 25842 25740 25848
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25516 23662 25544 24754
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25596 23588 25648 23594
rect 25596 23530 25648 23536
rect 25608 23254 25636 23530
rect 25596 23248 25648 23254
rect 25596 23190 25648 23196
rect 25608 23118 25636 23190
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25412 22636 25464 22642
rect 25412 22578 25464 22584
rect 25424 22030 25452 22578
rect 25596 22500 25648 22506
rect 25596 22442 25648 22448
rect 25608 22166 25636 22442
rect 25596 22160 25648 22166
rect 25596 22102 25648 22108
rect 25412 22024 25464 22030
rect 25412 21966 25464 21972
rect 25410 21856 25466 21865
rect 25700 21842 25728 25842
rect 25792 24206 25820 31214
rect 25872 30592 25924 30598
rect 25872 30534 25924 30540
rect 25884 30258 25912 30534
rect 25872 30252 25924 30258
rect 25872 30194 25924 30200
rect 25976 28626 26004 37742
rect 26160 37466 26188 37742
rect 26424 37664 26476 37670
rect 26424 37606 26476 37612
rect 26148 37460 26200 37466
rect 26148 37402 26200 37408
rect 26240 37324 26292 37330
rect 26240 37266 26292 37272
rect 26056 36168 26108 36174
rect 26056 36110 26108 36116
rect 26068 35698 26096 36110
rect 26148 36032 26200 36038
rect 26148 35974 26200 35980
rect 26160 35766 26188 35974
rect 26148 35760 26200 35766
rect 26148 35702 26200 35708
rect 26056 35692 26108 35698
rect 26056 35634 26108 35640
rect 26148 35624 26200 35630
rect 26148 35566 26200 35572
rect 26160 34406 26188 35566
rect 26252 34746 26280 37266
rect 26436 35562 26464 37606
rect 26712 37466 26740 37810
rect 26700 37460 26752 37466
rect 26700 37402 26752 37408
rect 26804 37330 26832 39442
rect 27620 39432 27672 39438
rect 27620 39374 27672 39380
rect 27344 38888 27396 38894
rect 27344 38830 27396 38836
rect 27356 38418 27384 38830
rect 27344 38412 27396 38418
rect 27344 38354 27396 38360
rect 26976 38344 27028 38350
rect 26976 38286 27028 38292
rect 26792 37324 26844 37330
rect 26712 37284 26792 37312
rect 26424 35556 26476 35562
rect 26424 35498 26476 35504
rect 26240 34740 26292 34746
rect 26240 34682 26292 34688
rect 26148 34400 26200 34406
rect 26148 34342 26200 34348
rect 26056 33516 26108 33522
rect 26056 33458 26108 33464
rect 26068 33114 26096 33458
rect 26516 33312 26568 33318
rect 26516 33254 26568 33260
rect 26056 33108 26108 33114
rect 26056 33050 26108 33056
rect 26528 32910 26556 33254
rect 26516 32904 26568 32910
rect 26516 32846 26568 32852
rect 26608 32836 26660 32842
rect 26608 32778 26660 32784
rect 26332 32428 26384 32434
rect 26332 32370 26384 32376
rect 26056 30660 26108 30666
rect 26056 30602 26108 30608
rect 25964 28620 26016 28626
rect 25964 28562 26016 28568
rect 25976 27146 26004 28562
rect 25884 27118 26004 27146
rect 25884 26042 25912 27118
rect 25962 27024 26018 27033
rect 25962 26959 25964 26968
rect 26016 26959 26018 26968
rect 25964 26930 26016 26936
rect 25962 26480 26018 26489
rect 25962 26415 26018 26424
rect 25872 26036 25924 26042
rect 25872 25978 25924 25984
rect 25976 25906 26004 26415
rect 26068 26382 26096 30602
rect 26240 30184 26292 30190
rect 26160 30132 26240 30138
rect 26160 30126 26292 30132
rect 26160 30110 26280 30126
rect 26160 29782 26188 30110
rect 26148 29776 26200 29782
rect 26148 29718 26200 29724
rect 26160 28558 26188 29718
rect 26148 28552 26200 28558
rect 26148 28494 26200 28500
rect 26344 27538 26372 32370
rect 26620 32366 26648 32778
rect 26712 32434 26740 37284
rect 26792 37266 26844 37272
rect 26988 36786 27016 38286
rect 27068 37664 27120 37670
rect 27068 37606 27120 37612
rect 27080 36854 27108 37606
rect 27068 36848 27120 36854
rect 27068 36790 27120 36796
rect 26976 36780 27028 36786
rect 26976 36722 27028 36728
rect 27356 35816 27384 38354
rect 27632 37874 27660 39374
rect 27816 38350 27844 41006
rect 27896 40452 27948 40458
rect 27896 40394 27948 40400
rect 27908 39642 27936 40394
rect 27896 39636 27948 39642
rect 27896 39578 27948 39584
rect 28000 39370 28028 41482
rect 28448 41064 28500 41070
rect 28448 41006 28500 41012
rect 28264 40384 28316 40390
rect 28264 40326 28316 40332
rect 28276 39438 28304 40326
rect 28460 40050 28488 41006
rect 28448 40044 28500 40050
rect 28448 39986 28500 39992
rect 28264 39432 28316 39438
rect 28264 39374 28316 39380
rect 27988 39364 28040 39370
rect 27988 39306 28040 39312
rect 28000 39030 28028 39306
rect 27988 39024 28040 39030
rect 27988 38966 28040 38972
rect 28460 38418 28488 39986
rect 28448 38412 28500 38418
rect 28448 38354 28500 38360
rect 27804 38344 27856 38350
rect 27804 38286 27856 38292
rect 28080 38276 28132 38282
rect 28080 38218 28132 38224
rect 27712 38208 27764 38214
rect 27712 38150 27764 38156
rect 27804 38208 27856 38214
rect 27804 38150 27856 38156
rect 27620 37868 27672 37874
rect 27620 37810 27672 37816
rect 27632 37330 27660 37810
rect 27620 37324 27672 37330
rect 27620 37266 27672 37272
rect 27724 37126 27752 38150
rect 27816 37942 27844 38150
rect 27804 37936 27856 37942
rect 27804 37878 27856 37884
rect 27896 37664 27948 37670
rect 27896 37606 27948 37612
rect 27908 37330 27936 37606
rect 28092 37398 28120 38218
rect 28172 38208 28224 38214
rect 28172 38150 28224 38156
rect 28184 37806 28212 38150
rect 28172 37800 28224 37806
rect 28172 37742 28224 37748
rect 28724 37800 28776 37806
rect 28724 37742 28776 37748
rect 28080 37392 28132 37398
rect 28080 37334 28132 37340
rect 27896 37324 27948 37330
rect 27896 37266 27948 37272
rect 27988 37324 28040 37330
rect 27988 37266 28040 37272
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 27526 36000 27582 36009
rect 27526 35935 27582 35944
rect 27172 35788 27384 35816
rect 26974 35728 27030 35737
rect 26974 35663 27030 35672
rect 26988 35630 27016 35663
rect 26976 35624 27028 35630
rect 26976 35566 27028 35572
rect 26884 35488 26936 35494
rect 26884 35430 26936 35436
rect 26896 35222 26924 35430
rect 26884 35216 26936 35222
rect 26790 35184 26846 35193
rect 26884 35158 26936 35164
rect 26790 35119 26846 35128
rect 26804 35086 26832 35119
rect 26792 35080 26844 35086
rect 26792 35022 26844 35028
rect 27172 32978 27200 35788
rect 27252 35692 27304 35698
rect 27252 35634 27304 35640
rect 27264 35290 27292 35634
rect 27342 35456 27398 35465
rect 27342 35391 27398 35400
rect 27252 35284 27304 35290
rect 27252 35226 27304 35232
rect 26792 32972 26844 32978
rect 26792 32914 26844 32920
rect 26884 32972 26936 32978
rect 26884 32914 26936 32920
rect 27160 32972 27212 32978
rect 27160 32914 27212 32920
rect 26804 32502 26832 32914
rect 26792 32496 26844 32502
rect 26792 32438 26844 32444
rect 26700 32428 26752 32434
rect 26700 32370 26752 32376
rect 26608 32360 26660 32366
rect 26608 32302 26660 32308
rect 26620 31890 26648 32302
rect 26608 31884 26660 31890
rect 26608 31826 26660 31832
rect 26700 31816 26752 31822
rect 26896 31804 26924 32914
rect 27160 32360 27212 32366
rect 27160 32302 27212 32308
rect 27172 32230 27200 32302
rect 27160 32224 27212 32230
rect 27160 32166 27212 32172
rect 27172 31890 27200 32166
rect 27356 31958 27384 35391
rect 27540 33368 27568 35935
rect 27896 35760 27948 35766
rect 27896 35702 27948 35708
rect 27908 35086 27936 35702
rect 28000 35465 28028 37266
rect 28092 36854 28120 37334
rect 28184 37312 28212 37742
rect 28736 37330 28764 37742
rect 28264 37324 28316 37330
rect 28184 37284 28264 37312
rect 28264 37266 28316 37272
rect 28356 37324 28408 37330
rect 28356 37266 28408 37272
rect 28724 37324 28776 37330
rect 28724 37266 28776 37272
rect 28276 36922 28304 37266
rect 28368 37126 28396 37266
rect 28540 37256 28592 37262
rect 28540 37198 28592 37204
rect 28356 37120 28408 37126
rect 28356 37062 28408 37068
rect 28264 36916 28316 36922
rect 28264 36858 28316 36864
rect 28080 36848 28132 36854
rect 28080 36790 28132 36796
rect 28552 36009 28580 37198
rect 28538 36000 28594 36009
rect 28538 35935 28594 35944
rect 27986 35456 28042 35465
rect 27986 35391 28042 35400
rect 27712 35080 27764 35086
rect 27712 35022 27764 35028
rect 27896 35080 27948 35086
rect 27896 35022 27948 35028
rect 28080 35080 28132 35086
rect 28080 35022 28132 35028
rect 28724 35080 28776 35086
rect 28724 35022 28776 35028
rect 27724 34950 27752 35022
rect 27804 35012 27856 35018
rect 27804 34954 27856 34960
rect 27712 34944 27764 34950
rect 27712 34886 27764 34892
rect 27620 34468 27672 34474
rect 27620 34410 27672 34416
rect 27632 33522 27660 34410
rect 27724 33658 27752 34886
rect 27816 34610 27844 34954
rect 27804 34604 27856 34610
rect 27804 34546 27856 34552
rect 27712 33652 27764 33658
rect 27712 33594 27764 33600
rect 27620 33516 27672 33522
rect 27620 33458 27672 33464
rect 27540 33340 27844 33368
rect 27528 32904 27580 32910
rect 27528 32846 27580 32852
rect 27540 32366 27568 32846
rect 27528 32360 27580 32366
rect 27528 32302 27580 32308
rect 27344 31952 27396 31958
rect 27344 31894 27396 31900
rect 27160 31884 27212 31890
rect 27160 31826 27212 31832
rect 26752 31776 26924 31804
rect 26700 31758 26752 31764
rect 26792 30252 26844 30258
rect 26792 30194 26844 30200
rect 26804 29850 26832 30194
rect 26792 29844 26844 29850
rect 26792 29786 26844 29792
rect 26608 28484 26660 28490
rect 26608 28426 26660 28432
rect 26620 28218 26648 28426
rect 26608 28212 26660 28218
rect 26608 28154 26660 28160
rect 26896 27946 26924 31776
rect 27356 30870 27384 31894
rect 27540 31890 27568 32302
rect 27620 32292 27672 32298
rect 27620 32234 27672 32240
rect 27632 32065 27660 32234
rect 27618 32056 27674 32065
rect 27618 31991 27674 32000
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 27816 31822 27844 33340
rect 27988 32564 28040 32570
rect 27988 32506 28040 32512
rect 28000 32434 28028 32506
rect 27988 32428 28040 32434
rect 27988 32370 28040 32376
rect 28000 31890 28028 32370
rect 27988 31884 28040 31890
rect 27988 31826 28040 31832
rect 27804 31816 27856 31822
rect 27856 31776 27936 31804
rect 27804 31758 27856 31764
rect 27528 31136 27580 31142
rect 27528 31078 27580 31084
rect 27540 30938 27568 31078
rect 27528 30932 27580 30938
rect 27528 30874 27580 30880
rect 27344 30864 27396 30870
rect 27344 30806 27396 30812
rect 27804 30796 27856 30802
rect 27804 30738 27856 30744
rect 27816 29850 27844 30738
rect 27344 29844 27396 29850
rect 27344 29786 27396 29792
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 27356 29714 27384 29786
rect 27344 29708 27396 29714
rect 27344 29650 27396 29656
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27252 28688 27304 28694
rect 27252 28630 27304 28636
rect 27264 28422 27292 28630
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 26884 27940 26936 27946
rect 26884 27882 26936 27888
rect 26332 27532 26384 27538
rect 26332 27474 26384 27480
rect 26146 26616 26202 26625
rect 26146 26551 26202 26560
rect 26160 26382 26188 26551
rect 26344 26518 26372 27474
rect 26516 27328 26568 27334
rect 26516 27270 26568 27276
rect 26608 27328 26660 27334
rect 26608 27270 26660 27276
rect 26528 27062 26556 27270
rect 26620 27130 26648 27270
rect 26608 27124 26660 27130
rect 26608 27066 26660 27072
rect 26516 27056 26568 27062
rect 26516 26998 26568 27004
rect 26896 26994 26924 27882
rect 26884 26988 26936 26994
rect 26884 26930 26936 26936
rect 26332 26512 26384 26518
rect 26332 26454 26384 26460
rect 26056 26376 26108 26382
rect 26056 26318 26108 26324
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26056 26240 26108 26246
rect 26056 26182 26108 26188
rect 25964 25900 26016 25906
rect 25964 25842 26016 25848
rect 26068 25226 26096 26182
rect 26252 25294 26280 26250
rect 26240 25288 26292 25294
rect 26240 25230 26292 25236
rect 26056 25220 26108 25226
rect 26056 25162 26108 25168
rect 26068 24970 26096 25162
rect 25884 24942 26096 24970
rect 25780 24200 25832 24206
rect 25780 24142 25832 24148
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 25792 22234 25820 22374
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 25410 21791 25466 21800
rect 25516 21814 25728 21842
rect 25424 17746 25452 21791
rect 25516 18222 25544 21814
rect 25686 21720 25742 21729
rect 25686 21655 25742 21664
rect 25700 21554 25728 21655
rect 25792 21554 25820 22170
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25780 21548 25832 21554
rect 25780 21490 25832 21496
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25688 19848 25740 19854
rect 25688 19790 25740 19796
rect 25608 19174 25636 19790
rect 25596 19168 25648 19174
rect 25596 19110 25648 19116
rect 25608 18834 25636 19110
rect 25700 18834 25728 19790
rect 25884 18834 25912 24942
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 26068 24410 26096 24754
rect 26056 24404 26108 24410
rect 26056 24346 26108 24352
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 26068 23730 26096 24006
rect 26056 23724 26108 23730
rect 26056 23666 26108 23672
rect 26068 22098 26096 23666
rect 26252 23254 26280 25230
rect 26976 25152 27028 25158
rect 26976 25094 27028 25100
rect 26988 24954 27016 25094
rect 26976 24948 27028 24954
rect 26976 24890 27028 24896
rect 26988 24750 27016 24890
rect 27252 24812 27304 24818
rect 27252 24754 27304 24760
rect 26976 24744 27028 24750
rect 27028 24692 27200 24698
rect 26976 24686 27200 24692
rect 26988 24670 27200 24686
rect 26608 24608 26660 24614
rect 26608 24550 26660 24556
rect 26700 24608 26752 24614
rect 26700 24550 26752 24556
rect 26976 24608 27028 24614
rect 26976 24550 27028 24556
rect 26620 24138 26648 24550
rect 26712 24342 26740 24550
rect 26988 24410 27016 24550
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 26700 24336 26752 24342
rect 26700 24278 26752 24284
rect 26712 24206 26740 24278
rect 26976 24268 27028 24274
rect 26976 24210 27028 24216
rect 26700 24200 26752 24206
rect 26700 24142 26752 24148
rect 26608 24132 26660 24138
rect 26608 24074 26660 24080
rect 26240 23248 26292 23254
rect 26240 23190 26292 23196
rect 26988 22506 27016 24210
rect 27068 24200 27120 24206
rect 27068 24142 27120 24148
rect 27080 23866 27108 24142
rect 27068 23860 27120 23866
rect 27068 23802 27120 23808
rect 27068 22568 27120 22574
rect 27068 22510 27120 22516
rect 26976 22500 27028 22506
rect 26976 22442 27028 22448
rect 26332 22228 26384 22234
rect 26332 22170 26384 22176
rect 25964 22092 26016 22098
rect 25964 22034 26016 22040
rect 26056 22092 26108 22098
rect 26056 22034 26108 22040
rect 25976 21865 26004 22034
rect 25962 21856 26018 21865
rect 25962 21791 26018 21800
rect 26068 21729 26096 22034
rect 26344 22030 26372 22170
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 26516 22024 26568 22030
rect 26516 21966 26568 21972
rect 26148 21888 26200 21894
rect 26148 21830 26200 21836
rect 26054 21720 26110 21729
rect 26054 21655 26110 21664
rect 25964 21548 26016 21554
rect 25964 21490 26016 21496
rect 25976 21146 26004 21490
rect 25964 21140 26016 21146
rect 25964 21082 26016 21088
rect 26056 21140 26108 21146
rect 26056 21082 26108 21088
rect 26068 20942 26096 21082
rect 26160 21078 26188 21830
rect 26528 21350 26556 21966
rect 26516 21344 26568 21350
rect 26516 21286 26568 21292
rect 26148 21072 26200 21078
rect 26148 21014 26200 21020
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 26240 20324 26292 20330
rect 26240 20266 26292 20272
rect 26252 19990 26280 20266
rect 26148 19984 26200 19990
rect 26148 19926 26200 19932
rect 26240 19984 26292 19990
rect 26240 19926 26292 19932
rect 25596 18828 25648 18834
rect 25596 18770 25648 18776
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25872 18828 25924 18834
rect 25872 18770 25924 18776
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 25884 18086 25912 18770
rect 26160 18086 26188 19926
rect 26332 19916 26384 19922
rect 26332 19858 26384 19864
rect 26344 18737 26372 19858
rect 26516 19848 26568 19854
rect 26516 19790 26568 19796
rect 26792 19848 26844 19854
rect 26844 19808 26924 19836
rect 26792 19790 26844 19796
rect 26424 18828 26476 18834
rect 26528 18816 26556 19790
rect 26792 19372 26844 19378
rect 26792 19314 26844 19320
rect 26476 18788 26556 18816
rect 26424 18770 26476 18776
rect 26330 18728 26386 18737
rect 26330 18663 26386 18672
rect 26240 18148 26292 18154
rect 26240 18090 26292 18096
rect 25872 18080 25924 18086
rect 25872 18022 25924 18028
rect 26148 18080 26200 18086
rect 26148 18022 26200 18028
rect 25412 17740 25464 17746
rect 25412 17682 25464 17688
rect 26252 17218 26280 18090
rect 26344 17338 26372 18663
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26332 17332 26384 17338
rect 26332 17274 26384 17280
rect 26436 17270 26464 17478
rect 26528 17338 26556 18788
rect 26608 18760 26660 18766
rect 26606 18728 26608 18737
rect 26700 18760 26752 18766
rect 26660 18728 26662 18737
rect 26700 18702 26752 18708
rect 26606 18663 26662 18672
rect 26712 18222 26740 18702
rect 26700 18216 26752 18222
rect 26700 18158 26752 18164
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26516 17332 26568 17338
rect 26516 17274 26568 17280
rect 26424 17264 26476 17270
rect 26252 17190 26372 17218
rect 26424 17206 26476 17212
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 25976 16590 26004 16934
rect 25964 16584 26016 16590
rect 25964 16526 26016 16532
rect 26344 16096 26372 17190
rect 26528 16590 26556 17274
rect 26620 16794 26648 17614
rect 26700 17536 26752 17542
rect 26700 17478 26752 17484
rect 26712 17134 26740 17478
rect 26804 17134 26832 19314
rect 26896 18154 26924 19808
rect 26884 18148 26936 18154
rect 26884 18090 26936 18096
rect 26884 17604 26936 17610
rect 26884 17546 26936 17552
rect 26896 17202 26924 17546
rect 26988 17542 27016 22442
rect 27080 22098 27108 22510
rect 27172 22506 27200 24670
rect 27264 24410 27292 24754
rect 27252 24404 27304 24410
rect 27252 24346 27304 24352
rect 27160 22500 27212 22506
rect 27160 22442 27212 22448
rect 27068 22092 27120 22098
rect 27356 22094 27384 29650
rect 27540 28626 27568 29650
rect 27528 28620 27580 28626
rect 27528 28562 27580 28568
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 27632 28082 27660 28358
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 27620 27464 27672 27470
rect 27620 27406 27672 27412
rect 27632 26994 27660 27406
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27908 24410 27936 31776
rect 27986 31240 28042 31249
rect 27986 31175 28042 31184
rect 28000 31142 28028 31175
rect 27988 31136 28040 31142
rect 27988 31078 28040 31084
rect 27988 30864 28040 30870
rect 27988 30806 28040 30812
rect 28000 30138 28028 30806
rect 28092 30258 28120 35022
rect 28356 34604 28408 34610
rect 28356 34546 28408 34552
rect 28540 34604 28592 34610
rect 28540 34546 28592 34552
rect 28368 32774 28396 34546
rect 28356 32768 28408 32774
rect 28356 32710 28408 32716
rect 28172 32360 28224 32366
rect 28172 32302 28224 32308
rect 28184 32026 28212 32302
rect 28172 32020 28224 32026
rect 28172 31962 28224 31968
rect 28368 31890 28396 32710
rect 28356 31884 28408 31890
rect 28356 31826 28408 31832
rect 28552 31754 28580 34546
rect 28736 34542 28764 35022
rect 28724 34536 28776 34542
rect 28724 34478 28776 34484
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 28460 31726 28580 31754
rect 28460 31346 28488 31726
rect 28264 31340 28316 31346
rect 28184 31300 28264 31328
rect 28080 30252 28132 30258
rect 28080 30194 28132 30200
rect 28000 30110 28120 30138
rect 27988 28212 28040 28218
rect 27988 28154 28040 28160
rect 28000 27946 28028 28154
rect 27988 27940 28040 27946
rect 27988 27882 28040 27888
rect 28000 27334 28028 27882
rect 27988 27328 28040 27334
rect 27988 27270 28040 27276
rect 27896 24404 27948 24410
rect 27896 24346 27948 24352
rect 27540 24274 27660 24290
rect 28092 24274 28120 30110
rect 28184 25226 28212 31300
rect 28264 31282 28316 31288
rect 28448 31340 28500 31346
rect 28448 31282 28500 31288
rect 28644 30734 28672 32166
rect 28632 30728 28684 30734
rect 28632 30670 28684 30676
rect 28264 30048 28316 30054
rect 28264 29990 28316 29996
rect 28356 30048 28408 30054
rect 28356 29990 28408 29996
rect 28276 29850 28304 29990
rect 28264 29844 28316 29850
rect 28264 29786 28316 29792
rect 28368 29510 28396 29990
rect 28356 29504 28408 29510
rect 28356 29446 28408 29452
rect 28540 28688 28592 28694
rect 28540 28630 28592 28636
rect 28262 28112 28318 28121
rect 28262 28047 28318 28056
rect 28448 28076 28500 28082
rect 28276 28014 28304 28047
rect 28448 28018 28500 28024
rect 28264 28008 28316 28014
rect 28264 27950 28316 27956
rect 28460 27674 28488 28018
rect 28448 27668 28500 27674
rect 28448 27610 28500 27616
rect 28552 27470 28580 28630
rect 28724 27872 28776 27878
rect 28724 27814 28776 27820
rect 28736 27470 28764 27814
rect 28540 27464 28592 27470
rect 28540 27406 28592 27412
rect 28724 27464 28776 27470
rect 28724 27406 28776 27412
rect 28540 26376 28592 26382
rect 28540 26318 28592 26324
rect 28172 25220 28224 25226
rect 28172 25162 28224 25168
rect 28356 24608 28408 24614
rect 28356 24550 28408 24556
rect 27528 24268 27660 24274
rect 27580 24262 27660 24268
rect 27528 24210 27580 24216
rect 27632 24188 27660 24262
rect 28080 24268 28132 24274
rect 28080 24210 28132 24216
rect 28368 24206 28396 24550
rect 27804 24200 27856 24206
rect 27632 24160 27752 24188
rect 27528 24132 27580 24138
rect 27580 24092 27660 24120
rect 27528 24074 27580 24080
rect 27632 23798 27660 24092
rect 27620 23792 27672 23798
rect 27620 23734 27672 23740
rect 27632 23610 27660 23734
rect 27724 23662 27752 24160
rect 27804 24142 27856 24148
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 27448 23582 27660 23610
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27816 23594 27844 24142
rect 28264 23724 28316 23730
rect 28368 23712 28396 24142
rect 28316 23684 28396 23712
rect 28264 23666 28316 23672
rect 27988 23656 28040 23662
rect 27986 23624 27988 23633
rect 28040 23624 28042 23633
rect 27448 23526 27476 23582
rect 27436 23520 27488 23526
rect 27436 23462 27488 23468
rect 27528 23520 27580 23526
rect 27528 23462 27580 23468
rect 27068 22034 27120 22040
rect 27172 22066 27384 22094
rect 27172 21418 27200 22066
rect 27344 21888 27396 21894
rect 27344 21830 27396 21836
rect 27356 21690 27384 21830
rect 27344 21684 27396 21690
rect 27344 21626 27396 21632
rect 27160 21412 27212 21418
rect 27160 21354 27212 21360
rect 27436 19712 27488 19718
rect 27436 19654 27488 19660
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 27172 18970 27200 19314
rect 27342 19000 27398 19009
rect 27160 18964 27212 18970
rect 27342 18935 27398 18944
rect 27160 18906 27212 18912
rect 27356 18834 27384 18935
rect 27344 18828 27396 18834
rect 27344 18770 27396 18776
rect 27448 18630 27476 19654
rect 27540 18698 27568 23462
rect 27632 22982 27660 23582
rect 27804 23588 27856 23594
rect 28552 23594 28580 26318
rect 28724 24812 28776 24818
rect 28724 24754 28776 24760
rect 28736 24410 28764 24754
rect 28632 24404 28684 24410
rect 28632 24346 28684 24352
rect 28724 24404 28776 24410
rect 28724 24346 28776 24352
rect 28644 24206 28672 24346
rect 28632 24200 28684 24206
rect 28632 24142 28684 24148
rect 27986 23559 28042 23568
rect 28540 23588 28592 23594
rect 27804 23530 27856 23536
rect 28540 23530 28592 23536
rect 28552 23497 28580 23530
rect 28538 23488 28594 23497
rect 28538 23423 28594 23432
rect 27712 23248 27764 23254
rect 27712 23190 27764 23196
rect 27620 22976 27672 22982
rect 27620 22918 27672 22924
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 27632 21894 27660 22578
rect 27620 21888 27672 21894
rect 27620 21830 27672 21836
rect 27620 19168 27672 19174
rect 27620 19110 27672 19116
rect 27632 18766 27660 19110
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27528 18692 27580 18698
rect 27528 18634 27580 18640
rect 27436 18624 27488 18630
rect 27436 18566 27488 18572
rect 26976 17536 27028 17542
rect 26976 17478 27028 17484
rect 26884 17196 26936 17202
rect 26884 17138 26936 17144
rect 26700 17128 26752 17134
rect 26700 17070 26752 17076
rect 26792 17128 26844 17134
rect 26792 17070 26844 17076
rect 26608 16788 26660 16794
rect 26608 16730 26660 16736
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26712 16250 26740 17070
rect 26700 16244 26752 16250
rect 26700 16186 26752 16192
rect 26516 16108 26568 16114
rect 26344 16068 26516 16096
rect 26516 16050 26568 16056
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 26056 15904 26108 15910
rect 26056 15846 26108 15852
rect 25228 14476 25280 14482
rect 25228 14418 25280 14424
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25412 14272 25464 14278
rect 25412 14214 25464 14220
rect 25424 14006 25452 14214
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 25608 13530 25636 14350
rect 25872 14340 25924 14346
rect 25872 14282 25924 14288
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 25504 13320 25556 13326
rect 25504 13262 25556 13268
rect 25148 12406 25268 12434
rect 24688 12294 24992 12322
rect 24688 12238 24716 12294
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 25044 12164 25096 12170
rect 25044 12106 25096 12112
rect 25056 11218 25084 12106
rect 25136 11280 25188 11286
rect 25136 11222 25188 11228
rect 25044 11212 25096 11218
rect 25044 11154 25096 11160
rect 25148 10742 25176 11222
rect 25136 10736 25188 10742
rect 25136 10678 25188 10684
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 24596 9574 24808 9602
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24596 9042 24624 9454
rect 24584 9036 24636 9042
rect 24584 8978 24636 8984
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 23664 8356 23716 8362
rect 23664 8298 23716 8304
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23400 5914 23428 7346
rect 23492 7342 23520 8230
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23940 7744 23992 7750
rect 23940 7686 23992 7692
rect 23664 7472 23716 7478
rect 23664 7414 23716 7420
rect 23480 7336 23532 7342
rect 23480 7278 23532 7284
rect 23676 6458 23704 7414
rect 23860 7410 23888 7686
rect 23952 7546 23980 7686
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 24228 6322 24256 7278
rect 24688 6866 24716 7346
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 23020 5908 23072 5914
rect 23020 5850 23072 5856
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22560 5704 22612 5710
rect 22664 5681 22692 5714
rect 22560 5646 22612 5652
rect 22650 5672 22706 5681
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 21732 4548 21784 4554
rect 21732 4490 21784 4496
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21100 3534 21128 3878
rect 21192 3738 21220 3878
rect 21180 3732 21232 3738
rect 21180 3674 21232 3680
rect 21376 3534 21404 4422
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 20916 3194 20944 3470
rect 21836 3466 21864 5102
rect 22572 4282 22600 5646
rect 22650 5607 22706 5616
rect 22652 5568 22704 5574
rect 22652 5510 22704 5516
rect 22192 4276 22244 4282
rect 22192 4218 22244 4224
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 22204 3738 22232 4218
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22376 3664 22428 3670
rect 22376 3606 22428 3612
rect 22388 3534 22416 3606
rect 22376 3528 22428 3534
rect 22376 3470 22428 3476
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21836 3058 21864 3402
rect 22480 3194 22508 4014
rect 22664 3398 22692 5510
rect 22836 5364 22888 5370
rect 22836 5306 22888 5312
rect 22848 4622 22876 5306
rect 23032 5098 23060 5850
rect 23480 5772 23532 5778
rect 23480 5714 23532 5720
rect 23492 5370 23520 5714
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23020 5092 23072 5098
rect 23020 5034 23072 5040
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 22744 3936 22796 3942
rect 22744 3878 22796 3884
rect 22756 3602 22784 3878
rect 23492 3738 23520 4082
rect 24032 4072 24084 4078
rect 24032 4014 24084 4020
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 22560 3392 22612 3398
rect 22560 3334 22612 3340
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 22572 2854 22600 3334
rect 22664 3194 22692 3334
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22848 2961 22876 3538
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 23124 3126 23152 3334
rect 23768 3126 23796 3878
rect 24044 3534 24072 4014
rect 24122 3632 24178 3641
rect 24122 3567 24124 3576
rect 24176 3567 24178 3576
rect 24124 3538 24176 3544
rect 24228 3534 24256 6258
rect 24504 5914 24532 6258
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24780 5370 24808 9574
rect 24952 9512 25004 9518
rect 24952 9454 25004 9460
rect 24964 9110 24992 9454
rect 24860 9104 24912 9110
rect 24860 9046 24912 9052
rect 24952 9104 25004 9110
rect 24952 9046 25004 9052
rect 25042 9072 25098 9081
rect 24872 6662 24900 9046
rect 25042 9007 25044 9016
rect 25096 9007 25098 9016
rect 25044 8978 25096 8984
rect 25148 8022 25176 9658
rect 25240 9586 25268 12406
rect 25516 12238 25544 13262
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25792 12442 25820 13126
rect 25780 12436 25832 12442
rect 25780 12378 25832 12384
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 25516 12102 25544 12174
rect 25884 12170 25912 14282
rect 25964 13388 26016 13394
rect 25964 13330 26016 13336
rect 25976 12850 26004 13330
rect 25964 12844 26016 12850
rect 25964 12786 26016 12792
rect 25964 12436 26016 12442
rect 25964 12378 26016 12384
rect 25872 12164 25924 12170
rect 25872 12106 25924 12112
rect 25504 12096 25556 12102
rect 25504 12038 25556 12044
rect 25976 11830 26004 12378
rect 25964 11824 26016 11830
rect 25964 11766 26016 11772
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25884 11286 25912 11494
rect 25872 11280 25924 11286
rect 25872 11222 25924 11228
rect 26068 11218 26096 15846
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 26344 15162 26372 15370
rect 26332 15156 26384 15162
rect 26332 15098 26384 15104
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26436 14618 26464 14962
rect 26528 14822 26556 16050
rect 26516 14816 26568 14822
rect 26516 14758 26568 14764
rect 26424 14612 26476 14618
rect 26424 14554 26476 14560
rect 26606 14512 26662 14521
rect 26606 14447 26608 14456
rect 26660 14447 26662 14456
rect 26608 14418 26660 14424
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 26160 13870 26188 14350
rect 26148 13864 26200 13870
rect 26148 13806 26200 13812
rect 26516 13728 26568 13734
rect 26516 13670 26568 13676
rect 26332 13456 26384 13462
rect 26332 13398 26384 13404
rect 26344 13190 26372 13398
rect 26528 13326 26556 13670
rect 26712 13394 26740 16186
rect 26804 15502 26832 17070
rect 26896 16658 26924 17138
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 27080 16114 27108 16390
rect 27724 16114 27752 23190
rect 28540 22704 28592 22710
rect 28540 22646 28592 22652
rect 28356 22568 28408 22574
rect 28356 22510 28408 22516
rect 28172 22500 28224 22506
rect 28172 22442 28224 22448
rect 27988 22432 28040 22438
rect 27988 22374 28040 22380
rect 27804 21956 27856 21962
rect 27804 21898 27856 21904
rect 27816 21690 27844 21898
rect 27804 21684 27856 21690
rect 27804 21626 27856 21632
rect 28000 21554 28028 22374
rect 28184 22234 28212 22442
rect 28172 22228 28224 22234
rect 28172 22170 28224 22176
rect 28080 22024 28132 22030
rect 28080 21966 28132 21972
rect 28092 21554 28120 21966
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 28080 21548 28132 21554
rect 28080 21490 28132 21496
rect 27896 20256 27948 20262
rect 27896 20198 27948 20204
rect 27908 19718 27936 20198
rect 27896 19712 27948 19718
rect 27896 19654 27948 19660
rect 27908 18834 27936 19654
rect 28184 19174 28212 22170
rect 28368 22030 28396 22510
rect 28356 22024 28408 22030
rect 28356 21966 28408 21972
rect 28552 21962 28580 22646
rect 28540 21956 28592 21962
rect 28540 21898 28592 21904
rect 28724 21888 28776 21894
rect 28724 21830 28776 21836
rect 28736 21622 28764 21830
rect 28724 21616 28776 21622
rect 28724 21558 28776 21564
rect 28540 19848 28592 19854
rect 28540 19790 28592 19796
rect 28172 19168 28224 19174
rect 28172 19110 28224 19116
rect 28184 18834 28212 19110
rect 27896 18828 27948 18834
rect 27896 18770 27948 18776
rect 28172 18828 28224 18834
rect 28172 18770 28224 18776
rect 28448 18692 28500 18698
rect 28448 18634 28500 18640
rect 28264 17740 28316 17746
rect 28264 17682 28316 17688
rect 28276 16114 28304 17682
rect 28460 16658 28488 18634
rect 28552 17134 28580 19790
rect 28632 19780 28684 19786
rect 28632 19722 28684 19728
rect 28644 19242 28672 19722
rect 28632 19236 28684 19242
rect 28632 19178 28684 19184
rect 28540 17128 28592 17134
rect 28540 17070 28592 17076
rect 28448 16652 28500 16658
rect 28448 16594 28500 16600
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 27712 16108 27764 16114
rect 27712 16050 27764 16056
rect 27896 16108 27948 16114
rect 27896 16050 27948 16056
rect 28264 16108 28316 16114
rect 28264 16050 28316 16056
rect 27712 15972 27764 15978
rect 27712 15914 27764 15920
rect 26792 15496 26844 15502
rect 26792 15438 26844 15444
rect 27344 15360 27396 15366
rect 27344 15302 27396 15308
rect 27356 15026 27384 15302
rect 27344 15020 27396 15026
rect 27344 14962 27396 14968
rect 26884 14952 26936 14958
rect 26884 14894 26936 14900
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 26896 14414 26924 14894
rect 26976 14476 27028 14482
rect 27028 14436 27108 14464
rect 26976 14418 27028 14424
rect 26884 14408 26936 14414
rect 26884 14350 26936 14356
rect 26896 13938 26924 14350
rect 26976 14272 27028 14278
rect 26976 14214 27028 14220
rect 26884 13932 26936 13938
rect 26884 13874 26936 13880
rect 26988 13870 27016 14214
rect 26976 13864 27028 13870
rect 26976 13806 27028 13812
rect 26700 13388 26752 13394
rect 26700 13330 26752 13336
rect 26516 13320 26568 13326
rect 26516 13262 26568 13268
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 26988 12152 27016 13806
rect 27080 13734 27108 14436
rect 27160 14408 27212 14414
rect 27158 14376 27160 14385
rect 27212 14376 27214 14385
rect 27158 14311 27214 14320
rect 27160 14272 27212 14278
rect 27160 14214 27212 14220
rect 27172 14006 27200 14214
rect 27160 14000 27212 14006
rect 27160 13942 27212 13948
rect 27160 13864 27212 13870
rect 27160 13806 27212 13812
rect 27068 13728 27120 13734
rect 27068 13670 27120 13676
rect 27172 13530 27200 13806
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 27448 13462 27476 14894
rect 27528 14476 27580 14482
rect 27528 14418 27580 14424
rect 27436 13456 27488 13462
rect 27436 13398 27488 13404
rect 27540 13326 27568 14418
rect 27724 13802 27752 15914
rect 27804 14884 27856 14890
rect 27804 14826 27856 14832
rect 27816 14618 27844 14826
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27712 13796 27764 13802
rect 27712 13738 27764 13744
rect 27528 13320 27580 13326
rect 27528 13262 27580 13268
rect 27252 12164 27304 12170
rect 26988 12124 27252 12152
rect 27252 12106 27304 12112
rect 26700 12096 26752 12102
rect 26700 12038 26752 12044
rect 26792 12096 26844 12102
rect 26792 12038 26844 12044
rect 26712 11898 26740 12038
rect 26700 11892 26752 11898
rect 26700 11834 26752 11840
rect 26804 11762 26832 12038
rect 27264 11812 27292 12106
rect 27264 11784 27384 11812
rect 26792 11756 26844 11762
rect 26792 11698 26844 11704
rect 27356 11558 27384 11784
rect 27540 11762 27568 13262
rect 27712 13252 27764 13258
rect 27632 13212 27712 13240
rect 27632 12714 27660 13212
rect 27712 13194 27764 13200
rect 27710 12880 27766 12889
rect 27710 12815 27712 12824
rect 27764 12815 27766 12824
rect 27712 12786 27764 12792
rect 27804 12776 27856 12782
rect 27804 12718 27856 12724
rect 27620 12708 27672 12714
rect 27620 12650 27672 12656
rect 27528 11756 27580 11762
rect 27528 11698 27580 11704
rect 27252 11552 27304 11558
rect 27252 11494 27304 11500
rect 27344 11552 27396 11558
rect 27344 11494 27396 11500
rect 26332 11280 26384 11286
rect 26332 11222 26384 11228
rect 26056 11212 26108 11218
rect 26056 11154 26108 11160
rect 25872 11144 25924 11150
rect 25410 11112 25466 11121
rect 25872 11086 25924 11092
rect 25410 11047 25412 11056
rect 25464 11047 25466 11056
rect 25412 11018 25464 11024
rect 25884 11014 25912 11086
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 26240 11008 26292 11014
rect 26240 10950 26292 10956
rect 26252 10198 26280 10950
rect 26240 10192 26292 10198
rect 26240 10134 26292 10140
rect 26344 9654 26372 11222
rect 26332 9648 26384 9654
rect 26332 9590 26384 9596
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 26792 9580 26844 9586
rect 26792 9522 26844 9528
rect 25412 9512 25464 9518
rect 25412 9454 25464 9460
rect 25424 8974 25452 9454
rect 26804 9178 26832 9522
rect 26792 9172 26844 9178
rect 26792 9114 26844 9120
rect 27264 9042 27292 11494
rect 27436 11076 27488 11082
rect 27436 11018 27488 11024
rect 25964 9036 26016 9042
rect 25964 8978 26016 8984
rect 27252 9036 27304 9042
rect 27252 8978 27304 8984
rect 25412 8968 25464 8974
rect 25596 8968 25648 8974
rect 25412 8910 25464 8916
rect 25594 8936 25596 8945
rect 25648 8936 25650 8945
rect 25136 8016 25188 8022
rect 25136 7958 25188 7964
rect 25424 7546 25452 8910
rect 25594 8871 25650 8880
rect 25976 8634 26004 8978
rect 26240 8832 26292 8838
rect 26240 8774 26292 8780
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 25608 6458 25636 8570
rect 26252 7886 26280 8774
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 26528 7478 26556 7890
rect 26792 7744 26844 7750
rect 26792 7686 26844 7692
rect 27160 7744 27212 7750
rect 27160 7686 27212 7692
rect 26516 7472 26568 7478
rect 26516 7414 26568 7420
rect 26240 7268 26292 7274
rect 26240 7210 26292 7216
rect 26148 6656 26200 6662
rect 26148 6598 26200 6604
rect 25596 6452 25648 6458
rect 25596 6394 25648 6400
rect 24860 5908 24912 5914
rect 24860 5850 24912 5856
rect 24872 5642 24900 5850
rect 24952 5840 25004 5846
rect 24952 5782 25004 5788
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 24964 5574 24992 5782
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 25044 5636 25096 5642
rect 25044 5578 25096 5584
rect 24952 5568 25004 5574
rect 24952 5510 25004 5516
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24952 5160 25004 5166
rect 24952 5102 25004 5108
rect 24964 4690 24992 5102
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 24860 4480 24912 4486
rect 24860 4422 24912 4428
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 23112 3120 23164 3126
rect 23112 3062 23164 3068
rect 23756 3120 23808 3126
rect 23756 3062 23808 3068
rect 24228 3058 24256 3470
rect 24872 3398 24900 4422
rect 25056 4078 25084 5578
rect 25148 4554 25176 5646
rect 25608 5642 25636 6394
rect 26160 6322 26188 6598
rect 25964 6316 26016 6322
rect 25964 6258 26016 6264
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 25780 5840 25832 5846
rect 25780 5782 25832 5788
rect 25596 5636 25648 5642
rect 25596 5578 25648 5584
rect 25792 4826 25820 5782
rect 25976 5574 26004 6258
rect 26252 5914 26280 7210
rect 26516 6724 26568 6730
rect 26516 6666 26568 6672
rect 26424 6656 26476 6662
rect 26424 6598 26476 6604
rect 26436 6458 26464 6598
rect 26528 6458 26556 6666
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 26516 6452 26568 6458
rect 26516 6394 26568 6400
rect 26700 6316 26752 6322
rect 26700 6258 26752 6264
rect 26712 6186 26740 6258
rect 26700 6180 26752 6186
rect 26700 6122 26752 6128
rect 26240 5908 26292 5914
rect 26240 5850 26292 5856
rect 25964 5568 26016 5574
rect 25964 5510 26016 5516
rect 26804 5370 26832 7686
rect 27172 7410 27200 7686
rect 27160 7404 27212 7410
rect 27160 7346 27212 7352
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 27080 6798 27108 7278
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 27264 6798 27292 7142
rect 27068 6792 27120 6798
rect 27068 6734 27120 6740
rect 27252 6792 27304 6798
rect 27252 6734 27304 6740
rect 27080 6458 27108 6734
rect 27068 6452 27120 6458
rect 27068 6394 27120 6400
rect 27344 6384 27396 6390
rect 27344 6326 27396 6332
rect 27356 6118 27384 6326
rect 27344 6112 27396 6118
rect 27344 6054 27396 6060
rect 26148 5364 26200 5370
rect 26148 5306 26200 5312
rect 26792 5364 26844 5370
rect 26792 5306 26844 5312
rect 26160 5234 26188 5306
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 25872 5160 25924 5166
rect 25872 5102 25924 5108
rect 26056 5160 26108 5166
rect 26056 5102 26108 5108
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 25884 4690 25912 5102
rect 25964 5024 26016 5030
rect 25964 4966 26016 4972
rect 25976 4758 26004 4966
rect 25964 4752 26016 4758
rect 25964 4694 26016 4700
rect 25596 4684 25648 4690
rect 25596 4626 25648 4632
rect 25872 4684 25924 4690
rect 25872 4626 25924 4632
rect 25136 4548 25188 4554
rect 25136 4490 25188 4496
rect 25044 4072 25096 4078
rect 25044 4014 25096 4020
rect 24952 3460 25004 3466
rect 24952 3402 25004 3408
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24872 3194 24900 3334
rect 24964 3194 24992 3402
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 24952 3188 25004 3194
rect 24952 3130 25004 3136
rect 24216 3052 24268 3058
rect 24216 2994 24268 3000
rect 25056 2990 25084 4014
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 25148 3058 25176 3878
rect 25608 3398 25636 4626
rect 25884 4282 25912 4626
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 25976 4282 26004 4558
rect 26068 4486 26096 5102
rect 27448 4758 27476 11018
rect 27816 10130 27844 12718
rect 27804 10124 27856 10130
rect 27804 10066 27856 10072
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27724 9722 27752 9998
rect 27712 9716 27764 9722
rect 27712 9658 27764 9664
rect 27528 9648 27580 9654
rect 27528 9590 27580 9596
rect 27540 9178 27568 9590
rect 27816 9466 27844 10066
rect 27724 9438 27844 9466
rect 27724 9382 27752 9438
rect 27712 9376 27764 9382
rect 27712 9318 27764 9324
rect 27908 9194 27936 16050
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 28184 15094 28212 15846
rect 28172 15088 28224 15094
rect 28172 15030 28224 15036
rect 28184 13938 28212 15030
rect 28172 13932 28224 13938
rect 28172 13874 28224 13880
rect 27988 13864 28040 13870
rect 27988 13806 28040 13812
rect 28000 13734 28028 13806
rect 27988 13728 28040 13734
rect 27988 13670 28040 13676
rect 28276 9450 28304 16050
rect 28460 15910 28488 16594
rect 28448 15904 28500 15910
rect 28448 15846 28500 15852
rect 28460 14958 28488 15846
rect 28632 15020 28684 15026
rect 28632 14962 28684 14968
rect 28448 14952 28500 14958
rect 28448 14894 28500 14900
rect 28644 14618 28672 14962
rect 28632 14612 28684 14618
rect 28632 14554 28684 14560
rect 28632 14272 28684 14278
rect 28632 14214 28684 14220
rect 28644 12782 28672 14214
rect 28724 13864 28776 13870
rect 28724 13806 28776 13812
rect 28736 13530 28764 13806
rect 28724 13524 28776 13530
rect 28724 13466 28776 13472
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 28632 12776 28684 12782
rect 28632 12718 28684 12724
rect 28736 11558 28764 13126
rect 28724 11552 28776 11558
rect 28724 11494 28776 11500
rect 28264 9444 28316 9450
rect 28264 9386 28316 9392
rect 27528 9172 27580 9178
rect 27528 9114 27580 9120
rect 27816 9166 27936 9194
rect 27540 9042 27568 9114
rect 27816 9042 27844 9166
rect 28276 9110 28304 9386
rect 28356 9376 28408 9382
rect 28356 9318 28408 9324
rect 28264 9104 28316 9110
rect 28264 9046 28316 9052
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27540 5914 27568 8774
rect 27816 7954 27844 8978
rect 28368 8974 28396 9318
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 27804 7948 27856 7954
rect 27804 7890 27856 7896
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28552 7002 28580 7822
rect 28540 6996 28592 7002
rect 28540 6938 28592 6944
rect 27528 5908 27580 5914
rect 27528 5850 27580 5856
rect 27540 5370 27568 5850
rect 28632 5772 28684 5778
rect 28632 5714 28684 5720
rect 27528 5364 27580 5370
rect 27528 5306 27580 5312
rect 27988 5160 28040 5166
rect 27988 5102 28040 5108
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27436 4752 27488 4758
rect 27436 4694 27488 4700
rect 26608 4616 26660 4622
rect 26608 4558 26660 4564
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 26620 4486 26648 4558
rect 26056 4480 26108 4486
rect 26056 4422 26108 4428
rect 26608 4480 26660 4486
rect 26608 4422 26660 4428
rect 27344 4480 27396 4486
rect 27344 4422 27396 4428
rect 25872 4276 25924 4282
rect 25872 4218 25924 4224
rect 25964 4276 26016 4282
rect 25964 4218 26016 4224
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25596 3392 25648 3398
rect 25596 3334 25648 3340
rect 25608 3126 25636 3334
rect 25792 3194 25820 4082
rect 25884 3738 25912 4218
rect 27356 4214 27384 4422
rect 27448 4214 27476 4558
rect 27344 4208 27396 4214
rect 27344 4150 27396 4156
rect 27436 4208 27488 4214
rect 27436 4150 27488 4156
rect 26056 3936 26108 3942
rect 26056 3878 26108 3884
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 26068 3534 26096 3878
rect 27448 3738 27476 4150
rect 27540 4146 27568 4966
rect 27620 4548 27672 4554
rect 27620 4490 27672 4496
rect 27528 4140 27580 4146
rect 27528 4082 27580 4088
rect 27632 4010 27660 4490
rect 28000 4282 28028 5102
rect 27988 4276 28040 4282
rect 27988 4218 28040 4224
rect 28644 4146 28672 5714
rect 28632 4140 28684 4146
rect 28632 4082 28684 4088
rect 27620 4004 27672 4010
rect 27620 3946 27672 3952
rect 27436 3732 27488 3738
rect 27436 3674 27488 3680
rect 26056 3528 26108 3534
rect 26056 3470 26108 3476
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 25780 3188 25832 3194
rect 25780 3130 25832 3136
rect 26332 3188 26384 3194
rect 26332 3130 26384 3136
rect 25596 3120 25648 3126
rect 25596 3062 25648 3068
rect 25136 3052 25188 3058
rect 25136 2994 25188 3000
rect 26344 2990 26372 3130
rect 27632 3126 27660 3470
rect 27620 3120 27672 3126
rect 27620 3062 27672 3068
rect 28644 3058 28672 4082
rect 28632 3052 28684 3058
rect 28632 2994 28684 3000
rect 25044 2984 25096 2990
rect 22834 2952 22890 2961
rect 26332 2984 26384 2990
rect 25044 2926 25096 2932
rect 26330 2952 26332 2961
rect 26384 2952 26386 2961
rect 22834 2887 22890 2896
rect 26330 2887 26386 2896
rect 22468 2848 22520 2854
rect 22468 2790 22520 2796
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 20732 2746 20852 2774
rect 20732 2514 20760 2746
rect 20994 2680 21050 2689
rect 22480 2666 22508 2790
rect 22848 2666 22876 2887
rect 28632 2848 28684 2854
rect 28828 2836 28856 42570
rect 29472 42294 29500 42638
rect 29932 42566 29960 43250
rect 30012 43172 30064 43178
rect 30012 43114 30064 43120
rect 30024 42906 30052 43114
rect 30012 42900 30064 42906
rect 30012 42842 30064 42848
rect 29552 42560 29604 42566
rect 29552 42502 29604 42508
rect 29920 42560 29972 42566
rect 29920 42502 29972 42508
rect 29460 42288 29512 42294
rect 29460 42230 29512 42236
rect 29564 42226 29592 42502
rect 30024 42294 30052 42842
rect 30208 42838 30236 43862
rect 30300 43772 30328 44338
rect 30472 43784 30524 43790
rect 30300 43744 30472 43772
rect 30472 43726 30524 43732
rect 30380 43648 30432 43654
rect 30380 43590 30432 43596
rect 30392 43450 30420 43590
rect 30288 43444 30340 43450
rect 30288 43386 30340 43392
rect 30380 43444 30432 43450
rect 30380 43386 30432 43392
rect 30300 43092 30328 43386
rect 30380 43104 30432 43110
rect 30300 43064 30380 43092
rect 30196 42832 30248 42838
rect 30196 42774 30248 42780
rect 30300 42702 30328 43064
rect 30380 43046 30432 43052
rect 30484 42770 30512 43726
rect 30668 43450 30696 44639
rect 30852 43722 30880 45902
rect 31116 45484 31168 45490
rect 31116 45426 31168 45432
rect 31024 45280 31076 45286
rect 31024 45222 31076 45228
rect 31036 45082 31064 45222
rect 31128 45082 31156 45426
rect 31576 45280 31628 45286
rect 31576 45222 31628 45228
rect 31024 45076 31076 45082
rect 31024 45018 31076 45024
rect 31116 45076 31168 45082
rect 31116 45018 31168 45024
rect 31588 45014 31616 45222
rect 31576 45008 31628 45014
rect 31576 44950 31628 44956
rect 31300 44872 31352 44878
rect 31300 44814 31352 44820
rect 31668 44872 31720 44878
rect 31720 44832 31800 44860
rect 31668 44814 31720 44820
rect 31312 44742 31340 44814
rect 31300 44736 31352 44742
rect 31300 44678 31352 44684
rect 31312 44334 31340 44678
rect 31772 44538 31800 44832
rect 31760 44532 31812 44538
rect 31760 44474 31812 44480
rect 31300 44328 31352 44334
rect 31300 44270 31352 44276
rect 32036 43784 32088 43790
rect 32036 43726 32088 43732
rect 30840 43716 30892 43722
rect 30840 43658 30892 43664
rect 30748 43648 30800 43654
rect 30748 43590 30800 43596
rect 30656 43444 30708 43450
rect 30656 43386 30708 43392
rect 30760 43314 30788 43590
rect 30838 43480 30894 43489
rect 30838 43415 30894 43424
rect 30852 43382 30880 43415
rect 30840 43376 30892 43382
rect 30840 43318 30892 43324
rect 32048 43314 32076 43726
rect 30748 43308 30800 43314
rect 30748 43250 30800 43256
rect 32036 43308 32088 43314
rect 32036 43250 32088 43256
rect 30472 42764 30524 42770
rect 30472 42706 30524 42712
rect 30288 42696 30340 42702
rect 30288 42638 30340 42644
rect 30196 42628 30248 42634
rect 30196 42570 30248 42576
rect 30012 42288 30064 42294
rect 30012 42230 30064 42236
rect 29552 42220 29604 42226
rect 29552 42162 29604 42168
rect 29920 42220 29972 42226
rect 29920 42162 29972 42168
rect 29932 41546 29960 42162
rect 30208 42090 30236 42570
rect 30840 42560 30892 42566
rect 30840 42502 30892 42508
rect 30852 42226 30880 42502
rect 31668 42356 31720 42362
rect 31588 42316 31668 42344
rect 30840 42220 30892 42226
rect 30840 42162 30892 42168
rect 30196 42084 30248 42090
rect 30196 42026 30248 42032
rect 29920 41540 29972 41546
rect 29920 41482 29972 41488
rect 30208 41478 30236 42026
rect 31588 41546 31616 42316
rect 31668 42298 31720 42304
rect 32048 42158 32076 43250
rect 32128 42696 32180 42702
rect 32128 42638 32180 42644
rect 32036 42152 32088 42158
rect 32036 42094 32088 42100
rect 31668 42016 31720 42022
rect 31668 41958 31720 41964
rect 31680 41546 31708 41958
rect 32140 41818 32168 42638
rect 32128 41812 32180 41818
rect 32128 41754 32180 41760
rect 31852 41608 31904 41614
rect 32036 41608 32088 41614
rect 31904 41556 32036 41562
rect 31852 41550 32088 41556
rect 31576 41540 31628 41546
rect 31576 41482 31628 41488
rect 31668 41540 31720 41546
rect 31864 41534 32076 41550
rect 31668 41482 31720 41488
rect 30196 41472 30248 41478
rect 30196 41414 30248 41420
rect 29368 40520 29420 40526
rect 29368 40462 29420 40468
rect 30932 40520 30984 40526
rect 30932 40462 30984 40468
rect 28908 40384 28960 40390
rect 28908 40326 28960 40332
rect 28920 40118 28948 40326
rect 29380 40186 29408 40462
rect 30564 40452 30616 40458
rect 30564 40394 30616 40400
rect 30576 40186 30604 40394
rect 29368 40180 29420 40186
rect 29368 40122 29420 40128
rect 30564 40180 30616 40186
rect 30564 40122 30616 40128
rect 28908 40112 28960 40118
rect 28908 40054 28960 40060
rect 29736 40044 29788 40050
rect 29736 39986 29788 39992
rect 29000 39908 29052 39914
rect 29000 39850 29052 39856
rect 29012 37754 29040 39850
rect 29748 39574 29776 39986
rect 30012 39976 30064 39982
rect 30012 39918 30064 39924
rect 30024 39642 30052 39918
rect 30012 39636 30064 39642
rect 30012 39578 30064 39584
rect 30840 39636 30892 39642
rect 30840 39578 30892 39584
rect 29736 39568 29788 39574
rect 29736 39510 29788 39516
rect 29092 39500 29144 39506
rect 29092 39442 29144 39448
rect 29104 39302 29132 39442
rect 29092 39296 29144 39302
rect 29092 39238 29144 39244
rect 29748 39030 29776 39510
rect 29736 39024 29788 39030
rect 29736 38966 29788 38972
rect 29920 38752 29972 38758
rect 29920 38694 29972 38700
rect 29828 38276 29880 38282
rect 29828 38218 29880 38224
rect 29840 38010 29868 38218
rect 29828 38004 29880 38010
rect 29828 37946 29880 37952
rect 29932 37874 29960 38694
rect 29920 37868 29972 37874
rect 29920 37810 29972 37816
rect 28920 37726 29040 37754
rect 28920 37670 28948 37726
rect 28908 37664 28960 37670
rect 28908 37606 28960 37612
rect 29000 37664 29052 37670
rect 29000 37606 29052 37612
rect 29920 37664 29972 37670
rect 29920 37606 29972 37612
rect 28908 35624 28960 35630
rect 29012 35612 29040 37606
rect 29184 37324 29236 37330
rect 29184 37266 29236 37272
rect 29092 36372 29144 36378
rect 29092 36314 29144 36320
rect 29104 35698 29132 36314
rect 29092 35692 29144 35698
rect 29092 35634 29144 35640
rect 28960 35584 29040 35612
rect 28908 35566 28960 35572
rect 29000 35488 29052 35494
rect 29000 35430 29052 35436
rect 28906 35184 28962 35193
rect 28906 35119 28962 35128
rect 28920 35086 28948 35119
rect 29012 35086 29040 35430
rect 29104 35290 29132 35634
rect 29092 35284 29144 35290
rect 29092 35226 29144 35232
rect 28908 35080 28960 35086
rect 28908 35022 28960 35028
rect 29000 35080 29052 35086
rect 29000 35022 29052 35028
rect 29092 35080 29144 35086
rect 29092 35022 29144 35028
rect 29104 34746 29132 35022
rect 29092 34740 29144 34746
rect 29092 34682 29144 34688
rect 29092 34604 29144 34610
rect 29092 34546 29144 34552
rect 29000 33040 29052 33046
rect 29000 32982 29052 32988
rect 29012 32065 29040 32982
rect 28998 32056 29054 32065
rect 28998 31991 29054 32000
rect 28908 31952 28960 31958
rect 28908 31894 28960 31900
rect 28920 29646 28948 31894
rect 29000 31680 29052 31686
rect 29000 31622 29052 31628
rect 29012 31210 29040 31622
rect 29104 31346 29132 34546
rect 29196 34474 29224 37266
rect 29932 37262 29960 37606
rect 29920 37256 29972 37262
rect 29920 37198 29972 37204
rect 29276 36644 29328 36650
rect 29276 36586 29328 36592
rect 29288 36174 29316 36586
rect 29276 36168 29328 36174
rect 29276 36110 29328 36116
rect 29460 36100 29512 36106
rect 29460 36042 29512 36048
rect 29276 35284 29328 35290
rect 29276 35226 29328 35232
rect 29184 34468 29236 34474
rect 29184 34410 29236 34416
rect 29288 33590 29316 35226
rect 29276 33584 29328 33590
rect 29276 33526 29328 33532
rect 29288 32858 29316 33526
rect 29196 32830 29316 32858
rect 29196 32570 29224 32830
rect 29276 32768 29328 32774
rect 29276 32710 29328 32716
rect 29368 32768 29420 32774
rect 29368 32710 29420 32716
rect 29184 32564 29236 32570
rect 29184 32506 29236 32512
rect 29184 32428 29236 32434
rect 29184 32370 29236 32376
rect 29196 32026 29224 32370
rect 29184 32020 29236 32026
rect 29184 31962 29236 31968
rect 29288 31890 29316 32710
rect 29276 31884 29328 31890
rect 29276 31826 29328 31832
rect 29380 31822 29408 32710
rect 29368 31816 29420 31822
rect 29368 31758 29420 31764
rect 29092 31340 29144 31346
rect 29092 31282 29144 31288
rect 29000 31204 29052 31210
rect 29000 31146 29052 31152
rect 29104 30666 29132 31282
rect 29092 30660 29144 30666
rect 29092 30602 29144 30608
rect 29472 29646 29500 36042
rect 29552 35692 29604 35698
rect 29552 35634 29604 35640
rect 29564 35290 29592 35634
rect 29736 35488 29788 35494
rect 29736 35430 29788 35436
rect 29552 35284 29604 35290
rect 29552 35226 29604 35232
rect 29748 35086 29776 35430
rect 29736 35080 29788 35086
rect 29736 35022 29788 35028
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 29552 34944 29604 34950
rect 29552 34886 29604 34892
rect 29736 34944 29788 34950
rect 29736 34886 29788 34892
rect 29564 34610 29592 34886
rect 29748 34746 29776 34886
rect 29736 34740 29788 34746
rect 29736 34682 29788 34688
rect 29932 34610 29960 35022
rect 29552 34604 29604 34610
rect 29552 34546 29604 34552
rect 29736 34604 29788 34610
rect 29736 34546 29788 34552
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 29748 34490 29776 34546
rect 29748 34462 29868 34490
rect 29734 33960 29790 33969
rect 29734 33895 29790 33904
rect 29644 32972 29696 32978
rect 29644 32914 29696 32920
rect 29552 32496 29604 32502
rect 29552 32438 29604 32444
rect 29564 31822 29592 32438
rect 29656 32230 29684 32914
rect 29644 32224 29696 32230
rect 29644 32166 29696 32172
rect 29552 31816 29604 31822
rect 29552 31758 29604 31764
rect 29748 31754 29776 33895
rect 29656 31726 29776 31754
rect 29656 30138 29684 31726
rect 29736 30592 29788 30598
rect 29736 30534 29788 30540
rect 29748 30258 29776 30534
rect 29736 30252 29788 30258
rect 29736 30194 29788 30200
rect 29656 30110 29776 30138
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 29092 29640 29144 29646
rect 29092 29582 29144 29588
rect 29460 29640 29512 29646
rect 29460 29582 29512 29588
rect 29104 28558 29132 29582
rect 29552 29504 29604 29510
rect 29552 29446 29604 29452
rect 29564 29170 29592 29446
rect 29368 29164 29420 29170
rect 29368 29106 29420 29112
rect 29552 29164 29604 29170
rect 29552 29106 29604 29112
rect 29644 29164 29696 29170
rect 29644 29106 29696 29112
rect 29380 29073 29408 29106
rect 29460 29096 29512 29102
rect 29366 29064 29422 29073
rect 29460 29038 29512 29044
rect 29366 28999 29422 29008
rect 29472 28762 29500 29038
rect 29460 28756 29512 28762
rect 29460 28698 29512 28704
rect 29092 28552 29144 28558
rect 29092 28494 29144 28500
rect 29000 28484 29052 28490
rect 29000 28426 29052 28432
rect 29184 28484 29236 28490
rect 29184 28426 29236 28432
rect 29012 28393 29040 28426
rect 28998 28384 29054 28393
rect 28998 28319 29054 28328
rect 29012 27985 29040 28319
rect 29196 28218 29224 28426
rect 29184 28212 29236 28218
rect 29184 28154 29236 28160
rect 28998 27976 29054 27985
rect 28998 27911 29054 27920
rect 29000 27872 29052 27878
rect 29000 27814 29052 27820
rect 29012 26790 29040 27814
rect 29092 27532 29144 27538
rect 29092 27474 29144 27480
rect 29104 26994 29132 27474
rect 29564 27470 29592 29106
rect 29656 28422 29684 29106
rect 29644 28416 29696 28422
rect 29644 28358 29696 28364
rect 29656 28218 29684 28358
rect 29644 28212 29696 28218
rect 29644 28154 29696 28160
rect 29644 27600 29696 27606
rect 29644 27542 29696 27548
rect 29552 27464 29604 27470
rect 29552 27406 29604 27412
rect 29184 27396 29236 27402
rect 29184 27338 29236 27344
rect 29196 27305 29224 27338
rect 29182 27296 29238 27305
rect 29182 27231 29238 27240
rect 29276 27124 29328 27130
rect 29276 27066 29328 27072
rect 29092 26988 29144 26994
rect 29092 26930 29144 26936
rect 29000 26784 29052 26790
rect 29000 26726 29052 26732
rect 28908 25492 28960 25498
rect 28908 25434 28960 25440
rect 28920 24426 28948 25434
rect 29092 24744 29144 24750
rect 29092 24686 29144 24692
rect 29104 24585 29132 24686
rect 29090 24576 29146 24585
rect 29090 24511 29146 24520
rect 28920 24398 29224 24426
rect 29092 24336 29144 24342
rect 29092 24278 29144 24284
rect 29000 24268 29052 24274
rect 29000 24210 29052 24216
rect 28908 23724 28960 23730
rect 29012 23712 29040 24210
rect 29104 23866 29132 24278
rect 29196 24274 29224 24398
rect 29184 24268 29236 24274
rect 29184 24210 29236 24216
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 28960 23684 29040 23712
rect 28908 23666 28960 23672
rect 29092 23656 29144 23662
rect 29144 23616 29224 23644
rect 29092 23598 29144 23604
rect 29092 22636 29144 22642
rect 29092 22578 29144 22584
rect 28908 22432 28960 22438
rect 28908 22374 28960 22380
rect 28920 22030 28948 22374
rect 28908 22024 28960 22030
rect 28908 21966 28960 21972
rect 28908 19984 28960 19990
rect 28908 19926 28960 19932
rect 28920 19378 28948 19926
rect 29104 19922 29132 22578
rect 29000 19916 29052 19922
rect 29000 19858 29052 19864
rect 29092 19916 29144 19922
rect 29092 19858 29144 19864
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 29012 17626 29040 19858
rect 29196 18329 29224 23616
rect 29288 21865 29316 27066
rect 29564 26874 29592 27406
rect 29656 26926 29684 27542
rect 29748 27130 29776 30110
rect 29840 27418 29868 34462
rect 30024 33114 30052 39578
rect 30196 39500 30248 39506
rect 30196 39442 30248 39448
rect 30208 34066 30236 39442
rect 30852 39438 30880 39578
rect 30944 39506 30972 40462
rect 31760 40384 31812 40390
rect 31760 40326 31812 40332
rect 31772 40186 31800 40326
rect 31760 40180 31812 40186
rect 31760 40122 31812 40128
rect 31482 40080 31538 40089
rect 31482 40015 31538 40024
rect 31392 39976 31444 39982
rect 31392 39918 31444 39924
rect 31300 39840 31352 39846
rect 31300 39782 31352 39788
rect 30932 39500 30984 39506
rect 30984 39460 31064 39488
rect 30932 39442 30984 39448
rect 30748 39432 30800 39438
rect 30748 39374 30800 39380
rect 30840 39432 30892 39438
rect 30840 39374 30892 39380
rect 30760 39302 30788 39374
rect 30748 39296 30800 39302
rect 30748 39238 30800 39244
rect 30288 39024 30340 39030
rect 30288 38966 30340 38972
rect 30300 38010 30328 38966
rect 30932 38956 30984 38962
rect 30932 38898 30984 38904
rect 30944 38554 30972 38898
rect 30932 38548 30984 38554
rect 30932 38490 30984 38496
rect 30288 38004 30340 38010
rect 30288 37946 30340 37952
rect 30300 36854 30328 37946
rect 30748 37868 30800 37874
rect 30748 37810 30800 37816
rect 30760 37466 30788 37810
rect 30748 37460 30800 37466
rect 30748 37402 30800 37408
rect 30288 36848 30340 36854
rect 30288 36790 30340 36796
rect 30300 35698 30328 36790
rect 30288 35692 30340 35698
rect 30288 35634 30340 35640
rect 30564 35556 30616 35562
rect 30564 35498 30616 35504
rect 30576 35154 30604 35498
rect 30656 35216 30708 35222
rect 30760 35204 30788 37402
rect 30944 36666 30972 38490
rect 31036 38418 31064 39460
rect 31312 39030 31340 39782
rect 31208 39024 31260 39030
rect 31208 38966 31260 38972
rect 31300 39024 31352 39030
rect 31300 38966 31352 38972
rect 31220 38758 31248 38966
rect 31208 38752 31260 38758
rect 31208 38694 31260 38700
rect 31024 38412 31076 38418
rect 31024 38354 31076 38360
rect 30708 35176 30788 35204
rect 30852 36638 30972 36666
rect 30656 35158 30708 35164
rect 30852 35154 30880 36638
rect 30932 35828 30984 35834
rect 30932 35770 30984 35776
rect 30944 35154 30972 35770
rect 31404 35630 31432 39918
rect 31496 39098 31524 40015
rect 31944 39500 31996 39506
rect 31944 39442 31996 39448
rect 31484 39092 31536 39098
rect 31484 39034 31536 39040
rect 31956 38962 31984 39442
rect 31944 38956 31996 38962
rect 31944 38898 31996 38904
rect 31668 38412 31720 38418
rect 31668 38354 31720 38360
rect 31576 38344 31628 38350
rect 31576 38286 31628 38292
rect 31588 38010 31616 38286
rect 31576 38004 31628 38010
rect 31576 37946 31628 37952
rect 31680 37330 31708 38354
rect 31668 37324 31720 37330
rect 31668 37266 31720 37272
rect 31680 36786 31708 37266
rect 31576 36780 31628 36786
rect 31576 36722 31628 36728
rect 31668 36780 31720 36786
rect 31668 36722 31720 36728
rect 31392 35624 31444 35630
rect 31392 35566 31444 35572
rect 30564 35148 30616 35154
rect 30564 35090 30616 35096
rect 30840 35148 30892 35154
rect 30840 35090 30892 35096
rect 30932 35148 30984 35154
rect 30932 35090 30984 35096
rect 30288 35080 30340 35086
rect 30340 35028 30512 35034
rect 30288 35022 30512 35028
rect 30300 35006 30512 35022
rect 30484 34542 30512 35006
rect 30472 34536 30524 34542
rect 30472 34478 30524 34484
rect 30196 34060 30248 34066
rect 30196 34002 30248 34008
rect 30484 33590 30512 34478
rect 30472 33584 30524 33590
rect 30472 33526 30524 33532
rect 30012 33108 30064 33114
rect 29932 33068 30012 33096
rect 29932 28778 29960 33068
rect 30012 33050 30064 33056
rect 30380 32904 30432 32910
rect 30380 32846 30432 32852
rect 30392 32570 30420 32846
rect 30380 32564 30432 32570
rect 30380 32506 30432 32512
rect 30196 32292 30248 32298
rect 30196 32234 30248 32240
rect 30012 29572 30064 29578
rect 30012 29514 30064 29520
rect 30024 29034 30052 29514
rect 30012 29028 30064 29034
rect 30012 28970 30064 28976
rect 29932 28750 30052 28778
rect 30208 28762 30236 32234
rect 30378 32056 30434 32065
rect 30378 31991 30434 32000
rect 30392 31822 30420 31991
rect 30380 31816 30432 31822
rect 30380 31758 30432 31764
rect 30576 31754 30604 35090
rect 30852 34610 30880 35090
rect 30944 34610 30972 35090
rect 31116 35080 31168 35086
rect 31116 35022 31168 35028
rect 30840 34604 30892 34610
rect 30840 34546 30892 34552
rect 30932 34604 30984 34610
rect 30932 34546 30984 34552
rect 30932 34128 30984 34134
rect 30932 34070 30984 34076
rect 30748 32836 30800 32842
rect 30748 32778 30800 32784
rect 30656 32768 30708 32774
rect 30656 32710 30708 32716
rect 30668 32366 30696 32710
rect 30760 32570 30788 32778
rect 30748 32564 30800 32570
rect 30748 32506 30800 32512
rect 30656 32360 30708 32366
rect 30656 32302 30708 32308
rect 30668 32026 30696 32302
rect 30760 32026 30788 32506
rect 30656 32020 30708 32026
rect 30656 31962 30708 31968
rect 30748 32020 30800 32026
rect 30748 31962 30800 31968
rect 30840 31884 30892 31890
rect 30840 31826 30892 31832
rect 30576 31726 30696 31754
rect 30562 30832 30618 30841
rect 30562 30767 30564 30776
rect 30616 30767 30618 30776
rect 30564 30738 30616 30744
rect 30576 30190 30604 30738
rect 30380 30184 30432 30190
rect 30380 30126 30432 30132
rect 30564 30184 30616 30190
rect 30564 30126 30616 30132
rect 29920 28416 29972 28422
rect 29920 28358 29972 28364
rect 29932 28218 29960 28358
rect 29920 28212 29972 28218
rect 29920 28154 29972 28160
rect 29932 27538 29960 28154
rect 30024 28014 30052 28750
rect 30196 28756 30248 28762
rect 30196 28698 30248 28704
rect 30012 28008 30064 28014
rect 30012 27950 30064 27956
rect 30024 27674 30052 27950
rect 30012 27668 30064 27674
rect 30012 27610 30064 27616
rect 29920 27532 29972 27538
rect 29920 27474 29972 27480
rect 30196 27532 30248 27538
rect 30196 27474 30248 27480
rect 29840 27390 30144 27418
rect 29920 27328 29972 27334
rect 29920 27270 29972 27276
rect 29736 27124 29788 27130
rect 29736 27066 29788 27072
rect 29828 26988 29880 26994
rect 29932 26976 29960 27270
rect 29880 26948 29960 26976
rect 30116 26976 30144 27390
rect 30208 27130 30236 27474
rect 30196 27124 30248 27130
rect 30196 27066 30248 27072
rect 30116 26948 30328 26976
rect 29828 26930 29880 26936
rect 29472 26858 29592 26874
rect 29644 26920 29696 26926
rect 30300 26874 30328 26948
rect 29644 26862 29696 26868
rect 29460 26852 29592 26858
rect 29512 26846 29592 26852
rect 30208 26846 30328 26874
rect 29460 26794 29512 26800
rect 29460 26036 29512 26042
rect 29460 25978 29512 25984
rect 29368 24676 29420 24682
rect 29368 24618 29420 24624
rect 29380 24070 29408 24618
rect 29368 24064 29420 24070
rect 29368 24006 29420 24012
rect 29472 23662 29500 25978
rect 29920 25288 29972 25294
rect 29920 25230 29972 25236
rect 29644 24676 29696 24682
rect 29644 24618 29696 24624
rect 29552 24132 29604 24138
rect 29552 24074 29604 24080
rect 29564 23769 29592 24074
rect 29656 23866 29684 24618
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29828 24608 29880 24614
rect 29828 24550 29880 24556
rect 29748 24206 29776 24550
rect 29840 24206 29868 24550
rect 29736 24200 29788 24206
rect 29736 24142 29788 24148
rect 29828 24200 29880 24206
rect 29828 24142 29880 24148
rect 29644 23860 29696 23866
rect 29644 23802 29696 23808
rect 29550 23760 29606 23769
rect 29550 23695 29606 23704
rect 29460 23656 29512 23662
rect 29460 23598 29512 23604
rect 29828 23656 29880 23662
rect 29828 23598 29880 23604
rect 29550 23488 29606 23497
rect 29550 23423 29606 23432
rect 29460 22568 29512 22574
rect 29460 22510 29512 22516
rect 29368 22500 29420 22506
rect 29368 22442 29420 22448
rect 29274 21856 29330 21865
rect 29274 21791 29330 21800
rect 29380 19990 29408 22442
rect 29472 21418 29500 22510
rect 29460 21412 29512 21418
rect 29460 21354 29512 21360
rect 29472 21078 29500 21354
rect 29460 21072 29512 21078
rect 29460 21014 29512 21020
rect 29368 19984 29420 19990
rect 29368 19926 29420 19932
rect 29368 19780 29420 19786
rect 29368 19722 29420 19728
rect 29276 19712 29328 19718
rect 29276 19654 29328 19660
rect 29288 19514 29316 19654
rect 29276 19508 29328 19514
rect 29276 19450 29328 19456
rect 29276 19372 29328 19378
rect 29276 19314 29328 19320
rect 29288 18970 29316 19314
rect 29276 18964 29328 18970
rect 29276 18906 29328 18912
rect 29380 18426 29408 19722
rect 29368 18420 29420 18426
rect 29368 18362 29420 18368
rect 29182 18320 29238 18329
rect 29182 18255 29238 18264
rect 29564 18170 29592 23423
rect 29840 23186 29868 23598
rect 29828 23180 29880 23186
rect 29828 23122 29880 23128
rect 29644 23112 29696 23118
rect 29644 23054 29696 23060
rect 29656 21049 29684 23054
rect 29736 22024 29788 22030
rect 29736 21966 29788 21972
rect 29748 21622 29776 21966
rect 29736 21616 29788 21622
rect 29736 21558 29788 21564
rect 29642 21040 29698 21049
rect 29642 20975 29698 20984
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 29748 20058 29776 20402
rect 29736 20052 29788 20058
rect 29736 19994 29788 20000
rect 29644 19168 29696 19174
rect 29644 19110 29696 19116
rect 29472 18154 29592 18170
rect 29460 18148 29592 18154
rect 29512 18142 29592 18148
rect 29460 18090 29512 18096
rect 29092 18080 29144 18086
rect 29092 18022 29144 18028
rect 29104 17746 29132 18022
rect 29092 17740 29144 17746
rect 29092 17682 29144 17688
rect 29184 17740 29236 17746
rect 29184 17682 29236 17688
rect 29012 17598 29132 17626
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 29012 17338 29040 17478
rect 29000 17332 29052 17338
rect 29000 17274 29052 17280
rect 29104 16590 29132 17598
rect 29092 16584 29144 16590
rect 29092 16526 29144 16532
rect 29196 16250 29224 17682
rect 29184 16244 29236 16250
rect 29184 16186 29236 16192
rect 28908 16176 28960 16182
rect 29092 16176 29144 16182
rect 28908 16118 28960 16124
rect 28998 16144 29054 16153
rect 28920 14618 28948 16118
rect 29092 16118 29144 16124
rect 28998 16079 29000 16088
rect 29052 16079 29054 16088
rect 29000 16050 29052 16056
rect 28908 14612 28960 14618
rect 28908 14554 28960 14560
rect 28908 13728 28960 13734
rect 28908 13670 28960 13676
rect 28920 12850 28948 13670
rect 28908 12844 28960 12850
rect 28908 12786 28960 12792
rect 29012 12434 29040 16050
rect 29104 15434 29132 16118
rect 29092 15428 29144 15434
rect 29092 15370 29144 15376
rect 29092 14816 29144 14822
rect 29092 14758 29144 14764
rect 29104 12850 29132 14758
rect 29196 14482 29224 16186
rect 29368 15496 29420 15502
rect 29368 15438 29420 15444
rect 29380 15162 29408 15438
rect 29368 15156 29420 15162
rect 29368 15098 29420 15104
rect 29184 14476 29236 14482
rect 29184 14418 29236 14424
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29092 12844 29144 12850
rect 29092 12786 29144 12792
rect 29012 12406 29132 12434
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 29012 10130 29040 10610
rect 29000 10124 29052 10130
rect 29000 10066 29052 10072
rect 29104 10010 29132 12406
rect 29288 12102 29316 13874
rect 29472 12434 29500 18090
rect 29552 17536 29604 17542
rect 29552 17478 29604 17484
rect 29564 17270 29592 17478
rect 29552 17264 29604 17270
rect 29552 17206 29604 17212
rect 29656 17066 29684 19110
rect 29736 18760 29788 18766
rect 29736 18702 29788 18708
rect 29748 18086 29776 18702
rect 29828 18216 29880 18222
rect 29828 18158 29880 18164
rect 29736 18080 29788 18086
rect 29736 18022 29788 18028
rect 29840 17746 29868 18158
rect 29828 17740 29880 17746
rect 29828 17682 29880 17688
rect 29840 17270 29868 17682
rect 29828 17264 29880 17270
rect 29828 17206 29880 17212
rect 29932 17134 29960 25230
rect 30208 24818 30236 26846
rect 30288 26784 30340 26790
rect 30392 26772 30420 30126
rect 30564 28756 30616 28762
rect 30564 28698 30616 28704
rect 30576 28200 30604 28698
rect 30484 28172 30604 28200
rect 30484 27946 30512 28172
rect 30564 28076 30616 28082
rect 30564 28018 30616 28024
rect 30472 27940 30524 27946
rect 30472 27882 30524 27888
rect 30576 27674 30604 28018
rect 30564 27668 30616 27674
rect 30564 27610 30616 27616
rect 30472 27464 30524 27470
rect 30472 27406 30524 27412
rect 30484 27334 30512 27406
rect 30472 27328 30524 27334
rect 30472 27270 30524 27276
rect 30564 26784 30616 26790
rect 30392 26744 30512 26772
rect 30288 26726 30340 26732
rect 30196 24812 30248 24818
rect 30116 24772 30196 24800
rect 30012 24744 30064 24750
rect 30012 24686 30064 24692
rect 30024 23118 30052 24686
rect 30012 23112 30064 23118
rect 30012 23054 30064 23060
rect 30012 22432 30064 22438
rect 30012 22374 30064 22380
rect 30024 22030 30052 22374
rect 30012 22024 30064 22030
rect 30012 21966 30064 21972
rect 30012 20392 30064 20398
rect 30010 20360 30012 20369
rect 30064 20360 30066 20369
rect 30010 20295 30066 20304
rect 30116 19334 30144 24772
rect 30196 24754 30248 24760
rect 30196 23520 30248 23526
rect 30196 23462 30248 23468
rect 30208 23118 30236 23462
rect 30196 23112 30248 23118
rect 30196 23054 30248 23060
rect 30196 19372 30248 19378
rect 30116 19320 30196 19334
rect 30116 19314 30248 19320
rect 30116 19306 30236 19314
rect 30104 18964 30156 18970
rect 30104 18906 30156 18912
rect 30012 18760 30064 18766
rect 30010 18728 30012 18737
rect 30064 18728 30066 18737
rect 30010 18663 30066 18672
rect 30012 18420 30064 18426
rect 30012 18362 30064 18368
rect 30024 17746 30052 18362
rect 30116 17814 30144 18906
rect 30104 17808 30156 17814
rect 30104 17750 30156 17756
rect 30012 17740 30064 17746
rect 30012 17682 30064 17688
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 29644 17060 29696 17066
rect 29644 17002 29696 17008
rect 29644 16584 29696 16590
rect 29644 16526 29696 16532
rect 29656 15910 29684 16526
rect 29644 15904 29696 15910
rect 29644 15846 29696 15852
rect 29552 14408 29604 14414
rect 29552 14350 29604 14356
rect 29564 13462 29592 14350
rect 29656 13802 29684 15846
rect 29932 15094 29960 17070
rect 30116 15978 30144 17750
rect 30104 15972 30156 15978
rect 30104 15914 30156 15920
rect 29920 15088 29972 15094
rect 29920 15030 29972 15036
rect 29736 14952 29788 14958
rect 29736 14894 29788 14900
rect 29748 14550 29776 14894
rect 29736 14544 29788 14550
rect 29736 14486 29788 14492
rect 30104 13864 30156 13870
rect 30104 13806 30156 13812
rect 29644 13796 29696 13802
rect 29644 13738 29696 13744
rect 30012 13796 30064 13802
rect 30012 13738 30064 13744
rect 29656 13530 29684 13738
rect 29644 13524 29696 13530
rect 29644 13466 29696 13472
rect 29552 13456 29604 13462
rect 29552 13398 29604 13404
rect 29380 12406 29500 12434
rect 29564 12434 29592 13398
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 29840 12714 29868 13330
rect 30024 13326 30052 13738
rect 30116 13394 30144 13806
rect 30104 13388 30156 13394
rect 30104 13330 30156 13336
rect 30012 13320 30064 13326
rect 30012 13262 30064 13268
rect 29920 12980 29972 12986
rect 29920 12922 29972 12928
rect 29932 12782 29960 12922
rect 29920 12776 29972 12782
rect 29920 12718 29972 12724
rect 29828 12708 29880 12714
rect 29828 12650 29880 12656
rect 29564 12406 29776 12434
rect 29276 12096 29328 12102
rect 29276 12038 29328 12044
rect 29276 11756 29328 11762
rect 29276 11698 29328 11704
rect 29288 11354 29316 11698
rect 29276 11348 29328 11354
rect 29276 11290 29328 11296
rect 29380 10606 29408 12406
rect 29472 10674 29684 10690
rect 29472 10668 29696 10674
rect 29472 10662 29644 10668
rect 29184 10600 29236 10606
rect 29184 10542 29236 10548
rect 29368 10600 29420 10606
rect 29368 10542 29420 10548
rect 29196 10062 29224 10542
rect 29012 9982 29132 10010
rect 29184 10056 29236 10062
rect 29184 9998 29236 10004
rect 29368 10056 29420 10062
rect 29368 9998 29420 10004
rect 28908 6792 28960 6798
rect 28908 6734 28960 6740
rect 28920 6322 28948 6734
rect 28908 6316 28960 6322
rect 28908 6258 28960 6264
rect 29012 6254 29040 9982
rect 29092 9920 29144 9926
rect 29092 9862 29144 9868
rect 29184 9920 29236 9926
rect 29184 9862 29236 9868
rect 29104 9722 29132 9862
rect 29092 9716 29144 9722
rect 29092 9658 29144 9664
rect 29196 9654 29224 9862
rect 29184 9648 29236 9654
rect 29184 9590 29236 9596
rect 29276 9444 29328 9450
rect 29276 9386 29328 9392
rect 29184 7812 29236 7818
rect 29184 7754 29236 7760
rect 29196 7546 29224 7754
rect 29184 7540 29236 7546
rect 29184 7482 29236 7488
rect 29288 7342 29316 9386
rect 29276 7336 29328 7342
rect 29276 7278 29328 7284
rect 29000 6248 29052 6254
rect 29000 6190 29052 6196
rect 29184 6248 29236 6254
rect 29184 6190 29236 6196
rect 29012 5234 29040 6190
rect 29196 5778 29224 6190
rect 29184 5772 29236 5778
rect 29184 5714 29236 5720
rect 28908 5228 28960 5234
rect 28908 5170 28960 5176
rect 29000 5228 29052 5234
rect 29000 5170 29052 5176
rect 28920 4758 28948 5170
rect 28908 4752 28960 4758
rect 28908 4694 28960 4700
rect 29000 4752 29052 4758
rect 29000 4694 29052 4700
rect 29012 4214 29040 4694
rect 29000 4208 29052 4214
rect 29000 4150 29052 4156
rect 29380 3602 29408 9998
rect 29472 9994 29500 10662
rect 29644 10610 29696 10616
rect 29552 10600 29604 10606
rect 29552 10542 29604 10548
rect 29564 10112 29592 10542
rect 29644 10124 29696 10130
rect 29564 10084 29644 10112
rect 29460 9988 29512 9994
rect 29460 9930 29512 9936
rect 29472 9382 29500 9930
rect 29564 9926 29592 10084
rect 29644 10066 29696 10072
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 29552 9648 29604 9654
rect 29552 9590 29604 9596
rect 29460 9376 29512 9382
rect 29460 9318 29512 9324
rect 29564 8498 29592 9590
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 29460 8424 29512 8430
rect 29460 8366 29512 8372
rect 29644 8424 29696 8430
rect 29644 8366 29696 8372
rect 29472 7954 29500 8366
rect 29460 7948 29512 7954
rect 29460 7890 29512 7896
rect 29656 7886 29684 8366
rect 29644 7880 29696 7886
rect 29644 7822 29696 7828
rect 29552 7404 29604 7410
rect 29552 7346 29604 7352
rect 29564 5710 29592 7346
rect 29656 5914 29684 7822
rect 29748 6866 29776 12406
rect 29918 12336 29974 12345
rect 29918 12271 29974 12280
rect 29932 12238 29960 12271
rect 29920 12232 29972 12238
rect 29920 12174 29972 12180
rect 29828 11756 29880 11762
rect 29828 11698 29880 11704
rect 29840 11286 29868 11698
rect 29932 11642 29960 12174
rect 30024 11830 30052 13262
rect 30104 12844 30156 12850
rect 30104 12786 30156 12792
rect 30012 11824 30064 11830
rect 30012 11766 30064 11772
rect 29932 11614 30052 11642
rect 29828 11280 29880 11286
rect 29828 11222 29880 11228
rect 29826 10976 29882 10985
rect 29826 10911 29882 10920
rect 29840 10674 29868 10911
rect 29828 10668 29880 10674
rect 29828 10610 29880 10616
rect 29920 10192 29972 10198
rect 29920 10134 29972 10140
rect 29828 7336 29880 7342
rect 29828 7278 29880 7284
rect 29840 6934 29868 7278
rect 29828 6928 29880 6934
rect 29828 6870 29880 6876
rect 29736 6860 29788 6866
rect 29736 6802 29788 6808
rect 29840 6186 29868 6870
rect 29828 6180 29880 6186
rect 29828 6122 29880 6128
rect 29644 5908 29696 5914
rect 29644 5850 29696 5856
rect 29552 5704 29604 5710
rect 29552 5646 29604 5652
rect 29656 5166 29684 5850
rect 29736 5704 29788 5710
rect 29736 5646 29788 5652
rect 29644 5160 29696 5166
rect 29644 5102 29696 5108
rect 29748 4690 29776 5646
rect 29840 5302 29868 6122
rect 29828 5296 29880 5302
rect 29828 5238 29880 5244
rect 29736 4684 29788 4690
rect 29736 4626 29788 4632
rect 29932 4622 29960 10134
rect 30024 7410 30052 11614
rect 30116 10198 30144 12786
rect 30208 11762 30236 19306
rect 30300 18970 30328 26726
rect 30484 24818 30512 26744
rect 30564 26726 30616 26732
rect 30576 26382 30604 26726
rect 30564 26376 30616 26382
rect 30564 26318 30616 26324
rect 30564 25832 30616 25838
rect 30564 25774 30616 25780
rect 30472 24812 30524 24818
rect 30472 24754 30524 24760
rect 30380 24676 30432 24682
rect 30380 24618 30432 24624
rect 30392 24154 30420 24618
rect 30484 24274 30512 24754
rect 30576 24750 30604 25774
rect 30668 25430 30696 31726
rect 30852 31482 30880 31826
rect 30840 31476 30892 31482
rect 30840 31418 30892 31424
rect 30840 31136 30892 31142
rect 30840 31078 30892 31084
rect 30852 30734 30880 31078
rect 30840 30728 30892 30734
rect 30840 30670 30892 30676
rect 30840 30592 30892 30598
rect 30840 30534 30892 30540
rect 30852 30326 30880 30534
rect 30840 30320 30892 30326
rect 30840 30262 30892 30268
rect 30748 28008 30800 28014
rect 30748 27950 30800 27956
rect 30656 25424 30708 25430
rect 30656 25366 30708 25372
rect 30656 24880 30708 24886
rect 30656 24822 30708 24828
rect 30564 24744 30616 24750
rect 30564 24686 30616 24692
rect 30472 24268 30524 24274
rect 30472 24210 30524 24216
rect 30392 24126 30604 24154
rect 30472 23724 30524 23730
rect 30472 23666 30524 23672
rect 30378 23624 30434 23633
rect 30378 23559 30434 23568
rect 30392 21894 30420 23559
rect 30484 22778 30512 23666
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30380 21888 30432 21894
rect 30380 21830 30432 21836
rect 30472 20256 30524 20262
rect 30472 20198 30524 20204
rect 30484 19310 30512 20198
rect 30576 19922 30604 24126
rect 30668 23905 30696 24822
rect 30654 23896 30710 23905
rect 30654 23831 30710 23840
rect 30656 22636 30708 22642
rect 30656 22578 30708 22584
rect 30668 22438 30696 22578
rect 30656 22432 30708 22438
rect 30656 22374 30708 22380
rect 30760 21554 30788 27950
rect 30944 27538 30972 34070
rect 31024 34060 31076 34066
rect 31024 34002 31076 34008
rect 31036 32366 31064 34002
rect 31024 32360 31076 32366
rect 31024 32302 31076 32308
rect 31024 32020 31076 32026
rect 31024 31962 31076 31968
rect 31036 31385 31064 31962
rect 31022 31376 31078 31385
rect 31022 31311 31078 31320
rect 30932 27532 30984 27538
rect 30932 27474 30984 27480
rect 30840 26920 30892 26926
rect 30840 26862 30892 26868
rect 30852 25294 30880 26862
rect 30840 25288 30892 25294
rect 30840 25230 30892 25236
rect 30840 25152 30892 25158
rect 30840 25094 30892 25100
rect 30852 24886 30880 25094
rect 30840 24880 30892 24886
rect 30840 24822 30892 24828
rect 30840 24268 30892 24274
rect 30840 24210 30892 24216
rect 30748 21548 30800 21554
rect 30748 21490 30800 21496
rect 30564 19916 30616 19922
rect 30564 19858 30616 19864
rect 30472 19304 30524 19310
rect 30472 19246 30524 19252
rect 30564 19168 30616 19174
rect 30564 19110 30616 19116
rect 30288 18964 30340 18970
rect 30288 18906 30340 18912
rect 30576 18698 30604 19110
rect 30564 18692 30616 18698
rect 30564 18634 30616 18640
rect 30286 18320 30342 18329
rect 30342 18290 30512 18306
rect 30342 18284 30524 18290
rect 30342 18278 30472 18284
rect 30286 18255 30342 18264
rect 30472 18226 30524 18232
rect 30288 18216 30340 18222
rect 30288 18158 30340 18164
rect 30300 17542 30328 18158
rect 30576 18086 30604 18634
rect 30564 18080 30616 18086
rect 30564 18022 30616 18028
rect 30656 18080 30708 18086
rect 30656 18022 30708 18028
rect 30576 17746 30604 18022
rect 30564 17740 30616 17746
rect 30564 17682 30616 17688
rect 30288 17536 30340 17542
rect 30668 17490 30696 18022
rect 30288 17478 30340 17484
rect 30300 17338 30328 17478
rect 30392 17462 30696 17490
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30392 17218 30420 17462
rect 30300 17190 30420 17218
rect 30300 16590 30328 17190
rect 30472 17060 30524 17066
rect 30472 17002 30524 17008
rect 30288 16584 30340 16590
rect 30288 16526 30340 16532
rect 30288 15972 30340 15978
rect 30288 15914 30340 15920
rect 30300 13462 30328 15914
rect 30378 13832 30434 13841
rect 30378 13767 30380 13776
rect 30432 13767 30434 13776
rect 30380 13738 30432 13744
rect 30288 13456 30340 13462
rect 30288 13398 30340 13404
rect 30300 12850 30328 13398
rect 30378 12880 30434 12889
rect 30288 12844 30340 12850
rect 30378 12815 30380 12824
rect 30288 12786 30340 12792
rect 30432 12815 30434 12824
rect 30380 12786 30432 12792
rect 30286 12744 30342 12753
rect 30286 12679 30342 12688
rect 30300 12306 30328 12679
rect 30484 12374 30512 17002
rect 30656 16720 30708 16726
rect 30656 16662 30708 16668
rect 30668 15314 30696 16662
rect 30760 15416 30788 21490
rect 30852 19378 30880 24210
rect 30944 22094 30972 27474
rect 31128 25702 31156 35022
rect 31300 31952 31352 31958
rect 31300 31894 31352 31900
rect 31312 31482 31340 31894
rect 31300 31476 31352 31482
rect 31300 31418 31352 31424
rect 31404 31278 31432 35566
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 31496 31521 31524 31758
rect 31482 31512 31538 31521
rect 31482 31447 31538 31456
rect 31392 31272 31444 31278
rect 31392 31214 31444 31220
rect 31208 31204 31260 31210
rect 31208 31146 31260 31152
rect 31220 30666 31248 31146
rect 31208 30660 31260 30666
rect 31208 30602 31260 30608
rect 31404 28994 31432 31214
rect 31482 30152 31538 30161
rect 31482 30087 31538 30096
rect 31496 29850 31524 30087
rect 31484 29844 31536 29850
rect 31484 29786 31536 29792
rect 31588 29578 31616 36722
rect 31760 34400 31812 34406
rect 31760 34342 31812 34348
rect 31852 34400 31904 34406
rect 31852 34342 31904 34348
rect 31668 33992 31720 33998
rect 31668 33934 31720 33940
rect 31680 33658 31708 33934
rect 31668 33652 31720 33658
rect 31668 33594 31720 33600
rect 31668 30864 31720 30870
rect 31668 30806 31720 30812
rect 31680 30394 31708 30806
rect 31772 30546 31800 34342
rect 31864 33998 31892 34342
rect 31852 33992 31904 33998
rect 31852 33934 31904 33940
rect 31852 33380 31904 33386
rect 31852 33322 31904 33328
rect 31864 31822 31892 33322
rect 31852 31816 31904 31822
rect 31852 31758 31904 31764
rect 31864 31385 31892 31758
rect 31956 31754 31984 38898
rect 32036 36848 32088 36854
rect 32036 36790 32088 36796
rect 32048 33454 32076 36790
rect 32128 36168 32180 36174
rect 32128 36110 32180 36116
rect 32140 35698 32168 36110
rect 32128 35692 32180 35698
rect 32128 35634 32180 35640
rect 32036 33448 32088 33454
rect 32036 33390 32088 33396
rect 32048 31958 32076 33390
rect 32128 32904 32180 32910
rect 32128 32846 32180 32852
rect 32140 32570 32168 32846
rect 32128 32564 32180 32570
rect 32128 32506 32180 32512
rect 32036 31952 32088 31958
rect 32036 31894 32088 31900
rect 31956 31726 32076 31754
rect 31850 31376 31906 31385
rect 31850 31311 31906 31320
rect 31944 31340 31996 31346
rect 31944 31282 31996 31288
rect 31852 31136 31904 31142
rect 31852 31078 31904 31084
rect 31864 30938 31892 31078
rect 31956 30938 31984 31282
rect 32048 31278 32076 31726
rect 32036 31272 32088 31278
rect 32036 31214 32088 31220
rect 31852 30932 31904 30938
rect 31852 30874 31904 30880
rect 31944 30932 31996 30938
rect 31944 30874 31996 30880
rect 32128 30796 32180 30802
rect 32128 30738 32180 30744
rect 31772 30518 32076 30546
rect 32048 30394 32076 30518
rect 31668 30388 31720 30394
rect 31668 30330 31720 30336
rect 32036 30388 32088 30394
rect 32036 30330 32088 30336
rect 32140 30258 32168 30738
rect 32232 30598 32260 46566
rect 32416 45529 32444 47534
rect 33508 47456 33560 47462
rect 33508 47398 33560 47404
rect 33324 47116 33376 47122
rect 33324 47058 33376 47064
rect 33336 46510 33364 47058
rect 33520 46986 33548 47398
rect 33508 46980 33560 46986
rect 33508 46922 33560 46928
rect 33324 46504 33376 46510
rect 33324 46446 33376 46452
rect 33232 46028 33284 46034
rect 33232 45970 33284 45976
rect 33138 45928 33194 45937
rect 33138 45863 33140 45872
rect 33192 45863 33194 45872
rect 33140 45834 33192 45840
rect 33140 45620 33192 45626
rect 33140 45562 33192 45568
rect 32402 45520 32458 45529
rect 33152 45506 33180 45562
rect 32968 45490 33180 45506
rect 32402 45455 32458 45464
rect 32588 45484 32640 45490
rect 32312 45280 32364 45286
rect 32312 45222 32364 45228
rect 32324 44878 32352 45222
rect 32312 44872 32364 44878
rect 32312 44814 32364 44820
rect 32416 44198 32444 45455
rect 32588 45426 32640 45432
rect 32956 45484 33180 45490
rect 33008 45478 33180 45484
rect 32956 45426 33008 45432
rect 32600 45082 32628 45426
rect 32588 45076 32640 45082
rect 32588 45018 32640 45024
rect 32680 44940 32732 44946
rect 32680 44882 32732 44888
rect 32404 44192 32456 44198
rect 32404 44134 32456 44140
rect 32692 43489 32720 44882
rect 32956 44872 33008 44878
rect 32956 44814 33008 44820
rect 32968 44538 32996 44814
rect 33244 44538 33272 45970
rect 33336 44962 33364 46446
rect 33416 45824 33468 45830
rect 33416 45766 33468 45772
rect 33428 45558 33456 45766
rect 33416 45552 33468 45558
rect 33416 45494 33468 45500
rect 33336 44934 33456 44962
rect 33324 44804 33376 44810
rect 33324 44746 33376 44752
rect 32956 44532 33008 44538
rect 32956 44474 33008 44480
rect 33232 44532 33284 44538
rect 33232 44474 33284 44480
rect 32678 43480 32734 43489
rect 32678 43415 32734 43424
rect 32968 42702 32996 44474
rect 33336 44402 33364 44746
rect 33324 44396 33376 44402
rect 33324 44338 33376 44344
rect 33336 43994 33364 44338
rect 33324 43988 33376 43994
rect 33324 43930 33376 43936
rect 33428 43314 33456 44934
rect 33416 43308 33468 43314
rect 33416 43250 33468 43256
rect 32956 42696 33008 42702
rect 32956 42638 33008 42644
rect 32588 42560 32640 42566
rect 32588 42502 32640 42508
rect 32600 42294 32628 42502
rect 32968 42362 32996 42638
rect 32956 42356 33008 42362
rect 32956 42298 33008 42304
rect 32588 42288 32640 42294
rect 32588 42230 32640 42236
rect 32864 41812 32916 41818
rect 32864 41754 32916 41760
rect 32876 41698 32904 41754
rect 32692 41682 32904 41698
rect 33140 41744 33192 41750
rect 33140 41686 33192 41692
rect 32680 41676 32904 41682
rect 32732 41670 32904 41676
rect 32680 41618 32732 41624
rect 32404 41472 32456 41478
rect 32588 41472 32640 41478
rect 32404 41414 32456 41420
rect 32586 41440 32588 41449
rect 32640 41440 32642 41449
rect 32416 36922 32444 41414
rect 32586 41375 32642 41384
rect 33048 40520 33100 40526
rect 33048 40462 33100 40468
rect 32772 40180 32824 40186
rect 32772 40122 32824 40128
rect 32680 39296 32732 39302
rect 32680 39238 32732 39244
rect 32496 38208 32548 38214
rect 32496 38150 32548 38156
rect 32508 38010 32536 38150
rect 32496 38004 32548 38010
rect 32496 37946 32548 37952
rect 32404 36916 32456 36922
rect 32404 36858 32456 36864
rect 32312 36372 32364 36378
rect 32312 36314 32364 36320
rect 32324 35698 32352 36314
rect 32508 36310 32536 37946
rect 32588 37800 32640 37806
rect 32588 37742 32640 37748
rect 32496 36304 32548 36310
rect 32496 36246 32548 36252
rect 32404 36236 32456 36242
rect 32404 36178 32456 36184
rect 32312 35692 32364 35698
rect 32312 35634 32364 35640
rect 32312 34400 32364 34406
rect 32312 34342 32364 34348
rect 32324 32910 32352 34342
rect 32416 33114 32444 36178
rect 32496 33856 32548 33862
rect 32496 33798 32548 33804
rect 32508 33658 32536 33798
rect 32496 33652 32548 33658
rect 32496 33594 32548 33600
rect 32404 33108 32456 33114
rect 32404 33050 32456 33056
rect 32312 32904 32364 32910
rect 32312 32846 32364 32852
rect 32496 32564 32548 32570
rect 32496 32506 32548 32512
rect 32312 31136 32364 31142
rect 32312 31078 32364 31084
rect 32324 30734 32352 31078
rect 32508 30802 32536 32506
rect 32600 32450 32628 37742
rect 32692 36242 32720 39238
rect 32784 36242 32812 40122
rect 32864 39296 32916 39302
rect 32864 39238 32916 39244
rect 32876 39030 32904 39238
rect 32864 39024 32916 39030
rect 32864 38966 32916 38972
rect 32876 38010 32904 38966
rect 33060 38894 33088 40462
rect 33152 40118 33180 41686
rect 33324 41608 33376 41614
rect 33324 41550 33376 41556
rect 33140 40112 33192 40118
rect 33140 40054 33192 40060
rect 33048 38888 33100 38894
rect 33048 38830 33100 38836
rect 33060 38706 33088 38830
rect 33060 38678 33180 38706
rect 32864 38004 32916 38010
rect 32864 37946 32916 37952
rect 33152 37262 33180 38678
rect 33232 38276 33284 38282
rect 33232 38218 33284 38224
rect 33244 37942 33272 38218
rect 33336 38010 33364 41550
rect 33416 40044 33468 40050
rect 33416 39986 33468 39992
rect 33324 38004 33376 38010
rect 33324 37946 33376 37952
rect 33232 37936 33284 37942
rect 33232 37878 33284 37884
rect 33140 37256 33192 37262
rect 33140 37198 33192 37204
rect 32864 36916 32916 36922
rect 32864 36858 32916 36864
rect 32680 36236 32732 36242
rect 32680 36178 32732 36184
rect 32772 36236 32824 36242
rect 32772 36178 32824 36184
rect 32692 35630 32720 36178
rect 32680 35624 32732 35630
rect 32680 35566 32732 35572
rect 32680 32768 32732 32774
rect 32680 32710 32732 32716
rect 32692 32570 32720 32710
rect 32680 32564 32732 32570
rect 32680 32506 32732 32512
rect 32600 32422 32720 32450
rect 32692 32366 32720 32422
rect 32680 32360 32732 32366
rect 32680 32302 32732 32308
rect 32588 31272 32640 31278
rect 32588 31214 32640 31220
rect 32496 30796 32548 30802
rect 32496 30738 32548 30744
rect 32312 30728 32364 30734
rect 32312 30670 32364 30676
rect 32220 30592 32272 30598
rect 32220 30534 32272 30540
rect 32128 30252 32180 30258
rect 32128 30194 32180 30200
rect 32324 30190 32352 30670
rect 32312 30184 32364 30190
rect 32312 30126 32364 30132
rect 31576 29572 31628 29578
rect 31576 29514 31628 29520
rect 32128 29164 32180 29170
rect 32128 29106 32180 29112
rect 31312 28966 31432 28994
rect 31312 27538 31340 28966
rect 31576 28620 31628 28626
rect 31576 28562 31628 28568
rect 31588 28218 31616 28562
rect 31944 28416 31996 28422
rect 31944 28358 31996 28364
rect 31576 28212 31628 28218
rect 31576 28154 31628 28160
rect 31300 27532 31352 27538
rect 31300 27474 31352 27480
rect 31312 26897 31340 27474
rect 31588 27402 31616 28154
rect 31956 28082 31984 28358
rect 31944 28076 31996 28082
rect 31944 28018 31996 28024
rect 32140 28014 32168 29106
rect 32496 28756 32548 28762
rect 32496 28698 32548 28704
rect 32508 28218 32536 28698
rect 32600 28626 32628 31214
rect 32692 28966 32720 32302
rect 32772 30796 32824 30802
rect 32772 30738 32824 30744
rect 32784 30394 32812 30738
rect 32876 30705 32904 36858
rect 33428 36310 33456 39986
rect 33520 36854 33548 46922
rect 33692 45960 33744 45966
rect 33690 45928 33692 45937
rect 33744 45928 33746 45937
rect 33690 45863 33746 45872
rect 33692 45824 33744 45830
rect 33692 45766 33744 45772
rect 33704 45626 33732 45766
rect 33692 45620 33744 45626
rect 33692 45562 33744 45568
rect 33968 45280 34020 45286
rect 33968 45222 34020 45228
rect 33980 44946 34008 45222
rect 33968 44940 34020 44946
rect 33968 44882 34020 44888
rect 34244 44532 34296 44538
rect 34244 44474 34296 44480
rect 33600 43716 33652 43722
rect 33600 43658 33652 43664
rect 33612 42362 33640 43658
rect 34152 42628 34204 42634
rect 34152 42570 34204 42576
rect 33600 42356 33652 42362
rect 33600 42298 33652 42304
rect 34164 42140 34192 42570
rect 34256 42294 34284 44474
rect 34244 42288 34296 42294
rect 34244 42230 34296 42236
rect 34244 42152 34296 42158
rect 34164 42112 34244 42140
rect 34244 42094 34296 42100
rect 34152 41200 34204 41206
rect 34152 41142 34204 41148
rect 33692 41132 33744 41138
rect 33692 41074 33744 41080
rect 33600 40384 33652 40390
rect 33600 40326 33652 40332
rect 33612 40050 33640 40326
rect 33704 40118 33732 41074
rect 34060 40452 34112 40458
rect 34060 40394 34112 40400
rect 34072 40186 34100 40394
rect 34060 40180 34112 40186
rect 34060 40122 34112 40128
rect 33692 40112 33744 40118
rect 33692 40054 33744 40060
rect 33784 40112 33836 40118
rect 33784 40054 33836 40060
rect 33600 40044 33652 40050
rect 33600 39986 33652 39992
rect 33508 36848 33560 36854
rect 33508 36790 33560 36796
rect 33416 36304 33468 36310
rect 33416 36246 33468 36252
rect 33140 36236 33192 36242
rect 33140 36178 33192 36184
rect 33508 36236 33560 36242
rect 33508 36178 33560 36184
rect 32956 36168 33008 36174
rect 32956 36110 33008 36116
rect 32968 32570 32996 36110
rect 33152 35698 33180 36178
rect 33140 35692 33192 35698
rect 33140 35634 33192 35640
rect 33324 35624 33376 35630
rect 33324 35566 33376 35572
rect 33336 35154 33364 35566
rect 33324 35148 33376 35154
rect 33324 35090 33376 35096
rect 33046 34912 33102 34921
rect 33046 34847 33102 34856
rect 33060 34610 33088 34847
rect 33048 34604 33100 34610
rect 33048 34546 33100 34552
rect 33324 34536 33376 34542
rect 33324 34478 33376 34484
rect 32956 32564 33008 32570
rect 32956 32506 33008 32512
rect 33048 31340 33100 31346
rect 33048 31282 33100 31288
rect 33060 30734 33088 31282
rect 33140 30932 33192 30938
rect 33140 30874 33192 30880
rect 33152 30734 33180 30874
rect 33336 30734 33364 34478
rect 33520 33454 33548 36178
rect 33612 35086 33640 39986
rect 33796 38350 33824 40054
rect 34164 39982 34192 41142
rect 34256 40934 34284 42094
rect 34244 40928 34296 40934
rect 34244 40870 34296 40876
rect 34152 39976 34204 39982
rect 34152 39918 34204 39924
rect 34152 39024 34204 39030
rect 34152 38966 34204 38972
rect 33784 38344 33836 38350
rect 33784 38286 33836 38292
rect 34060 36576 34112 36582
rect 34060 36518 34112 36524
rect 34072 36378 34100 36518
rect 34060 36372 34112 36378
rect 34060 36314 34112 36320
rect 34072 36106 34100 36314
rect 34060 36100 34112 36106
rect 34060 36042 34112 36048
rect 34164 36038 34192 38966
rect 34256 38944 34284 40870
rect 34348 39302 34376 47602
rect 36452 47592 36504 47598
rect 36452 47534 36504 47540
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34980 47048 35032 47054
rect 34980 46990 35032 46996
rect 34796 46912 34848 46918
rect 34796 46854 34848 46860
rect 34808 46646 34836 46854
rect 34992 46714 35020 46990
rect 35440 46980 35492 46986
rect 35440 46922 35492 46928
rect 34980 46708 35032 46714
rect 34980 46650 35032 46656
rect 34796 46640 34848 46646
rect 34796 46582 34848 46588
rect 35452 46510 35480 46922
rect 35594 46812 35902 46821
rect 35594 46810 35600 46812
rect 35656 46810 35680 46812
rect 35736 46810 35760 46812
rect 35816 46810 35840 46812
rect 35896 46810 35902 46812
rect 35656 46758 35658 46810
rect 35838 46758 35840 46810
rect 35594 46756 35600 46758
rect 35656 46756 35680 46758
rect 35736 46756 35760 46758
rect 35816 46756 35840 46758
rect 35896 46756 35902 46758
rect 35594 46747 35902 46756
rect 35716 46572 35768 46578
rect 35716 46514 35768 46520
rect 35808 46572 35860 46578
rect 35808 46514 35860 46520
rect 35440 46504 35492 46510
rect 35440 46446 35492 46452
rect 35348 46368 35400 46374
rect 35348 46310 35400 46316
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 35360 45966 35388 46310
rect 35728 46034 35756 46514
rect 35440 46028 35492 46034
rect 35440 45970 35492 45976
rect 35716 46028 35768 46034
rect 35716 45970 35768 45976
rect 34796 45960 34848 45966
rect 34796 45902 34848 45908
rect 35348 45960 35400 45966
rect 35348 45902 35400 45908
rect 34428 45824 34480 45830
rect 34428 45766 34480 45772
rect 34440 44441 34468 45766
rect 34808 45558 34836 45902
rect 34796 45552 34848 45558
rect 34796 45494 34848 45500
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34796 45008 34848 45014
rect 34796 44950 34848 44956
rect 34426 44432 34482 44441
rect 34808 44402 34836 44950
rect 35452 44470 35480 45970
rect 35820 45830 35848 46514
rect 36360 46368 36412 46374
rect 36360 46310 36412 46316
rect 36372 45966 36400 46310
rect 36360 45960 36412 45966
rect 36360 45902 36412 45908
rect 35808 45824 35860 45830
rect 35808 45766 35860 45772
rect 35594 45724 35902 45733
rect 35594 45722 35600 45724
rect 35656 45722 35680 45724
rect 35736 45722 35760 45724
rect 35816 45722 35840 45724
rect 35896 45722 35902 45724
rect 35656 45670 35658 45722
rect 35838 45670 35840 45722
rect 35594 45668 35600 45670
rect 35656 45668 35680 45670
rect 35736 45668 35760 45670
rect 35816 45668 35840 45670
rect 35896 45668 35902 45670
rect 35594 45659 35902 45668
rect 35594 44636 35902 44645
rect 35594 44634 35600 44636
rect 35656 44634 35680 44636
rect 35736 44634 35760 44636
rect 35816 44634 35840 44636
rect 35896 44634 35902 44636
rect 35656 44582 35658 44634
rect 35838 44582 35840 44634
rect 35594 44580 35600 44582
rect 35656 44580 35680 44582
rect 35736 44580 35760 44582
rect 35816 44580 35840 44582
rect 35896 44580 35902 44582
rect 35594 44571 35902 44580
rect 36464 44538 36492 47534
rect 36728 45824 36780 45830
rect 36728 45766 36780 45772
rect 36740 45558 36768 45766
rect 36728 45552 36780 45558
rect 36728 45494 36780 45500
rect 36452 44532 36504 44538
rect 36452 44474 36504 44480
rect 35348 44464 35400 44470
rect 35348 44406 35400 44412
rect 35440 44464 35492 44470
rect 35440 44406 35492 44412
rect 34426 44367 34482 44376
rect 34796 44396 34848 44402
rect 34440 41596 34468 44367
rect 34796 44338 34848 44344
rect 34520 44328 34572 44334
rect 34520 44270 34572 44276
rect 34532 43246 34560 44270
rect 34704 43716 34756 43722
rect 34704 43658 34756 43664
rect 34716 43314 34744 43658
rect 34808 43450 34836 44338
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 35360 43994 35388 44406
rect 36464 43994 36492 44474
rect 35348 43988 35400 43994
rect 35348 43930 35400 43936
rect 36452 43988 36504 43994
rect 36452 43930 36504 43936
rect 34888 43920 34940 43926
rect 34888 43862 34940 43868
rect 34900 43450 34928 43862
rect 35992 43852 36044 43858
rect 36044 43812 36308 43840
rect 35992 43794 36044 43800
rect 35348 43784 35400 43790
rect 35348 43726 35400 43732
rect 34796 43444 34848 43450
rect 34796 43386 34848 43392
rect 34888 43444 34940 43450
rect 34888 43386 34940 43392
rect 34900 43330 34928 43386
rect 34704 43308 34756 43314
rect 34704 43250 34756 43256
rect 34808 43302 34928 43330
rect 35072 43308 35124 43314
rect 34520 43240 34572 43246
rect 34716 43217 34744 43250
rect 34520 43182 34572 43188
rect 34702 43208 34758 43217
rect 34612 43172 34664 43178
rect 34702 43143 34758 43152
rect 34612 43114 34664 43120
rect 34520 43104 34572 43110
rect 34520 43046 34572 43052
rect 34532 41750 34560 43046
rect 34520 41744 34572 41750
rect 34520 41686 34572 41692
rect 34440 41568 34560 41596
rect 34428 41472 34480 41478
rect 34428 41414 34480 41420
rect 34440 41138 34468 41414
rect 34428 41132 34480 41138
rect 34428 41074 34480 41080
rect 34428 40996 34480 41002
rect 34428 40938 34480 40944
rect 34440 40118 34468 40938
rect 34532 40769 34560 41568
rect 34624 41546 34652 43114
rect 34704 42220 34756 42226
rect 34704 42162 34756 42168
rect 34612 41540 34664 41546
rect 34612 41482 34664 41488
rect 34612 41268 34664 41274
rect 34612 41210 34664 41216
rect 34518 40760 34574 40769
rect 34518 40695 34574 40704
rect 34428 40112 34480 40118
rect 34428 40054 34480 40060
rect 34428 39976 34480 39982
rect 34428 39918 34480 39924
rect 34336 39296 34388 39302
rect 34336 39238 34388 39244
rect 34348 39098 34376 39238
rect 34440 39114 34468 39918
rect 34440 39098 34560 39114
rect 34336 39092 34388 39098
rect 34336 39034 34388 39040
rect 34440 39092 34572 39098
rect 34440 39086 34520 39092
rect 34336 38956 34388 38962
rect 34256 38916 34336 38944
rect 34336 38898 34388 38904
rect 34440 38418 34468 39086
rect 34520 39034 34572 39040
rect 34428 38412 34480 38418
rect 34428 38354 34480 38360
rect 34624 38350 34652 41210
rect 34716 40882 34744 42162
rect 34808 41682 34836 43302
rect 35072 43250 35124 43256
rect 35084 43194 35112 43250
rect 35360 43194 35388 43726
rect 35440 43716 35492 43722
rect 35440 43658 35492 43664
rect 35992 43716 36044 43722
rect 35992 43658 36044 43664
rect 35452 43432 35480 43658
rect 35594 43548 35902 43557
rect 35594 43546 35600 43548
rect 35656 43546 35680 43548
rect 35736 43546 35760 43548
rect 35816 43546 35840 43548
rect 35896 43546 35902 43548
rect 35656 43494 35658 43546
rect 35838 43494 35840 43546
rect 35594 43492 35600 43494
rect 35656 43492 35680 43494
rect 35736 43492 35760 43494
rect 35816 43492 35840 43494
rect 35896 43492 35902 43494
rect 35594 43483 35902 43492
rect 36004 43450 36032 43658
rect 35992 43444 36044 43450
rect 35452 43404 35572 43432
rect 35440 43308 35492 43314
rect 35440 43250 35492 43256
rect 35084 43166 35388 43194
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 35360 42786 35388 43166
rect 35452 42906 35480 43250
rect 35544 43246 35572 43404
rect 35992 43386 36044 43392
rect 36084 43444 36136 43450
rect 36084 43386 36136 43392
rect 36096 43330 36124 43386
rect 36004 43314 36124 43330
rect 36280 43314 36308 43812
rect 35992 43308 36124 43314
rect 36044 43302 36124 43308
rect 36268 43308 36320 43314
rect 35992 43250 36044 43256
rect 36268 43250 36320 43256
rect 35532 43240 35584 43246
rect 35532 43182 35584 43188
rect 36004 43110 36032 43250
rect 35992 43104 36044 43110
rect 35992 43046 36044 43052
rect 35440 42900 35492 42906
rect 35440 42842 35492 42848
rect 35360 42758 35480 42786
rect 35072 42696 35124 42702
rect 35072 42638 35124 42644
rect 35084 42158 35112 42638
rect 35452 42276 35480 42758
rect 35992 42628 36044 42634
rect 35992 42570 36044 42576
rect 35594 42460 35902 42469
rect 35594 42458 35600 42460
rect 35656 42458 35680 42460
rect 35736 42458 35760 42460
rect 35816 42458 35840 42460
rect 35896 42458 35902 42460
rect 35656 42406 35658 42458
rect 35838 42406 35840 42458
rect 35594 42404 35600 42406
rect 35656 42404 35680 42406
rect 35736 42404 35760 42406
rect 35816 42404 35840 42406
rect 35896 42404 35902 42406
rect 35594 42395 35902 42404
rect 35452 42248 35572 42276
rect 35348 42220 35400 42226
rect 35348 42162 35400 42168
rect 35072 42152 35124 42158
rect 35072 42094 35124 42100
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34888 41812 34940 41818
rect 34888 41754 34940 41760
rect 35164 41812 35216 41818
rect 35164 41754 35216 41760
rect 34900 41721 34928 41754
rect 34886 41712 34942 41721
rect 34796 41676 34848 41682
rect 34886 41647 34942 41656
rect 34796 41618 34848 41624
rect 34796 41540 34848 41546
rect 34796 41482 34848 41488
rect 34808 41070 34836 41482
rect 34900 41274 34928 41647
rect 34980 41608 35032 41614
rect 35176 41585 35204 41754
rect 35360 41682 35388 42162
rect 35440 42016 35492 42022
rect 35440 41958 35492 41964
rect 35452 41818 35480 41958
rect 35440 41812 35492 41818
rect 35440 41754 35492 41760
rect 35348 41676 35400 41682
rect 35348 41618 35400 41624
rect 34980 41550 35032 41556
rect 35162 41576 35218 41585
rect 34888 41268 34940 41274
rect 34888 41210 34940 41216
rect 34992 41138 35020 41550
rect 35072 41540 35124 41546
rect 35360 41562 35388 41618
rect 35162 41511 35218 41520
rect 35268 41534 35388 41562
rect 35440 41608 35492 41614
rect 35440 41550 35492 41556
rect 35072 41482 35124 41488
rect 35084 41274 35112 41482
rect 35072 41268 35124 41274
rect 35072 41210 35124 41216
rect 34980 41132 35032 41138
rect 34980 41074 35032 41080
rect 34796 41064 34848 41070
rect 34796 41006 34848 41012
rect 34796 40928 34848 40934
rect 34716 40876 34796 40882
rect 34716 40870 34848 40876
rect 35268 40882 35296 41534
rect 35348 41472 35400 41478
rect 35348 41414 35400 41420
rect 35360 41274 35388 41414
rect 35348 41268 35400 41274
rect 35348 41210 35400 41216
rect 35452 41154 35480 41550
rect 35544 41478 35572 42248
rect 35624 42152 35676 42158
rect 35624 42094 35676 42100
rect 35636 41478 35664 42094
rect 35714 41712 35770 41721
rect 35714 41647 35770 41656
rect 35728 41614 35756 41647
rect 35716 41608 35768 41614
rect 35716 41550 35768 41556
rect 36004 41478 36032 42570
rect 36280 41585 36308 43250
rect 36544 43104 36596 43110
rect 36544 43046 36596 43052
rect 36556 42838 36584 43046
rect 36544 42832 36596 42838
rect 36544 42774 36596 42780
rect 36728 41812 36780 41818
rect 36728 41754 36780 41760
rect 36360 41676 36412 41682
rect 36360 41618 36412 41624
rect 36266 41576 36322 41585
rect 36266 41511 36322 41520
rect 35532 41472 35584 41478
rect 35532 41414 35584 41420
rect 35624 41472 35676 41478
rect 35624 41414 35676 41420
rect 35992 41472 36044 41478
rect 35992 41414 36044 41420
rect 35594 41372 35902 41381
rect 35594 41370 35600 41372
rect 35656 41370 35680 41372
rect 35736 41370 35760 41372
rect 35816 41370 35840 41372
rect 35896 41370 35902 41372
rect 35656 41318 35658 41370
rect 35838 41318 35840 41370
rect 35594 41316 35600 41318
rect 35656 41316 35680 41318
rect 35736 41316 35760 41318
rect 35816 41316 35840 41318
rect 35896 41316 35902 41318
rect 35594 41307 35902 41316
rect 36084 41200 36136 41206
rect 35452 41138 35572 41154
rect 36136 41148 36216 41154
rect 36084 41142 36216 41148
rect 35348 41132 35400 41138
rect 35348 41074 35400 41080
rect 35452 41132 35584 41138
rect 35452 41126 35532 41132
rect 35360 41002 35388 41074
rect 35348 40996 35400 41002
rect 35348 40938 35400 40944
rect 34716 40854 34836 40870
rect 35268 40854 35388 40882
rect 34702 40760 34758 40769
rect 34702 40695 34758 40704
rect 34612 38344 34664 38350
rect 34612 38286 34664 38292
rect 34336 38208 34388 38214
rect 34336 38150 34388 38156
rect 34244 36848 34296 36854
rect 34244 36790 34296 36796
rect 34152 36032 34204 36038
rect 34152 35974 34204 35980
rect 33600 35080 33652 35086
rect 33600 35022 33652 35028
rect 33508 33448 33560 33454
rect 33508 33390 33560 33396
rect 33508 33108 33560 33114
rect 33508 33050 33560 33056
rect 33416 32904 33468 32910
rect 33416 32846 33468 32852
rect 33428 31278 33456 32846
rect 33520 31754 33548 33050
rect 33520 31726 33732 31754
rect 33416 31272 33468 31278
rect 33416 31214 33468 31220
rect 33428 30841 33456 31214
rect 33414 30832 33470 30841
rect 33414 30767 33470 30776
rect 33048 30728 33100 30734
rect 32862 30696 32918 30705
rect 33048 30670 33100 30676
rect 33140 30728 33192 30734
rect 33140 30670 33192 30676
rect 33324 30728 33376 30734
rect 33324 30670 33376 30676
rect 32862 30631 32918 30640
rect 32772 30388 32824 30394
rect 32772 30330 32824 30336
rect 32680 28960 32732 28966
rect 32680 28902 32732 28908
rect 32692 28762 32720 28902
rect 32680 28756 32732 28762
rect 32680 28698 32732 28704
rect 32588 28620 32640 28626
rect 32588 28562 32640 28568
rect 32496 28212 32548 28218
rect 32496 28154 32548 28160
rect 32600 28150 32628 28562
rect 32680 28484 32732 28490
rect 32680 28426 32732 28432
rect 32588 28144 32640 28150
rect 32588 28086 32640 28092
rect 32128 28008 32180 28014
rect 32128 27950 32180 27956
rect 31576 27396 31628 27402
rect 31576 27338 31628 27344
rect 31852 27328 31904 27334
rect 31852 27270 31904 27276
rect 31864 26994 31892 27270
rect 31852 26988 31904 26994
rect 32140 26976 32168 27950
rect 32692 27538 32720 28426
rect 32680 27532 32732 27538
rect 32680 27474 32732 27480
rect 32692 26994 32720 27474
rect 31852 26930 31904 26936
rect 31956 26948 32168 26976
rect 32680 26988 32732 26994
rect 31298 26888 31354 26897
rect 31298 26823 31354 26832
rect 31956 26466 31984 26948
rect 32680 26930 32732 26936
rect 32036 26784 32088 26790
rect 32036 26726 32088 26732
rect 31576 26444 31628 26450
rect 31576 26386 31628 26392
rect 31864 26438 31984 26466
rect 31116 25696 31168 25702
rect 31116 25638 31168 25644
rect 31024 25288 31076 25294
rect 31024 25230 31076 25236
rect 31036 24410 31064 25230
rect 31024 24404 31076 24410
rect 31024 24346 31076 24352
rect 31392 24268 31444 24274
rect 31392 24210 31444 24216
rect 31208 24200 31260 24206
rect 31260 24160 31340 24188
rect 31208 24142 31260 24148
rect 31312 23798 31340 24160
rect 31300 23792 31352 23798
rect 31300 23734 31352 23740
rect 31208 23588 31260 23594
rect 31208 23530 31260 23536
rect 31220 23322 31248 23530
rect 31208 23316 31260 23322
rect 31208 23258 31260 23264
rect 31024 23180 31076 23186
rect 31024 23122 31076 23128
rect 31036 22982 31064 23122
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 31220 22778 31248 23258
rect 31208 22772 31260 22778
rect 31208 22714 31260 22720
rect 31312 22642 31340 23734
rect 31404 23662 31432 24210
rect 31392 23656 31444 23662
rect 31392 23598 31444 23604
rect 31404 23322 31432 23598
rect 31392 23316 31444 23322
rect 31392 23258 31444 23264
rect 31300 22636 31352 22642
rect 31300 22578 31352 22584
rect 31208 22432 31260 22438
rect 31208 22374 31260 22380
rect 31220 22234 31248 22374
rect 31208 22228 31260 22234
rect 31208 22170 31260 22176
rect 31312 22098 31340 22578
rect 31588 22137 31616 26386
rect 31864 26382 31892 26438
rect 32048 26382 32076 26726
rect 32784 26382 32812 30330
rect 33060 30190 33088 30670
rect 33152 30258 33180 30670
rect 33336 30394 33364 30670
rect 33324 30388 33376 30394
rect 33324 30330 33376 30336
rect 33140 30252 33192 30258
rect 33140 30194 33192 30200
rect 33048 30184 33100 30190
rect 33048 30126 33100 30132
rect 33324 30184 33376 30190
rect 33324 30126 33376 30132
rect 32864 30116 32916 30122
rect 32864 30058 32916 30064
rect 32876 29102 32904 30058
rect 32864 29096 32916 29102
rect 32864 29038 32916 29044
rect 33232 29096 33284 29102
rect 33232 29038 33284 29044
rect 32864 28416 32916 28422
rect 32864 28358 32916 28364
rect 32876 28150 32904 28358
rect 32864 28144 32916 28150
rect 32864 28086 32916 28092
rect 33244 27538 33272 29038
rect 33336 28626 33364 30126
rect 33600 29504 33652 29510
rect 33600 29446 33652 29452
rect 33612 29170 33640 29446
rect 33600 29164 33652 29170
rect 33600 29106 33652 29112
rect 33416 28960 33468 28966
rect 33416 28902 33468 28908
rect 33324 28620 33376 28626
rect 33324 28562 33376 28568
rect 33428 28490 33456 28902
rect 33508 28620 33560 28626
rect 33508 28562 33560 28568
rect 33416 28484 33468 28490
rect 33416 28426 33468 28432
rect 33520 27878 33548 28562
rect 33600 28144 33652 28150
rect 33600 28086 33652 28092
rect 33508 27872 33560 27878
rect 33508 27814 33560 27820
rect 33232 27532 33284 27538
rect 33232 27474 33284 27480
rect 32864 27464 32916 27470
rect 33244 27418 33272 27474
rect 33612 27470 33640 28086
rect 32864 27406 32916 27412
rect 32876 27130 32904 27406
rect 33152 27390 33272 27418
rect 33600 27464 33652 27470
rect 33600 27406 33652 27412
rect 32864 27124 32916 27130
rect 32864 27066 32916 27072
rect 31852 26376 31904 26382
rect 31852 26318 31904 26324
rect 32036 26376 32088 26382
rect 32036 26318 32088 26324
rect 32772 26376 32824 26382
rect 32772 26318 32824 26324
rect 33048 25900 33100 25906
rect 33048 25842 33100 25848
rect 33060 25294 33088 25842
rect 31760 25288 31812 25294
rect 31760 25230 31812 25236
rect 33048 25288 33100 25294
rect 33048 25230 33100 25236
rect 31668 24608 31720 24614
rect 31668 24550 31720 24556
rect 31680 24070 31708 24550
rect 31772 24206 31800 25230
rect 33152 24834 33180 27390
rect 33612 26926 33640 27406
rect 33600 26920 33652 26926
rect 33600 26862 33652 26868
rect 33704 26858 33732 31726
rect 33968 31680 34020 31686
rect 33968 31622 34020 31628
rect 33980 31414 34008 31622
rect 33784 31408 33836 31414
rect 33784 31350 33836 31356
rect 33968 31408 34020 31414
rect 33968 31350 34020 31356
rect 33796 30938 33824 31350
rect 33784 30932 33836 30938
rect 33784 30874 33836 30880
rect 34060 30048 34112 30054
rect 34060 29990 34112 29996
rect 34072 29578 34100 29990
rect 34060 29572 34112 29578
rect 34060 29514 34112 29520
rect 34164 29238 34192 35974
rect 34256 35170 34284 36790
rect 34348 36632 34376 38150
rect 34428 37800 34480 37806
rect 34428 37742 34480 37748
rect 34440 37262 34468 37742
rect 34428 37256 34480 37262
rect 34428 37198 34480 37204
rect 34520 37188 34572 37194
rect 34520 37130 34572 37136
rect 34532 36922 34560 37130
rect 34520 36916 34572 36922
rect 34520 36858 34572 36864
rect 34612 36780 34664 36786
rect 34612 36722 34664 36728
rect 34520 36644 34572 36650
rect 34348 36604 34520 36632
rect 34520 36586 34572 36592
rect 34256 35142 34376 35170
rect 34244 35080 34296 35086
rect 34244 35022 34296 35028
rect 34256 34542 34284 35022
rect 34244 34536 34296 34542
rect 34244 34478 34296 34484
rect 34244 32564 34296 32570
rect 34244 32506 34296 32512
rect 34152 29232 34204 29238
rect 34152 29174 34204 29180
rect 33876 29164 33928 29170
rect 33876 29106 33928 29112
rect 33888 28762 33916 29106
rect 33876 28756 33928 28762
rect 33876 28698 33928 28704
rect 33876 28552 33928 28558
rect 33876 28494 33928 28500
rect 33888 27470 33916 28494
rect 34060 27532 34112 27538
rect 34060 27474 34112 27480
rect 33876 27464 33928 27470
rect 33876 27406 33928 27412
rect 33692 26852 33744 26858
rect 33692 26794 33744 26800
rect 33324 26784 33376 26790
rect 33324 26726 33376 26732
rect 33336 26314 33364 26726
rect 33324 26308 33376 26314
rect 33324 26250 33376 26256
rect 33508 25832 33560 25838
rect 33508 25774 33560 25780
rect 33232 25220 33284 25226
rect 33232 25162 33284 25168
rect 33244 24954 33272 25162
rect 33232 24948 33284 24954
rect 33232 24890 33284 24896
rect 32404 24812 32456 24818
rect 32404 24754 32456 24760
rect 33060 24806 33180 24834
rect 33324 24812 33376 24818
rect 32220 24608 32272 24614
rect 32220 24550 32272 24556
rect 32232 24206 32260 24550
rect 31760 24200 31812 24206
rect 31760 24142 31812 24148
rect 32220 24200 32272 24206
rect 32220 24142 32272 24148
rect 31668 24064 31720 24070
rect 31668 24006 31720 24012
rect 31574 22128 31630 22137
rect 30944 22066 31064 22094
rect 31036 21350 31064 22066
rect 31300 22092 31352 22098
rect 31574 22063 31630 22072
rect 31300 22034 31352 22040
rect 31024 21344 31076 21350
rect 31024 21286 31076 21292
rect 31036 20074 31064 21286
rect 31392 20460 31444 20466
rect 31392 20402 31444 20408
rect 31036 20046 31248 20074
rect 31404 20058 31432 20402
rect 31116 19984 31168 19990
rect 31116 19926 31168 19932
rect 31024 19916 31076 19922
rect 31024 19858 31076 19864
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 31036 19242 31064 19858
rect 31024 19236 31076 19242
rect 31024 19178 31076 19184
rect 31128 18426 31156 19926
rect 31116 18420 31168 18426
rect 31116 18362 31168 18368
rect 30840 17672 30892 17678
rect 30840 17614 30892 17620
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 30852 17542 30880 17614
rect 30840 17536 30892 17542
rect 30840 17478 30892 17484
rect 31036 17134 31064 17614
rect 31024 17128 31076 17134
rect 31024 17070 31076 17076
rect 31116 16516 31168 16522
rect 31116 16458 31168 16464
rect 31128 16250 31156 16458
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 30760 15388 30880 15416
rect 30668 15286 30788 15314
rect 30656 15156 30708 15162
rect 30656 15098 30708 15104
rect 30564 14476 30616 14482
rect 30564 14418 30616 14424
rect 30576 12866 30604 14418
rect 30668 13938 30696 15098
rect 30760 14618 30788 15286
rect 30748 14612 30800 14618
rect 30748 14554 30800 14560
rect 30852 14482 30880 15388
rect 30932 15360 30984 15366
rect 30932 15302 30984 15308
rect 30944 15162 30972 15302
rect 30932 15156 30984 15162
rect 30932 15098 30984 15104
rect 30840 14476 30892 14482
rect 30840 14418 30892 14424
rect 30748 14340 30800 14346
rect 30748 14282 30800 14288
rect 30760 13938 30788 14282
rect 31024 14272 31076 14278
rect 31024 14214 31076 14220
rect 31036 14074 31064 14214
rect 31024 14068 31076 14074
rect 31024 14010 31076 14016
rect 31220 13954 31248 20046
rect 31392 20052 31444 20058
rect 31392 19994 31444 20000
rect 31300 19372 31352 19378
rect 31300 19314 31352 19320
rect 31312 17082 31340 19314
rect 31588 19310 31616 22063
rect 31772 21622 31800 24142
rect 32416 23866 32444 24754
rect 32956 24676 33008 24682
rect 32956 24618 33008 24624
rect 32772 24064 32824 24070
rect 32772 24006 32824 24012
rect 32784 23866 32812 24006
rect 32404 23860 32456 23866
rect 32404 23802 32456 23808
rect 32772 23860 32824 23866
rect 32772 23802 32824 23808
rect 32036 23316 32088 23322
rect 32036 23258 32088 23264
rect 31760 21616 31812 21622
rect 31760 21558 31812 21564
rect 31772 20754 31800 21558
rect 31944 20936 31996 20942
rect 31944 20878 31996 20884
rect 31956 20754 31984 20878
rect 31680 20726 31984 20754
rect 31680 20602 31708 20726
rect 31668 20596 31720 20602
rect 31668 20538 31720 20544
rect 31852 20256 31904 20262
rect 31852 20198 31904 20204
rect 31864 19961 31892 20198
rect 31850 19952 31906 19961
rect 31850 19887 31906 19896
rect 31864 19854 31892 19887
rect 31956 19854 31984 20726
rect 32048 19922 32076 23258
rect 32968 23254 32996 24618
rect 33060 24154 33088 24806
rect 33324 24754 33376 24760
rect 33232 24608 33284 24614
rect 33232 24550 33284 24556
rect 33244 24410 33272 24550
rect 33336 24410 33364 24754
rect 33416 24744 33468 24750
rect 33416 24686 33468 24692
rect 33232 24404 33284 24410
rect 33232 24346 33284 24352
rect 33324 24404 33376 24410
rect 33324 24346 33376 24352
rect 33060 24126 33180 24154
rect 33048 23656 33100 23662
rect 33048 23598 33100 23604
rect 32956 23248 33008 23254
rect 32956 23190 33008 23196
rect 32968 23118 32996 23190
rect 32956 23112 33008 23118
rect 32956 23054 33008 23060
rect 32864 23044 32916 23050
rect 32864 22986 32916 22992
rect 32876 22438 32904 22986
rect 32956 22772 33008 22778
rect 32956 22714 33008 22720
rect 32864 22432 32916 22438
rect 32864 22374 32916 22380
rect 32404 21956 32456 21962
rect 32404 21898 32456 21904
rect 32416 21690 32444 21898
rect 32968 21690 32996 22714
rect 32404 21684 32456 21690
rect 32404 21626 32456 21632
rect 32956 21684 33008 21690
rect 32956 21626 33008 21632
rect 32968 21418 32996 21626
rect 33060 21486 33088 23598
rect 33048 21480 33100 21486
rect 33048 21422 33100 21428
rect 32956 21412 33008 21418
rect 32956 21354 33008 21360
rect 32220 21344 32272 21350
rect 32220 21286 32272 21292
rect 32232 20942 32260 21286
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 33152 20398 33180 24126
rect 33324 23792 33376 23798
rect 33324 23734 33376 23740
rect 33336 23186 33364 23734
rect 33428 23662 33456 24686
rect 33520 24342 33548 25774
rect 33600 25696 33652 25702
rect 33600 25638 33652 25644
rect 33508 24336 33560 24342
rect 33508 24278 33560 24284
rect 33508 24200 33560 24206
rect 33508 24142 33560 24148
rect 33416 23656 33468 23662
rect 33416 23598 33468 23604
rect 33324 23180 33376 23186
rect 33324 23122 33376 23128
rect 33520 22094 33548 24142
rect 33612 23866 33640 25638
rect 33600 23860 33652 23866
rect 33600 23802 33652 23808
rect 33428 22066 33548 22094
rect 33704 22094 33732 26794
rect 33888 25673 33916 27406
rect 34072 26994 34100 27474
rect 34060 26988 34112 26994
rect 34060 26930 34112 26936
rect 34072 26586 34100 26930
rect 34256 26926 34284 32506
rect 34348 30938 34376 35142
rect 34428 34944 34480 34950
rect 34428 34886 34480 34892
rect 34440 33454 34468 34886
rect 34532 34202 34560 36586
rect 34624 36378 34652 36722
rect 34612 36372 34664 36378
rect 34612 36314 34664 36320
rect 34612 36236 34664 36242
rect 34612 36178 34664 36184
rect 34624 34202 34652 36178
rect 34520 34196 34572 34202
rect 34520 34138 34572 34144
rect 34612 34196 34664 34202
rect 34612 34138 34664 34144
rect 34532 33998 34560 34138
rect 34624 34066 34652 34138
rect 34612 34060 34664 34066
rect 34612 34002 34664 34008
rect 34520 33992 34572 33998
rect 34520 33934 34572 33940
rect 34428 33448 34480 33454
rect 34428 33390 34480 33396
rect 34440 32910 34468 33390
rect 34428 32904 34480 32910
rect 34428 32846 34480 32852
rect 34612 31816 34664 31822
rect 34612 31758 34664 31764
rect 34520 31748 34572 31754
rect 34520 31690 34572 31696
rect 34336 30932 34388 30938
rect 34336 30874 34388 30880
rect 34532 30870 34560 31690
rect 34624 31482 34652 31758
rect 34612 31476 34664 31482
rect 34612 31418 34664 31424
rect 34520 30864 34572 30870
rect 34716 30818 34744 40695
rect 34808 40610 34836 40854
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35360 40610 35388 40854
rect 34808 40582 34928 40610
rect 34900 40526 34928 40582
rect 35268 40582 35388 40610
rect 34888 40520 34940 40526
rect 34888 40462 34940 40468
rect 34796 40384 34848 40390
rect 34796 40326 34848 40332
rect 34808 40118 34836 40326
rect 34900 40118 34928 40462
rect 34796 40112 34848 40118
rect 34796 40054 34848 40060
rect 34888 40112 34940 40118
rect 34888 40054 34940 40060
rect 35268 40050 35296 40582
rect 35348 40520 35400 40526
rect 35348 40462 35400 40468
rect 35256 40044 35308 40050
rect 35256 39986 35308 39992
rect 34796 39976 34848 39982
rect 34796 39918 34848 39924
rect 34808 38962 34836 39918
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35164 39296 35216 39302
rect 35164 39238 35216 39244
rect 35176 38962 35204 39238
rect 35360 38962 35388 40462
rect 35452 39982 35480 41126
rect 36096 41126 36216 41142
rect 35532 41074 35584 41080
rect 35808 41064 35860 41070
rect 35808 41006 35860 41012
rect 35820 40526 35848 41006
rect 35808 40520 35860 40526
rect 35808 40462 35860 40468
rect 35594 40284 35902 40293
rect 35594 40282 35600 40284
rect 35656 40282 35680 40284
rect 35736 40282 35760 40284
rect 35816 40282 35840 40284
rect 35896 40282 35902 40284
rect 35656 40230 35658 40282
rect 35838 40230 35840 40282
rect 35594 40228 35600 40230
rect 35656 40228 35680 40230
rect 35736 40228 35760 40230
rect 35816 40228 35840 40230
rect 35896 40228 35902 40230
rect 35594 40219 35902 40228
rect 35992 40112 36044 40118
rect 35992 40054 36044 40060
rect 35440 39976 35492 39982
rect 35440 39918 35492 39924
rect 36004 39370 36032 40054
rect 35440 39364 35492 39370
rect 35440 39306 35492 39312
rect 35992 39364 36044 39370
rect 35992 39306 36044 39312
rect 34796 38956 34848 38962
rect 34796 38898 34848 38904
rect 34888 38956 34940 38962
rect 34888 38898 34940 38904
rect 35164 38956 35216 38962
rect 35164 38898 35216 38904
rect 35348 38956 35400 38962
rect 35348 38898 35400 38904
rect 34900 38842 34928 38898
rect 34808 38814 34928 38842
rect 34808 38418 34836 38814
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34796 38412 34848 38418
rect 34796 38354 34848 38360
rect 34808 36786 34836 38354
rect 35360 38350 35388 38898
rect 35452 38554 35480 39306
rect 35594 39196 35902 39205
rect 35594 39194 35600 39196
rect 35656 39194 35680 39196
rect 35736 39194 35760 39196
rect 35816 39194 35840 39196
rect 35896 39194 35902 39196
rect 35656 39142 35658 39194
rect 35838 39142 35840 39194
rect 35594 39140 35600 39142
rect 35656 39140 35680 39142
rect 35736 39140 35760 39142
rect 35816 39140 35840 39142
rect 35896 39140 35902 39142
rect 35594 39131 35902 39140
rect 36188 38962 36216 41126
rect 36268 40996 36320 41002
rect 36268 40938 36320 40944
rect 36280 40458 36308 40938
rect 36372 40934 36400 41618
rect 36452 41472 36504 41478
rect 36452 41414 36504 41420
rect 36360 40928 36412 40934
rect 36360 40870 36412 40876
rect 36372 40594 36400 40870
rect 36360 40588 36412 40594
rect 36360 40530 36412 40536
rect 36268 40452 36320 40458
rect 36268 40394 36320 40400
rect 36176 38956 36228 38962
rect 36176 38898 36228 38904
rect 35532 38888 35584 38894
rect 35532 38830 35584 38836
rect 35808 38888 35860 38894
rect 35808 38830 35860 38836
rect 35440 38548 35492 38554
rect 35440 38490 35492 38496
rect 35348 38344 35400 38350
rect 35348 38286 35400 38292
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34886 37360 34942 37369
rect 34886 37295 34942 37304
rect 34796 36780 34848 36786
rect 34796 36722 34848 36728
rect 34900 36666 34928 37295
rect 35452 36786 35480 38490
rect 35544 38214 35572 38830
rect 35820 38486 35848 38830
rect 35808 38480 35860 38486
rect 35808 38422 35860 38428
rect 35992 38276 36044 38282
rect 35992 38218 36044 38224
rect 35532 38208 35584 38214
rect 35532 38150 35584 38156
rect 35594 38108 35902 38117
rect 35594 38106 35600 38108
rect 35656 38106 35680 38108
rect 35736 38106 35760 38108
rect 35816 38106 35840 38108
rect 35896 38106 35902 38108
rect 35656 38054 35658 38106
rect 35838 38054 35840 38106
rect 35594 38052 35600 38054
rect 35656 38052 35680 38054
rect 35736 38052 35760 38054
rect 35816 38052 35840 38054
rect 35896 38052 35902 38054
rect 35594 38043 35902 38052
rect 36004 37992 36032 38218
rect 36188 38010 36216 38898
rect 35820 37964 36032 37992
rect 36176 38004 36228 38010
rect 35820 37913 35848 37964
rect 36176 37946 36228 37952
rect 35806 37904 35862 37913
rect 35806 37839 35862 37848
rect 35820 37398 35848 37839
rect 36176 37664 36228 37670
rect 36176 37606 36228 37612
rect 35808 37392 35860 37398
rect 35806 37360 35808 37369
rect 35860 37360 35862 37369
rect 35806 37295 35862 37304
rect 36084 37120 36136 37126
rect 36082 37088 36084 37097
rect 36136 37088 36138 37097
rect 35594 37020 35902 37029
rect 36082 37023 36138 37032
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 36096 36922 36124 37023
rect 36084 36916 36136 36922
rect 36084 36858 36136 36864
rect 36188 36786 36216 37606
rect 35440 36780 35492 36786
rect 35440 36722 35492 36728
rect 36176 36780 36228 36786
rect 36176 36722 36228 36728
rect 34520 30806 34572 30812
rect 34624 30790 34744 30818
rect 34808 36638 34928 36666
rect 35992 36644 36044 36650
rect 34808 30818 34836 36638
rect 35992 36586 36044 36592
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 36004 36174 36032 36586
rect 36188 36378 36216 36722
rect 36176 36372 36228 36378
rect 36176 36314 36228 36320
rect 36280 36258 36308 40394
rect 36372 40390 36400 40530
rect 36360 40384 36412 40390
rect 36360 40326 36412 40332
rect 36372 40050 36400 40326
rect 36360 40044 36412 40050
rect 36360 39986 36412 39992
rect 36372 39438 36400 39986
rect 36464 39574 36492 41414
rect 36740 41206 36768 41754
rect 36728 41200 36780 41206
rect 36728 41142 36780 41148
rect 36544 40996 36596 41002
rect 36544 40938 36596 40944
rect 36556 40594 36584 40938
rect 36740 40730 36768 41142
rect 36820 41064 36872 41070
rect 36820 41006 36872 41012
rect 36728 40724 36780 40730
rect 36728 40666 36780 40672
rect 36544 40588 36596 40594
rect 36544 40530 36596 40536
rect 36832 40526 36860 41006
rect 36728 40520 36780 40526
rect 36728 40462 36780 40468
rect 36820 40520 36872 40526
rect 36820 40462 36872 40468
rect 36740 40050 36768 40462
rect 36728 40044 36780 40050
rect 36728 39986 36780 39992
rect 36452 39568 36504 39574
rect 36452 39510 36504 39516
rect 36360 39432 36412 39438
rect 36360 39374 36412 39380
rect 36544 39432 36596 39438
rect 36544 39374 36596 39380
rect 36636 39432 36688 39438
rect 36832 39409 36860 40462
rect 36924 40390 36952 47602
rect 37280 46572 37332 46578
rect 37280 46514 37332 46520
rect 37292 45354 37320 46514
rect 37372 46436 37424 46442
rect 37372 46378 37424 46384
rect 37384 45558 37412 46378
rect 38108 45620 38160 45626
rect 38108 45562 38160 45568
rect 37372 45552 37424 45558
rect 37372 45494 37424 45500
rect 37280 45348 37332 45354
rect 37280 45290 37332 45296
rect 37384 44538 37412 45494
rect 38120 45286 38148 45562
rect 38108 45280 38160 45286
rect 38108 45222 38160 45228
rect 37372 44532 37424 44538
rect 37372 44474 37424 44480
rect 37280 44396 37332 44402
rect 37280 44338 37332 44344
rect 37292 43994 37320 44338
rect 37280 43988 37332 43994
rect 37280 43930 37332 43936
rect 37280 43784 37332 43790
rect 37280 43726 37332 43732
rect 37292 42702 37320 43726
rect 37384 43450 37412 44474
rect 37646 43752 37702 43761
rect 37646 43687 37702 43696
rect 37832 43716 37884 43722
rect 37660 43450 37688 43687
rect 37832 43658 37884 43664
rect 37372 43444 37424 43450
rect 37372 43386 37424 43392
rect 37648 43444 37700 43450
rect 37648 43386 37700 43392
rect 37384 43314 37412 43386
rect 37372 43308 37424 43314
rect 37372 43250 37424 43256
rect 37740 43240 37792 43246
rect 37740 43182 37792 43188
rect 37752 42945 37780 43182
rect 37738 42936 37794 42945
rect 37738 42871 37794 42880
rect 37280 42696 37332 42702
rect 37280 42638 37332 42644
rect 37096 42016 37148 42022
rect 37096 41958 37148 41964
rect 37004 41200 37056 41206
rect 37004 41142 37056 41148
rect 36912 40384 36964 40390
rect 36912 40326 36964 40332
rect 36912 39976 36964 39982
rect 36912 39918 36964 39924
rect 36924 39506 36952 39918
rect 36912 39500 36964 39506
rect 36912 39442 36964 39448
rect 36636 39374 36688 39380
rect 36818 39400 36874 39409
rect 36556 39273 36584 39374
rect 36648 39302 36676 39374
rect 36818 39335 36874 39344
rect 36912 39364 36964 39370
rect 36912 39306 36964 39312
rect 36636 39296 36688 39302
rect 36542 39264 36598 39273
rect 36636 39238 36688 39244
rect 36728 39296 36780 39302
rect 36728 39238 36780 39244
rect 36542 39199 36598 39208
rect 36556 39030 36584 39199
rect 36544 39024 36596 39030
rect 36544 38966 36596 38972
rect 36544 38888 36596 38894
rect 36544 38830 36596 38836
rect 36556 37874 36584 38830
rect 36544 37868 36596 37874
rect 36544 37810 36596 37816
rect 36544 37120 36596 37126
rect 36544 37062 36596 37068
rect 36452 36916 36504 36922
rect 36452 36858 36504 36864
rect 36188 36230 36308 36258
rect 35992 36168 36044 36174
rect 35992 36110 36044 36116
rect 35992 36032 36044 36038
rect 35992 35974 36044 35980
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 36004 35494 36032 35974
rect 35992 35488 36044 35494
rect 35992 35430 36044 35436
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 36004 35086 36032 35430
rect 34980 35080 35032 35086
rect 34978 35048 34980 35057
rect 35992 35080 36044 35086
rect 35032 35048 35034 35057
rect 35992 35022 36044 35028
rect 34978 34983 35034 34992
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 35808 34536 35860 34542
rect 35808 34478 35860 34484
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35820 33862 35848 34478
rect 36004 33998 36032 35022
rect 36084 34604 36136 34610
rect 36084 34546 36136 34552
rect 36096 34202 36124 34546
rect 36084 34196 36136 34202
rect 36084 34138 36136 34144
rect 35992 33992 36044 33998
rect 35992 33934 36044 33940
rect 35808 33856 35860 33862
rect 35808 33798 35860 33804
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 36004 33522 36032 33934
rect 35992 33516 36044 33522
rect 35992 33458 36044 33464
rect 36188 33454 36216 36230
rect 36268 36168 36320 36174
rect 36268 36110 36320 36116
rect 36280 35834 36308 36110
rect 36360 36032 36412 36038
rect 36360 35974 36412 35980
rect 36268 35828 36320 35834
rect 36268 35770 36320 35776
rect 36372 35766 36400 35974
rect 36360 35760 36412 35766
rect 36360 35702 36412 35708
rect 36464 34218 36492 36858
rect 36556 36310 36584 37062
rect 36648 36582 36676 39238
rect 36740 38350 36768 39238
rect 36924 38962 36952 39306
rect 36912 38956 36964 38962
rect 36912 38898 36964 38904
rect 37016 38758 37044 41142
rect 37108 40934 37136 41958
rect 37648 41812 37700 41818
rect 37648 41754 37700 41760
rect 37660 41138 37688 41754
rect 37280 41132 37332 41138
rect 37280 41074 37332 41080
rect 37648 41132 37700 41138
rect 37648 41074 37700 41080
rect 37096 40928 37148 40934
rect 37096 40870 37148 40876
rect 37108 40610 37136 40870
rect 37108 40582 37228 40610
rect 37200 40526 37228 40582
rect 37188 40520 37240 40526
rect 37188 40462 37240 40468
rect 37096 40384 37148 40390
rect 37096 40326 37148 40332
rect 37004 38752 37056 38758
rect 37004 38694 37056 38700
rect 37016 38418 37044 38694
rect 37004 38412 37056 38418
rect 37004 38354 37056 38360
rect 36728 38344 36780 38350
rect 36728 38286 36780 38292
rect 36820 38276 36872 38282
rect 36820 38218 36872 38224
rect 36728 37936 36780 37942
rect 36728 37878 36780 37884
rect 36740 37262 36768 37878
rect 36832 37874 36860 38218
rect 36912 38208 36964 38214
rect 36912 38150 36964 38156
rect 36820 37868 36872 37874
rect 36820 37810 36872 37816
rect 36728 37256 36780 37262
rect 36728 37198 36780 37204
rect 36924 36854 36952 38150
rect 37016 37942 37044 38354
rect 37004 37936 37056 37942
rect 37004 37878 37056 37884
rect 36912 36848 36964 36854
rect 36912 36790 36964 36796
rect 36636 36576 36688 36582
rect 36636 36518 36688 36524
rect 36544 36304 36596 36310
rect 36544 36246 36596 36252
rect 36820 36168 36872 36174
rect 36820 36110 36872 36116
rect 36544 36032 36596 36038
rect 36544 35974 36596 35980
rect 36556 35086 36584 35974
rect 36832 35834 36860 36110
rect 36636 35828 36688 35834
rect 36636 35770 36688 35776
rect 36820 35828 36872 35834
rect 36820 35770 36872 35776
rect 36544 35080 36596 35086
rect 36544 35022 36596 35028
rect 36648 35018 36676 35770
rect 36636 35012 36688 35018
rect 36636 34954 36688 34960
rect 36372 34190 36492 34218
rect 36176 33448 36228 33454
rect 36176 33390 36228 33396
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35992 32904 36044 32910
rect 35992 32846 36044 32852
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 35348 32360 35400 32366
rect 36004 32337 36032 32846
rect 36084 32836 36136 32842
rect 36084 32778 36136 32784
rect 35348 32302 35400 32308
rect 35990 32328 36046 32337
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34886 31920 34942 31929
rect 34886 31855 34942 31864
rect 34900 31822 34928 31855
rect 35360 31822 35388 32302
rect 35990 32263 36046 32272
rect 36096 32212 36124 32778
rect 36004 32184 36124 32212
rect 36004 31822 36032 32184
rect 34888 31816 34940 31822
rect 34888 31758 34940 31764
rect 35256 31816 35308 31822
rect 35256 31758 35308 31764
rect 35348 31816 35400 31822
rect 35348 31758 35400 31764
rect 35992 31816 36044 31822
rect 35992 31758 36044 31764
rect 36084 31816 36136 31822
rect 36084 31758 36136 31764
rect 35164 31680 35216 31686
rect 35164 31622 35216 31628
rect 35176 31142 35204 31622
rect 35268 31249 35296 31758
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35438 31512 35494 31521
rect 35594 31515 35902 31524
rect 35438 31447 35440 31456
rect 35492 31447 35494 31456
rect 35440 31418 35492 31424
rect 35346 31376 35402 31385
rect 35346 31311 35402 31320
rect 35254 31240 35310 31249
rect 35254 31175 35310 31184
rect 35164 31136 35216 31142
rect 35164 31078 35216 31084
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35072 30932 35124 30938
rect 35072 30874 35124 30880
rect 34808 30790 35020 30818
rect 34428 30388 34480 30394
rect 34428 30330 34480 30336
rect 34440 28994 34468 30330
rect 34624 29102 34652 30790
rect 34704 30728 34756 30734
rect 34704 30670 34756 30676
rect 34716 30394 34744 30670
rect 34704 30388 34756 30394
rect 34704 30330 34756 30336
rect 34704 30252 34756 30258
rect 34704 30194 34756 30200
rect 34612 29096 34664 29102
rect 34612 29038 34664 29044
rect 34440 28966 34652 28994
rect 34520 27940 34572 27946
rect 34520 27882 34572 27888
rect 34532 27606 34560 27882
rect 34520 27600 34572 27606
rect 34520 27542 34572 27548
rect 34244 26920 34296 26926
rect 34244 26862 34296 26868
rect 34060 26580 34112 26586
rect 34060 26522 34112 26528
rect 34256 26466 34284 26862
rect 34072 26438 34284 26466
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 33874 25664 33930 25673
rect 33874 25599 33930 25608
rect 33876 25492 33928 25498
rect 33876 25434 33928 25440
rect 33784 24744 33836 24750
rect 33784 24686 33836 24692
rect 33796 24410 33824 24686
rect 33784 24404 33836 24410
rect 33784 24346 33836 24352
rect 33796 23594 33824 24346
rect 33888 24206 33916 25434
rect 33980 24750 34008 26318
rect 33968 24744 34020 24750
rect 33968 24686 34020 24692
rect 33876 24200 33928 24206
rect 33876 24142 33928 24148
rect 33888 23594 33916 24142
rect 34072 23882 34100 26438
rect 34152 26376 34204 26382
rect 34152 26318 34204 26324
rect 34164 25974 34192 26318
rect 34152 25968 34204 25974
rect 34152 25910 34204 25916
rect 34428 25832 34480 25838
rect 34428 25774 34480 25780
rect 34336 25152 34388 25158
rect 34336 25094 34388 25100
rect 34348 24818 34376 25094
rect 34336 24812 34388 24818
rect 34336 24754 34388 24760
rect 34152 24744 34204 24750
rect 34152 24686 34204 24692
rect 34164 24138 34192 24686
rect 34244 24268 34296 24274
rect 34244 24210 34296 24216
rect 34152 24132 34204 24138
rect 34152 24074 34204 24080
rect 33980 23854 34100 23882
rect 33784 23588 33836 23594
rect 33784 23530 33836 23536
rect 33876 23588 33928 23594
rect 33876 23530 33928 23536
rect 33704 22066 33916 22094
rect 33324 21548 33376 21554
rect 33324 21490 33376 21496
rect 33232 21480 33284 21486
rect 33232 21422 33284 21428
rect 33140 20392 33192 20398
rect 33140 20334 33192 20340
rect 32036 19916 32088 19922
rect 32036 19858 32088 19864
rect 31852 19848 31904 19854
rect 31852 19790 31904 19796
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 31668 19372 31720 19378
rect 31668 19314 31720 19320
rect 31576 19304 31628 19310
rect 31576 19246 31628 19252
rect 31576 18828 31628 18834
rect 31576 18770 31628 18776
rect 31392 17740 31444 17746
rect 31392 17682 31444 17688
rect 31404 17202 31432 17682
rect 31392 17196 31444 17202
rect 31392 17138 31444 17144
rect 31312 17054 31432 17082
rect 31300 16992 31352 16998
rect 31300 16934 31352 16940
rect 31312 16114 31340 16934
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 31300 15088 31352 15094
rect 31300 15030 31352 15036
rect 30656 13932 30708 13938
rect 30656 13874 30708 13880
rect 30748 13932 30800 13938
rect 30748 13874 30800 13880
rect 31128 13926 31248 13954
rect 30668 13394 30696 13874
rect 30656 13388 30708 13394
rect 30656 13330 30708 13336
rect 30760 13376 30788 13874
rect 31128 13870 31156 13926
rect 31116 13864 31168 13870
rect 31116 13806 31168 13812
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 30932 13388 30984 13394
rect 30760 13348 30932 13376
rect 30760 12986 30788 13348
rect 30932 13330 30984 13336
rect 30748 12980 30800 12986
rect 30748 12922 30800 12928
rect 31036 12918 31064 13466
rect 31024 12912 31076 12918
rect 30576 12838 30880 12866
rect 31024 12854 31076 12860
rect 30472 12368 30524 12374
rect 30472 12310 30524 12316
rect 30288 12300 30340 12306
rect 30288 12242 30340 12248
rect 30196 11756 30248 11762
rect 30196 11698 30248 11704
rect 30380 11756 30432 11762
rect 30380 11698 30432 11704
rect 30392 11150 30420 11698
rect 30484 11676 30512 12310
rect 30564 11688 30616 11694
rect 30484 11648 30564 11676
rect 30564 11630 30616 11636
rect 30472 11280 30524 11286
rect 30472 11222 30524 11228
rect 30380 11144 30432 11150
rect 30380 11086 30432 11092
rect 30484 10810 30512 11222
rect 30472 10804 30524 10810
rect 30472 10746 30524 10752
rect 30104 10192 30156 10198
rect 30104 10134 30156 10140
rect 30116 8430 30144 10134
rect 30748 10124 30800 10130
rect 30668 10084 30748 10112
rect 30564 10056 30616 10062
rect 30564 9998 30616 10004
rect 30576 9926 30604 9998
rect 30564 9920 30616 9926
rect 30564 9862 30616 9868
rect 30668 8498 30696 10084
rect 30748 10066 30800 10072
rect 30852 9042 30880 12838
rect 31128 12730 31156 13806
rect 31312 13394 31340 15030
rect 31300 13388 31352 13394
rect 31300 13330 31352 13336
rect 31036 12702 31156 12730
rect 31036 12458 31064 12702
rect 31312 12594 31340 13330
rect 30944 12430 31064 12458
rect 31128 12566 31340 12594
rect 30840 9036 30892 9042
rect 30840 8978 30892 8984
rect 30748 8832 30800 8838
rect 30748 8774 30800 8780
rect 30656 8492 30708 8498
rect 30656 8434 30708 8440
rect 30104 8424 30156 8430
rect 30104 8366 30156 8372
rect 30380 8424 30432 8430
rect 30380 8366 30432 8372
rect 30564 8424 30616 8430
rect 30564 8366 30616 8372
rect 30194 7984 30250 7993
rect 30104 7948 30156 7954
rect 30392 7970 30420 8366
rect 30250 7942 30328 7970
rect 30392 7942 30512 7970
rect 30576 7954 30604 8366
rect 30760 8090 30788 8774
rect 30852 8294 30880 8978
rect 30840 8288 30892 8294
rect 30840 8230 30892 8236
rect 30748 8084 30800 8090
rect 30748 8026 30800 8032
rect 30944 7970 30972 12430
rect 31128 10130 31156 12566
rect 31404 11762 31432 17054
rect 31588 16590 31616 18770
rect 31680 17814 31708 19314
rect 31852 19304 31904 19310
rect 31852 19246 31904 19252
rect 31760 18760 31812 18766
rect 31760 18702 31812 18708
rect 31772 18426 31800 18702
rect 31760 18420 31812 18426
rect 31760 18362 31812 18368
rect 31668 17808 31720 17814
rect 31668 17750 31720 17756
rect 31576 16584 31628 16590
rect 31576 16526 31628 16532
rect 31588 16114 31616 16526
rect 31576 16108 31628 16114
rect 31576 16050 31628 16056
rect 31864 14482 31892 19246
rect 31944 16176 31996 16182
rect 31944 16118 31996 16124
rect 31956 15366 31984 16118
rect 32048 15570 32076 19858
rect 32496 19712 32548 19718
rect 32496 19654 32548 19660
rect 32508 18698 32536 19654
rect 32496 18692 32548 18698
rect 32496 18634 32548 18640
rect 32508 18426 32536 18634
rect 32588 18624 32640 18630
rect 32588 18566 32640 18572
rect 32600 18426 32628 18566
rect 32496 18420 32548 18426
rect 32496 18362 32548 18368
rect 32588 18420 32640 18426
rect 32588 18362 32640 18368
rect 33140 18148 33192 18154
rect 33140 18090 33192 18096
rect 32128 17264 32180 17270
rect 32128 17206 32180 17212
rect 32140 16794 32168 17206
rect 32864 16992 32916 16998
rect 32864 16934 32916 16940
rect 32128 16788 32180 16794
rect 32128 16730 32180 16736
rect 32876 16590 32904 16934
rect 32864 16584 32916 16590
rect 32864 16526 32916 16532
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 32416 15706 32444 16050
rect 32404 15700 32456 15706
rect 32404 15642 32456 15648
rect 32036 15564 32088 15570
rect 32036 15506 32088 15512
rect 31944 15360 31996 15366
rect 31944 15302 31996 15308
rect 32496 15360 32548 15366
rect 32496 15302 32548 15308
rect 32508 14482 32536 15302
rect 33152 15178 33180 18090
rect 33244 17202 33272 21422
rect 33336 21078 33364 21490
rect 33324 21072 33376 21078
rect 33324 21014 33376 21020
rect 33428 20890 33456 22066
rect 33784 22024 33836 22030
rect 33784 21966 33836 21972
rect 33600 21684 33652 21690
rect 33600 21626 33652 21632
rect 33508 21344 33560 21350
rect 33508 21286 33560 21292
rect 33520 21146 33548 21286
rect 33508 21140 33560 21146
rect 33508 21082 33560 21088
rect 33336 20862 33456 20890
rect 33506 20904 33562 20913
rect 33336 18154 33364 20862
rect 33506 20839 33562 20848
rect 33416 20800 33468 20806
rect 33416 20742 33468 20748
rect 33428 19854 33456 20742
rect 33520 20346 33548 20839
rect 33612 20466 33640 21626
rect 33692 21480 33744 21486
rect 33692 21422 33744 21428
rect 33704 20602 33732 21422
rect 33692 20596 33744 20602
rect 33692 20538 33744 20544
rect 33600 20460 33652 20466
rect 33600 20402 33652 20408
rect 33520 20318 33640 20346
rect 33416 19848 33468 19854
rect 33416 19790 33468 19796
rect 33508 19304 33560 19310
rect 33508 19246 33560 19252
rect 33520 18222 33548 19246
rect 33508 18216 33560 18222
rect 33508 18158 33560 18164
rect 33612 18170 33640 20318
rect 33692 19304 33744 19310
rect 33796 19281 33824 21966
rect 33888 21593 33916 22066
rect 33980 22030 34008 23854
rect 34164 23662 34192 24074
rect 34152 23656 34204 23662
rect 34152 23598 34204 23604
rect 34060 23248 34112 23254
rect 34060 23190 34112 23196
rect 33968 22024 34020 22030
rect 33968 21966 34020 21972
rect 33968 21888 34020 21894
rect 33968 21830 34020 21836
rect 33874 21584 33930 21593
rect 33874 21519 33930 21528
rect 33888 19310 33916 21519
rect 33980 21418 34008 21830
rect 34072 21486 34100 23190
rect 34060 21480 34112 21486
rect 34060 21422 34112 21428
rect 33968 21412 34020 21418
rect 33968 21354 34020 21360
rect 33980 21146 34008 21354
rect 33968 21140 34020 21146
rect 33968 21082 34020 21088
rect 33980 21010 34008 21082
rect 34150 21040 34206 21049
rect 33968 21004 34020 21010
rect 34256 21010 34284 24210
rect 34336 24132 34388 24138
rect 34336 24074 34388 24080
rect 34348 23730 34376 24074
rect 34336 23724 34388 23730
rect 34336 23666 34388 23672
rect 34440 21706 34468 25774
rect 34520 25152 34572 25158
rect 34520 25094 34572 25100
rect 34532 24206 34560 25094
rect 34624 24857 34652 28966
rect 34716 28257 34744 30194
rect 34992 30138 35020 30790
rect 35084 30734 35112 30874
rect 35162 30832 35218 30841
rect 35162 30767 35218 30776
rect 35176 30734 35204 30767
rect 35072 30728 35124 30734
rect 35072 30670 35124 30676
rect 35164 30728 35216 30734
rect 35164 30670 35216 30676
rect 35084 30258 35112 30670
rect 35072 30252 35124 30258
rect 35072 30194 35124 30200
rect 34808 30110 35020 30138
rect 34702 28248 34758 28257
rect 34702 28183 34758 28192
rect 34716 25838 34744 28183
rect 34704 25832 34756 25838
rect 34704 25774 34756 25780
rect 34610 24848 34666 24857
rect 34610 24783 34612 24792
rect 34664 24783 34666 24792
rect 34612 24754 34664 24760
rect 34808 24698 34836 30110
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35164 27464 35216 27470
rect 35164 27406 35216 27412
rect 35176 27130 35204 27406
rect 35164 27124 35216 27130
rect 35164 27066 35216 27072
rect 35360 26926 35388 31311
rect 35452 30938 35480 31418
rect 35714 31376 35770 31385
rect 35714 31311 35770 31320
rect 35728 31278 35756 31311
rect 35716 31272 35768 31278
rect 35716 31214 35768 31220
rect 35624 31204 35676 31210
rect 35624 31146 35676 31152
rect 35440 30932 35492 30938
rect 35440 30874 35492 30880
rect 35636 30598 35664 31146
rect 36004 30818 36032 31758
rect 36096 31414 36124 31758
rect 36372 31754 36400 34190
rect 36544 32224 36596 32230
rect 36544 32166 36596 32172
rect 36280 31726 36400 31754
rect 36084 31408 36136 31414
rect 36084 31350 36136 31356
rect 36004 30790 36216 30818
rect 35992 30728 36044 30734
rect 35992 30670 36044 30676
rect 36084 30728 36136 30734
rect 36084 30670 36136 30676
rect 35624 30592 35676 30598
rect 35624 30534 35676 30540
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 35624 30116 35676 30122
rect 35624 30058 35676 30064
rect 35438 29744 35494 29753
rect 35438 29679 35494 29688
rect 35452 29646 35480 29679
rect 35636 29646 35664 30058
rect 36004 29646 36032 30670
rect 35440 29640 35492 29646
rect 35440 29582 35492 29588
rect 35624 29640 35676 29646
rect 35624 29582 35676 29588
rect 35992 29640 36044 29646
rect 35992 29582 36044 29588
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 35992 29096 36044 29102
rect 35806 29064 35862 29073
rect 35992 29038 36044 29044
rect 35806 28999 35862 29008
rect 35820 28762 35848 28999
rect 35808 28756 35860 28762
rect 35808 28698 35860 28704
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 35440 28008 35492 28014
rect 35440 27950 35492 27956
rect 35452 27384 35480 27950
rect 35624 27396 35676 27402
rect 35452 27356 35624 27384
rect 35452 26994 35480 27356
rect 35624 27338 35676 27344
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35440 26988 35492 26994
rect 35440 26930 35492 26936
rect 35348 26920 35400 26926
rect 35348 26862 35400 26868
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35360 26586 35388 26862
rect 35348 26580 35400 26586
rect 35348 26522 35400 26528
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35348 25288 35400 25294
rect 35348 25230 35400 25236
rect 34716 24670 34836 24698
rect 34520 24200 34572 24206
rect 34520 24142 34572 24148
rect 34716 24154 34744 24670
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34716 24126 34836 24154
rect 34704 24064 34756 24070
rect 34704 24006 34756 24012
rect 34612 23860 34664 23866
rect 34612 23802 34664 23808
rect 34624 23662 34652 23802
rect 34612 23656 34664 23662
rect 34612 23598 34664 23604
rect 34624 22166 34652 23598
rect 34716 23186 34744 24006
rect 34704 23180 34756 23186
rect 34704 23122 34756 23128
rect 34612 22160 34664 22166
rect 34612 22102 34664 22108
rect 34612 21956 34664 21962
rect 34612 21898 34664 21904
rect 34624 21842 34652 21898
rect 34624 21814 34744 21842
rect 34440 21678 34652 21706
rect 34336 21480 34388 21486
rect 34520 21480 34572 21486
rect 34388 21440 34468 21468
rect 34336 21422 34388 21428
rect 34150 20975 34206 20984
rect 34244 21004 34296 21010
rect 33968 20946 34020 20952
rect 34164 20806 34192 20975
rect 34244 20946 34296 20952
rect 34336 21004 34388 21010
rect 34336 20946 34388 20952
rect 34256 20913 34284 20946
rect 34242 20904 34298 20913
rect 34242 20839 34298 20848
rect 34152 20800 34204 20806
rect 34152 20742 34204 20748
rect 34348 20602 34376 20946
rect 34440 20874 34468 21440
rect 34520 21422 34572 21428
rect 34532 21078 34560 21422
rect 34520 21072 34572 21078
rect 34520 21014 34572 21020
rect 34428 20868 34480 20874
rect 34428 20810 34480 20816
rect 34336 20596 34388 20602
rect 34336 20538 34388 20544
rect 34440 20398 34468 20810
rect 34532 20466 34560 21014
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34428 20392 34480 20398
rect 34428 20334 34480 20340
rect 33968 20324 34020 20330
rect 33968 20266 34020 20272
rect 33876 19304 33928 19310
rect 33692 19246 33744 19252
rect 33782 19272 33838 19281
rect 33704 18426 33732 19246
rect 33876 19246 33928 19252
rect 33782 19207 33838 19216
rect 33784 18760 33836 18766
rect 33782 18728 33784 18737
rect 33836 18728 33838 18737
rect 33782 18663 33838 18672
rect 33692 18420 33744 18426
rect 33692 18362 33744 18368
rect 33704 18290 33732 18362
rect 33692 18284 33744 18290
rect 33692 18226 33744 18232
rect 33876 18216 33928 18222
rect 33324 18148 33376 18154
rect 33612 18142 33732 18170
rect 33876 18158 33928 18164
rect 33324 18090 33376 18096
rect 33232 17196 33284 17202
rect 33232 17138 33284 17144
rect 33600 17128 33652 17134
rect 33600 17070 33652 17076
rect 33060 15150 33180 15178
rect 31852 14476 31904 14482
rect 31852 14418 31904 14424
rect 32036 14476 32088 14482
rect 32036 14418 32088 14424
rect 32496 14476 32548 14482
rect 32496 14418 32548 14424
rect 31852 14272 31904 14278
rect 31852 14214 31904 14220
rect 31864 13530 31892 14214
rect 31944 13728 31996 13734
rect 31944 13670 31996 13676
rect 31852 13524 31904 13530
rect 31852 13466 31904 13472
rect 31668 13388 31720 13394
rect 31668 13330 31720 13336
rect 31484 12640 31536 12646
rect 31482 12608 31484 12617
rect 31536 12608 31538 12617
rect 31482 12543 31538 12552
rect 31576 11824 31628 11830
rect 31576 11766 31628 11772
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 31392 11552 31444 11558
rect 31392 11494 31444 11500
rect 31208 11076 31260 11082
rect 31208 11018 31260 11024
rect 31220 10810 31248 11018
rect 31208 10804 31260 10810
rect 31208 10746 31260 10752
rect 31404 10674 31432 11494
rect 31588 11354 31616 11766
rect 31576 11348 31628 11354
rect 31576 11290 31628 11296
rect 31680 11150 31708 13330
rect 31956 13326 31984 13670
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31852 11892 31904 11898
rect 31852 11834 31904 11840
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 31392 10668 31444 10674
rect 31392 10610 31444 10616
rect 31484 10464 31536 10470
rect 31484 10406 31536 10412
rect 31496 10198 31524 10406
rect 31484 10192 31536 10198
rect 31484 10134 31536 10140
rect 31116 10124 31168 10130
rect 31116 10066 31168 10072
rect 31300 9580 31352 9586
rect 31300 9522 31352 9528
rect 31024 8968 31076 8974
rect 31024 8910 31076 8916
rect 30194 7919 30196 7928
rect 30104 7890 30156 7896
rect 30248 7919 30250 7928
rect 30196 7890 30248 7896
rect 30116 7834 30144 7890
rect 30116 7806 30236 7834
rect 30208 7478 30236 7806
rect 30196 7472 30248 7478
rect 30196 7414 30248 7420
rect 30012 7404 30064 7410
rect 30012 7346 30064 7352
rect 30208 6458 30236 7414
rect 30300 6662 30328 7942
rect 30484 7886 30512 7942
rect 30564 7948 30616 7954
rect 30564 7890 30616 7896
rect 30760 7942 30972 7970
rect 30760 7886 30788 7942
rect 30472 7880 30524 7886
rect 30472 7822 30524 7828
rect 30748 7880 30800 7886
rect 30748 7822 30800 7828
rect 30484 7274 30512 7822
rect 30472 7268 30524 7274
rect 30472 7210 30524 7216
rect 30760 6730 30788 7822
rect 30840 7200 30892 7206
rect 30840 7142 30892 7148
rect 30852 6798 30880 7142
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30748 6724 30800 6730
rect 30748 6666 30800 6672
rect 30288 6656 30340 6662
rect 30288 6598 30340 6604
rect 30656 6656 30708 6662
rect 30656 6598 30708 6604
rect 30196 6452 30248 6458
rect 30196 6394 30248 6400
rect 30668 6390 30696 6598
rect 30656 6384 30708 6390
rect 30656 6326 30708 6332
rect 31036 5642 31064 8910
rect 31312 8634 31340 9522
rect 31300 8628 31352 8634
rect 31300 8570 31352 8576
rect 31208 7744 31260 7750
rect 31208 7686 31260 7692
rect 31220 7206 31248 7686
rect 31208 7200 31260 7206
rect 31208 7142 31260 7148
rect 31484 6316 31536 6322
rect 31484 6258 31536 6264
rect 31300 6112 31352 6118
rect 31300 6054 31352 6060
rect 31312 5710 31340 6054
rect 31300 5704 31352 5710
rect 31300 5646 31352 5652
rect 31024 5636 31076 5642
rect 31024 5578 31076 5584
rect 31496 5370 31524 6258
rect 31484 5364 31536 5370
rect 31484 5306 31536 5312
rect 30196 5160 30248 5166
rect 30196 5102 30248 5108
rect 29920 4616 29972 4622
rect 29920 4558 29972 4564
rect 29828 4480 29880 4486
rect 29828 4422 29880 4428
rect 29368 3596 29420 3602
rect 29368 3538 29420 3544
rect 29840 3534 29868 4422
rect 29932 4010 29960 4558
rect 29920 4004 29972 4010
rect 29920 3946 29972 3952
rect 30208 3602 30236 5102
rect 31864 4826 31892 11834
rect 32048 10130 32076 14418
rect 32508 14074 32536 14418
rect 32496 14068 32548 14074
rect 32496 14010 32548 14016
rect 32680 13864 32732 13870
rect 32680 13806 32732 13812
rect 32692 12918 32720 13806
rect 32680 12912 32732 12918
rect 32680 12854 32732 12860
rect 33060 12434 33088 15150
rect 33508 14612 33560 14618
rect 33508 14554 33560 14560
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 33324 13932 33376 13938
rect 33324 13874 33376 13880
rect 33244 13530 33272 13874
rect 33232 13524 33284 13530
rect 33232 13466 33284 13472
rect 33140 13456 33192 13462
rect 33140 13398 33192 13404
rect 33152 12986 33180 13398
rect 33140 12980 33192 12986
rect 33140 12922 33192 12928
rect 33336 12866 33364 13874
rect 33520 13870 33548 14554
rect 33508 13864 33560 13870
rect 33508 13806 33560 13812
rect 33416 13728 33468 13734
rect 33416 13670 33468 13676
rect 33428 13190 33456 13670
rect 33416 13184 33468 13190
rect 33416 13126 33468 13132
rect 32876 12406 33088 12434
rect 33152 12838 33364 12866
rect 32772 12232 32824 12238
rect 32772 12174 32824 12180
rect 32496 11756 32548 11762
rect 32548 11716 32628 11744
rect 32496 11698 32548 11704
rect 32036 10124 32088 10130
rect 32036 10066 32088 10072
rect 31944 9648 31996 9654
rect 31944 9590 31996 9596
rect 31956 9178 31984 9590
rect 32048 9518 32076 10066
rect 32036 9512 32088 9518
rect 32036 9454 32088 9460
rect 32128 9512 32180 9518
rect 32128 9454 32180 9460
rect 32312 9512 32364 9518
rect 32312 9454 32364 9460
rect 31944 9172 31996 9178
rect 31944 9114 31996 9120
rect 31944 7404 31996 7410
rect 31944 7346 31996 7352
rect 31956 7002 31984 7346
rect 31944 6996 31996 7002
rect 31944 6938 31996 6944
rect 32140 6390 32168 9454
rect 32220 8968 32272 8974
rect 32324 8956 32352 9454
rect 32272 8928 32352 8956
rect 32220 8910 32272 8916
rect 32232 7410 32260 8910
rect 32404 8900 32456 8906
rect 32404 8842 32456 8848
rect 32416 8634 32444 8842
rect 32404 8628 32456 8634
rect 32404 8570 32456 8576
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 32508 8090 32536 8434
rect 32496 8084 32548 8090
rect 32496 8026 32548 8032
rect 32220 7404 32272 7410
rect 32220 7346 32272 7352
rect 32128 6384 32180 6390
rect 32128 6326 32180 6332
rect 32128 5160 32180 5166
rect 32128 5102 32180 5108
rect 31852 4820 31904 4826
rect 31852 4762 31904 4768
rect 32140 4690 32168 5102
rect 32128 4684 32180 4690
rect 32128 4626 32180 4632
rect 32036 4616 32088 4622
rect 32036 4558 32088 4564
rect 31852 4480 31904 4486
rect 31852 4422 31904 4428
rect 31864 4214 31892 4422
rect 31852 4208 31904 4214
rect 31852 4150 31904 4156
rect 31024 4140 31076 4146
rect 31024 4082 31076 4088
rect 31944 4140 31996 4146
rect 31944 4082 31996 4088
rect 30748 3936 30800 3942
rect 30748 3878 30800 3884
rect 30012 3596 30064 3602
rect 30012 3538 30064 3544
rect 30196 3596 30248 3602
rect 30196 3538 30248 3544
rect 29828 3528 29880 3534
rect 29828 3470 29880 3476
rect 29368 3392 29420 3398
rect 29368 3334 29420 3340
rect 29184 3052 29236 3058
rect 29184 2994 29236 3000
rect 28684 2808 28856 2836
rect 28632 2790 28684 2796
rect 22480 2638 22876 2666
rect 20994 2615 21050 2624
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 21008 2446 21036 2615
rect 28644 2446 28672 2790
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 16132 800 16160 2382
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18708 800 18736 2246
rect 20640 800 20668 2314
rect 23216 800 23244 2382
rect 25148 800 25176 2382
rect 29196 2310 29224 2994
rect 29380 2446 29408 3334
rect 30024 3194 30052 3538
rect 30760 3534 30788 3878
rect 30564 3528 30616 3534
rect 30564 3470 30616 3476
rect 30748 3528 30800 3534
rect 30748 3470 30800 3476
rect 30012 3188 30064 3194
rect 30012 3130 30064 3136
rect 30576 3126 30604 3470
rect 31036 3194 31064 4082
rect 31956 3738 31984 4082
rect 32048 3738 32076 4558
rect 32140 3942 32168 4626
rect 32232 4146 32260 7346
rect 32600 6866 32628 11716
rect 32680 11552 32732 11558
rect 32680 11494 32732 11500
rect 32692 11150 32720 11494
rect 32680 11144 32732 11150
rect 32680 11086 32732 11092
rect 32680 8424 32732 8430
rect 32680 8366 32732 8372
rect 32692 7886 32720 8366
rect 32784 7954 32812 12174
rect 32772 7948 32824 7954
rect 32772 7890 32824 7896
rect 32680 7880 32732 7886
rect 32680 7822 32732 7828
rect 32692 7410 32720 7822
rect 32680 7404 32732 7410
rect 32680 7346 32732 7352
rect 32588 6860 32640 6866
rect 32588 6802 32640 6808
rect 32312 5160 32364 5166
rect 32312 5102 32364 5108
rect 32324 4622 32352 5102
rect 32312 4616 32364 4622
rect 32312 4558 32364 4564
rect 32220 4140 32272 4146
rect 32220 4082 32272 4088
rect 32128 3936 32180 3942
rect 32128 3878 32180 3884
rect 31944 3732 31996 3738
rect 31944 3674 31996 3680
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 31852 3664 31904 3670
rect 31852 3606 31904 3612
rect 31760 3596 31812 3602
rect 31760 3538 31812 3544
rect 31666 3496 31722 3505
rect 31484 3460 31536 3466
rect 31666 3431 31722 3440
rect 31484 3402 31536 3408
rect 31024 3188 31076 3194
rect 31024 3130 31076 3136
rect 31496 3126 31524 3402
rect 30564 3120 30616 3126
rect 30564 3062 30616 3068
rect 31484 3120 31536 3126
rect 31484 3062 31536 3068
rect 31680 2854 31708 3431
rect 31772 3398 31800 3538
rect 31760 3392 31812 3398
rect 31760 3334 31812 3340
rect 31772 2990 31800 3334
rect 31864 3194 31892 3606
rect 31956 3482 31984 3674
rect 31956 3454 32076 3482
rect 31944 3392 31996 3398
rect 31944 3334 31996 3340
rect 31852 3188 31904 3194
rect 31852 3130 31904 3136
rect 31956 3126 31984 3334
rect 31944 3120 31996 3126
rect 31944 3062 31996 3068
rect 32048 3058 32076 3454
rect 32140 3398 32168 3878
rect 32600 3602 32628 6802
rect 32678 4720 32734 4729
rect 32678 4655 32680 4664
rect 32732 4655 32734 4664
rect 32680 4626 32732 4632
rect 32784 4010 32812 7890
rect 32876 4758 32904 12406
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 32956 8288 33008 8294
rect 32956 8230 33008 8236
rect 32968 7954 32996 8230
rect 33060 8090 33088 8774
rect 33152 8129 33180 12838
rect 33520 12782 33548 13806
rect 33508 12776 33560 12782
rect 33508 12718 33560 12724
rect 33232 12708 33284 12714
rect 33284 12668 33456 12696
rect 33232 12650 33284 12656
rect 33232 11076 33284 11082
rect 33232 11018 33284 11024
rect 33244 10674 33272 11018
rect 33232 10668 33284 10674
rect 33232 10610 33284 10616
rect 33324 9920 33376 9926
rect 33324 9862 33376 9868
rect 33138 8120 33194 8129
rect 33048 8084 33100 8090
rect 33138 8055 33194 8064
rect 33048 8026 33100 8032
rect 32956 7948 33008 7954
rect 32956 7890 33008 7896
rect 33048 7880 33100 7886
rect 33152 7834 33180 8055
rect 33100 7828 33180 7834
rect 33048 7822 33180 7828
rect 33060 7806 33180 7822
rect 33140 7744 33192 7750
rect 33140 7686 33192 7692
rect 33048 6996 33100 7002
rect 33048 6938 33100 6944
rect 33060 6390 33088 6938
rect 33152 6934 33180 7686
rect 33232 7200 33284 7206
rect 33232 7142 33284 7148
rect 33140 6928 33192 6934
rect 33140 6870 33192 6876
rect 33244 6866 33272 7142
rect 33232 6860 33284 6866
rect 33232 6802 33284 6808
rect 33048 6384 33100 6390
rect 33048 6326 33100 6332
rect 33336 5370 33364 9862
rect 33428 8362 33456 12668
rect 33612 12170 33640 17070
rect 33704 15570 33732 18142
rect 33888 17610 33916 18158
rect 33876 17604 33928 17610
rect 33876 17546 33928 17552
rect 33692 15564 33744 15570
rect 33692 15506 33744 15512
rect 33704 12442 33732 15506
rect 33784 15020 33836 15026
rect 33784 14962 33836 14968
rect 33796 13841 33824 14962
rect 33980 13870 34008 20266
rect 34440 20058 34468 20334
rect 34428 20052 34480 20058
rect 34428 19994 34480 20000
rect 34060 19508 34112 19514
rect 34060 19450 34112 19456
rect 34072 18086 34100 19450
rect 34244 19304 34296 19310
rect 34520 19304 34572 19310
rect 34244 19246 34296 19252
rect 34440 19264 34520 19292
rect 34152 18760 34204 18766
rect 34152 18702 34204 18708
rect 34060 18080 34112 18086
rect 34060 18022 34112 18028
rect 34164 17134 34192 18702
rect 34256 18222 34284 19246
rect 34336 18760 34388 18766
rect 34336 18702 34388 18708
rect 34244 18216 34296 18222
rect 34244 18158 34296 18164
rect 34152 17128 34204 17134
rect 34152 17070 34204 17076
rect 34152 16992 34204 16998
rect 34152 16934 34204 16940
rect 34060 16516 34112 16522
rect 34060 16458 34112 16464
rect 34072 16250 34100 16458
rect 34060 16244 34112 16250
rect 34060 16186 34112 16192
rect 34164 14822 34192 16934
rect 34256 16454 34284 18158
rect 34348 17202 34376 18702
rect 34440 18272 34468 19264
rect 34520 19246 34572 19252
rect 34520 18284 34572 18290
rect 34440 18244 34520 18272
rect 34440 17338 34468 18244
rect 34520 18226 34572 18232
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 34428 17332 34480 17338
rect 34428 17274 34480 17280
rect 34336 17196 34388 17202
rect 34336 17138 34388 17144
rect 34336 17060 34388 17066
rect 34336 17002 34388 17008
rect 34348 16590 34376 17002
rect 34440 16794 34468 17274
rect 34428 16788 34480 16794
rect 34428 16730 34480 16736
rect 34336 16584 34388 16590
rect 34336 16526 34388 16532
rect 34244 16448 34296 16454
rect 34244 16390 34296 16396
rect 34348 16114 34376 16526
rect 34428 16448 34480 16454
rect 34428 16390 34480 16396
rect 34244 16108 34296 16114
rect 34244 16050 34296 16056
rect 34336 16108 34388 16114
rect 34336 16050 34388 16056
rect 34256 15706 34284 16050
rect 34244 15700 34296 15706
rect 34244 15642 34296 15648
rect 34440 15502 34468 16390
rect 34532 15994 34560 17614
rect 34624 17082 34652 21678
rect 34716 20602 34744 21814
rect 34704 20596 34756 20602
rect 34704 20538 34756 20544
rect 34702 20496 34758 20505
rect 34702 20431 34704 20440
rect 34756 20431 34758 20440
rect 34704 20402 34756 20408
rect 34716 17678 34744 20402
rect 34704 17672 34756 17678
rect 34704 17614 34756 17620
rect 34704 17536 34756 17542
rect 34704 17478 34756 17484
rect 34716 17202 34744 17478
rect 34704 17196 34756 17202
rect 34704 17138 34756 17144
rect 34624 17054 34744 17082
rect 34612 16584 34664 16590
rect 34612 16526 34664 16532
rect 34624 16182 34652 16526
rect 34612 16176 34664 16182
rect 34612 16118 34664 16124
rect 34532 15966 34652 15994
rect 34428 15496 34480 15502
rect 34428 15438 34480 15444
rect 34152 14816 34204 14822
rect 34152 14758 34204 14764
rect 34336 14816 34388 14822
rect 34336 14758 34388 14764
rect 34244 14476 34296 14482
rect 34244 14418 34296 14424
rect 33968 13864 34020 13870
rect 33782 13832 33838 13841
rect 33968 13806 34020 13812
rect 34152 13864 34204 13870
rect 34152 13806 34204 13812
rect 33782 13767 33838 13776
rect 33876 13796 33928 13802
rect 33876 13738 33928 13744
rect 33888 13258 33916 13738
rect 33876 13252 33928 13258
rect 33876 13194 33928 13200
rect 33888 12986 33916 13194
rect 33968 13184 34020 13190
rect 33968 13126 34020 13132
rect 33876 12980 33928 12986
rect 33876 12922 33928 12928
rect 33980 12866 34008 13126
rect 33796 12838 34008 12866
rect 34164 12850 34192 13806
rect 34256 13394 34284 14418
rect 34348 13394 34376 14758
rect 34520 14272 34572 14278
rect 34520 14214 34572 14220
rect 34428 13864 34480 13870
rect 34428 13806 34480 13812
rect 34244 13388 34296 13394
rect 34244 13330 34296 13336
rect 34336 13388 34388 13394
rect 34336 13330 34388 13336
rect 34152 12844 34204 12850
rect 33796 12782 33824 12838
rect 34152 12786 34204 12792
rect 33784 12776 33836 12782
rect 33784 12718 33836 12724
rect 33968 12776 34020 12782
rect 33968 12718 34020 12724
rect 33980 12594 34008 12718
rect 34058 12608 34114 12617
rect 33980 12566 34058 12594
rect 34058 12543 34114 12552
rect 33692 12436 33744 12442
rect 33692 12378 33744 12384
rect 33600 12164 33652 12170
rect 33600 12106 33652 12112
rect 33612 11694 33640 12106
rect 33704 12102 33732 12378
rect 33692 12096 33744 12102
rect 33692 12038 33744 12044
rect 33704 11694 33732 12038
rect 33600 11688 33652 11694
rect 33600 11630 33652 11636
rect 33692 11688 33744 11694
rect 33692 11630 33744 11636
rect 33600 8832 33652 8838
rect 33600 8774 33652 8780
rect 33612 8378 33640 8774
rect 34072 8650 34100 12543
rect 34164 11762 34192 12786
rect 34256 11898 34284 13330
rect 34348 13190 34376 13330
rect 34336 13184 34388 13190
rect 34336 13126 34388 13132
rect 34440 12866 34468 13806
rect 34532 12986 34560 14214
rect 34624 13938 34652 15966
rect 34612 13932 34664 13938
rect 34612 13874 34664 13880
rect 34520 12980 34572 12986
rect 34520 12922 34572 12928
rect 34348 12850 34468 12866
rect 34336 12844 34468 12850
rect 34388 12838 34468 12844
rect 34336 12786 34388 12792
rect 34440 12434 34468 12838
rect 34624 12434 34652 13874
rect 34348 12406 34468 12434
rect 34532 12406 34652 12434
rect 34244 11892 34296 11898
rect 34244 11834 34296 11840
rect 34348 11830 34376 12406
rect 34336 11824 34388 11830
rect 34336 11766 34388 11772
rect 34152 11756 34204 11762
rect 34152 11698 34204 11704
rect 34164 10810 34192 11698
rect 34348 11354 34376 11766
rect 34428 11552 34480 11558
rect 34428 11494 34480 11500
rect 34336 11348 34388 11354
rect 34336 11290 34388 11296
rect 34440 11150 34468 11494
rect 34428 11144 34480 11150
rect 34428 11086 34480 11092
rect 34244 11008 34296 11014
rect 34244 10950 34296 10956
rect 34152 10804 34204 10810
rect 34152 10746 34204 10752
rect 34256 10742 34284 10950
rect 34244 10736 34296 10742
rect 34244 10678 34296 10684
rect 34072 8622 34192 8650
rect 34164 8498 34192 8622
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 33692 8424 33744 8430
rect 33612 8372 33692 8378
rect 33612 8366 33744 8372
rect 33968 8424 34020 8430
rect 33968 8366 34020 8372
rect 33416 8356 33468 8362
rect 33416 8298 33468 8304
rect 33612 8350 33732 8366
rect 33324 5364 33376 5370
rect 33324 5306 33376 5312
rect 33060 5222 33272 5250
rect 33060 5166 33088 5222
rect 33048 5160 33100 5166
rect 33048 5102 33100 5108
rect 33140 5160 33192 5166
rect 33140 5102 33192 5108
rect 32864 4752 32916 4758
rect 32864 4694 32916 4700
rect 33152 4622 33180 5102
rect 33140 4616 33192 4622
rect 33140 4558 33192 4564
rect 32772 4004 32824 4010
rect 32772 3946 32824 3952
rect 32784 3738 32812 3946
rect 32772 3732 32824 3738
rect 32772 3674 32824 3680
rect 33152 3670 33180 4558
rect 33244 4434 33272 5222
rect 33428 5030 33456 8298
rect 33612 7954 33640 8350
rect 33980 7970 34008 8366
rect 33600 7948 33652 7954
rect 33600 7890 33652 7896
rect 33704 7942 34008 7970
rect 33704 7886 33732 7942
rect 33692 7880 33744 7886
rect 33520 7828 33692 7834
rect 33520 7822 33744 7828
rect 33856 7880 33908 7886
rect 33908 7828 33916 7868
rect 33856 7822 33916 7828
rect 33520 7806 33732 7822
rect 33520 7206 33548 7806
rect 33508 7200 33560 7206
rect 33508 7142 33560 7148
rect 33520 6798 33548 7142
rect 33508 6792 33560 6798
rect 33508 6734 33560 6740
rect 33888 6186 33916 7822
rect 34060 7336 34112 7342
rect 34060 7278 34112 7284
rect 34072 6934 34100 7278
rect 34060 6928 34112 6934
rect 34060 6870 34112 6876
rect 33876 6180 33928 6186
rect 33876 6122 33928 6128
rect 34164 5166 34192 8434
rect 34336 8288 34388 8294
rect 34336 8230 34388 8236
rect 34348 8022 34376 8230
rect 34336 8016 34388 8022
rect 34336 7958 34388 7964
rect 34532 7954 34560 12406
rect 34612 10668 34664 10674
rect 34612 10610 34664 10616
rect 34624 8362 34652 10610
rect 34612 8356 34664 8362
rect 34612 8298 34664 8304
rect 34520 7948 34572 7954
rect 34520 7890 34572 7896
rect 34612 7948 34664 7954
rect 34612 7890 34664 7896
rect 34624 7562 34652 7890
rect 34440 7534 34652 7562
rect 34242 7440 34298 7449
rect 34440 7410 34468 7534
rect 34242 7375 34298 7384
rect 34428 7404 34480 7410
rect 34256 7342 34284 7375
rect 34428 7346 34480 7352
rect 34520 7404 34572 7410
rect 34520 7346 34572 7352
rect 34244 7336 34296 7342
rect 34244 7278 34296 7284
rect 34152 5160 34204 5166
rect 34152 5102 34204 5108
rect 33416 5024 33468 5030
rect 33416 4966 33468 4972
rect 33508 5024 33560 5030
rect 33508 4966 33560 4972
rect 33520 4842 33548 4966
rect 33336 4814 33548 4842
rect 33336 4729 33364 4814
rect 33322 4720 33378 4729
rect 33322 4655 33378 4664
rect 33508 4684 33560 4690
rect 33336 4622 33364 4655
rect 33508 4626 33560 4632
rect 33324 4616 33376 4622
rect 33324 4558 33376 4564
rect 33520 4434 33548 4626
rect 33244 4406 33548 4434
rect 33244 3754 33272 4406
rect 33244 3726 33364 3754
rect 33140 3664 33192 3670
rect 33046 3632 33102 3641
rect 32588 3596 32640 3602
rect 33140 3606 33192 3612
rect 33046 3567 33102 3576
rect 33232 3596 33284 3602
rect 32588 3538 32640 3544
rect 33060 3466 33088 3567
rect 33232 3538 33284 3544
rect 33048 3460 33100 3466
rect 33048 3402 33100 3408
rect 32128 3392 32180 3398
rect 32128 3334 32180 3340
rect 32036 3052 32088 3058
rect 32036 2994 32088 3000
rect 31760 2984 31812 2990
rect 31760 2926 31812 2932
rect 33244 2854 33272 3538
rect 33336 3482 33364 3726
rect 34256 3670 34284 7278
rect 34336 7200 34388 7206
rect 34336 7142 34388 7148
rect 34348 6798 34376 7142
rect 34336 6792 34388 6798
rect 34336 6734 34388 6740
rect 34532 6662 34560 7346
rect 34624 7002 34652 7534
rect 34612 6996 34664 7002
rect 34612 6938 34664 6944
rect 34520 6656 34572 6662
rect 34520 6598 34572 6604
rect 34624 5166 34652 6938
rect 34612 5160 34664 5166
rect 34612 5102 34664 5108
rect 34244 3664 34296 3670
rect 33874 3632 33930 3641
rect 34244 3606 34296 3612
rect 33874 3567 33876 3576
rect 33928 3567 33930 3576
rect 33876 3538 33928 3544
rect 34716 3534 34744 17054
rect 34808 9625 34836 24126
rect 35254 23896 35310 23905
rect 35360 23866 35388 25230
rect 35440 25152 35492 25158
rect 35440 25094 35492 25100
rect 35452 24206 35480 25094
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 35440 24200 35492 24206
rect 35440 24142 35492 24148
rect 35440 24064 35492 24070
rect 35440 24006 35492 24012
rect 35452 23866 35480 24006
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 35254 23831 35256 23840
rect 35308 23831 35310 23840
rect 35348 23860 35400 23866
rect 35256 23802 35308 23808
rect 35348 23802 35400 23808
rect 35440 23860 35492 23866
rect 35440 23802 35492 23808
rect 35348 23588 35400 23594
rect 35348 23530 35400 23536
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35360 22250 35388 23530
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 35268 22222 35388 22250
rect 35716 22228 35768 22234
rect 35072 22160 35124 22166
rect 35072 22102 35124 22108
rect 34978 21992 35034 22001
rect 34978 21927 35034 21936
rect 34992 21486 35020 21927
rect 34980 21480 35032 21486
rect 34980 21422 35032 21428
rect 35084 21434 35112 22102
rect 35268 22098 35296 22222
rect 35716 22170 35768 22176
rect 35256 22092 35308 22098
rect 35256 22034 35308 22040
rect 35348 22092 35400 22098
rect 35348 22034 35400 22040
rect 35164 22024 35216 22030
rect 35216 21972 35296 21978
rect 35164 21966 35296 21972
rect 35176 21950 35296 21966
rect 35268 21690 35296 21950
rect 35256 21684 35308 21690
rect 35256 21626 35308 21632
rect 35360 21554 35388 22034
rect 35728 22030 35756 22170
rect 35440 22024 35492 22030
rect 35440 21966 35492 21972
rect 35716 22024 35768 22030
rect 35716 21966 35768 21972
rect 35452 21672 35480 21966
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 35452 21644 35572 21672
rect 35348 21548 35400 21554
rect 35348 21490 35400 21496
rect 35084 21406 35480 21434
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35256 21140 35308 21146
rect 35256 21082 35308 21088
rect 35268 20244 35296 21082
rect 35268 20216 35388 20244
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34888 19304 34940 19310
rect 34886 19272 34888 19281
rect 34940 19272 34942 19281
rect 34886 19207 34942 19216
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18850 35388 20216
rect 35268 18822 35388 18850
rect 35268 18426 35296 18822
rect 35256 18420 35308 18426
rect 35256 18362 35308 18368
rect 35452 18222 35480 21406
rect 35544 21146 35572 21644
rect 35532 21140 35584 21146
rect 35532 21082 35584 21088
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 36004 19514 36032 29038
rect 36096 27470 36124 30670
rect 36084 27464 36136 27470
rect 36084 27406 36136 27412
rect 36188 27282 36216 30790
rect 36280 28665 36308 31726
rect 36556 31346 36584 32166
rect 36360 31340 36412 31346
rect 36360 31282 36412 31288
rect 36544 31340 36596 31346
rect 36544 31282 36596 31288
rect 36372 30802 36400 31282
rect 36544 31136 36596 31142
rect 36542 31104 36544 31113
rect 36596 31104 36598 31113
rect 36542 31039 36598 31048
rect 36360 30796 36412 30802
rect 36360 30738 36412 30744
rect 36452 30728 36504 30734
rect 36450 30696 36452 30705
rect 36504 30696 36506 30705
rect 36360 30660 36412 30666
rect 36450 30631 36506 30640
rect 36360 30602 36412 30608
rect 36372 30122 36400 30602
rect 36452 30592 36504 30598
rect 36452 30534 36504 30540
rect 36464 30258 36492 30534
rect 36452 30252 36504 30258
rect 36452 30194 36504 30200
rect 36360 30116 36412 30122
rect 36360 30058 36412 30064
rect 36452 30048 36504 30054
rect 36452 29990 36504 29996
rect 36360 29164 36412 29170
rect 36464 29152 36492 29990
rect 36648 29578 36676 34954
rect 36832 32978 36860 35770
rect 37108 34746 37136 40326
rect 37200 39846 37228 40462
rect 37292 40089 37320 41074
rect 37844 40662 37872 43658
rect 38120 43654 38148 45222
rect 38292 44736 38344 44742
rect 38292 44678 38344 44684
rect 38304 44402 38332 44678
rect 38396 44538 38424 47670
rect 38672 47666 38700 49624
rect 41340 47818 41368 49694
rect 43166 49694 43300 49722
rect 43166 49624 43222 49694
rect 41340 47802 41460 47818
rect 41340 47796 41472 47802
rect 41340 47790 41420 47796
rect 41420 47738 41472 47744
rect 43272 47666 43300 49694
rect 45742 49694 45876 49722
rect 45742 49624 45798 49694
rect 45848 47666 45876 49694
rect 47674 49624 47730 50424
rect 45926 47696 45982 47705
rect 38660 47660 38712 47666
rect 38660 47602 38712 47608
rect 43260 47660 43312 47666
rect 43260 47602 43312 47608
rect 45836 47660 45888 47666
rect 45926 47631 45928 47640
rect 45836 47602 45888 47608
rect 45980 47631 45982 47640
rect 45928 47602 45980 47608
rect 42892 47592 42944 47598
rect 42892 47534 42944 47540
rect 46204 47592 46256 47598
rect 46204 47534 46256 47540
rect 38844 47456 38896 47462
rect 38844 47398 38896 47404
rect 38856 44878 38884 47398
rect 38844 44872 38896 44878
rect 38844 44814 38896 44820
rect 38384 44532 38436 44538
rect 38384 44474 38436 44480
rect 38292 44396 38344 44402
rect 38292 44338 38344 44344
rect 38396 44334 38424 44474
rect 38844 44464 38896 44470
rect 38844 44406 38896 44412
rect 38476 44396 38528 44402
rect 38476 44338 38528 44344
rect 38384 44328 38436 44334
rect 38384 44270 38436 44276
rect 38108 43648 38160 43654
rect 38108 43590 38160 43596
rect 37832 40656 37884 40662
rect 37832 40598 37884 40604
rect 38016 40520 38068 40526
rect 38016 40462 38068 40468
rect 37464 40384 37516 40390
rect 37464 40326 37516 40332
rect 37476 40118 37504 40326
rect 37556 40180 37608 40186
rect 37556 40122 37608 40128
rect 37464 40112 37516 40118
rect 37278 40080 37334 40089
rect 37464 40054 37516 40060
rect 37278 40015 37334 40024
rect 37188 39840 37240 39846
rect 37188 39782 37240 39788
rect 37280 39840 37332 39846
rect 37280 39782 37332 39788
rect 37188 39568 37240 39574
rect 37188 39510 37240 39516
rect 37200 38418 37228 39510
rect 37292 39098 37320 39782
rect 37476 39642 37504 40054
rect 37464 39636 37516 39642
rect 37464 39578 37516 39584
rect 37462 39264 37518 39273
rect 37462 39199 37518 39208
rect 37280 39092 37332 39098
rect 37280 39034 37332 39040
rect 37292 38418 37320 39034
rect 37476 38962 37504 39199
rect 37464 38956 37516 38962
rect 37464 38898 37516 38904
rect 37464 38752 37516 38758
rect 37464 38694 37516 38700
rect 37188 38412 37240 38418
rect 37188 38354 37240 38360
rect 37280 38412 37332 38418
rect 37280 38354 37332 38360
rect 37372 38412 37424 38418
rect 37372 38354 37424 38360
rect 37200 37194 37228 38354
rect 37292 37942 37320 38354
rect 37280 37936 37332 37942
rect 37280 37878 37332 37884
rect 37384 37262 37412 38354
rect 37476 38010 37504 38694
rect 37464 38004 37516 38010
rect 37464 37946 37516 37952
rect 37372 37256 37424 37262
rect 37372 37198 37424 37204
rect 37188 37188 37240 37194
rect 37188 37130 37240 37136
rect 37384 36258 37412 37198
rect 37384 36230 37504 36258
rect 37372 36168 37424 36174
rect 37372 36110 37424 36116
rect 37384 35290 37412 36110
rect 37372 35284 37424 35290
rect 37372 35226 37424 35232
rect 37096 34740 37148 34746
rect 37096 34682 37148 34688
rect 37004 33312 37056 33318
rect 37004 33254 37056 33260
rect 36820 32972 36872 32978
rect 36820 32914 36872 32920
rect 36832 32298 36860 32914
rect 36820 32292 36872 32298
rect 36820 32234 36872 32240
rect 37016 31754 37044 33254
rect 37108 32910 37136 34682
rect 37188 33856 37240 33862
rect 37188 33798 37240 33804
rect 37200 33590 37228 33798
rect 37188 33584 37240 33590
rect 37188 33526 37240 33532
rect 37188 33448 37240 33454
rect 37188 33390 37240 33396
rect 37096 32904 37148 32910
rect 37096 32846 37148 32852
rect 37108 32366 37136 32846
rect 37096 32360 37148 32366
rect 37096 32302 37148 32308
rect 37016 31726 37136 31754
rect 36728 31136 36780 31142
rect 36728 31078 36780 31084
rect 36912 31136 36964 31142
rect 36912 31078 36964 31084
rect 36636 29572 36688 29578
rect 36636 29514 36688 29520
rect 36544 29504 36596 29510
rect 36544 29446 36596 29452
rect 36412 29124 36492 29152
rect 36360 29106 36412 29112
rect 36266 28656 36322 28665
rect 36266 28591 36322 28600
rect 36096 27254 36216 27282
rect 36096 25770 36124 27254
rect 36360 26988 36412 26994
rect 36360 26930 36412 26936
rect 36372 26518 36400 26930
rect 36360 26512 36412 26518
rect 36360 26454 36412 26460
rect 36358 25936 36414 25945
rect 36358 25871 36414 25880
rect 36084 25764 36136 25770
rect 36084 25706 36136 25712
rect 36096 24834 36124 25706
rect 36176 25696 36228 25702
rect 36176 25638 36228 25644
rect 36188 24954 36216 25638
rect 36268 25356 36320 25362
rect 36268 25298 36320 25304
rect 36280 24954 36308 25298
rect 36176 24948 36228 24954
rect 36176 24890 36228 24896
rect 36268 24948 36320 24954
rect 36268 24890 36320 24896
rect 36096 24806 36308 24834
rect 36372 24818 36400 25871
rect 36176 24744 36228 24750
rect 36176 24686 36228 24692
rect 36084 24064 36136 24070
rect 36084 24006 36136 24012
rect 36096 23730 36124 24006
rect 36084 23724 36136 23730
rect 36084 23666 36136 23672
rect 36084 21888 36136 21894
rect 36084 21830 36136 21836
rect 36096 21622 36124 21830
rect 36084 21616 36136 21622
rect 36084 21558 36136 21564
rect 35992 19508 36044 19514
rect 35992 19450 36044 19456
rect 35992 19372 36044 19378
rect 35992 19314 36044 19320
rect 35716 19168 35768 19174
rect 35716 19110 35768 19116
rect 35728 18766 35756 19110
rect 35716 18760 35768 18766
rect 35716 18702 35768 18708
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 36004 18426 36032 19314
rect 36188 18737 36216 24686
rect 36280 22642 36308 24806
rect 36360 24812 36412 24818
rect 36360 24754 36412 24760
rect 36464 24274 36492 29124
rect 36556 25906 36584 29446
rect 36648 27674 36676 29514
rect 36740 29170 36768 31078
rect 36924 30054 36952 31078
rect 37004 30252 37056 30258
rect 37004 30194 37056 30200
rect 36912 30048 36964 30054
rect 36912 29990 36964 29996
rect 36818 29336 36874 29345
rect 36818 29271 36874 29280
rect 36832 29238 36860 29271
rect 36820 29232 36872 29238
rect 36820 29174 36872 29180
rect 36728 29164 36780 29170
rect 36728 29106 36780 29112
rect 37016 28490 37044 30194
rect 37108 29646 37136 31726
rect 37096 29640 37148 29646
rect 37096 29582 37148 29588
rect 37004 28484 37056 28490
rect 37004 28426 37056 28432
rect 36636 27668 36688 27674
rect 36636 27610 36688 27616
rect 36912 27396 36964 27402
rect 36912 27338 36964 27344
rect 36636 27328 36688 27334
rect 36636 27270 36688 27276
rect 36648 27130 36676 27270
rect 36636 27124 36688 27130
rect 36636 27066 36688 27072
rect 36924 27062 36952 27338
rect 36912 27056 36964 27062
rect 36912 26998 36964 27004
rect 37016 25906 37044 28426
rect 37096 27600 37148 27606
rect 37096 27542 37148 27548
rect 37108 27470 37136 27542
rect 37096 27464 37148 27470
rect 37096 27406 37148 27412
rect 37096 26784 37148 26790
rect 37096 26726 37148 26732
rect 37108 26314 37136 26726
rect 37096 26308 37148 26314
rect 37096 26250 37148 26256
rect 36544 25900 36596 25906
rect 36544 25842 36596 25848
rect 37004 25900 37056 25906
rect 37004 25842 37056 25848
rect 36544 25288 36596 25294
rect 37096 25288 37148 25294
rect 36544 25230 36596 25236
rect 37002 25256 37058 25265
rect 36452 24268 36504 24274
rect 36452 24210 36504 24216
rect 36360 24132 36412 24138
rect 36360 24074 36412 24080
rect 36372 23662 36400 24074
rect 36556 23730 36584 25230
rect 37096 25230 37148 25236
rect 37002 25191 37058 25200
rect 36912 24948 36964 24954
rect 36912 24890 36964 24896
rect 36820 24404 36872 24410
rect 36820 24346 36872 24352
rect 36728 24268 36780 24274
rect 36728 24210 36780 24216
rect 36636 24132 36688 24138
rect 36636 24074 36688 24080
rect 36544 23724 36596 23730
rect 36464 23684 36544 23712
rect 36360 23656 36412 23662
rect 36360 23598 36412 23604
rect 36268 22636 36320 22642
rect 36268 22578 36320 22584
rect 36268 22160 36320 22166
rect 36268 22102 36320 22108
rect 36174 18728 36230 18737
rect 36174 18663 36230 18672
rect 36084 18624 36136 18630
rect 36084 18566 36136 18572
rect 35532 18420 35584 18426
rect 35532 18362 35584 18368
rect 35992 18420 36044 18426
rect 35992 18362 36044 18368
rect 35440 18216 35492 18222
rect 35440 18158 35492 18164
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35544 17746 35572 18362
rect 36096 18358 36124 18566
rect 36188 18426 36216 18663
rect 36176 18420 36228 18426
rect 36176 18362 36228 18368
rect 36084 18352 36136 18358
rect 36084 18294 36136 18300
rect 36280 18222 36308 22102
rect 36372 22098 36400 23598
rect 36360 22092 36412 22098
rect 36360 22034 36412 22040
rect 36360 21888 36412 21894
rect 36360 21830 36412 21836
rect 36372 21554 36400 21830
rect 36360 21548 36412 21554
rect 36360 21490 36412 21496
rect 36464 21486 36492 23684
rect 36544 23666 36596 23672
rect 36544 23588 36596 23594
rect 36544 23530 36596 23536
rect 36452 21480 36504 21486
rect 36452 21422 36504 21428
rect 36360 19508 36412 19514
rect 36360 19450 36412 19456
rect 36176 18216 36228 18222
rect 36176 18158 36228 18164
rect 36268 18216 36320 18222
rect 36268 18158 36320 18164
rect 35532 17740 35584 17746
rect 35532 17682 35584 17688
rect 34980 17672 35032 17678
rect 34980 17614 35032 17620
rect 34992 16998 35020 17614
rect 35348 17604 35400 17610
rect 35348 17546 35400 17552
rect 35164 17536 35216 17542
rect 35164 17478 35216 17484
rect 35176 17134 35204 17478
rect 35164 17128 35216 17134
rect 35164 17070 35216 17076
rect 34980 16992 35032 16998
rect 34980 16934 35032 16940
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35360 16250 35388 17546
rect 35992 17536 36044 17542
rect 35992 17478 36044 17484
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 35532 16992 35584 16998
rect 35532 16934 35584 16940
rect 35544 16590 35572 16934
rect 35532 16584 35584 16590
rect 35532 16526 35584 16532
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 35348 16244 35400 16250
rect 35348 16186 35400 16192
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 36004 15502 36032 17478
rect 36084 17196 36136 17202
rect 36084 17138 36136 17144
rect 36096 15910 36124 17138
rect 36084 15904 36136 15910
rect 36084 15846 36136 15852
rect 35992 15496 36044 15502
rect 35992 15438 36044 15444
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 35348 15020 35400 15026
rect 35348 14962 35400 14968
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35256 14340 35308 14346
rect 35256 14282 35308 14288
rect 35268 14074 35296 14282
rect 35256 14068 35308 14074
rect 35256 14010 35308 14016
rect 35360 13734 35388 14962
rect 35900 14952 35952 14958
rect 35900 14894 35952 14900
rect 35912 14414 35940 14894
rect 35900 14408 35952 14414
rect 35952 14356 36032 14362
rect 35900 14350 36032 14356
rect 35912 14334 36032 14350
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 35716 13864 35768 13870
rect 36004 13818 36032 14334
rect 36084 14340 36136 14346
rect 36084 14282 36136 14288
rect 35768 13812 36032 13818
rect 35716 13806 36032 13812
rect 35728 13790 36032 13806
rect 35348 13728 35400 13734
rect 35348 13670 35400 13676
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 36004 12434 36032 13790
rect 36096 12986 36124 14282
rect 36084 12980 36136 12986
rect 36084 12922 36136 12928
rect 36004 12406 36124 12434
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 35900 11620 35952 11626
rect 35900 11562 35952 11568
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35348 11212 35400 11218
rect 35348 11154 35400 11160
rect 35360 10674 35388 11154
rect 35912 11150 35940 11562
rect 35900 11144 35952 11150
rect 35900 11086 35952 11092
rect 35990 11112 36046 11121
rect 35990 11047 36046 11056
rect 35440 11008 35492 11014
rect 35440 10950 35492 10956
rect 35348 10668 35400 10674
rect 35348 10610 35400 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35256 9716 35308 9722
rect 35256 9658 35308 9664
rect 34794 9616 34850 9625
rect 34794 9551 34850 9560
rect 34796 9444 34848 9450
rect 34796 9386 34848 9392
rect 34808 8634 34836 9386
rect 35268 9330 35296 9658
rect 35360 9518 35388 10610
rect 35452 10062 35480 10950
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 36004 10674 36032 11047
rect 35992 10668 36044 10674
rect 35992 10610 36044 10616
rect 35440 10056 35492 10062
rect 35440 9998 35492 10004
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 35992 9648 36044 9654
rect 35992 9590 36044 9596
rect 35348 9512 35400 9518
rect 35348 9454 35400 9460
rect 35808 9512 35860 9518
rect 35808 9454 35860 9460
rect 35268 9302 35480 9330
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 8628 34848 8634
rect 34796 8570 34848 8576
rect 35348 8356 35400 8362
rect 35348 8298 35400 8304
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35360 8106 35388 8298
rect 35268 8078 35388 8106
rect 35268 7954 35296 8078
rect 35256 7948 35308 7954
rect 35256 7890 35308 7896
rect 35164 7880 35216 7886
rect 35164 7822 35216 7828
rect 35176 7546 35204 7822
rect 35164 7540 35216 7546
rect 35164 7482 35216 7488
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35348 5704 35400 5710
rect 35348 5646 35400 5652
rect 35072 5568 35124 5574
rect 35072 5510 35124 5516
rect 35084 5302 35112 5510
rect 35072 5296 35124 5302
rect 35072 5238 35124 5244
rect 34796 5160 34848 5166
rect 34796 5102 34848 5108
rect 34808 4146 34836 5102
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35360 4826 35388 5646
rect 35452 5234 35480 9302
rect 35820 8838 35848 9454
rect 35808 8832 35860 8838
rect 35808 8774 35860 8780
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 35440 5228 35492 5234
rect 35440 5170 35492 5176
rect 35440 5024 35492 5030
rect 35440 4966 35492 4972
rect 35348 4820 35400 4826
rect 35348 4762 35400 4768
rect 35452 4622 35480 4966
rect 36004 4622 36032 9590
rect 36096 8566 36124 12406
rect 36188 9722 36216 18158
rect 36280 15706 36308 18158
rect 36268 15700 36320 15706
rect 36268 15642 36320 15648
rect 36268 13932 36320 13938
rect 36268 13874 36320 13880
rect 36280 13530 36308 13874
rect 36372 13530 36400 19450
rect 36556 15502 36584 23530
rect 36648 23322 36676 24074
rect 36636 23316 36688 23322
rect 36636 23258 36688 23264
rect 36636 21888 36688 21894
rect 36636 21830 36688 21836
rect 36648 21350 36676 21830
rect 36636 21344 36688 21350
rect 36636 21286 36688 21292
rect 36648 20806 36676 21286
rect 36636 20800 36688 20806
rect 36636 20742 36688 20748
rect 36636 18692 36688 18698
rect 36636 18634 36688 18640
rect 36648 18426 36676 18634
rect 36636 18420 36688 18426
rect 36636 18362 36688 18368
rect 36544 15496 36596 15502
rect 36544 15438 36596 15444
rect 36268 13524 36320 13530
rect 36268 13466 36320 13472
rect 36360 13524 36412 13530
rect 36360 13466 36412 13472
rect 36556 12434 36584 15438
rect 36636 13184 36688 13190
rect 36636 13126 36688 13132
rect 36648 12646 36676 13126
rect 36636 12640 36688 12646
rect 36636 12582 36688 12588
rect 36556 12406 36676 12434
rect 36452 12368 36504 12374
rect 36452 12310 36504 12316
rect 36176 9716 36228 9722
rect 36176 9658 36228 9664
rect 36464 9654 36492 12310
rect 36544 12232 36596 12238
rect 36544 12174 36596 12180
rect 36452 9648 36504 9654
rect 36452 9590 36504 9596
rect 36556 8974 36584 12174
rect 36452 8968 36504 8974
rect 36452 8910 36504 8916
rect 36544 8968 36596 8974
rect 36544 8910 36596 8916
rect 36084 8560 36136 8566
rect 36084 8502 36136 8508
rect 36268 8084 36320 8090
rect 36268 8026 36320 8032
rect 36280 7478 36308 8026
rect 36268 7472 36320 7478
rect 36268 7414 36320 7420
rect 36084 4684 36136 4690
rect 36084 4626 36136 4632
rect 35440 4616 35492 4622
rect 35440 4558 35492 4564
rect 35992 4616 36044 4622
rect 35992 4558 36044 4564
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 36096 4282 36124 4626
rect 36084 4276 36136 4282
rect 36084 4218 36136 4224
rect 34796 4140 34848 4146
rect 34796 4082 34848 4088
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35256 3596 35308 3602
rect 35256 3538 35308 3544
rect 33508 3528 33560 3534
rect 33336 3476 33508 3482
rect 33336 3470 33560 3476
rect 34704 3528 34756 3534
rect 35268 3505 35296 3538
rect 34704 3470 34756 3476
rect 35254 3496 35310 3505
rect 33336 3454 33548 3470
rect 33336 3194 33364 3454
rect 35254 3431 35310 3440
rect 34704 3392 34756 3398
rect 34704 3334 34756 3340
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 33324 3188 33376 3194
rect 33324 3130 33376 3136
rect 34612 3188 34664 3194
rect 34612 3130 34664 3136
rect 33416 3052 33468 3058
rect 33416 2994 33468 3000
rect 31668 2848 31720 2854
rect 31668 2790 31720 2796
rect 33232 2848 33284 2854
rect 33232 2790 33284 2796
rect 29368 2440 29420 2446
rect 29368 2382 29420 2388
rect 33428 2310 33456 2994
rect 34624 2378 34652 3130
rect 34716 2446 34744 3334
rect 35176 3194 35204 3334
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 35164 3188 35216 3194
rect 35164 3130 35216 3136
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 36464 2650 36492 8910
rect 36648 7834 36676 12406
rect 36740 12238 36768 24210
rect 36832 24070 36860 24346
rect 36924 24290 36952 24890
rect 37016 24410 37044 25191
rect 37108 24721 37136 25230
rect 37094 24712 37150 24721
rect 37094 24647 37150 24656
rect 37004 24404 37056 24410
rect 37004 24346 37056 24352
rect 36924 24262 37136 24290
rect 36820 24064 36872 24070
rect 36820 24006 36872 24012
rect 36832 23118 36860 24006
rect 36912 23180 36964 23186
rect 36912 23122 36964 23128
rect 36820 23112 36872 23118
rect 36820 23054 36872 23060
rect 36924 22166 36952 23122
rect 36912 22160 36964 22166
rect 36912 22102 36964 22108
rect 36912 22024 36964 22030
rect 36912 21966 36964 21972
rect 36924 21690 36952 21966
rect 36912 21684 36964 21690
rect 36912 21626 36964 21632
rect 36820 21480 36872 21486
rect 36820 21422 36872 21428
rect 36832 18766 36860 21422
rect 36924 21010 36952 21626
rect 36912 21004 36964 21010
rect 36912 20946 36964 20952
rect 36912 20052 36964 20058
rect 36912 19994 36964 20000
rect 36820 18760 36872 18766
rect 36820 18702 36872 18708
rect 36924 15502 36952 19994
rect 37004 15700 37056 15706
rect 37004 15642 37056 15648
rect 36912 15496 36964 15502
rect 36912 15438 36964 15444
rect 36728 12232 36780 12238
rect 36728 12174 36780 12180
rect 36924 11354 36952 15438
rect 37016 13802 37044 15642
rect 37108 15026 37136 24262
rect 37096 15020 37148 15026
rect 37096 14962 37148 14968
rect 37004 13796 37056 13802
rect 37004 13738 37056 13744
rect 37016 13394 37044 13738
rect 37096 13728 37148 13734
rect 37096 13670 37148 13676
rect 37004 13388 37056 13394
rect 37004 13330 37056 13336
rect 37108 13326 37136 13670
rect 37096 13320 37148 13326
rect 37096 13262 37148 13268
rect 36912 11348 36964 11354
rect 36912 11290 36964 11296
rect 36556 7806 36676 7834
rect 36556 7342 36584 7806
rect 36544 7336 36596 7342
rect 36544 7278 36596 7284
rect 36556 4690 36584 7278
rect 36544 4684 36596 4690
rect 36544 4626 36596 4632
rect 36452 2644 36504 2650
rect 36452 2586 36504 2592
rect 34886 2544 34942 2553
rect 37200 2514 37228 33390
rect 37384 33046 37412 35226
rect 37476 34610 37504 36230
rect 37568 34746 37596 40122
rect 37832 39908 37884 39914
rect 37832 39850 37884 39856
rect 37648 39840 37700 39846
rect 37648 39782 37700 39788
rect 37660 39574 37688 39782
rect 37648 39568 37700 39574
rect 37648 39510 37700 39516
rect 37660 38962 37688 39510
rect 37844 39370 37872 39850
rect 37924 39432 37976 39438
rect 37924 39374 37976 39380
rect 37832 39364 37884 39370
rect 37832 39306 37884 39312
rect 37740 39296 37792 39302
rect 37740 39238 37792 39244
rect 37752 39098 37780 39238
rect 37740 39092 37792 39098
rect 37740 39034 37792 39040
rect 37648 38956 37700 38962
rect 37648 38898 37700 38904
rect 37936 37738 37964 39374
rect 38028 38962 38056 40462
rect 38016 38956 38068 38962
rect 38016 38898 38068 38904
rect 38016 38752 38068 38758
rect 38016 38694 38068 38700
rect 38028 38350 38056 38694
rect 38016 38344 38068 38350
rect 38016 38286 38068 38292
rect 38028 37806 38056 38286
rect 38016 37800 38068 37806
rect 38016 37742 38068 37748
rect 37924 37732 37976 37738
rect 37924 37674 37976 37680
rect 37648 37664 37700 37670
rect 37648 37606 37700 37612
rect 37660 36786 37688 37606
rect 38028 36786 38056 37742
rect 37648 36780 37700 36786
rect 37648 36722 37700 36728
rect 38016 36780 38068 36786
rect 38016 36722 38068 36728
rect 37660 36378 37688 36722
rect 37648 36372 37700 36378
rect 37648 36314 37700 36320
rect 37832 34944 37884 34950
rect 37832 34886 37884 34892
rect 37844 34746 37872 34886
rect 37556 34740 37608 34746
rect 37556 34682 37608 34688
rect 37832 34740 37884 34746
rect 37832 34682 37884 34688
rect 38016 34740 38068 34746
rect 38016 34682 38068 34688
rect 37464 34604 37516 34610
rect 37464 34546 37516 34552
rect 37832 34604 37884 34610
rect 37832 34546 37884 34552
rect 37924 34604 37976 34610
rect 37924 34546 37976 34552
rect 37476 33998 37504 34546
rect 37464 33992 37516 33998
rect 37464 33934 37516 33940
rect 37740 33924 37792 33930
rect 37740 33866 37792 33872
rect 37372 33040 37424 33046
rect 37372 32982 37424 32988
rect 37280 32768 37332 32774
rect 37280 32710 37332 32716
rect 37292 31346 37320 32710
rect 37384 32570 37412 32982
rect 37648 32768 37700 32774
rect 37648 32710 37700 32716
rect 37372 32564 37424 32570
rect 37372 32506 37424 32512
rect 37556 32360 37608 32366
rect 37556 32302 37608 32308
rect 37568 32026 37596 32302
rect 37660 32230 37688 32710
rect 37648 32224 37700 32230
rect 37648 32166 37700 32172
rect 37556 32020 37608 32026
rect 37556 31962 37608 31968
rect 37648 31884 37700 31890
rect 37752 31872 37780 33866
rect 37844 32910 37872 34546
rect 37832 32904 37884 32910
rect 37832 32846 37884 32852
rect 37700 31844 37780 31872
rect 37648 31826 37700 31832
rect 37464 31816 37516 31822
rect 37464 31758 37516 31764
rect 37280 31340 37332 31346
rect 37280 31282 37332 31288
rect 37292 30734 37320 31282
rect 37372 31136 37424 31142
rect 37372 31078 37424 31084
rect 37384 30734 37412 31078
rect 37280 30728 37332 30734
rect 37280 30670 37332 30676
rect 37372 30728 37424 30734
rect 37372 30670 37424 30676
rect 37292 30326 37320 30670
rect 37280 30320 37332 30326
rect 37280 30262 37332 30268
rect 37280 30048 37332 30054
rect 37280 29990 37332 29996
rect 37292 29306 37320 29990
rect 37280 29300 37332 29306
rect 37280 29242 37332 29248
rect 37280 29164 37332 29170
rect 37280 29106 37332 29112
rect 37292 29073 37320 29106
rect 37278 29064 37334 29073
rect 37278 28999 37334 29008
rect 37384 26994 37412 30670
rect 37476 30326 37504 31758
rect 37660 31754 37688 31826
rect 37568 31726 37688 31754
rect 37568 31346 37596 31726
rect 37556 31340 37608 31346
rect 37556 31282 37608 31288
rect 37464 30320 37516 30326
rect 37464 30262 37516 30268
rect 37464 29504 37516 29510
rect 37464 29446 37516 29452
rect 37476 27538 37504 29446
rect 37464 27532 37516 27538
rect 37464 27474 37516 27480
rect 37372 26988 37424 26994
rect 37372 26930 37424 26936
rect 37372 26376 37424 26382
rect 37372 26318 37424 26324
rect 37278 25392 37334 25401
rect 37278 25327 37280 25336
rect 37332 25327 37334 25336
rect 37280 25298 37332 25304
rect 37292 24886 37320 25298
rect 37280 24880 37332 24886
rect 37280 24822 37332 24828
rect 37384 23594 37412 26318
rect 37372 23588 37424 23594
rect 37372 23530 37424 23536
rect 37372 22568 37424 22574
rect 37372 22510 37424 22516
rect 37384 22030 37412 22510
rect 37372 22024 37424 22030
rect 37372 21966 37424 21972
rect 37280 20936 37332 20942
rect 37384 20890 37412 21966
rect 37332 20884 37412 20890
rect 37280 20878 37412 20884
rect 37292 20862 37412 20878
rect 37278 17232 37334 17241
rect 37278 17167 37334 17176
rect 37292 16590 37320 17167
rect 37280 16584 37332 16590
rect 37280 16526 37332 16532
rect 37280 16040 37332 16046
rect 37384 15994 37412 20862
rect 37476 20602 37504 27474
rect 37568 22030 37596 31282
rect 37936 31142 37964 34546
rect 38028 32502 38056 34682
rect 38016 32496 38068 32502
rect 38016 32438 38068 32444
rect 37924 31136 37976 31142
rect 37924 31078 37976 31084
rect 37648 30728 37700 30734
rect 37648 30670 37700 30676
rect 37660 30161 37688 30670
rect 37740 30592 37792 30598
rect 37740 30534 37792 30540
rect 37646 30152 37702 30161
rect 37646 30087 37702 30096
rect 37752 29782 37780 30534
rect 38016 30048 38068 30054
rect 38016 29990 38068 29996
rect 37740 29776 37792 29782
rect 37740 29718 37792 29724
rect 37752 29578 37780 29718
rect 37740 29572 37792 29578
rect 37740 29514 37792 29520
rect 37740 29028 37792 29034
rect 37740 28970 37792 28976
rect 37648 28756 37700 28762
rect 37648 28698 37700 28704
rect 37660 27674 37688 28698
rect 37752 28370 37780 28970
rect 37832 28960 37884 28966
rect 37832 28902 37884 28908
rect 37844 28558 37872 28902
rect 37832 28552 37884 28558
rect 37832 28494 37884 28500
rect 37752 28342 37872 28370
rect 37648 27668 37700 27674
rect 37648 27610 37700 27616
rect 37660 26586 37688 27610
rect 37648 26580 37700 26586
rect 37648 26522 37700 26528
rect 37844 24342 37872 28342
rect 37924 25900 37976 25906
rect 37924 25842 37976 25848
rect 37832 24336 37884 24342
rect 37832 24278 37884 24284
rect 37830 23216 37886 23225
rect 37830 23151 37886 23160
rect 37556 22024 37608 22030
rect 37556 21966 37608 21972
rect 37464 20596 37516 20602
rect 37464 20538 37516 20544
rect 37464 20460 37516 20466
rect 37464 20402 37516 20408
rect 37476 17678 37504 20402
rect 37740 19984 37792 19990
rect 37740 19926 37792 19932
rect 37556 19848 37608 19854
rect 37556 19790 37608 19796
rect 37568 19514 37596 19790
rect 37556 19508 37608 19514
rect 37556 19450 37608 19456
rect 37648 18964 37700 18970
rect 37648 18906 37700 18912
rect 37660 18426 37688 18906
rect 37648 18420 37700 18426
rect 37648 18362 37700 18368
rect 37752 18306 37780 19926
rect 37844 19854 37872 23151
rect 37936 20466 37964 25842
rect 38028 22094 38056 29990
rect 38120 29306 38148 43590
rect 38488 42702 38516 44338
rect 38856 43994 38884 44406
rect 39028 44328 39080 44334
rect 39028 44270 39080 44276
rect 38844 43988 38896 43994
rect 38844 43930 38896 43936
rect 38752 43716 38804 43722
rect 38752 43658 38804 43664
rect 38764 43450 38792 43658
rect 38568 43444 38620 43450
rect 38568 43386 38620 43392
rect 38752 43444 38804 43450
rect 38752 43386 38804 43392
rect 38292 42696 38344 42702
rect 38292 42638 38344 42644
rect 38476 42696 38528 42702
rect 38476 42638 38528 42644
rect 38304 39506 38332 42638
rect 38382 41168 38438 41177
rect 38382 41103 38384 41112
rect 38436 41103 38438 41112
rect 38384 41074 38436 41080
rect 38476 40996 38528 41002
rect 38476 40938 38528 40944
rect 38488 40730 38516 40938
rect 38476 40724 38528 40730
rect 38476 40666 38528 40672
rect 38580 40610 38608 43386
rect 38856 43246 38884 43930
rect 38844 43240 38896 43246
rect 38844 43182 38896 43188
rect 38844 42560 38896 42566
rect 38844 42502 38896 42508
rect 38856 41818 38884 42502
rect 38844 41812 38896 41818
rect 38844 41754 38896 41760
rect 38660 41472 38712 41478
rect 38660 41414 38712 41420
rect 38672 41138 38700 41414
rect 38856 41138 38884 41754
rect 38936 41472 38988 41478
rect 38936 41414 38988 41420
rect 38660 41132 38712 41138
rect 38660 41074 38712 41080
rect 38844 41132 38896 41138
rect 38844 41074 38896 41080
rect 38488 40582 38608 40610
rect 38292 39500 38344 39506
rect 38292 39442 38344 39448
rect 38200 39296 38252 39302
rect 38200 39238 38252 39244
rect 38212 38554 38240 39238
rect 38304 39030 38332 39442
rect 38292 39024 38344 39030
rect 38292 38966 38344 38972
rect 38488 38570 38516 40582
rect 38672 40526 38700 41074
rect 38856 40662 38884 41074
rect 38948 41070 38976 41414
rect 38936 41064 38988 41070
rect 38936 41006 38988 41012
rect 38844 40656 38896 40662
rect 38844 40598 38896 40604
rect 38660 40520 38712 40526
rect 38660 40462 38712 40468
rect 38672 40186 38700 40462
rect 38660 40180 38712 40186
rect 38660 40122 38712 40128
rect 38856 40118 38884 40598
rect 38936 40452 38988 40458
rect 38936 40394 38988 40400
rect 38844 40112 38896 40118
rect 38844 40054 38896 40060
rect 38948 39982 38976 40394
rect 38936 39976 38988 39982
rect 38936 39918 38988 39924
rect 38568 38956 38620 38962
rect 38568 38898 38620 38904
rect 38580 38706 38608 38898
rect 38580 38678 38700 38706
rect 38672 38654 38700 38678
rect 38672 38626 38792 38654
rect 38200 38548 38252 38554
rect 38488 38542 38608 38570
rect 38200 38490 38252 38496
rect 38580 37126 38608 38542
rect 38764 37874 38792 38626
rect 38752 37868 38804 37874
rect 38752 37810 38804 37816
rect 38568 37120 38620 37126
rect 38568 37062 38620 37068
rect 38384 34944 38436 34950
rect 38384 34886 38436 34892
rect 38396 34406 38424 34886
rect 38384 34400 38436 34406
rect 38384 34342 38436 34348
rect 38200 32904 38252 32910
rect 38200 32846 38252 32852
rect 38212 29646 38240 32846
rect 38580 32298 38608 37062
rect 38660 36712 38712 36718
rect 38660 36654 38712 36660
rect 38672 36378 38700 36654
rect 38660 36372 38712 36378
rect 38660 36314 38712 36320
rect 38660 33992 38712 33998
rect 38660 33934 38712 33940
rect 38672 33114 38700 33934
rect 38660 33108 38712 33114
rect 38660 33050 38712 33056
rect 38568 32292 38620 32298
rect 38568 32234 38620 32240
rect 38476 32224 38528 32230
rect 38476 32166 38528 32172
rect 38384 30252 38436 30258
rect 38384 30194 38436 30200
rect 38200 29640 38252 29646
rect 38200 29582 38252 29588
rect 38108 29300 38160 29306
rect 38108 29242 38160 29248
rect 38120 29209 38148 29242
rect 38106 29200 38162 29209
rect 38106 29135 38108 29144
rect 38160 29135 38162 29144
rect 38108 29106 38160 29112
rect 38212 27878 38240 29582
rect 38396 29510 38424 30194
rect 38384 29504 38436 29510
rect 38384 29446 38436 29452
rect 38290 29336 38346 29345
rect 38290 29271 38292 29280
rect 38344 29271 38346 29280
rect 38292 29242 38344 29248
rect 38384 28008 38436 28014
rect 38384 27950 38436 27956
rect 38200 27872 38252 27878
rect 38200 27814 38252 27820
rect 38212 27674 38240 27814
rect 38200 27668 38252 27674
rect 38200 27610 38252 27616
rect 38108 26988 38160 26994
rect 38108 26930 38160 26936
rect 38120 23730 38148 26930
rect 38212 26382 38240 27610
rect 38292 27328 38344 27334
rect 38292 27270 38344 27276
rect 38304 26994 38332 27270
rect 38396 27130 38424 27950
rect 38384 27124 38436 27130
rect 38384 27066 38436 27072
rect 38292 26988 38344 26994
rect 38292 26930 38344 26936
rect 38384 26512 38436 26518
rect 38384 26454 38436 26460
rect 38200 26376 38252 26382
rect 38200 26318 38252 26324
rect 38396 25498 38424 26454
rect 38384 25492 38436 25498
rect 38384 25434 38436 25440
rect 38488 25294 38516 32166
rect 38672 29866 38700 33050
rect 38580 29850 38700 29866
rect 38568 29844 38700 29850
rect 38620 29838 38700 29844
rect 38568 29786 38620 29792
rect 38672 28762 38700 29838
rect 38764 28994 38792 37810
rect 38844 37120 38896 37126
rect 38844 37062 38896 37068
rect 38856 36922 38884 37062
rect 38844 36916 38896 36922
rect 38844 36858 38896 36864
rect 39040 36378 39068 44270
rect 39212 43648 39264 43654
rect 39212 43590 39264 43596
rect 39856 43648 39908 43654
rect 39856 43590 39908 43596
rect 39224 41070 39252 43590
rect 39868 43382 39896 43590
rect 40408 43444 40460 43450
rect 40408 43386 40460 43392
rect 39856 43376 39908 43382
rect 40420 43353 40448 43386
rect 39856 43318 39908 43324
rect 40406 43344 40462 43353
rect 39580 43308 39632 43314
rect 40406 43279 40462 43288
rect 39580 43250 39632 43256
rect 39592 42906 39620 43250
rect 40420 43110 40448 43279
rect 40408 43104 40460 43110
rect 40408 43046 40460 43052
rect 39580 42900 39632 42906
rect 39580 42842 39632 42848
rect 39396 41540 39448 41546
rect 39396 41482 39448 41488
rect 39408 41206 39436 41482
rect 39396 41200 39448 41206
rect 39396 41142 39448 41148
rect 39212 41064 39264 41070
rect 39212 41006 39264 41012
rect 39224 40526 39252 41006
rect 39212 40520 39264 40526
rect 39212 40462 39264 40468
rect 39408 40390 39436 41142
rect 40132 41064 40184 41070
rect 40132 41006 40184 41012
rect 40144 40594 40172 41006
rect 40132 40588 40184 40594
rect 40132 40530 40184 40536
rect 39396 40384 39448 40390
rect 39396 40326 39448 40332
rect 39580 40384 39632 40390
rect 39580 40326 39632 40332
rect 39856 40384 39908 40390
rect 39856 40326 39908 40332
rect 40408 40384 40460 40390
rect 40408 40326 40460 40332
rect 39408 40186 39436 40326
rect 39396 40180 39448 40186
rect 39396 40122 39448 40128
rect 39408 38554 39436 40122
rect 39592 40089 39620 40326
rect 39578 40080 39634 40089
rect 39868 40050 39896 40326
rect 40420 40118 40448 40326
rect 40408 40112 40460 40118
rect 40408 40054 40460 40060
rect 39578 40015 39634 40024
rect 39856 40044 39908 40050
rect 39856 39986 39908 39992
rect 39580 39976 39632 39982
rect 39580 39918 39632 39924
rect 39396 38548 39448 38554
rect 39396 38490 39448 38496
rect 39592 38010 39620 39918
rect 39868 39914 39896 39986
rect 39856 39908 39908 39914
rect 39856 39850 39908 39856
rect 39868 39642 39896 39850
rect 39856 39636 39908 39642
rect 39856 39578 39908 39584
rect 39580 38004 39632 38010
rect 39580 37946 39632 37952
rect 39212 37120 39264 37126
rect 39212 37062 39264 37068
rect 39224 36854 39252 37062
rect 39212 36848 39264 36854
rect 39212 36790 39264 36796
rect 39028 36372 39080 36378
rect 39028 36314 39080 36320
rect 39040 35086 39068 36314
rect 42904 35894 42932 47534
rect 45652 47456 45704 47462
rect 45652 47398 45704 47404
rect 45664 46510 45692 47398
rect 45652 46504 45704 46510
rect 45652 46446 45704 46452
rect 45836 43308 45888 43314
rect 45836 43250 45888 43256
rect 45560 40520 45612 40526
rect 45560 40462 45612 40468
rect 44180 37868 44232 37874
rect 44180 37810 44232 37816
rect 44192 36922 44220 37810
rect 44180 36916 44232 36922
rect 44180 36858 44232 36864
rect 42904 35866 43300 35894
rect 39854 35728 39910 35737
rect 39854 35663 39910 35672
rect 40040 35692 40092 35698
rect 39764 35624 39816 35630
rect 39764 35566 39816 35572
rect 39776 35086 39804 35566
rect 39028 35080 39080 35086
rect 39028 35022 39080 35028
rect 39764 35080 39816 35086
rect 39764 35022 39816 35028
rect 39580 34740 39632 34746
rect 39580 34682 39632 34688
rect 39304 33516 39356 33522
rect 39304 33458 39356 33464
rect 39212 33312 39264 33318
rect 39212 33254 39264 33260
rect 39028 32836 39080 32842
rect 39028 32778 39080 32784
rect 38936 30116 38988 30122
rect 38936 30058 38988 30064
rect 38844 29504 38896 29510
rect 38844 29446 38896 29452
rect 38856 29306 38884 29446
rect 38844 29300 38896 29306
rect 38844 29242 38896 29248
rect 38844 29164 38896 29170
rect 38948 29152 38976 30058
rect 39040 29510 39068 32778
rect 39120 30796 39172 30802
rect 39120 30738 39172 30744
rect 39132 30258 39160 30738
rect 39120 30252 39172 30258
rect 39120 30194 39172 30200
rect 39120 30116 39172 30122
rect 39120 30058 39172 30064
rect 39028 29504 39080 29510
rect 39028 29446 39080 29452
rect 39132 29322 39160 30058
rect 38896 29124 38976 29152
rect 38844 29106 38896 29112
rect 38764 28966 38884 28994
rect 38660 28756 38712 28762
rect 38660 28698 38712 28704
rect 38752 28076 38804 28082
rect 38752 28018 38804 28024
rect 38568 27872 38620 27878
rect 38568 27814 38620 27820
rect 38660 27872 38712 27878
rect 38660 27814 38712 27820
rect 38580 27402 38608 27814
rect 38672 27674 38700 27814
rect 38660 27668 38712 27674
rect 38660 27610 38712 27616
rect 38568 27396 38620 27402
rect 38568 27338 38620 27344
rect 38764 27130 38792 28018
rect 38752 27124 38804 27130
rect 38752 27066 38804 27072
rect 38568 26920 38620 26926
rect 38568 26862 38620 26868
rect 38580 26450 38608 26862
rect 38752 26784 38804 26790
rect 38752 26726 38804 26732
rect 38568 26444 38620 26450
rect 38568 26386 38620 26392
rect 38476 25288 38528 25294
rect 38476 25230 38528 25236
rect 38580 24818 38608 26386
rect 38764 25378 38792 26726
rect 38856 25430 38884 28966
rect 38672 25350 38792 25378
rect 38844 25424 38896 25430
rect 38844 25366 38896 25372
rect 38568 24812 38620 24818
rect 38568 24754 38620 24760
rect 38568 24336 38620 24342
rect 38568 24278 38620 24284
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 38476 24200 38528 24206
rect 38476 24142 38528 24148
rect 38304 23866 38332 24142
rect 38384 24064 38436 24070
rect 38384 24006 38436 24012
rect 38292 23860 38344 23866
rect 38292 23802 38344 23808
rect 38290 23760 38346 23769
rect 38108 23724 38160 23730
rect 38290 23695 38292 23704
rect 38108 23666 38160 23672
rect 38344 23695 38346 23704
rect 38292 23666 38344 23672
rect 38396 22982 38424 24006
rect 38488 23497 38516 24142
rect 38474 23488 38530 23497
rect 38474 23423 38530 23432
rect 38580 23066 38608 24278
rect 38672 23186 38700 25350
rect 38752 25220 38804 25226
rect 38752 25162 38804 25168
rect 38660 23180 38712 23186
rect 38660 23122 38712 23128
rect 38580 23038 38700 23066
rect 38384 22976 38436 22982
rect 38384 22918 38436 22924
rect 38200 22704 38252 22710
rect 38200 22646 38252 22652
rect 38028 22066 38148 22094
rect 38016 20936 38068 20942
rect 38016 20878 38068 20884
rect 37924 20460 37976 20466
rect 37924 20402 37976 20408
rect 37924 20324 37976 20330
rect 37924 20266 37976 20272
rect 37936 19854 37964 20266
rect 37832 19848 37884 19854
rect 37832 19790 37884 19796
rect 37924 19848 37976 19854
rect 37924 19790 37976 19796
rect 37832 19712 37884 19718
rect 37832 19654 37884 19660
rect 37844 19378 37872 19654
rect 37832 19372 37884 19378
rect 37832 19314 37884 19320
rect 37832 19236 37884 19242
rect 37832 19178 37884 19184
rect 37844 18698 37872 19178
rect 37832 18692 37884 18698
rect 37832 18634 37884 18640
rect 37936 18630 37964 19790
rect 37924 18624 37976 18630
rect 37924 18566 37976 18572
rect 37752 18278 37872 18306
rect 37740 18216 37792 18222
rect 37740 18158 37792 18164
rect 37752 17814 37780 18158
rect 37740 17808 37792 17814
rect 37740 17750 37792 17756
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37332 15988 37412 15994
rect 37280 15982 37412 15988
rect 37292 15966 37412 15982
rect 37280 13728 37332 13734
rect 37280 13670 37332 13676
rect 37292 12850 37320 13670
rect 37280 12844 37332 12850
rect 37280 12786 37332 12792
rect 37384 10266 37412 15966
rect 37476 13190 37504 17614
rect 37556 16108 37608 16114
rect 37556 16050 37608 16056
rect 37568 16017 37596 16050
rect 37554 16008 37610 16017
rect 37554 15943 37610 15952
rect 37648 14612 37700 14618
rect 37648 14554 37700 14560
rect 37660 14074 37688 14554
rect 37740 14476 37792 14482
rect 37740 14418 37792 14424
rect 37648 14068 37700 14074
rect 37648 14010 37700 14016
rect 37556 13320 37608 13326
rect 37556 13262 37608 13268
rect 37464 13184 37516 13190
rect 37464 13126 37516 13132
rect 37476 12102 37504 13126
rect 37464 12096 37516 12102
rect 37464 12038 37516 12044
rect 37372 10260 37424 10266
rect 37372 10202 37424 10208
rect 37372 9920 37424 9926
rect 37372 9862 37424 9868
rect 37384 9042 37412 9862
rect 37372 9036 37424 9042
rect 37372 8978 37424 8984
rect 37568 8922 37596 13262
rect 37752 11257 37780 14418
rect 37844 14278 37872 18278
rect 37936 17678 37964 18566
rect 37924 17672 37976 17678
rect 37924 17614 37976 17620
rect 37936 16522 37964 17614
rect 38028 16998 38056 20878
rect 38120 18766 38148 22066
rect 38108 18760 38160 18766
rect 38108 18702 38160 18708
rect 38108 17604 38160 17610
rect 38108 17546 38160 17552
rect 38016 16992 38068 16998
rect 38016 16934 38068 16940
rect 38120 16697 38148 17546
rect 38106 16688 38162 16697
rect 38016 16652 38068 16658
rect 38106 16623 38162 16632
rect 38016 16594 38068 16600
rect 37924 16516 37976 16522
rect 37924 16458 37976 16464
rect 37832 14272 37884 14278
rect 37832 14214 37884 14220
rect 37844 14074 37872 14214
rect 37832 14068 37884 14074
rect 37832 14010 37884 14016
rect 37832 11824 37884 11830
rect 37832 11766 37884 11772
rect 37738 11248 37794 11257
rect 37738 11183 37794 11192
rect 37752 11150 37780 11183
rect 37740 11144 37792 11150
rect 37740 11086 37792 11092
rect 37844 10674 37872 11766
rect 37936 11234 37964 16458
rect 38028 13258 38056 16594
rect 38108 15632 38160 15638
rect 38108 15574 38160 15580
rect 38120 14346 38148 15574
rect 38212 14618 38240 22646
rect 38476 22636 38528 22642
rect 38476 22578 38528 22584
rect 38488 22234 38516 22578
rect 38476 22228 38528 22234
rect 38476 22170 38528 22176
rect 38672 22094 38700 23038
rect 38764 22778 38792 25162
rect 38948 25158 38976 29124
rect 39040 29294 39160 29322
rect 39040 29034 39068 29294
rect 39120 29164 39172 29170
rect 39120 29106 39172 29112
rect 39028 29028 39080 29034
rect 39028 28970 39080 28976
rect 39040 28490 39068 28970
rect 39028 28484 39080 28490
rect 39028 28426 39080 28432
rect 38844 25152 38896 25158
rect 38844 25094 38896 25100
rect 38936 25152 38988 25158
rect 38936 25094 38988 25100
rect 38856 24886 38884 25094
rect 38844 24880 38896 24886
rect 38844 24822 38896 24828
rect 38856 23322 38884 24822
rect 38844 23316 38896 23322
rect 38844 23258 38896 23264
rect 38752 22772 38804 22778
rect 38752 22714 38804 22720
rect 38750 22672 38806 22681
rect 38750 22607 38752 22616
rect 38804 22607 38806 22616
rect 38752 22578 38804 22584
rect 38752 22432 38804 22438
rect 38752 22374 38804 22380
rect 38764 22234 38792 22374
rect 38948 22273 38976 25094
rect 39040 23338 39068 28426
rect 39132 28218 39160 29106
rect 39120 28212 39172 28218
rect 39120 28154 39172 28160
rect 39224 28150 39252 33254
rect 39316 33114 39344 33458
rect 39304 33108 39356 33114
rect 39304 33050 39356 33056
rect 39396 30592 39448 30598
rect 39396 30534 39448 30540
rect 39408 30258 39436 30534
rect 39304 30252 39356 30258
rect 39304 30194 39356 30200
rect 39396 30252 39448 30258
rect 39396 30194 39448 30200
rect 39316 29782 39344 30194
rect 39488 30184 39540 30190
rect 39488 30126 39540 30132
rect 39304 29776 39356 29782
rect 39304 29718 39356 29724
rect 39316 29238 39344 29718
rect 39500 29306 39528 30126
rect 39488 29300 39540 29306
rect 39488 29242 39540 29248
rect 39304 29232 39356 29238
rect 39304 29174 39356 29180
rect 39212 28144 39264 28150
rect 39212 28086 39264 28092
rect 39224 27606 39252 28086
rect 39120 27600 39172 27606
rect 39120 27542 39172 27548
rect 39212 27600 39264 27606
rect 39212 27542 39264 27548
rect 39132 27470 39160 27542
rect 39120 27464 39172 27470
rect 39316 27418 39344 29174
rect 39120 27406 39172 27412
rect 39132 26790 39160 27406
rect 39224 27390 39344 27418
rect 39396 27396 39448 27402
rect 39120 26784 39172 26790
rect 39120 26726 39172 26732
rect 39120 26240 39172 26246
rect 39120 26182 39172 26188
rect 39132 25294 39160 26182
rect 39120 25288 39172 25294
rect 39120 25230 39172 25236
rect 39224 25106 39252 27390
rect 39396 27338 39448 27344
rect 39408 26994 39436 27338
rect 39396 26988 39448 26994
rect 39316 26948 39396 26976
rect 39316 25226 39344 26948
rect 39396 26930 39448 26936
rect 39304 25220 39356 25226
rect 39304 25162 39356 25168
rect 39132 25078 39252 25106
rect 39132 23508 39160 25078
rect 39212 24812 39264 24818
rect 39212 24754 39264 24760
rect 39224 24721 39252 24754
rect 39316 24732 39344 25162
rect 39592 24818 39620 34682
rect 39776 34610 39804 35022
rect 39868 34610 39896 35663
rect 40040 35634 40092 35640
rect 40052 35601 40080 35634
rect 40038 35592 40094 35601
rect 40038 35527 40094 35536
rect 41236 35488 41288 35494
rect 41236 35430 41288 35436
rect 40130 35184 40186 35193
rect 40130 35119 40186 35128
rect 40144 35086 40172 35119
rect 40132 35080 40184 35086
rect 40132 35022 40184 35028
rect 41248 34610 41276 35430
rect 41420 34944 41472 34950
rect 41420 34886 41472 34892
rect 39764 34604 39816 34610
rect 39764 34546 39816 34552
rect 39856 34604 39908 34610
rect 39856 34546 39908 34552
rect 41236 34604 41288 34610
rect 41236 34546 41288 34552
rect 41052 33992 41104 33998
rect 41052 33934 41104 33940
rect 40316 33856 40368 33862
rect 40316 33798 40368 33804
rect 40328 33522 40356 33798
rect 41064 33658 41092 33934
rect 41144 33924 41196 33930
rect 41144 33866 41196 33872
rect 41052 33652 41104 33658
rect 41052 33594 41104 33600
rect 40316 33516 40368 33522
rect 40316 33458 40368 33464
rect 41156 33318 41184 33866
rect 41328 33516 41380 33522
rect 41328 33458 41380 33464
rect 40040 33312 40092 33318
rect 40040 33254 40092 33260
rect 41144 33312 41196 33318
rect 41144 33254 41196 33260
rect 41236 33312 41288 33318
rect 41236 33254 41288 33260
rect 40052 30734 40080 33254
rect 40500 32836 40552 32842
rect 40500 32778 40552 32784
rect 40776 32836 40828 32842
rect 40776 32778 40828 32784
rect 40512 32434 40540 32778
rect 40500 32428 40552 32434
rect 40500 32370 40552 32376
rect 40224 32360 40276 32366
rect 40224 32302 40276 32308
rect 40236 31822 40264 32302
rect 40224 31816 40276 31822
rect 40224 31758 40276 31764
rect 40236 30802 40264 31758
rect 40408 31136 40460 31142
rect 40408 31078 40460 31084
rect 40224 30796 40276 30802
rect 40224 30738 40276 30744
rect 40420 30734 40448 31078
rect 40512 30938 40540 32370
rect 40788 32366 40816 32778
rect 40776 32360 40828 32366
rect 40776 32302 40828 32308
rect 40592 31816 40644 31822
rect 40592 31758 40644 31764
rect 40500 30932 40552 30938
rect 40500 30874 40552 30880
rect 40040 30728 40092 30734
rect 40040 30670 40092 30676
rect 40316 30728 40368 30734
rect 40316 30670 40368 30676
rect 40408 30728 40460 30734
rect 40408 30670 40460 30676
rect 40328 30258 40356 30670
rect 40408 30592 40460 30598
rect 40408 30534 40460 30540
rect 40040 30252 40092 30258
rect 40316 30252 40368 30258
rect 40040 30194 40092 30200
rect 40236 30212 40316 30240
rect 39672 30184 39724 30190
rect 39672 30126 39724 30132
rect 39684 29850 39712 30126
rect 39948 30048 40000 30054
rect 39948 29990 40000 29996
rect 39960 29850 39988 29990
rect 39672 29844 39724 29850
rect 39672 29786 39724 29792
rect 39948 29844 40000 29850
rect 39948 29786 40000 29792
rect 40052 29782 40080 30194
rect 40040 29776 40092 29782
rect 40040 29718 40092 29724
rect 40052 29102 40080 29718
rect 40236 29646 40264 30212
rect 40420 30240 40448 30534
rect 40500 30252 40552 30258
rect 40420 30212 40500 30240
rect 40316 30194 40368 30200
rect 40500 30194 40552 30200
rect 40224 29640 40276 29646
rect 40224 29582 40276 29588
rect 40132 29504 40184 29510
rect 40132 29446 40184 29452
rect 40144 29238 40172 29446
rect 40132 29232 40184 29238
rect 40132 29174 40184 29180
rect 40040 29096 40092 29102
rect 40040 29038 40092 29044
rect 40144 28200 40172 29174
rect 40052 28172 40172 28200
rect 39948 28076 40000 28082
rect 39948 28018 40000 28024
rect 39764 27940 39816 27946
rect 39764 27882 39816 27888
rect 39776 26994 39804 27882
rect 39960 27713 39988 28018
rect 39946 27704 40002 27713
rect 39946 27639 40002 27648
rect 39948 27396 40000 27402
rect 39948 27338 40000 27344
rect 39960 26994 39988 27338
rect 40052 27334 40080 28172
rect 40236 28082 40264 29582
rect 40512 28150 40540 30194
rect 40500 28144 40552 28150
rect 40500 28086 40552 28092
rect 40132 28076 40184 28082
rect 40132 28018 40184 28024
rect 40224 28076 40276 28082
rect 40276 28036 40356 28064
rect 40224 28018 40276 28024
rect 40040 27328 40092 27334
rect 40040 27270 40092 27276
rect 39764 26988 39816 26994
rect 39948 26988 40000 26994
rect 39816 26948 39896 26976
rect 39764 26930 39816 26936
rect 39672 26240 39724 26246
rect 39672 26182 39724 26188
rect 39684 25906 39712 26182
rect 39672 25900 39724 25906
rect 39672 25842 39724 25848
rect 39580 24812 39632 24818
rect 39580 24754 39632 24760
rect 39396 24744 39448 24750
rect 39210 24712 39266 24721
rect 39210 24647 39266 24656
rect 39316 24704 39396 24732
rect 39212 24608 39264 24614
rect 39212 24550 39264 24556
rect 39224 24052 39252 24550
rect 39316 24206 39344 24704
rect 39396 24686 39448 24692
rect 39488 24608 39540 24614
rect 39488 24550 39540 24556
rect 39304 24200 39356 24206
rect 39304 24142 39356 24148
rect 39224 24024 39436 24052
rect 39408 23594 39436 24024
rect 39500 23730 39528 24550
rect 39488 23724 39540 23730
rect 39488 23666 39540 23672
rect 39396 23588 39448 23594
rect 39396 23530 39448 23536
rect 39304 23520 39356 23526
rect 39132 23480 39304 23508
rect 39304 23462 39356 23468
rect 39040 23310 39252 23338
rect 39028 23180 39080 23186
rect 39028 23122 39080 23128
rect 38934 22264 38990 22273
rect 38752 22228 38804 22234
rect 38934 22199 38990 22208
rect 38752 22170 38804 22176
rect 38672 22066 38976 22094
rect 38752 22024 38804 22030
rect 38752 21966 38804 21972
rect 38568 21888 38620 21894
rect 38568 21830 38620 21836
rect 38580 20942 38608 21830
rect 38764 21622 38792 21966
rect 38844 21956 38896 21962
rect 38844 21898 38896 21904
rect 38856 21690 38884 21898
rect 38844 21684 38896 21690
rect 38844 21626 38896 21632
rect 38752 21616 38804 21622
rect 38752 21558 38804 21564
rect 38568 20936 38620 20942
rect 38568 20878 38620 20884
rect 38384 20596 38436 20602
rect 38384 20538 38436 20544
rect 38396 19378 38424 20538
rect 38660 20392 38712 20398
rect 38660 20334 38712 20340
rect 38568 20052 38620 20058
rect 38568 19994 38620 20000
rect 38384 19372 38436 19378
rect 38304 19332 38384 19360
rect 38304 16674 38332 19332
rect 38384 19314 38436 19320
rect 38580 19310 38608 19994
rect 38568 19304 38620 19310
rect 38568 19246 38620 19252
rect 38672 18970 38700 20334
rect 38764 19854 38792 21558
rect 38844 21480 38896 21486
rect 38844 21422 38896 21428
rect 38856 20330 38884 21422
rect 38844 20324 38896 20330
rect 38844 20266 38896 20272
rect 38752 19848 38804 19854
rect 38752 19790 38804 19796
rect 38752 19508 38804 19514
rect 38752 19450 38804 19456
rect 38764 19378 38792 19450
rect 38752 19372 38804 19378
rect 38752 19314 38804 19320
rect 38660 18964 38712 18970
rect 38660 18906 38712 18912
rect 38764 18902 38792 19314
rect 38752 18896 38804 18902
rect 38658 18864 38714 18873
rect 38752 18838 38804 18844
rect 38658 18799 38714 18808
rect 38672 18766 38700 18799
rect 38384 18760 38436 18766
rect 38384 18702 38436 18708
rect 38660 18760 38712 18766
rect 38660 18702 38712 18708
rect 38396 17270 38424 18702
rect 38672 17678 38700 18702
rect 38660 17672 38712 17678
rect 38660 17614 38712 17620
rect 38844 17672 38896 17678
rect 38844 17614 38896 17620
rect 38856 17338 38884 17614
rect 38844 17332 38896 17338
rect 38844 17274 38896 17280
rect 38384 17264 38436 17270
rect 38384 17206 38436 17212
rect 38844 17196 38896 17202
rect 38948 17184 38976 22066
rect 38896 17156 38976 17184
rect 38844 17138 38896 17144
rect 38936 17060 38988 17066
rect 38936 17002 38988 17008
rect 38476 16992 38528 16998
rect 38476 16934 38528 16940
rect 38304 16646 38424 16674
rect 38292 16584 38344 16590
rect 38292 16526 38344 16532
rect 38304 16250 38332 16526
rect 38292 16244 38344 16250
rect 38292 16186 38344 16192
rect 38200 14612 38252 14618
rect 38200 14554 38252 14560
rect 38108 14340 38160 14346
rect 38108 14282 38160 14288
rect 38016 13252 38068 13258
rect 38016 13194 38068 13200
rect 38120 13138 38148 14282
rect 38396 13326 38424 16646
rect 38488 16590 38516 16934
rect 38476 16584 38528 16590
rect 38476 16526 38528 16532
rect 38844 16584 38896 16590
rect 38844 16526 38896 16532
rect 38856 15978 38884 16526
rect 38948 16454 38976 17002
rect 38936 16448 38988 16454
rect 38936 16390 38988 16396
rect 38948 16182 38976 16390
rect 38936 16176 38988 16182
rect 38936 16118 38988 16124
rect 39040 15978 39068 23122
rect 39120 22636 39172 22642
rect 39120 22578 39172 22584
rect 39132 22409 39160 22578
rect 39118 22400 39174 22409
rect 39118 22335 39174 22344
rect 39118 22264 39174 22273
rect 39118 22199 39174 22208
rect 39132 18698 39160 22199
rect 39224 19174 39252 23310
rect 39212 19168 39264 19174
rect 39212 19110 39264 19116
rect 39120 18692 39172 18698
rect 39120 18634 39172 18640
rect 39132 18290 39160 18634
rect 39120 18284 39172 18290
rect 39120 18226 39172 18232
rect 38844 15972 38896 15978
rect 38844 15914 38896 15920
rect 39028 15972 39080 15978
rect 39028 15914 39080 15920
rect 39224 15570 39252 19110
rect 39212 15564 39264 15570
rect 39212 15506 39264 15512
rect 38476 15020 38528 15026
rect 38476 14962 38528 14968
rect 38488 14482 38516 14962
rect 39224 14890 39252 15506
rect 39316 15026 39344 23462
rect 39408 16114 39436 23530
rect 39500 23225 39528 23666
rect 39486 23216 39542 23225
rect 39486 23151 39542 23160
rect 39488 22092 39540 22098
rect 39488 22034 39540 22040
rect 39500 20641 39528 22034
rect 39592 21350 39620 24754
rect 39764 24064 39816 24070
rect 39764 24006 39816 24012
rect 39776 23730 39804 24006
rect 39764 23724 39816 23730
rect 39764 23666 39816 23672
rect 39868 23610 39896 26948
rect 39948 26930 40000 26936
rect 40040 25152 40092 25158
rect 40040 25094 40092 25100
rect 40052 24206 40080 25094
rect 40144 24682 40172 28018
rect 40328 27470 40356 28036
rect 40316 27464 40368 27470
rect 40316 27406 40368 27412
rect 40328 26858 40356 27406
rect 40316 26852 40368 26858
rect 40316 26794 40368 26800
rect 40316 25696 40368 25702
rect 40316 25638 40368 25644
rect 40328 25294 40356 25638
rect 40316 25288 40368 25294
rect 40316 25230 40368 25236
rect 40132 24676 40184 24682
rect 40132 24618 40184 24624
rect 40040 24200 40092 24206
rect 40604 24154 40632 31758
rect 40960 30592 41012 30598
rect 40960 30534 41012 30540
rect 40868 30048 40920 30054
rect 40696 29996 40868 30002
rect 40696 29990 40920 29996
rect 40696 29974 40908 29990
rect 40696 29850 40724 29974
rect 40684 29844 40736 29850
rect 40684 29786 40736 29792
rect 40972 29714 41000 30534
rect 41052 30116 41104 30122
rect 41052 30058 41104 30064
rect 40960 29708 41012 29714
rect 40960 29650 41012 29656
rect 40972 29594 41000 29650
rect 40880 29578 41000 29594
rect 40868 29572 41000 29578
rect 40920 29566 41000 29572
rect 40868 29514 40920 29520
rect 40960 29504 41012 29510
rect 40960 29446 41012 29452
rect 40972 29170 41000 29446
rect 40960 29164 41012 29170
rect 40960 29106 41012 29112
rect 40776 28756 40828 28762
rect 40776 28698 40828 28704
rect 40788 27402 40816 28698
rect 40960 27872 41012 27878
rect 40960 27814 41012 27820
rect 40776 27396 40828 27402
rect 40776 27338 40828 27344
rect 40684 27328 40736 27334
rect 40684 27270 40736 27276
rect 40696 27062 40724 27270
rect 40684 27056 40736 27062
rect 40684 26998 40736 27004
rect 40684 24812 40736 24818
rect 40788 24800 40816 27338
rect 40972 26518 41000 27814
rect 41064 27402 41092 30058
rect 41156 29782 41184 33254
rect 41248 32434 41276 33254
rect 41236 32428 41288 32434
rect 41236 32370 41288 32376
rect 41340 32298 41368 33458
rect 41328 32292 41380 32298
rect 41328 32234 41380 32240
rect 41236 30184 41288 30190
rect 41236 30126 41288 30132
rect 41144 29776 41196 29782
rect 41144 29718 41196 29724
rect 41156 29646 41184 29718
rect 41144 29640 41196 29646
rect 41144 29582 41196 29588
rect 41144 29504 41196 29510
rect 41144 29446 41196 29452
rect 41156 29170 41184 29446
rect 41248 29238 41276 30126
rect 41328 29300 41380 29306
rect 41328 29242 41380 29248
rect 41236 29232 41288 29238
rect 41236 29174 41288 29180
rect 41144 29164 41196 29170
rect 41144 29106 41196 29112
rect 41156 29073 41184 29106
rect 41142 29064 41198 29073
rect 41142 28999 41198 29008
rect 41248 27826 41276 29174
rect 41340 29102 41368 29242
rect 41328 29096 41380 29102
rect 41328 29038 41380 29044
rect 41340 28014 41368 29038
rect 41432 28966 41460 34886
rect 41788 34604 41840 34610
rect 41788 34546 41840 34552
rect 42156 34604 42208 34610
rect 42156 34546 42208 34552
rect 41696 34400 41748 34406
rect 41696 34342 41748 34348
rect 41604 33924 41656 33930
rect 41604 33866 41656 33872
rect 41616 33402 41644 33866
rect 41708 33862 41736 34342
rect 41800 34134 41828 34546
rect 42168 34474 42196 34546
rect 42156 34468 42208 34474
rect 42156 34410 42208 34416
rect 42708 34468 42760 34474
rect 42708 34410 42760 34416
rect 41972 34400 42024 34406
rect 42168 34377 42196 34410
rect 41972 34342 42024 34348
rect 42154 34368 42210 34377
rect 41788 34128 41840 34134
rect 41788 34070 41840 34076
rect 41984 33930 42012 34342
rect 42154 34303 42210 34312
rect 42248 34128 42300 34134
rect 42248 34070 42300 34076
rect 42064 34060 42116 34066
rect 42064 34002 42116 34008
rect 41972 33924 42024 33930
rect 41972 33866 42024 33872
rect 41696 33856 41748 33862
rect 41696 33798 41748 33804
rect 41708 33522 41736 33798
rect 41972 33652 42024 33658
rect 41972 33594 42024 33600
rect 41696 33516 41748 33522
rect 41696 33458 41748 33464
rect 41880 33448 41932 33454
rect 41616 33374 41736 33402
rect 41880 33390 41932 33396
rect 41708 33318 41736 33374
rect 41696 33312 41748 33318
rect 41696 33254 41748 33260
rect 41604 33040 41656 33046
rect 41604 32982 41656 32988
rect 41616 32609 41644 32982
rect 41708 32892 41736 33254
rect 41892 33114 41920 33390
rect 41880 33108 41932 33114
rect 41880 33050 41932 33056
rect 41984 32978 42012 33594
rect 42076 33522 42104 34002
rect 42064 33516 42116 33522
rect 42064 33458 42116 33464
rect 42154 33008 42210 33017
rect 41972 32972 42024 32978
rect 42154 32943 42210 32952
rect 41972 32914 42024 32920
rect 41788 32904 41840 32910
rect 41708 32864 41788 32892
rect 41788 32846 41840 32852
rect 42064 32904 42116 32910
rect 42064 32846 42116 32852
rect 41696 32768 41748 32774
rect 41694 32736 41696 32745
rect 41748 32736 41750 32745
rect 41694 32671 41750 32680
rect 41602 32600 41658 32609
rect 41602 32535 41658 32544
rect 41512 32224 41564 32230
rect 41512 32166 41564 32172
rect 41604 32224 41656 32230
rect 41604 32166 41656 32172
rect 41524 31890 41552 32166
rect 41512 31884 41564 31890
rect 41512 31826 41564 31832
rect 41524 31482 41552 31826
rect 41512 31476 41564 31482
rect 41512 31418 41564 31424
rect 41616 30258 41644 32166
rect 41800 30258 41828 32846
rect 42076 32570 42104 32846
rect 42064 32564 42116 32570
rect 42064 32506 42116 32512
rect 42168 32434 42196 32943
rect 42260 32910 42288 34070
rect 42432 33856 42484 33862
rect 42432 33798 42484 33804
rect 42524 33856 42576 33862
rect 42524 33798 42576 33804
rect 42444 33590 42472 33798
rect 42432 33584 42484 33590
rect 42432 33526 42484 33532
rect 42340 33312 42392 33318
rect 42340 33254 42392 33260
rect 42352 33114 42380 33254
rect 42340 33108 42392 33114
rect 42340 33050 42392 33056
rect 42248 32904 42300 32910
rect 42444 32858 42472 33526
rect 42536 33522 42564 33798
rect 42720 33522 42748 34410
rect 42524 33516 42576 33522
rect 42708 33516 42760 33522
rect 42576 33476 42656 33504
rect 42524 33458 42576 33464
rect 42524 33040 42576 33046
rect 42522 33008 42524 33017
rect 42576 33008 42578 33017
rect 42522 32943 42578 32952
rect 42628 32910 42656 33476
rect 42708 33458 42760 33464
rect 42248 32846 42300 32852
rect 42352 32830 42472 32858
rect 42616 32904 42668 32910
rect 42616 32846 42668 32852
rect 42524 32836 42576 32842
rect 42156 32428 42208 32434
rect 42156 32370 42208 32376
rect 42352 32366 42380 32830
rect 42524 32778 42576 32784
rect 42432 32768 42484 32774
rect 42432 32710 42484 32716
rect 42444 32570 42472 32710
rect 42432 32564 42484 32570
rect 42432 32506 42484 32512
rect 42340 32360 42392 32366
rect 42536 32314 42564 32778
rect 42628 32434 42656 32846
rect 42720 32502 42748 33458
rect 42892 32904 42944 32910
rect 42892 32846 42944 32852
rect 42800 32768 42852 32774
rect 42798 32736 42800 32745
rect 42852 32736 42854 32745
rect 42798 32671 42854 32680
rect 42708 32496 42760 32502
rect 42708 32438 42760 32444
rect 42616 32428 42668 32434
rect 42616 32370 42668 32376
rect 42340 32302 42392 32308
rect 42352 32026 42380 32302
rect 42444 32286 42564 32314
rect 41972 32020 42024 32026
rect 41972 31962 42024 31968
rect 42340 32020 42392 32026
rect 42340 31962 42392 31968
rect 41604 30252 41656 30258
rect 41604 30194 41656 30200
rect 41788 30252 41840 30258
rect 41788 30194 41840 30200
rect 41696 29572 41748 29578
rect 41696 29514 41748 29520
rect 41880 29572 41932 29578
rect 41880 29514 41932 29520
rect 41512 29164 41564 29170
rect 41564 29124 41644 29152
rect 41512 29106 41564 29112
rect 41510 29064 41566 29073
rect 41510 28999 41566 29008
rect 41420 28960 41472 28966
rect 41420 28902 41472 28908
rect 41432 28064 41460 28902
rect 41524 28234 41552 28999
rect 41616 28966 41644 29124
rect 41604 28960 41656 28966
rect 41604 28902 41656 28908
rect 41524 28206 41644 28234
rect 41512 28076 41564 28082
rect 41432 28036 41512 28064
rect 41512 28018 41564 28024
rect 41328 28008 41380 28014
rect 41328 27950 41380 27956
rect 41418 27840 41474 27849
rect 41248 27798 41368 27826
rect 41052 27396 41104 27402
rect 41052 27338 41104 27344
rect 41144 27396 41196 27402
rect 41144 27338 41196 27344
rect 41156 27130 41184 27338
rect 41144 27124 41196 27130
rect 41144 27066 41196 27072
rect 41236 26784 41288 26790
rect 41236 26726 41288 26732
rect 40960 26512 41012 26518
rect 40960 26454 41012 26460
rect 41144 25968 41196 25974
rect 41144 25910 41196 25916
rect 40868 25152 40920 25158
rect 40868 25094 40920 25100
rect 40880 24818 40908 25094
rect 41156 24954 41184 25910
rect 41144 24948 41196 24954
rect 41144 24890 41196 24896
rect 40736 24772 40816 24800
rect 40868 24812 40920 24818
rect 40684 24754 40736 24760
rect 40868 24754 40920 24760
rect 40040 24142 40092 24148
rect 40512 24126 40632 24154
rect 40512 23730 40540 24126
rect 40592 24064 40644 24070
rect 40592 24006 40644 24012
rect 40604 23730 40632 24006
rect 39948 23724 40000 23730
rect 39948 23666 40000 23672
rect 40500 23724 40552 23730
rect 40500 23666 40552 23672
rect 40592 23724 40644 23730
rect 40592 23666 40644 23672
rect 39776 23594 39896 23610
rect 39764 23588 39896 23594
rect 39816 23582 39896 23588
rect 39764 23530 39816 23536
rect 39672 23112 39724 23118
rect 39672 23054 39724 23060
rect 39684 22778 39712 23054
rect 39672 22772 39724 22778
rect 39672 22714 39724 22720
rect 39580 21344 39632 21350
rect 39580 21286 39632 21292
rect 39684 21146 39712 22714
rect 39776 21554 39804 23530
rect 39960 23526 39988 23666
rect 39948 23520 40000 23526
rect 39948 23462 40000 23468
rect 39856 22500 39908 22506
rect 39856 22442 39908 22448
rect 39868 22166 39896 22442
rect 39856 22160 39908 22166
rect 39856 22102 39908 22108
rect 39764 21548 39816 21554
rect 39764 21490 39816 21496
rect 39672 21140 39724 21146
rect 39672 21082 39724 21088
rect 39486 20632 39542 20641
rect 39486 20567 39542 20576
rect 39396 16108 39448 16114
rect 39396 16050 39448 16056
rect 39408 15026 39436 16050
rect 39776 15434 39804 21490
rect 39868 19334 39896 22102
rect 40512 22094 40540 23666
rect 40420 22066 40540 22094
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 39948 21888 40000 21894
rect 39948 21830 40000 21836
rect 39960 21622 39988 21830
rect 39948 21616 40000 21622
rect 39948 21558 40000 21564
rect 40052 20262 40080 21966
rect 40316 21684 40368 21690
rect 40316 21626 40368 21632
rect 40130 21448 40186 21457
rect 40130 21383 40186 21392
rect 40144 20942 40172 21383
rect 40132 20936 40184 20942
rect 40132 20878 40184 20884
rect 40224 20392 40276 20398
rect 40224 20334 40276 20340
rect 40040 20256 40092 20262
rect 40040 20198 40092 20204
rect 39868 19306 39988 19334
rect 39960 17678 39988 19306
rect 40040 18760 40092 18766
rect 40040 18702 40092 18708
rect 40052 18426 40080 18702
rect 40040 18420 40092 18426
rect 40040 18362 40092 18368
rect 40132 18284 40184 18290
rect 40132 18226 40184 18232
rect 39948 17672 40000 17678
rect 39948 17614 40000 17620
rect 39960 17338 39988 17614
rect 39948 17332 40000 17338
rect 39948 17274 40000 17280
rect 39856 17128 39908 17134
rect 39856 17070 39908 17076
rect 39868 16794 39896 17070
rect 39856 16788 39908 16794
rect 39856 16730 39908 16736
rect 39868 15706 39896 16730
rect 39960 16590 39988 17274
rect 40040 17196 40092 17202
rect 40040 17138 40092 17144
rect 39948 16584 40000 16590
rect 39948 16526 40000 16532
rect 40052 16454 40080 17138
rect 40040 16448 40092 16454
rect 40040 16390 40092 16396
rect 39856 15700 39908 15706
rect 39856 15642 39908 15648
rect 39764 15428 39816 15434
rect 39764 15370 39816 15376
rect 39304 15020 39356 15026
rect 39304 14962 39356 14968
rect 39396 15020 39448 15026
rect 39396 14962 39448 14968
rect 39212 14884 39264 14890
rect 39212 14826 39264 14832
rect 38660 14816 38712 14822
rect 38660 14758 38712 14764
rect 39672 14816 39724 14822
rect 39672 14758 39724 14764
rect 38476 14476 38528 14482
rect 38476 14418 38528 14424
rect 38568 14408 38620 14414
rect 38568 14350 38620 14356
rect 38476 14272 38528 14278
rect 38476 14214 38528 14220
rect 38384 13320 38436 13326
rect 38384 13262 38436 13268
rect 38120 13110 38424 13138
rect 38396 12434 38424 13110
rect 38304 12406 38424 12434
rect 38016 12300 38068 12306
rect 38016 12242 38068 12248
rect 38028 11898 38056 12242
rect 38016 11892 38068 11898
rect 38016 11834 38068 11840
rect 38108 11620 38160 11626
rect 38108 11562 38160 11568
rect 37936 11206 38056 11234
rect 37924 11144 37976 11150
rect 37924 11086 37976 11092
rect 37936 10810 37964 11086
rect 37924 10804 37976 10810
rect 37924 10746 37976 10752
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 37844 10198 37872 10610
rect 37832 10192 37884 10198
rect 37832 10134 37884 10140
rect 37740 9444 37792 9450
rect 37740 9386 37792 9392
rect 37752 8974 37780 9386
rect 37384 8906 37596 8922
rect 37740 8968 37792 8974
rect 37740 8910 37792 8916
rect 37372 8900 37596 8906
rect 37424 8894 37596 8900
rect 37372 8842 37424 8848
rect 37568 8566 37596 8894
rect 37924 8900 37976 8906
rect 37924 8842 37976 8848
rect 37936 8634 37964 8842
rect 37924 8628 37976 8634
rect 37924 8570 37976 8576
rect 37556 8560 37608 8566
rect 37556 8502 37608 8508
rect 38028 8498 38056 11206
rect 38120 10674 38148 11562
rect 38108 10668 38160 10674
rect 38108 10610 38160 10616
rect 38120 9382 38148 10610
rect 38304 10470 38332 12406
rect 38488 11762 38516 14214
rect 38580 12209 38608 14350
rect 38566 12200 38622 12209
rect 38566 12135 38622 12144
rect 38476 11756 38528 11762
rect 38476 11698 38528 11704
rect 38568 11552 38620 11558
rect 38568 11494 38620 11500
rect 38580 11286 38608 11494
rect 38568 11280 38620 11286
rect 38382 11248 38438 11257
rect 38568 11222 38620 11228
rect 38382 11183 38438 11192
rect 38396 11150 38424 11183
rect 38384 11144 38436 11150
rect 38384 11086 38436 11092
rect 38384 11008 38436 11014
rect 38384 10950 38436 10956
rect 38396 10674 38424 10950
rect 38384 10668 38436 10674
rect 38384 10610 38436 10616
rect 38672 10606 38700 14758
rect 39684 14618 39712 14758
rect 39672 14612 39724 14618
rect 39672 14554 39724 14560
rect 39212 12844 39264 12850
rect 39212 12786 39264 12792
rect 39580 12844 39632 12850
rect 39580 12786 39632 12792
rect 39224 12442 39252 12786
rect 38752 12436 38804 12442
rect 38752 12378 38804 12384
rect 38844 12436 38896 12442
rect 38844 12378 38896 12384
rect 39212 12436 39264 12442
rect 39592 12434 39620 12786
rect 39212 12378 39264 12384
rect 39500 12406 39620 12434
rect 38764 11801 38792 12378
rect 38856 12238 38884 12378
rect 39500 12374 39528 12406
rect 39488 12368 39540 12374
rect 39488 12310 39540 12316
rect 39776 12238 39804 15370
rect 40144 15094 40172 18226
rect 40236 16998 40264 20334
rect 40328 18358 40356 21626
rect 40420 21350 40448 22066
rect 40408 21344 40460 21350
rect 40408 21286 40460 21292
rect 40696 20874 40724 24754
rect 41248 24750 41276 26726
rect 41236 24744 41288 24750
rect 41236 24686 41288 24692
rect 41248 24041 41276 24686
rect 41234 24032 41290 24041
rect 41234 23967 41290 23976
rect 40960 21344 41012 21350
rect 40960 21286 41012 21292
rect 40684 20868 40736 20874
rect 40684 20810 40736 20816
rect 40972 20466 41000 21286
rect 41052 20800 41104 20806
rect 41052 20742 41104 20748
rect 40684 20460 40736 20466
rect 40684 20402 40736 20408
rect 40960 20460 41012 20466
rect 40960 20402 41012 20408
rect 40590 19816 40646 19825
rect 40590 19751 40646 19760
rect 40604 19378 40632 19751
rect 40500 19372 40552 19378
rect 40420 19320 40500 19334
rect 40420 19314 40552 19320
rect 40592 19372 40644 19378
rect 40592 19314 40644 19320
rect 40420 19306 40540 19314
rect 40420 18834 40448 19306
rect 40592 19236 40644 19242
rect 40592 19178 40644 19184
rect 40408 18828 40460 18834
rect 40408 18770 40460 18776
rect 40316 18352 40368 18358
rect 40316 18294 40368 18300
rect 40328 17338 40356 18294
rect 40420 17746 40448 18770
rect 40604 18766 40632 19178
rect 40500 18760 40552 18766
rect 40500 18702 40552 18708
rect 40592 18760 40644 18766
rect 40592 18702 40644 18708
rect 40512 18222 40540 18702
rect 40592 18624 40644 18630
rect 40696 18612 40724 20402
rect 40868 20256 40920 20262
rect 40868 20198 40920 20204
rect 40880 19922 40908 20198
rect 40868 19916 40920 19922
rect 40868 19858 40920 19864
rect 40644 18584 40724 18612
rect 40592 18566 40644 18572
rect 40500 18216 40552 18222
rect 40500 18158 40552 18164
rect 40408 17740 40460 17746
rect 40408 17682 40460 17688
rect 40316 17332 40368 17338
rect 40316 17274 40368 17280
rect 40224 16992 40276 16998
rect 40224 16934 40276 16940
rect 40236 16114 40264 16934
rect 40316 16516 40368 16522
rect 40316 16458 40368 16464
rect 40224 16108 40276 16114
rect 40224 16050 40276 16056
rect 40132 15088 40184 15094
rect 40132 15030 40184 15036
rect 40144 14498 40172 15030
rect 40236 14600 40264 16050
rect 40328 16046 40356 16458
rect 40316 16040 40368 16046
rect 40316 15982 40368 15988
rect 40604 15994 40632 18566
rect 40776 18420 40828 18426
rect 40776 18362 40828 18368
rect 40684 16720 40736 16726
rect 40788 16674 40816 18362
rect 41064 17814 41092 20742
rect 41340 20466 41368 27798
rect 41418 27775 41474 27784
rect 41432 27606 41460 27775
rect 41420 27600 41472 27606
rect 41420 27542 41472 27548
rect 41524 27470 41552 28018
rect 41512 27464 41564 27470
rect 41512 27406 41564 27412
rect 41616 26926 41644 28206
rect 41604 26920 41656 26926
rect 41604 26862 41656 26868
rect 41708 26382 41736 29514
rect 41892 29170 41920 29514
rect 41984 29306 42012 31962
rect 42248 31816 42300 31822
rect 42444 31804 42472 32286
rect 42524 32224 42576 32230
rect 42524 32166 42576 32172
rect 42300 31776 42472 31804
rect 42248 31758 42300 31764
rect 42340 30320 42392 30326
rect 42340 30262 42392 30268
rect 42156 30048 42208 30054
rect 42156 29990 42208 29996
rect 42168 29850 42196 29990
rect 42156 29844 42208 29850
rect 42156 29786 42208 29792
rect 42064 29640 42116 29646
rect 42064 29582 42116 29588
rect 41972 29300 42024 29306
rect 41972 29242 42024 29248
rect 42076 29170 42104 29582
rect 41880 29164 41932 29170
rect 41800 29124 41880 29152
rect 41800 28558 41828 29124
rect 41880 29106 41932 29112
rect 42064 29164 42116 29170
rect 42064 29106 42116 29112
rect 42156 29164 42208 29170
rect 42156 29106 42208 29112
rect 42168 29034 42196 29106
rect 42156 29028 42208 29034
rect 42156 28970 42208 28976
rect 41972 28960 42024 28966
rect 41972 28902 42024 28908
rect 41984 28558 42012 28902
rect 42064 28620 42116 28626
rect 42064 28562 42116 28568
rect 41788 28552 41840 28558
rect 41788 28494 41840 28500
rect 41972 28552 42024 28558
rect 41972 28494 42024 28500
rect 41800 28218 41828 28494
rect 41788 28212 41840 28218
rect 41788 28154 41840 28160
rect 41800 27996 41828 28154
rect 41880 28008 41932 28014
rect 41800 27968 41880 27996
rect 41880 27950 41932 27956
rect 41984 27946 42012 28494
rect 41972 27940 42024 27946
rect 41972 27882 42024 27888
rect 42076 27878 42104 28562
rect 41788 27872 41840 27878
rect 41788 27814 41840 27820
rect 42064 27872 42116 27878
rect 42064 27814 42116 27820
rect 41800 27674 41828 27814
rect 41788 27668 41840 27674
rect 41788 27610 41840 27616
rect 41800 27538 42012 27554
rect 41788 27532 42024 27538
rect 41840 27526 41972 27532
rect 41788 27474 41840 27480
rect 41972 27474 42024 27480
rect 41972 27396 42024 27402
rect 41972 27338 42024 27344
rect 41880 27328 41932 27334
rect 41880 27270 41932 27276
rect 41788 27056 41840 27062
rect 41788 26998 41840 27004
rect 41696 26376 41748 26382
rect 41696 26318 41748 26324
rect 41696 24948 41748 24954
rect 41696 24890 41748 24896
rect 41420 24812 41472 24818
rect 41420 24754 41472 24760
rect 41432 23730 41460 24754
rect 41512 24744 41564 24750
rect 41512 24686 41564 24692
rect 41524 24410 41552 24686
rect 41512 24404 41564 24410
rect 41512 24346 41564 24352
rect 41604 24200 41656 24206
rect 41602 24168 41604 24177
rect 41656 24168 41658 24177
rect 41602 24103 41658 24112
rect 41708 23769 41736 24890
rect 41800 24886 41828 26998
rect 41892 26858 41920 27270
rect 41880 26852 41932 26858
rect 41880 26794 41932 26800
rect 41984 26382 42012 27338
rect 42076 27130 42104 27814
rect 42064 27124 42116 27130
rect 42064 27066 42116 27072
rect 42076 26858 42104 27066
rect 42064 26852 42116 26858
rect 42064 26794 42116 26800
rect 41972 26376 42024 26382
rect 41972 26318 42024 26324
rect 42076 25838 42104 26794
rect 42064 25832 42116 25838
rect 42064 25774 42116 25780
rect 41788 24880 41840 24886
rect 41788 24822 41840 24828
rect 41694 23760 41750 23769
rect 41420 23724 41472 23730
rect 41420 23666 41472 23672
rect 41604 23724 41656 23730
rect 41694 23695 41696 23704
rect 41604 23666 41656 23672
rect 41748 23695 41750 23704
rect 41696 23666 41748 23672
rect 41616 21894 41644 23666
rect 41800 22094 41828 24822
rect 42168 24426 42196 28970
rect 42248 27464 42300 27470
rect 42248 27406 42300 27412
rect 42260 26994 42288 27406
rect 42248 26988 42300 26994
rect 42248 26930 42300 26936
rect 42260 26382 42288 26930
rect 42248 26376 42300 26382
rect 42248 26318 42300 26324
rect 42076 24398 42196 24426
rect 41878 24304 41934 24313
rect 41878 24239 41934 24248
rect 41892 24206 41920 24239
rect 41880 24200 41932 24206
rect 41880 24142 41932 24148
rect 41972 24200 42024 24206
rect 41972 24142 42024 24148
rect 41984 23882 42012 24142
rect 41892 23854 42012 23882
rect 41892 23798 41920 23854
rect 41880 23792 41932 23798
rect 41880 23734 41932 23740
rect 41892 23322 41920 23734
rect 41880 23316 41932 23322
rect 41880 23258 41932 23264
rect 42076 23254 42104 24398
rect 42156 24336 42208 24342
rect 42156 24278 42208 24284
rect 42168 24154 42196 24278
rect 42168 24126 42288 24154
rect 42156 24064 42208 24070
rect 42156 24006 42208 24012
rect 42168 23866 42196 24006
rect 42156 23860 42208 23866
rect 42156 23802 42208 23808
rect 42260 23594 42288 24126
rect 42352 23866 42380 30262
rect 42536 29714 42564 32166
rect 42720 31822 42748 32438
rect 42904 32366 42932 32846
rect 43166 32600 43222 32609
rect 43166 32535 43222 32544
rect 43180 32502 43208 32535
rect 43168 32496 43220 32502
rect 43168 32438 43220 32444
rect 42892 32360 42944 32366
rect 42892 32302 42944 32308
rect 43076 32224 43128 32230
rect 43076 32166 43128 32172
rect 42708 31816 42760 31822
rect 42708 31758 42760 31764
rect 43088 31346 43116 32166
rect 43076 31340 43128 31346
rect 43076 31282 43128 31288
rect 42708 31272 42760 31278
rect 42708 31214 42760 31220
rect 42720 29866 42748 31214
rect 43180 30258 43208 32438
rect 43272 32314 43300 35866
rect 44180 34740 44232 34746
rect 44180 34682 44232 34688
rect 43812 34400 43864 34406
rect 43812 34342 43864 34348
rect 43824 34066 43852 34342
rect 44192 34066 44220 34682
rect 43812 34060 43864 34066
rect 43812 34002 43864 34008
rect 44180 34060 44232 34066
rect 44180 34002 44232 34008
rect 45192 34060 45244 34066
rect 45192 34002 45244 34008
rect 43824 33590 43852 34002
rect 44456 33992 44508 33998
rect 44456 33934 44508 33940
rect 43812 33584 43864 33590
rect 43812 33526 43864 33532
rect 44468 33522 44496 33934
rect 45008 33924 45060 33930
rect 45008 33866 45060 33872
rect 45020 33522 45048 33866
rect 43904 33516 43956 33522
rect 43904 33458 43956 33464
rect 44456 33516 44508 33522
rect 44456 33458 44508 33464
rect 44548 33516 44600 33522
rect 44548 33458 44600 33464
rect 44916 33516 44968 33522
rect 44916 33458 44968 33464
rect 45008 33516 45060 33522
rect 45008 33458 45060 33464
rect 43444 33312 43496 33318
rect 43444 33254 43496 33260
rect 43456 32434 43484 33254
rect 43812 33108 43864 33114
rect 43812 33050 43864 33056
rect 43444 32428 43496 32434
rect 43444 32370 43496 32376
rect 43272 32286 43484 32314
rect 43168 30252 43220 30258
rect 43168 30194 43220 30200
rect 42720 29838 42932 29866
rect 42616 29776 42668 29782
rect 42616 29718 42668 29724
rect 42524 29708 42576 29714
rect 42524 29650 42576 29656
rect 42628 29170 42656 29718
rect 42708 29708 42760 29714
rect 42708 29650 42760 29656
rect 42616 29164 42668 29170
rect 42616 29106 42668 29112
rect 42432 28620 42484 28626
rect 42432 28562 42484 28568
rect 42444 28014 42472 28562
rect 42616 28416 42668 28422
rect 42616 28358 42668 28364
rect 42628 28218 42656 28358
rect 42616 28212 42668 28218
rect 42616 28154 42668 28160
rect 42432 28008 42484 28014
rect 42432 27950 42484 27956
rect 42444 27062 42472 27950
rect 42524 27940 42576 27946
rect 42524 27882 42576 27888
rect 42432 27056 42484 27062
rect 42432 26998 42484 27004
rect 42432 26920 42484 26926
rect 42432 26862 42484 26868
rect 42444 26382 42472 26862
rect 42432 26376 42484 26382
rect 42432 26318 42484 26324
rect 42536 25906 42564 27882
rect 42616 27872 42668 27878
rect 42614 27840 42616 27849
rect 42668 27840 42670 27849
rect 42614 27775 42670 27784
rect 42616 26988 42668 26994
rect 42616 26930 42668 26936
rect 42628 26586 42656 26930
rect 42616 26580 42668 26586
rect 42616 26522 42668 26528
rect 42628 26450 42656 26522
rect 42616 26444 42668 26450
rect 42616 26386 42668 26392
rect 42524 25900 42576 25906
rect 42524 25842 42576 25848
rect 42616 25832 42668 25838
rect 42616 25774 42668 25780
rect 42524 25696 42576 25702
rect 42524 25638 42576 25644
rect 42536 24818 42564 25638
rect 42524 24812 42576 24818
rect 42524 24754 42576 24760
rect 42522 24304 42578 24313
rect 42432 24268 42484 24274
rect 42522 24239 42524 24248
rect 42432 24210 42484 24216
rect 42576 24239 42578 24248
rect 42524 24210 42576 24216
rect 42444 24177 42472 24210
rect 42430 24168 42486 24177
rect 42430 24103 42486 24112
rect 42340 23860 42392 23866
rect 42340 23802 42392 23808
rect 42248 23588 42300 23594
rect 42248 23530 42300 23536
rect 42064 23248 42116 23254
rect 42064 23190 42116 23196
rect 41708 22066 41828 22094
rect 41604 21888 41656 21894
rect 41604 21830 41656 21836
rect 41604 21548 41656 21554
rect 41604 21490 41656 21496
rect 41616 20466 41644 21490
rect 41708 21486 41736 22066
rect 42352 22012 42380 23802
rect 42432 23316 42484 23322
rect 42432 23258 42484 23264
rect 42444 23118 42472 23258
rect 42524 23180 42576 23186
rect 42524 23122 42576 23128
rect 42432 23112 42484 23118
rect 42432 23054 42484 23060
rect 42536 22166 42564 23122
rect 42628 22982 42656 25774
rect 42616 22976 42668 22982
rect 42616 22918 42668 22924
rect 42720 22642 42748 29650
rect 42904 29578 42932 29838
rect 43180 29782 43208 30194
rect 43168 29776 43220 29782
rect 43168 29718 43220 29724
rect 43076 29640 43128 29646
rect 43076 29582 43128 29588
rect 42892 29572 42944 29578
rect 42892 29514 42944 29520
rect 42904 27946 42932 29514
rect 43088 29238 43116 29582
rect 43076 29232 43128 29238
rect 43076 29174 43128 29180
rect 43180 29170 43208 29718
rect 43168 29164 43220 29170
rect 43168 29106 43220 29112
rect 42892 27940 42944 27946
rect 42892 27882 42944 27888
rect 42800 27872 42852 27878
rect 42800 27814 42852 27820
rect 42812 27538 42840 27814
rect 42800 27532 42852 27538
rect 42800 27474 42852 27480
rect 43352 27056 43404 27062
rect 43352 26998 43404 27004
rect 43260 26988 43312 26994
rect 43260 26930 43312 26936
rect 42984 26920 43036 26926
rect 42984 26862 43036 26868
rect 42800 26512 42852 26518
rect 42800 26454 42852 26460
rect 42812 25838 42840 26454
rect 42996 26382 43024 26862
rect 43168 26580 43220 26586
rect 43168 26522 43220 26528
rect 43180 26382 43208 26522
rect 43272 26450 43300 26930
rect 43260 26444 43312 26450
rect 43260 26386 43312 26392
rect 43364 26382 43392 26998
rect 42984 26376 43036 26382
rect 42984 26318 43036 26324
rect 43168 26376 43220 26382
rect 43168 26318 43220 26324
rect 43352 26376 43404 26382
rect 43352 26318 43404 26324
rect 42892 26036 42944 26042
rect 42892 25978 42944 25984
rect 42800 25832 42852 25838
rect 42800 25774 42852 25780
rect 42812 23798 42840 25774
rect 42800 23792 42852 23798
rect 42800 23734 42852 23740
rect 42904 23118 42932 25978
rect 42996 24177 43024 26318
rect 43180 25838 43208 26318
rect 43260 26240 43312 26246
rect 43364 26194 43392 26318
rect 43312 26188 43392 26194
rect 43260 26182 43392 26188
rect 43272 26166 43392 26182
rect 43272 25906 43300 26166
rect 43260 25900 43312 25906
rect 43260 25842 43312 25848
rect 43168 25832 43220 25838
rect 43168 25774 43220 25780
rect 43272 25702 43300 25842
rect 43260 25696 43312 25702
rect 43260 25638 43312 25644
rect 43352 24268 43404 24274
rect 43352 24210 43404 24216
rect 43076 24200 43128 24206
rect 42982 24168 43038 24177
rect 43260 24200 43312 24206
rect 43076 24142 43128 24148
rect 43258 24168 43260 24177
rect 43312 24168 43314 24177
rect 42982 24103 43038 24112
rect 42982 24032 43038 24041
rect 42982 23967 43038 23976
rect 42892 23112 42944 23118
rect 42892 23054 42944 23060
rect 42892 22976 42944 22982
rect 42892 22918 42944 22924
rect 42904 22642 42932 22918
rect 42708 22636 42760 22642
rect 42708 22578 42760 22584
rect 42892 22636 42944 22642
rect 42892 22578 42944 22584
rect 42616 22568 42668 22574
rect 42616 22510 42668 22516
rect 42524 22160 42576 22166
rect 42524 22102 42576 22108
rect 42628 22094 42656 22510
rect 42892 22160 42944 22166
rect 42892 22102 42944 22108
rect 42628 22066 42840 22094
rect 42628 22030 42656 22066
rect 42812 22030 42840 22066
rect 42432 22024 42484 22030
rect 42352 21984 42432 22012
rect 42432 21966 42484 21972
rect 42616 22024 42668 22030
rect 42616 21966 42668 21972
rect 42708 22024 42760 22030
rect 42708 21966 42760 21972
rect 42800 22024 42852 22030
rect 42800 21966 42852 21972
rect 42156 21888 42208 21894
rect 42156 21830 42208 21836
rect 42168 21554 42196 21830
rect 42720 21622 42748 21966
rect 42708 21616 42760 21622
rect 42708 21558 42760 21564
rect 42156 21548 42208 21554
rect 42156 21490 42208 21496
rect 41696 21480 41748 21486
rect 41696 21422 41748 21428
rect 41328 20460 41380 20466
rect 41328 20402 41380 20408
rect 41420 20460 41472 20466
rect 41420 20402 41472 20408
rect 41604 20460 41656 20466
rect 41604 20402 41656 20408
rect 41432 20058 41460 20402
rect 41604 20324 41656 20330
rect 41604 20266 41656 20272
rect 41512 20256 41564 20262
rect 41512 20198 41564 20204
rect 41420 20052 41472 20058
rect 41420 19994 41472 20000
rect 41524 19854 41552 20198
rect 41616 20058 41644 20266
rect 41604 20052 41656 20058
rect 41604 19994 41656 20000
rect 41512 19848 41564 19854
rect 41512 19790 41564 19796
rect 41616 19666 41644 19994
rect 41524 19638 41644 19666
rect 41328 19304 41380 19310
rect 41328 19246 41380 19252
rect 41340 18970 41368 19246
rect 41420 19236 41472 19242
rect 41420 19178 41472 19184
rect 41328 18964 41380 18970
rect 41328 18906 41380 18912
rect 41144 18760 41196 18766
rect 41144 18702 41196 18708
rect 41156 18222 41184 18702
rect 41340 18272 41368 18906
rect 41432 18834 41460 19178
rect 41420 18828 41472 18834
rect 41420 18770 41472 18776
rect 41524 18630 41552 19638
rect 41708 19530 41736 21422
rect 42616 21412 42668 21418
rect 42616 21354 42668 21360
rect 41880 21344 41932 21350
rect 41880 21286 41932 21292
rect 41616 19502 41736 19530
rect 41512 18624 41564 18630
rect 41512 18566 41564 18572
rect 41420 18284 41472 18290
rect 41340 18244 41420 18272
rect 41420 18226 41472 18232
rect 41524 18222 41552 18566
rect 41144 18216 41196 18222
rect 41144 18158 41196 18164
rect 41512 18216 41564 18222
rect 41512 18158 41564 18164
rect 41052 17808 41104 17814
rect 41052 17750 41104 17756
rect 40868 17060 40920 17066
rect 40868 17002 40920 17008
rect 40880 16726 40908 17002
rect 40736 16668 40816 16674
rect 40684 16662 40816 16668
rect 40868 16720 40920 16726
rect 40868 16662 40920 16668
rect 40696 16646 40816 16662
rect 41064 16658 41092 17750
rect 41156 17134 41184 18158
rect 41236 18080 41288 18086
rect 41236 18022 41288 18028
rect 41248 17882 41276 18022
rect 41236 17876 41288 17882
rect 41236 17818 41288 17824
rect 41328 17672 41380 17678
rect 41328 17614 41380 17620
rect 41340 17338 41368 17614
rect 41236 17332 41288 17338
rect 41236 17274 41288 17280
rect 41328 17332 41380 17338
rect 41328 17274 41380 17280
rect 41248 17134 41276 17274
rect 41144 17128 41196 17134
rect 41144 17070 41196 17076
rect 41236 17128 41288 17134
rect 41236 17070 41288 17076
rect 40788 16590 40816 16646
rect 41052 16652 41104 16658
rect 41052 16594 41104 16600
rect 41248 16590 41276 17070
rect 40776 16584 40828 16590
rect 40776 16526 40828 16532
rect 40960 16584 41012 16590
rect 40960 16526 41012 16532
rect 41236 16584 41288 16590
rect 41236 16526 41288 16532
rect 40972 16454 41000 16526
rect 41616 16454 41644 19502
rect 41788 18828 41840 18834
rect 41788 18770 41840 18776
rect 41696 18216 41748 18222
rect 41696 18158 41748 18164
rect 41708 18086 41736 18158
rect 41800 18154 41828 18770
rect 41788 18148 41840 18154
rect 41788 18090 41840 18096
rect 41696 18080 41748 18086
rect 41696 18022 41748 18028
rect 41708 17202 41736 18022
rect 41892 17542 41920 21286
rect 42524 21004 42576 21010
rect 42524 20946 42576 20952
rect 42340 20460 42392 20466
rect 42340 20402 42392 20408
rect 42352 20330 42380 20402
rect 42340 20324 42392 20330
rect 42340 20266 42392 20272
rect 42352 19310 42380 20266
rect 42432 20256 42484 20262
rect 42432 20198 42484 20204
rect 42444 19854 42472 20198
rect 42432 19848 42484 19854
rect 42432 19790 42484 19796
rect 42340 19304 42392 19310
rect 42340 19246 42392 19252
rect 42064 18760 42116 18766
rect 42064 18702 42116 18708
rect 42076 18222 42104 18702
rect 42064 18216 42116 18222
rect 42116 18176 42288 18204
rect 42064 18158 42116 18164
rect 41880 17536 41932 17542
rect 41880 17478 41932 17484
rect 42260 17338 42288 18176
rect 42156 17332 42208 17338
rect 42156 17274 42208 17280
rect 42248 17332 42300 17338
rect 42248 17274 42300 17280
rect 42064 17264 42116 17270
rect 42064 17206 42116 17212
rect 41696 17196 41748 17202
rect 41696 17138 41748 17144
rect 42076 16794 42104 17206
rect 42064 16788 42116 16794
rect 42064 16730 42116 16736
rect 42168 16590 42196 17274
rect 42260 17066 42288 17274
rect 42248 17060 42300 17066
rect 42248 17002 42300 17008
rect 42340 16992 42392 16998
rect 42340 16934 42392 16940
rect 42352 16590 42380 16934
rect 42536 16590 42564 20946
rect 42628 20448 42656 21354
rect 42904 21010 42932 22102
rect 42892 21004 42944 21010
rect 42892 20946 42944 20952
rect 42892 20868 42944 20874
rect 42892 20810 42944 20816
rect 42708 20460 42760 20466
rect 42628 20420 42708 20448
rect 42628 20058 42656 20420
rect 42708 20402 42760 20408
rect 42616 20052 42668 20058
rect 42616 19994 42668 20000
rect 42800 19780 42852 19786
rect 42800 19722 42852 19728
rect 42812 19446 42840 19722
rect 42800 19440 42852 19446
rect 42800 19382 42852 19388
rect 42812 19174 42840 19382
rect 42800 19168 42852 19174
rect 42800 19110 42852 19116
rect 42904 17882 42932 20810
rect 42996 20806 43024 23967
rect 43088 23866 43116 24142
rect 43258 24103 43314 24112
rect 43076 23860 43128 23866
rect 43076 23802 43128 23808
rect 43364 23798 43392 24210
rect 43352 23792 43404 23798
rect 43352 23734 43404 23740
rect 43076 23656 43128 23662
rect 43076 23598 43128 23604
rect 43088 23254 43116 23598
rect 43076 23248 43128 23254
rect 43076 23190 43128 23196
rect 43260 22976 43312 22982
rect 43260 22918 43312 22924
rect 43272 22574 43300 22918
rect 43260 22568 43312 22574
rect 43260 22510 43312 22516
rect 43260 22432 43312 22438
rect 43260 22374 43312 22380
rect 43272 21554 43300 22374
rect 43352 22228 43404 22234
rect 43352 22170 43404 22176
rect 43168 21548 43220 21554
rect 43168 21490 43220 21496
rect 43260 21548 43312 21554
rect 43260 21490 43312 21496
rect 42984 20800 43036 20806
rect 42984 20742 43036 20748
rect 42984 20460 43036 20466
rect 42984 20402 43036 20408
rect 42996 20058 43024 20402
rect 43180 20262 43208 21490
rect 43364 20942 43392 22170
rect 43352 20936 43404 20942
rect 43352 20878 43404 20884
rect 43168 20256 43220 20262
rect 43168 20198 43220 20204
rect 42984 20052 43036 20058
rect 42984 19994 43036 20000
rect 42892 17876 42944 17882
rect 42892 17818 42944 17824
rect 42800 17604 42852 17610
rect 42800 17546 42852 17552
rect 42812 17338 42840 17546
rect 42800 17332 42852 17338
rect 42800 17274 42852 17280
rect 42812 16794 42840 17274
rect 42708 16788 42760 16794
rect 42708 16730 42760 16736
rect 42800 16788 42852 16794
rect 42800 16730 42852 16736
rect 42616 16652 42668 16658
rect 42616 16594 42668 16600
rect 42156 16584 42208 16590
rect 42156 16526 42208 16532
rect 42340 16584 42392 16590
rect 42340 16526 42392 16532
rect 42524 16584 42576 16590
rect 42524 16526 42576 16532
rect 40776 16448 40828 16454
rect 40776 16390 40828 16396
rect 40960 16448 41012 16454
rect 40960 16390 41012 16396
rect 41328 16448 41380 16454
rect 41328 16390 41380 16396
rect 41604 16448 41656 16454
rect 41604 16390 41656 16396
rect 40788 16114 40816 16390
rect 40776 16108 40828 16114
rect 40776 16050 40828 16056
rect 40604 15966 40816 15994
rect 40316 14612 40368 14618
rect 40236 14572 40316 14600
rect 40316 14554 40368 14560
rect 40144 14470 40264 14498
rect 40236 14414 40264 14470
rect 40592 14476 40644 14482
rect 40592 14418 40644 14424
rect 39856 14408 39908 14414
rect 39856 14350 39908 14356
rect 40132 14408 40184 14414
rect 40132 14350 40184 14356
rect 40224 14408 40276 14414
rect 40224 14350 40276 14356
rect 39868 12986 39896 14350
rect 40144 14074 40172 14350
rect 40500 14272 40552 14278
rect 40500 14214 40552 14220
rect 40132 14068 40184 14074
rect 40132 14010 40184 14016
rect 40512 14006 40540 14214
rect 40500 14000 40552 14006
rect 40500 13942 40552 13948
rect 39856 12980 39908 12986
rect 39856 12922 39908 12928
rect 39948 12844 40000 12850
rect 39948 12786 40000 12792
rect 39960 12714 39988 12786
rect 39948 12708 40000 12714
rect 39948 12650 40000 12656
rect 38844 12232 38896 12238
rect 39764 12232 39816 12238
rect 39210 12200 39266 12209
rect 38896 12180 39068 12186
rect 38844 12174 39068 12180
rect 38856 12158 39068 12174
rect 38844 12096 38896 12102
rect 38844 12038 38896 12044
rect 38936 12096 38988 12102
rect 38936 12038 38988 12044
rect 38856 11830 38884 12038
rect 38844 11824 38896 11830
rect 38750 11792 38806 11801
rect 38844 11766 38896 11772
rect 38750 11727 38806 11736
rect 38844 11688 38896 11694
rect 38948 11676 38976 12038
rect 38896 11648 38976 11676
rect 38844 11630 38896 11636
rect 39040 11354 39068 12158
rect 39120 12164 39172 12170
rect 39764 12174 39816 12180
rect 39210 12135 39266 12144
rect 39120 12106 39172 12112
rect 38752 11348 38804 11354
rect 38752 11290 38804 11296
rect 39028 11348 39080 11354
rect 39028 11290 39080 11296
rect 38764 10674 38792 11290
rect 39132 11150 39160 12106
rect 38844 11144 38896 11150
rect 38844 11086 38896 11092
rect 39120 11144 39172 11150
rect 39120 11086 39172 11092
rect 38856 10810 38884 11086
rect 39132 11014 39160 11086
rect 39120 11008 39172 11014
rect 39120 10950 39172 10956
rect 38844 10804 38896 10810
rect 38844 10746 38896 10752
rect 39132 10674 39160 10950
rect 38752 10668 38804 10674
rect 38752 10610 38804 10616
rect 39120 10668 39172 10674
rect 39120 10610 39172 10616
rect 38660 10600 38712 10606
rect 38660 10542 38712 10548
rect 38384 10532 38436 10538
rect 38384 10474 38436 10480
rect 38292 10464 38344 10470
rect 38292 10406 38344 10412
rect 38304 9994 38332 10406
rect 38292 9988 38344 9994
rect 38292 9930 38344 9936
rect 38396 9586 38424 10474
rect 39224 10130 39252 12135
rect 39396 11756 39448 11762
rect 39396 11698 39448 11704
rect 39304 11144 39356 11150
rect 39304 11086 39356 11092
rect 39316 10810 39344 11086
rect 39408 11014 39436 11698
rect 39960 11540 39988 12650
rect 40040 12640 40092 12646
rect 40040 12582 40092 12588
rect 40052 12442 40080 12582
rect 40040 12436 40092 12442
rect 40040 12378 40092 12384
rect 40408 12232 40460 12238
rect 40408 12174 40460 12180
rect 40224 12096 40276 12102
rect 40224 12038 40276 12044
rect 40040 11552 40092 11558
rect 39960 11512 40040 11540
rect 40040 11494 40092 11500
rect 39488 11280 39540 11286
rect 39488 11222 39540 11228
rect 39396 11008 39448 11014
rect 39396 10950 39448 10956
rect 39304 10804 39356 10810
rect 39304 10746 39356 10752
rect 39500 10554 39528 11222
rect 39580 11008 39632 11014
rect 39580 10950 39632 10956
rect 39592 10742 39620 10950
rect 39580 10736 39632 10742
rect 39580 10678 39632 10684
rect 40052 10674 40080 11494
rect 40040 10668 40092 10674
rect 40040 10610 40092 10616
rect 39408 10538 39528 10554
rect 39854 10568 39910 10577
rect 39408 10532 39540 10538
rect 39408 10526 39488 10532
rect 39212 10124 39264 10130
rect 39212 10066 39264 10072
rect 39408 10062 39436 10526
rect 39854 10503 39910 10512
rect 39488 10474 39540 10480
rect 39396 10056 39448 10062
rect 39396 9998 39448 10004
rect 39488 10056 39540 10062
rect 39488 9998 39540 10004
rect 38384 9580 38436 9586
rect 38384 9522 38436 9528
rect 38660 9580 38712 9586
rect 38660 9522 38712 9528
rect 38108 9376 38160 9382
rect 38108 9318 38160 9324
rect 38384 9376 38436 9382
rect 38384 9318 38436 9324
rect 38396 9178 38424 9318
rect 38384 9172 38436 9178
rect 38384 9114 38436 9120
rect 38476 8832 38528 8838
rect 38476 8774 38528 8780
rect 37648 8492 37700 8498
rect 37648 8434 37700 8440
rect 38016 8492 38068 8498
rect 38016 8434 38068 8440
rect 37464 8288 37516 8294
rect 37464 8230 37516 8236
rect 37476 7546 37504 8230
rect 37464 7540 37516 7546
rect 37464 7482 37516 7488
rect 37476 6934 37504 7482
rect 37464 6928 37516 6934
rect 37464 6870 37516 6876
rect 37462 2680 37518 2689
rect 37462 2615 37518 2624
rect 34886 2479 34942 2488
rect 37188 2508 37240 2514
rect 34900 2446 34928 2479
rect 37188 2450 37240 2456
rect 37476 2446 37504 2615
rect 37660 2582 37688 8434
rect 38028 7886 38056 8434
rect 38488 8430 38516 8774
rect 38476 8424 38528 8430
rect 38476 8366 38528 8372
rect 38672 8090 38700 9522
rect 39500 9518 39528 9998
rect 39764 9920 39816 9926
rect 39764 9862 39816 9868
rect 39488 9512 39540 9518
rect 39488 9454 39540 9460
rect 39672 8968 39724 8974
rect 39672 8910 39724 8916
rect 39684 8566 39712 8910
rect 39776 8634 39804 9862
rect 39868 9722 39896 10503
rect 39856 9716 39908 9722
rect 39856 9658 39908 9664
rect 39868 8634 39896 9658
rect 40052 9586 40080 10610
rect 40040 9580 40092 9586
rect 40040 9522 40092 9528
rect 39764 8628 39816 8634
rect 39764 8570 39816 8576
rect 39856 8628 39908 8634
rect 39856 8570 39908 8576
rect 39672 8560 39724 8566
rect 39672 8502 39724 8508
rect 40236 8498 40264 12038
rect 40420 11762 40448 12174
rect 40408 11756 40460 11762
rect 40408 11698 40460 11704
rect 40420 10810 40448 11698
rect 40408 10804 40460 10810
rect 40408 10746 40460 10752
rect 40500 10736 40552 10742
rect 40500 10678 40552 10684
rect 40408 10668 40460 10674
rect 40408 10610 40460 10616
rect 40316 10532 40368 10538
rect 40316 10474 40368 10480
rect 40328 9586 40356 10474
rect 40420 10266 40448 10610
rect 40408 10260 40460 10266
rect 40408 10202 40460 10208
rect 40512 9654 40540 10678
rect 40604 10130 40632 14418
rect 40684 14272 40736 14278
rect 40684 14214 40736 14220
rect 40696 13938 40724 14214
rect 40684 13932 40736 13938
rect 40684 13874 40736 13880
rect 40788 12434 40816 15966
rect 41236 15496 41288 15502
rect 41236 15438 41288 15444
rect 41144 14816 41196 14822
rect 41144 14758 41196 14764
rect 40960 14408 41012 14414
rect 40960 14350 41012 14356
rect 40972 14074 41000 14350
rect 40960 14068 41012 14074
rect 40960 14010 41012 14016
rect 41156 13938 41184 14758
rect 41248 14618 41276 15438
rect 41236 14612 41288 14618
rect 41236 14554 41288 14560
rect 41144 13932 41196 13938
rect 41144 13874 41196 13880
rect 40960 13864 41012 13870
rect 40960 13806 41012 13812
rect 40972 12782 41000 13806
rect 40960 12776 41012 12782
rect 40960 12718 41012 12724
rect 41052 12776 41104 12782
rect 41052 12718 41104 12724
rect 40696 12406 40816 12434
rect 40592 10124 40644 10130
rect 40592 10066 40644 10072
rect 40500 9648 40552 9654
rect 40500 9590 40552 9596
rect 40696 9586 40724 12406
rect 40868 12368 40920 12374
rect 40868 12310 40920 12316
rect 40774 11656 40830 11665
rect 40774 11591 40830 11600
rect 40788 11150 40816 11591
rect 40776 11144 40828 11150
rect 40776 11086 40828 11092
rect 40776 10668 40828 10674
rect 40880 10656 40908 12310
rect 41064 12170 41092 12718
rect 41052 12164 41104 12170
rect 41052 12106 41104 12112
rect 41340 11665 41368 16390
rect 42168 16114 42196 16526
rect 42156 16108 42208 16114
rect 42156 16050 42208 16056
rect 42524 15972 42576 15978
rect 42524 15914 42576 15920
rect 42536 15026 42564 15914
rect 42156 15020 42208 15026
rect 42156 14962 42208 14968
rect 42524 15020 42576 15026
rect 42524 14962 42576 14968
rect 42168 14618 42196 14962
rect 42156 14612 42208 14618
rect 42156 14554 42208 14560
rect 42248 13932 42300 13938
rect 42248 13874 42300 13880
rect 41604 12708 41656 12714
rect 41604 12650 41656 12656
rect 41616 12442 41644 12650
rect 41604 12436 41656 12442
rect 41604 12378 41656 12384
rect 41696 12436 41748 12442
rect 41696 12378 41748 12384
rect 41708 12238 41736 12378
rect 42260 12238 42288 13874
rect 42536 13326 42564 14962
rect 42524 13320 42576 13326
rect 42524 13262 42576 13268
rect 41696 12232 41748 12238
rect 41696 12174 41748 12180
rect 42248 12232 42300 12238
rect 42300 12192 42564 12220
rect 42248 12174 42300 12180
rect 41420 12096 41472 12102
rect 41420 12038 41472 12044
rect 41432 11898 41460 12038
rect 41708 11898 41736 12174
rect 41420 11892 41472 11898
rect 41420 11834 41472 11840
rect 41696 11892 41748 11898
rect 41696 11834 41748 11840
rect 42064 11756 42116 11762
rect 42064 11698 42116 11704
rect 41326 11656 41382 11665
rect 42076 11642 42104 11698
rect 42432 11688 42484 11694
rect 42076 11636 42432 11642
rect 42076 11630 42484 11636
rect 42076 11614 42472 11630
rect 41326 11591 41382 11600
rect 42444 10810 42472 11614
rect 42536 11354 42564 12192
rect 42524 11348 42576 11354
rect 42524 11290 42576 11296
rect 42628 11150 42656 16594
rect 42720 16590 42748 16730
rect 42708 16584 42760 16590
rect 42708 16526 42760 16532
rect 42708 16448 42760 16454
rect 42708 16390 42760 16396
rect 42720 16114 42748 16390
rect 42708 16108 42760 16114
rect 42708 16050 42760 16056
rect 42904 13818 42932 17818
rect 43076 17196 43128 17202
rect 43076 17138 43128 17144
rect 43088 16590 43116 17138
rect 43180 17134 43208 20198
rect 43364 19854 43392 20878
rect 43456 20602 43484 32286
rect 43720 31816 43772 31822
rect 43720 31758 43772 31764
rect 43732 30258 43760 31758
rect 43720 30252 43772 30258
rect 43720 30194 43772 30200
rect 43720 29096 43772 29102
rect 43720 29038 43772 29044
rect 43732 28558 43760 29038
rect 43720 28552 43772 28558
rect 43720 28494 43772 28500
rect 43536 28076 43588 28082
rect 43536 28018 43588 28024
rect 43548 27946 43576 28018
rect 43536 27940 43588 27946
rect 43536 27882 43588 27888
rect 43720 25356 43772 25362
rect 43720 25298 43772 25304
rect 43732 24682 43760 25298
rect 43720 24676 43772 24682
rect 43720 24618 43772 24624
rect 43536 24132 43588 24138
rect 43536 24074 43588 24080
rect 43548 23118 43576 24074
rect 43718 23760 43774 23769
rect 43718 23695 43720 23704
rect 43772 23695 43774 23704
rect 43720 23666 43772 23672
rect 43720 23520 43772 23526
rect 43720 23462 43772 23468
rect 43626 23216 43682 23225
rect 43732 23186 43760 23462
rect 43626 23151 43682 23160
rect 43720 23180 43772 23186
rect 43640 23118 43668 23151
rect 43720 23122 43772 23128
rect 43536 23112 43588 23118
rect 43536 23054 43588 23060
rect 43628 23112 43680 23118
rect 43628 23054 43680 23060
rect 43732 23050 43760 23122
rect 43720 23044 43772 23050
rect 43720 22986 43772 22992
rect 43824 22506 43852 33050
rect 43916 32570 43944 33458
rect 44560 33114 44588 33458
rect 44732 33312 44784 33318
rect 44732 33254 44784 33260
rect 44364 33108 44416 33114
rect 44364 33050 44416 33056
rect 44548 33108 44600 33114
rect 44548 33050 44600 33056
rect 44640 33108 44692 33114
rect 44640 33050 44692 33056
rect 43904 32564 43956 32570
rect 43904 32506 43956 32512
rect 44180 32496 44232 32502
rect 44180 32438 44232 32444
rect 44192 30274 44220 32438
rect 44376 32434 44404 33050
rect 44652 32842 44680 33050
rect 44640 32836 44692 32842
rect 44640 32778 44692 32784
rect 44364 32428 44416 32434
rect 44364 32370 44416 32376
rect 44640 32360 44692 32366
rect 44640 32302 44692 32308
rect 44652 32026 44680 32302
rect 44640 32020 44692 32026
rect 44640 31962 44692 31968
rect 44744 31278 44772 33254
rect 44928 32774 44956 33458
rect 45008 32904 45060 32910
rect 45008 32846 45060 32852
rect 44916 32768 44968 32774
rect 44916 32710 44968 32716
rect 44928 32502 44956 32710
rect 44916 32496 44968 32502
rect 44916 32438 44968 32444
rect 44824 32360 44876 32366
rect 44824 32302 44876 32308
rect 44836 31482 44864 32302
rect 44928 31822 44956 32438
rect 45020 32434 45048 32846
rect 45100 32836 45152 32842
rect 45100 32778 45152 32784
rect 45008 32428 45060 32434
rect 45008 32370 45060 32376
rect 45020 31958 45048 32370
rect 45112 32230 45140 32778
rect 45100 32224 45152 32230
rect 45100 32166 45152 32172
rect 45008 31952 45060 31958
rect 45008 31894 45060 31900
rect 44916 31816 44968 31822
rect 44916 31758 44968 31764
rect 44824 31476 44876 31482
rect 44824 31418 44876 31424
rect 44732 31272 44784 31278
rect 44732 31214 44784 31220
rect 44100 30258 44220 30274
rect 44088 30252 44220 30258
rect 44140 30246 44220 30252
rect 44088 30194 44140 30200
rect 43904 30048 43956 30054
rect 43904 29990 43956 29996
rect 43916 29714 43944 29990
rect 44192 29782 44220 30246
rect 44272 30252 44324 30258
rect 44272 30194 44324 30200
rect 44456 30252 44508 30258
rect 44456 30194 44508 30200
rect 44284 29850 44312 30194
rect 44272 29844 44324 29850
rect 44272 29786 44324 29792
rect 44180 29776 44232 29782
rect 44180 29718 44232 29724
rect 43904 29708 43956 29714
rect 43904 29650 43956 29656
rect 44192 28558 44220 29718
rect 44180 28552 44232 28558
rect 44180 28494 44232 28500
rect 43996 28416 44048 28422
rect 43996 28358 44048 28364
rect 44008 28150 44036 28358
rect 43996 28144 44048 28150
rect 43996 28086 44048 28092
rect 44088 28144 44140 28150
rect 44088 28086 44140 28092
rect 43996 27872 44048 27878
rect 44100 27860 44128 28086
rect 44468 28082 44496 30194
rect 44744 29646 44772 31214
rect 44928 30190 44956 31758
rect 45008 31204 45060 31210
rect 45008 31146 45060 31152
rect 44916 30184 44968 30190
rect 44916 30126 44968 30132
rect 45020 29714 45048 31146
rect 45112 30104 45140 32166
rect 45204 31210 45232 34002
rect 45376 33992 45428 33998
rect 45428 33940 45508 33946
rect 45376 33934 45508 33940
rect 45388 33918 45508 33934
rect 45376 33856 45428 33862
rect 45376 33798 45428 33804
rect 45388 33590 45416 33798
rect 45376 33584 45428 33590
rect 45376 33526 45428 33532
rect 45480 33522 45508 33918
rect 45468 33516 45520 33522
rect 45468 33458 45520 33464
rect 45480 33114 45508 33458
rect 45468 33108 45520 33114
rect 45468 33050 45520 33056
rect 45480 32570 45508 33050
rect 45468 32564 45520 32570
rect 45468 32506 45520 32512
rect 45376 32292 45428 32298
rect 45376 32234 45428 32240
rect 45192 31204 45244 31210
rect 45192 31146 45244 31152
rect 45388 30802 45416 32234
rect 45468 31476 45520 31482
rect 45468 31418 45520 31424
rect 45376 30796 45428 30802
rect 45376 30738 45428 30744
rect 45388 30394 45416 30738
rect 45480 30734 45508 31418
rect 45468 30728 45520 30734
rect 45468 30670 45520 30676
rect 45376 30388 45428 30394
rect 45376 30330 45428 30336
rect 45376 30252 45428 30258
rect 45376 30194 45428 30200
rect 45284 30116 45336 30122
rect 45112 30076 45284 30104
rect 45112 29850 45140 30076
rect 45284 30058 45336 30064
rect 45100 29844 45152 29850
rect 45100 29786 45152 29792
rect 45008 29708 45060 29714
rect 45060 29668 45140 29696
rect 45008 29650 45060 29656
rect 44732 29640 44784 29646
rect 44732 29582 44784 29588
rect 44744 29102 44772 29582
rect 44732 29096 44784 29102
rect 44732 29038 44784 29044
rect 45008 29096 45060 29102
rect 45008 29038 45060 29044
rect 44548 28756 44600 28762
rect 44548 28698 44600 28704
rect 44560 28150 44588 28698
rect 45020 28558 45048 29038
rect 45112 28558 45140 29668
rect 45388 29578 45416 30194
rect 45468 30048 45520 30054
rect 45468 29990 45520 29996
rect 45480 29646 45508 29990
rect 45468 29640 45520 29646
rect 45468 29582 45520 29588
rect 45376 29572 45428 29578
rect 45376 29514 45428 29520
rect 45468 29504 45520 29510
rect 45468 29446 45520 29452
rect 45480 28626 45508 29446
rect 45468 28620 45520 28626
rect 45468 28562 45520 28568
rect 44916 28552 44968 28558
rect 44916 28494 44968 28500
rect 45008 28552 45060 28558
rect 45008 28494 45060 28500
rect 45100 28552 45152 28558
rect 45100 28494 45152 28500
rect 44928 28218 44956 28494
rect 45192 28416 45244 28422
rect 45192 28358 45244 28364
rect 44916 28212 44968 28218
rect 44916 28154 44968 28160
rect 44548 28144 44600 28150
rect 44548 28086 44600 28092
rect 45204 28082 45232 28358
rect 44456 28076 44508 28082
rect 44456 28018 44508 28024
rect 44640 28076 44692 28082
rect 44640 28018 44692 28024
rect 45192 28076 45244 28082
rect 45192 28018 45244 28024
rect 44048 27832 44128 27860
rect 43996 27814 44048 27820
rect 44652 26790 44680 28018
rect 45468 27872 45520 27878
rect 45468 27814 45520 27820
rect 45480 27538 45508 27814
rect 45468 27532 45520 27538
rect 45468 27474 45520 27480
rect 45572 27112 45600 40462
rect 45744 34060 45796 34066
rect 45744 34002 45796 34008
rect 45756 33522 45784 34002
rect 45744 33516 45796 33522
rect 45744 33458 45796 33464
rect 45848 33046 45876 43250
rect 46020 33924 46072 33930
rect 46020 33866 46072 33872
rect 46032 33114 46060 33866
rect 46112 33312 46164 33318
rect 46112 33254 46164 33260
rect 46020 33108 46072 33114
rect 46020 33050 46072 33056
rect 45836 33040 45888 33046
rect 45836 32982 45888 32988
rect 45834 30968 45890 30977
rect 45834 30903 45890 30912
rect 45744 30796 45796 30802
rect 45744 30738 45796 30744
rect 45650 27704 45706 27713
rect 45650 27639 45652 27648
rect 45704 27639 45706 27648
rect 45652 27610 45704 27616
rect 45652 27464 45704 27470
rect 45652 27406 45704 27412
rect 45664 27130 45692 27406
rect 45480 27084 45600 27112
rect 45652 27124 45704 27130
rect 44640 26784 44692 26790
rect 44640 26726 44692 26732
rect 43996 26308 44048 26314
rect 43996 26250 44048 26256
rect 44008 25974 44036 26250
rect 44088 26036 44140 26042
rect 44088 25978 44140 25984
rect 43996 25968 44048 25974
rect 43996 25910 44048 25916
rect 43904 25696 43956 25702
rect 43904 25638 43956 25644
rect 43916 25362 43944 25638
rect 43904 25356 43956 25362
rect 43904 25298 43956 25304
rect 44008 25294 44036 25910
rect 44100 25770 44128 25978
rect 45480 25922 45508 27084
rect 45652 27066 45704 27072
rect 45756 26994 45784 30738
rect 45560 26988 45612 26994
rect 45560 26930 45612 26936
rect 45744 26988 45796 26994
rect 45744 26930 45796 26936
rect 45572 26042 45600 26930
rect 45744 26376 45796 26382
rect 45744 26318 45796 26324
rect 45560 26036 45612 26042
rect 45560 25978 45612 25984
rect 45480 25894 45600 25922
rect 45756 25906 45784 26318
rect 44088 25764 44140 25770
rect 44088 25706 44140 25712
rect 44100 25514 44128 25706
rect 45284 25696 45336 25702
rect 45284 25638 45336 25644
rect 44100 25486 44220 25514
rect 43996 25288 44048 25294
rect 43996 25230 44048 25236
rect 44192 24954 44220 25486
rect 45296 25430 45324 25638
rect 45284 25424 45336 25430
rect 45284 25366 45336 25372
rect 44456 25288 44508 25294
rect 44456 25230 44508 25236
rect 44548 25288 44600 25294
rect 44548 25230 44600 25236
rect 44180 24948 44232 24954
rect 44180 24890 44232 24896
rect 44468 24818 44496 25230
rect 44560 24886 44588 25230
rect 44732 25152 44784 25158
rect 44732 25094 44784 25100
rect 44548 24880 44600 24886
rect 44548 24822 44600 24828
rect 44744 24818 44772 25094
rect 43996 24812 44048 24818
rect 43996 24754 44048 24760
rect 44456 24812 44508 24818
rect 44456 24754 44508 24760
rect 44732 24812 44784 24818
rect 44732 24754 44784 24760
rect 44008 23866 44036 24754
rect 44468 24342 44496 24754
rect 44456 24336 44508 24342
rect 45572 24290 45600 25894
rect 45744 25900 45796 25906
rect 45744 25842 45796 25848
rect 45848 25362 45876 30903
rect 45928 30592 45980 30598
rect 45928 30534 45980 30540
rect 45940 30258 45968 30534
rect 45928 30252 45980 30258
rect 45928 30194 45980 30200
rect 46032 29850 46060 33050
rect 46124 30734 46152 33254
rect 46216 30870 46244 47534
rect 47688 47054 47716 49624
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 46572 46912 46624 46918
rect 46572 46854 46624 46860
rect 46584 43790 46612 46854
rect 46756 45484 46808 45490
rect 46756 45426 46808 45432
rect 46768 44985 46796 45426
rect 46754 44976 46810 44985
rect 46754 44911 46810 44920
rect 46572 43784 46624 43790
rect 46572 43726 46624 43732
rect 46480 43104 46532 43110
rect 46480 43046 46532 43052
rect 46664 43104 46716 43110
rect 46664 43046 46716 43052
rect 46204 30864 46256 30870
rect 46204 30806 46256 30812
rect 46112 30728 46164 30734
rect 46112 30670 46164 30676
rect 46204 30184 46256 30190
rect 46204 30126 46256 30132
rect 46020 29844 46072 29850
rect 46020 29786 46072 29792
rect 46032 29646 46060 29786
rect 46020 29640 46072 29646
rect 46020 29582 46072 29588
rect 46020 28144 46072 28150
rect 46020 28086 46072 28092
rect 46032 26858 46060 28086
rect 46216 27606 46244 30126
rect 46112 27600 46164 27606
rect 46112 27542 46164 27548
rect 46204 27600 46256 27606
rect 46204 27542 46256 27548
rect 46020 26852 46072 26858
rect 46020 26794 46072 26800
rect 46020 26580 46072 26586
rect 46020 26522 46072 26528
rect 46032 25702 46060 26522
rect 46020 25696 46072 25702
rect 46020 25638 46072 25644
rect 45836 25356 45888 25362
rect 45836 25298 45888 25304
rect 45928 25288 45980 25294
rect 45926 25256 45928 25265
rect 45980 25256 45982 25265
rect 45744 25220 45796 25226
rect 45926 25191 45982 25200
rect 45744 25162 45796 25168
rect 45756 24290 45784 25162
rect 44456 24278 44508 24284
rect 44468 23866 44496 24278
rect 45388 24262 45600 24290
rect 45664 24262 45784 24290
rect 45928 24268 45980 24274
rect 44916 24200 44968 24206
rect 44914 24168 44916 24177
rect 45192 24200 45244 24206
rect 44968 24168 44970 24177
rect 45192 24142 45244 24148
rect 44914 24103 44970 24112
rect 43996 23860 44048 23866
rect 43996 23802 44048 23808
rect 44456 23860 44508 23866
rect 44456 23802 44508 23808
rect 44178 23760 44234 23769
rect 44178 23695 44234 23704
rect 44272 23724 44324 23730
rect 44192 23526 44220 23695
rect 44272 23666 44324 23672
rect 44180 23520 44232 23526
rect 44180 23462 44232 23468
rect 44192 23118 44220 23462
rect 44284 23118 44312 23666
rect 44456 23656 44508 23662
rect 44456 23598 44508 23604
rect 44180 23112 44232 23118
rect 44180 23054 44232 23060
rect 44272 23112 44324 23118
rect 44272 23054 44324 23060
rect 44468 22778 44496 23598
rect 44640 23248 44692 23254
rect 44640 23190 44692 23196
rect 44456 22772 44508 22778
rect 44456 22714 44508 22720
rect 43812 22500 43864 22506
rect 43812 22442 43864 22448
rect 43904 21480 43956 21486
rect 43904 21422 43956 21428
rect 43916 21146 43944 21422
rect 43904 21140 43956 21146
rect 43904 21082 43956 21088
rect 44652 21010 44680 23190
rect 44928 23186 44956 24103
rect 45204 23866 45232 24142
rect 45192 23860 45244 23866
rect 45192 23802 45244 23808
rect 44916 23180 44968 23186
rect 44916 23122 44968 23128
rect 45204 23050 45232 23802
rect 45388 23662 45416 24262
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 45468 24132 45520 24138
rect 45468 24074 45520 24080
rect 45480 23798 45508 24074
rect 45468 23792 45520 23798
rect 45468 23734 45520 23740
rect 45376 23656 45428 23662
rect 45572 23644 45600 24142
rect 45664 24138 45692 24262
rect 45928 24210 45980 24216
rect 45940 24138 45968 24210
rect 46020 24200 46072 24206
rect 46018 24168 46020 24177
rect 46072 24168 46074 24177
rect 45652 24132 45704 24138
rect 45652 24074 45704 24080
rect 45928 24132 45980 24138
rect 46018 24103 46074 24112
rect 45928 24074 45980 24080
rect 45664 23798 45692 24074
rect 45652 23792 45704 23798
rect 45652 23734 45704 23740
rect 45940 23730 45968 24074
rect 45928 23724 45980 23730
rect 45928 23666 45980 23672
rect 45744 23656 45796 23662
rect 45572 23616 45744 23644
rect 45376 23598 45428 23604
rect 45744 23598 45796 23604
rect 45756 23050 45784 23598
rect 45940 23118 45968 23666
rect 45928 23112 45980 23118
rect 45928 23054 45980 23060
rect 45192 23044 45244 23050
rect 45192 22986 45244 22992
rect 45744 23044 45796 23050
rect 45744 22986 45796 22992
rect 45744 21344 45796 21350
rect 45744 21286 45796 21292
rect 45756 21010 45784 21286
rect 46020 21140 46072 21146
rect 46020 21082 46072 21088
rect 44640 21004 44692 21010
rect 44640 20946 44692 20952
rect 45744 21004 45796 21010
rect 45744 20946 45796 20952
rect 43628 20868 43680 20874
rect 43628 20810 43680 20816
rect 44548 20868 44600 20874
rect 44548 20810 44600 20816
rect 43444 20596 43496 20602
rect 43444 20538 43496 20544
rect 43536 20460 43588 20466
rect 43536 20402 43588 20408
rect 43548 20058 43576 20402
rect 43536 20052 43588 20058
rect 43536 19994 43588 20000
rect 43352 19848 43404 19854
rect 43352 19790 43404 19796
rect 43364 19378 43392 19790
rect 43352 19372 43404 19378
rect 43352 19314 43404 19320
rect 43168 17128 43220 17134
rect 43168 17070 43220 17076
rect 43536 17128 43588 17134
rect 43536 17070 43588 17076
rect 43352 17060 43404 17066
rect 43352 17002 43404 17008
rect 43364 16658 43392 17002
rect 43352 16652 43404 16658
rect 43352 16594 43404 16600
rect 43076 16584 43128 16590
rect 43076 16526 43128 16532
rect 43548 16522 43576 17070
rect 43536 16516 43588 16522
rect 43536 16458 43588 16464
rect 43260 16448 43312 16454
rect 43640 16402 43668 20810
rect 44560 20602 44588 20810
rect 44548 20596 44600 20602
rect 44548 20538 44600 20544
rect 44560 19854 44588 20538
rect 44652 19854 44680 20946
rect 46032 20890 46060 21082
rect 45560 20868 45612 20874
rect 45560 20810 45612 20816
rect 45940 20862 46060 20890
rect 45284 20392 45336 20398
rect 45284 20334 45336 20340
rect 44548 19848 44600 19854
rect 44548 19790 44600 19796
rect 44640 19848 44692 19854
rect 44640 19790 44692 19796
rect 44180 19712 44232 19718
rect 44180 19654 44232 19660
rect 44364 19712 44416 19718
rect 44364 19654 44416 19660
rect 44192 19514 44220 19654
rect 43812 19508 43864 19514
rect 43812 19450 43864 19456
rect 44180 19508 44232 19514
rect 44180 19450 44232 19456
rect 43824 18290 43852 19450
rect 44272 19372 44324 19378
rect 44272 19314 44324 19320
rect 44284 18834 44312 19314
rect 44376 19310 44404 19654
rect 44364 19304 44416 19310
rect 44364 19246 44416 19252
rect 44272 18828 44324 18834
rect 44272 18770 44324 18776
rect 44560 18766 44588 19790
rect 44548 18760 44600 18766
rect 44548 18702 44600 18708
rect 44652 18698 44680 19790
rect 45296 19310 45324 20334
rect 45572 19854 45600 20810
rect 45940 20058 45968 20862
rect 45928 20052 45980 20058
rect 45928 19994 45980 20000
rect 45560 19848 45612 19854
rect 45560 19790 45612 19796
rect 45284 19304 45336 19310
rect 45284 19246 45336 19252
rect 44732 18760 44784 18766
rect 44732 18702 44784 18708
rect 44272 18692 44324 18698
rect 44272 18634 44324 18640
rect 44640 18692 44692 18698
rect 44640 18634 44692 18640
rect 43812 18284 43864 18290
rect 43812 18226 43864 18232
rect 44180 18284 44232 18290
rect 44180 18226 44232 18232
rect 43812 18080 43864 18086
rect 43812 18022 43864 18028
rect 43824 17610 43852 18022
rect 44088 17808 44140 17814
rect 44088 17750 44140 17756
rect 43812 17604 43864 17610
rect 43812 17546 43864 17552
rect 44100 16998 44128 17750
rect 44192 17678 44220 18226
rect 44180 17672 44232 17678
rect 44180 17614 44232 17620
rect 44088 16992 44140 16998
rect 44088 16934 44140 16940
rect 44100 16726 44128 16934
rect 44088 16720 44140 16726
rect 44088 16662 44140 16668
rect 43812 16584 43864 16590
rect 43812 16526 43864 16532
rect 43260 16390 43312 16396
rect 43272 15026 43300 16390
rect 43548 16374 43668 16402
rect 43260 15020 43312 15026
rect 43260 14962 43312 14968
rect 42984 14816 43036 14822
rect 42984 14758 43036 14764
rect 42996 14074 43024 14758
rect 43076 14272 43128 14278
rect 43076 14214 43128 14220
rect 42984 14068 43036 14074
rect 42984 14010 43036 14016
rect 43088 13938 43116 14214
rect 43076 13932 43128 13938
rect 43076 13874 43128 13880
rect 43168 13864 43220 13870
rect 42904 13790 43116 13818
rect 43168 13806 43220 13812
rect 42800 13728 42852 13734
rect 42800 13670 42852 13676
rect 42812 12782 42840 13670
rect 43088 13190 43116 13790
rect 43076 13184 43128 13190
rect 43076 13126 43128 13132
rect 43180 12986 43208 13806
rect 43260 13728 43312 13734
rect 43260 13670 43312 13676
rect 43272 13326 43300 13670
rect 43260 13320 43312 13326
rect 43260 13262 43312 13268
rect 43260 13184 43312 13190
rect 43260 13126 43312 13132
rect 43168 12980 43220 12986
rect 43168 12922 43220 12928
rect 42800 12776 42852 12782
rect 42800 12718 42852 12724
rect 43076 12776 43128 12782
rect 43076 12718 43128 12724
rect 43168 12776 43220 12782
rect 43168 12718 43220 12724
rect 43088 12442 43116 12718
rect 43076 12436 43128 12442
rect 43076 12378 43128 12384
rect 42708 12232 42760 12238
rect 42706 12200 42708 12209
rect 42760 12200 42762 12209
rect 43180 12170 43208 12718
rect 43272 12170 43300 13126
rect 43548 12646 43576 16374
rect 43824 16250 43852 16526
rect 43812 16244 43864 16250
rect 43812 16186 43864 16192
rect 43720 15904 43772 15910
rect 43720 15846 43772 15852
rect 43732 15026 43760 15846
rect 44284 15094 44312 18634
rect 44744 18426 44772 18702
rect 44824 18624 44876 18630
rect 44824 18566 44876 18572
rect 44732 18420 44784 18426
rect 44732 18362 44784 18368
rect 44836 18222 44864 18566
rect 45008 18284 45060 18290
rect 44928 18244 45008 18272
rect 44364 18216 44416 18222
rect 44364 18158 44416 18164
rect 44824 18216 44876 18222
rect 44824 18158 44876 18164
rect 44376 17678 44404 18158
rect 44364 17672 44416 17678
rect 44364 17614 44416 17620
rect 44548 17672 44600 17678
rect 44548 17614 44600 17620
rect 44560 17338 44588 17614
rect 44548 17332 44600 17338
rect 44548 17274 44600 17280
rect 44836 17270 44864 18158
rect 44824 17264 44876 17270
rect 44824 17206 44876 17212
rect 44364 17196 44416 17202
rect 44364 17138 44416 17144
rect 44732 17196 44784 17202
rect 44732 17138 44784 17144
rect 44376 16522 44404 17138
rect 44744 16794 44772 17138
rect 44928 17066 44956 18244
rect 45008 18226 45060 18232
rect 45572 17678 45600 19790
rect 45836 18624 45888 18630
rect 45836 18566 45888 18572
rect 45848 18290 45876 18566
rect 45836 18284 45888 18290
rect 45836 18226 45888 18232
rect 45836 17876 45888 17882
rect 45940 17864 45968 19994
rect 46124 18850 46152 27542
rect 46204 27464 46256 27470
rect 46204 27406 46256 27412
rect 46216 26586 46244 27406
rect 46204 26580 46256 26586
rect 46204 26522 46256 26528
rect 46204 25900 46256 25906
rect 46204 25842 46256 25848
rect 46216 20942 46244 25842
rect 46296 25696 46348 25702
rect 46296 25638 46348 25644
rect 46308 21146 46336 25638
rect 46388 24812 46440 24818
rect 46388 24754 46440 24760
rect 46400 23594 46428 24754
rect 46388 23588 46440 23594
rect 46388 23530 46440 23536
rect 46400 23254 46428 23530
rect 46388 23248 46440 23254
rect 46388 23190 46440 23196
rect 46296 21140 46348 21146
rect 46296 21082 46348 21088
rect 46204 20936 46256 20942
rect 46204 20878 46256 20884
rect 46492 20466 46520 43046
rect 46676 42945 46704 43046
rect 46662 42936 46718 42945
rect 46662 42871 46718 42880
rect 46664 40384 46716 40390
rect 46664 40326 46716 40332
rect 46676 40225 46704 40326
rect 46662 40216 46718 40225
rect 46662 40151 46718 40160
rect 46664 37664 46716 37670
rect 46664 37606 46716 37612
rect 46676 37505 46704 37606
rect 46662 37496 46718 37505
rect 46662 37431 46718 37440
rect 46848 36576 46900 36582
rect 46848 36518 46900 36524
rect 46860 35894 46888 36518
rect 46860 35866 46980 35894
rect 46848 35692 46900 35698
rect 46848 35634 46900 35640
rect 46664 35488 46716 35494
rect 46662 35456 46664 35465
rect 46716 35456 46718 35465
rect 46662 35391 46718 35400
rect 46664 32768 46716 32774
rect 46662 32736 46664 32745
rect 46716 32736 46718 32745
rect 46662 32671 46718 32680
rect 46662 30016 46718 30025
rect 46662 29951 46718 29960
rect 46676 29306 46704 29951
rect 46664 29300 46716 29306
rect 46664 29242 46716 29248
rect 46662 28520 46718 28529
rect 46662 28455 46718 28464
rect 46676 28218 46704 28455
rect 46664 28212 46716 28218
rect 46664 28154 46716 28160
rect 46572 28076 46624 28082
rect 46572 28018 46624 28024
rect 46584 27985 46612 28018
rect 46570 27976 46626 27985
rect 46570 27911 46626 27920
rect 46756 26988 46808 26994
rect 46756 26930 46808 26936
rect 46768 26586 46796 26930
rect 46756 26580 46808 26586
rect 46756 26522 46808 26528
rect 46572 24608 46624 24614
rect 46572 24550 46624 24556
rect 46584 24206 46612 24550
rect 46664 24268 46716 24274
rect 46664 24210 46716 24216
rect 46572 24200 46624 24206
rect 46572 24142 46624 24148
rect 46676 23866 46704 24210
rect 46664 23860 46716 23866
rect 46664 23802 46716 23808
rect 46570 23216 46626 23225
rect 46570 23151 46626 23160
rect 46584 23118 46612 23151
rect 46572 23112 46624 23118
rect 46572 23054 46624 23060
rect 46756 21548 46808 21554
rect 46756 21490 46808 21496
rect 46768 21146 46796 21490
rect 46756 21140 46808 21146
rect 46756 21082 46808 21088
rect 46664 20596 46716 20602
rect 46664 20538 46716 20544
rect 46676 20505 46704 20538
rect 46662 20496 46718 20505
rect 46204 20460 46256 20466
rect 46204 20402 46256 20408
rect 46480 20460 46532 20466
rect 46662 20431 46718 20440
rect 46480 20402 46532 20408
rect 46216 20058 46244 20402
rect 46204 20052 46256 20058
rect 46204 19994 46256 20000
rect 46124 18822 46244 18850
rect 46112 18760 46164 18766
rect 46112 18702 46164 18708
rect 46124 17882 46152 18702
rect 45888 17836 45968 17864
rect 46112 17876 46164 17882
rect 45836 17818 45888 17824
rect 46112 17818 46164 17824
rect 45560 17672 45612 17678
rect 45560 17614 45612 17620
rect 45008 17536 45060 17542
rect 45008 17478 45060 17484
rect 44916 17060 44968 17066
rect 44916 17002 44968 17008
rect 44732 16788 44784 16794
rect 44732 16730 44784 16736
rect 44824 16788 44876 16794
rect 44824 16730 44876 16736
rect 44836 16674 44864 16730
rect 44744 16646 44864 16674
rect 44916 16720 44968 16726
rect 44916 16662 44968 16668
rect 44364 16516 44416 16522
rect 44364 16458 44416 16464
rect 44272 15088 44324 15094
rect 44272 15030 44324 15036
rect 43720 15020 43772 15026
rect 43720 14962 43772 14968
rect 43628 14884 43680 14890
rect 43628 14826 43680 14832
rect 43536 12640 43588 12646
rect 43536 12582 43588 12588
rect 43352 12300 43404 12306
rect 43352 12242 43404 12248
rect 42706 12135 42762 12144
rect 43168 12164 43220 12170
rect 43168 12106 43220 12112
rect 43260 12164 43312 12170
rect 43260 12106 43312 12112
rect 43180 11898 43208 12106
rect 43168 11892 43220 11898
rect 43168 11834 43220 11840
rect 43074 11792 43130 11801
rect 43074 11727 43130 11736
rect 43168 11756 43220 11762
rect 42984 11688 43036 11694
rect 42984 11630 43036 11636
rect 42708 11552 42760 11558
rect 42708 11494 42760 11500
rect 42616 11144 42668 11150
rect 42614 11112 42616 11121
rect 42720 11132 42748 11494
rect 42800 11144 42852 11150
rect 42668 11112 42670 11121
rect 42720 11104 42800 11132
rect 42800 11086 42852 11092
rect 42890 11112 42946 11121
rect 42614 11047 42670 11056
rect 42890 11047 42946 11056
rect 41052 10804 41104 10810
rect 41052 10746 41104 10752
rect 42432 10804 42484 10810
rect 42432 10746 42484 10752
rect 40828 10628 40908 10656
rect 40776 10610 40828 10616
rect 40880 10130 40908 10628
rect 40868 10124 40920 10130
rect 40868 10066 40920 10072
rect 40880 9674 40908 10066
rect 41064 10062 41092 10746
rect 42444 10062 42472 10746
rect 42904 10674 42932 11047
rect 42996 10724 43024 11630
rect 43088 11558 43116 11727
rect 43168 11698 43220 11704
rect 43076 11552 43128 11558
rect 43076 11494 43128 11500
rect 43180 11150 43208 11698
rect 43260 11688 43312 11694
rect 43258 11656 43260 11665
rect 43312 11656 43314 11665
rect 43364 11626 43392 12242
rect 43640 12238 43668 14826
rect 43732 14482 43760 14962
rect 43720 14476 43772 14482
rect 43720 14418 43772 14424
rect 44180 14272 44232 14278
rect 44180 14214 44232 14220
rect 44192 13938 44220 14214
rect 44180 13932 44232 13938
rect 44180 13874 44232 13880
rect 43720 13456 43772 13462
rect 43720 13398 43772 13404
rect 43628 12232 43680 12238
rect 43626 12200 43628 12209
rect 43680 12200 43682 12209
rect 43626 12135 43682 12144
rect 43536 12096 43588 12102
rect 43536 12038 43588 12044
rect 43548 11762 43576 12038
rect 43640 11762 43668 12135
rect 43536 11756 43588 11762
rect 43536 11698 43588 11704
rect 43628 11756 43680 11762
rect 43628 11698 43680 11704
rect 43444 11688 43496 11694
rect 43444 11630 43496 11636
rect 43258 11591 43314 11600
rect 43352 11620 43404 11626
rect 43352 11562 43404 11568
rect 43364 11234 43392 11562
rect 43456 11354 43484 11630
rect 43444 11348 43496 11354
rect 43444 11290 43496 11296
rect 43364 11206 43484 11234
rect 43168 11144 43220 11150
rect 43220 11092 43300 11098
rect 43168 11086 43300 11092
rect 43180 11070 43300 11086
rect 43168 11008 43220 11014
rect 43168 10950 43220 10956
rect 43076 10736 43128 10742
rect 42996 10696 43076 10724
rect 42892 10668 42944 10674
rect 42892 10610 42944 10616
rect 42996 10062 43024 10696
rect 43076 10678 43128 10684
rect 43076 10192 43128 10198
rect 43076 10134 43128 10140
rect 41052 10056 41104 10062
rect 41052 9998 41104 10004
rect 42432 10056 42484 10062
rect 42432 9998 42484 10004
rect 42984 10056 43036 10062
rect 42984 9998 43036 10004
rect 40788 9646 40908 9674
rect 41064 9654 41092 9998
rect 42800 9988 42852 9994
rect 42800 9930 42852 9936
rect 41052 9648 41104 9654
rect 40316 9580 40368 9586
rect 40316 9522 40368 9528
rect 40684 9580 40736 9586
rect 40684 9522 40736 9528
rect 40788 9518 40816 9646
rect 41052 9590 41104 9596
rect 40776 9512 40828 9518
rect 40776 9454 40828 9460
rect 40788 9178 40816 9454
rect 41064 9450 41092 9590
rect 41144 9580 41196 9586
rect 41144 9522 41196 9528
rect 41052 9444 41104 9450
rect 41052 9386 41104 9392
rect 41156 9330 41184 9522
rect 42708 9444 42760 9450
rect 42708 9386 42760 9392
rect 41420 9376 41472 9382
rect 41156 9324 41420 9330
rect 41156 9318 41472 9324
rect 41156 9302 41460 9318
rect 40776 9172 40828 9178
rect 40776 9114 40828 9120
rect 42720 8974 42748 9386
rect 42812 9178 42840 9930
rect 42892 9580 42944 9586
rect 42892 9522 42944 9528
rect 42800 9172 42852 9178
rect 42800 9114 42852 9120
rect 42904 8974 42932 9522
rect 43088 9518 43116 10134
rect 43180 9926 43208 10950
rect 43168 9920 43220 9926
rect 43168 9862 43220 9868
rect 43180 9586 43208 9862
rect 43168 9580 43220 9586
rect 43168 9522 43220 9528
rect 43272 9518 43300 11070
rect 43352 11076 43404 11082
rect 43352 11018 43404 11024
rect 43364 10810 43392 11018
rect 43352 10804 43404 10810
rect 43352 10746 43404 10752
rect 43364 10470 43392 10746
rect 43456 10742 43484 11206
rect 43628 11212 43680 11218
rect 43628 11154 43680 11160
rect 43536 11144 43588 11150
rect 43534 11112 43536 11121
rect 43588 11112 43590 11121
rect 43534 11047 43590 11056
rect 43640 11014 43668 11154
rect 43628 11008 43680 11014
rect 43628 10950 43680 10956
rect 43640 10810 43668 10950
rect 43628 10804 43680 10810
rect 43628 10746 43680 10752
rect 43444 10736 43496 10742
rect 43444 10678 43496 10684
rect 43352 10464 43404 10470
rect 43352 10406 43404 10412
rect 43352 9648 43404 9654
rect 43456 9636 43484 10678
rect 43732 10130 43760 13398
rect 44088 12640 44140 12646
rect 44088 12582 44140 12588
rect 44100 12374 44128 12582
rect 44088 12368 44140 12374
rect 44088 12310 44140 12316
rect 43812 12232 43864 12238
rect 43812 12174 43864 12180
rect 43996 12232 44048 12238
rect 43996 12174 44048 12180
rect 44180 12232 44232 12238
rect 44180 12174 44232 12180
rect 43824 11642 43852 12174
rect 44008 11830 44036 12174
rect 43996 11824 44048 11830
rect 43996 11766 44048 11772
rect 43996 11688 44048 11694
rect 43824 11636 43996 11642
rect 43824 11630 44048 11636
rect 43824 11614 44036 11630
rect 44008 11286 44036 11614
rect 43996 11280 44048 11286
rect 43996 11222 44048 11228
rect 44192 10674 44220 12174
rect 44180 10668 44232 10674
rect 44180 10610 44232 10616
rect 43720 10124 43772 10130
rect 43720 10066 43772 10072
rect 44192 10062 44220 10610
rect 44180 10056 44232 10062
rect 44180 9998 44232 10004
rect 43404 9608 43484 9636
rect 43352 9590 43404 9596
rect 43076 9512 43128 9518
rect 43076 9454 43128 9460
rect 43260 9512 43312 9518
rect 43260 9454 43312 9460
rect 43272 8974 43300 9454
rect 42708 8968 42760 8974
rect 42708 8910 42760 8916
rect 42892 8968 42944 8974
rect 42892 8910 42944 8916
rect 43260 8968 43312 8974
rect 43260 8910 43312 8916
rect 40224 8492 40276 8498
rect 40224 8434 40276 8440
rect 38660 8084 38712 8090
rect 38660 8026 38712 8032
rect 38016 7880 38068 7886
rect 38016 7822 38068 7828
rect 38752 7880 38804 7886
rect 38752 7822 38804 7828
rect 38292 4616 38344 4622
rect 38292 4558 38344 4564
rect 38304 4214 38332 4558
rect 38292 4208 38344 4214
rect 38292 4150 38344 4156
rect 38764 2650 38792 7822
rect 44376 5710 44404 16458
rect 44744 16454 44772 16646
rect 44732 16448 44784 16454
rect 44732 16390 44784 16396
rect 44824 16448 44876 16454
rect 44824 16390 44876 16396
rect 44744 16114 44772 16390
rect 44732 16108 44784 16114
rect 44732 16050 44784 16056
rect 44836 16046 44864 16390
rect 44824 16040 44876 16046
rect 44824 15982 44876 15988
rect 44928 15978 44956 16662
rect 45020 16590 45048 17478
rect 45100 16992 45152 16998
rect 45100 16934 45152 16940
rect 45008 16584 45060 16590
rect 45008 16526 45060 16532
rect 45112 16046 45140 16934
rect 45376 16652 45428 16658
rect 45376 16594 45428 16600
rect 45388 16250 45416 16594
rect 45376 16244 45428 16250
rect 45376 16186 45428 16192
rect 45100 16040 45152 16046
rect 45100 15982 45152 15988
rect 45468 16040 45520 16046
rect 45468 15982 45520 15988
rect 44916 15972 44968 15978
rect 44916 15914 44968 15920
rect 45192 15496 45244 15502
rect 45192 15438 45244 15444
rect 45204 15162 45232 15438
rect 45192 15156 45244 15162
rect 45192 15098 45244 15104
rect 45204 15026 45232 15098
rect 45192 15020 45244 15026
rect 45192 14962 45244 14968
rect 45204 14414 45232 14962
rect 45480 14822 45508 15982
rect 45572 15570 45600 17614
rect 45744 16516 45796 16522
rect 45744 16458 45796 16464
rect 45756 15706 45784 16458
rect 45848 16114 45876 17818
rect 45836 16108 45888 16114
rect 45836 16050 45888 16056
rect 45744 15700 45796 15706
rect 45744 15642 45796 15648
rect 45560 15564 45612 15570
rect 45560 15506 45612 15512
rect 45468 14816 45520 14822
rect 45388 14776 45468 14804
rect 45388 14618 45416 14776
rect 45468 14758 45520 14764
rect 45376 14612 45428 14618
rect 45376 14554 45428 14560
rect 45192 14408 45244 14414
rect 45192 14350 45244 14356
rect 45204 13938 45232 14350
rect 45192 13932 45244 13938
rect 45192 13874 45244 13880
rect 45388 13734 45416 14554
rect 45376 13728 45428 13734
rect 45376 13670 45428 13676
rect 45468 13728 45520 13734
rect 45468 13670 45520 13676
rect 45480 13326 45508 13670
rect 46112 13524 46164 13530
rect 46112 13466 46164 13472
rect 45468 13320 45520 13326
rect 45468 13262 45520 13268
rect 45100 13184 45152 13190
rect 45100 13126 45152 13132
rect 45112 12850 45140 13126
rect 45100 12844 45152 12850
rect 45100 12786 45152 12792
rect 44916 12776 44968 12782
rect 44916 12718 44968 12724
rect 44548 12640 44600 12646
rect 44548 12582 44600 12588
rect 44560 12238 44588 12582
rect 44548 12232 44600 12238
rect 44548 12174 44600 12180
rect 44928 11694 44956 12718
rect 44916 11688 44968 11694
rect 44916 11630 44968 11636
rect 46124 8498 46152 13466
rect 46216 13326 46244 18822
rect 46386 17776 46442 17785
rect 46386 17711 46442 17720
rect 46754 17776 46810 17785
rect 46754 17711 46810 17720
rect 46400 17678 46428 17711
rect 46768 17678 46796 17711
rect 46388 17672 46440 17678
rect 46388 17614 46440 17620
rect 46756 17672 46808 17678
rect 46756 17614 46808 17620
rect 46480 16108 46532 16114
rect 46480 16050 46532 16056
rect 46492 15638 46520 16050
rect 46664 15904 46716 15910
rect 46664 15846 46716 15852
rect 46676 15745 46704 15846
rect 46662 15736 46718 15745
rect 46662 15671 46718 15680
rect 46480 15632 46532 15638
rect 46480 15574 46532 15580
rect 46388 15496 46440 15502
rect 46388 15438 46440 15444
rect 46400 15162 46428 15438
rect 46388 15156 46440 15162
rect 46388 15098 46440 15104
rect 46860 13870 46888 35634
rect 46952 23254 46980 35866
rect 46940 23248 46992 23254
rect 46940 23190 46992 23196
rect 46848 13864 46900 13870
rect 46848 13806 46900 13812
rect 46204 13320 46256 13326
rect 46204 13262 46256 13268
rect 46664 13184 46716 13190
rect 46664 13126 46716 13132
rect 46676 13025 46704 13126
rect 46662 13016 46718 13025
rect 46662 12951 46718 12960
rect 46480 10668 46532 10674
rect 46480 10610 46532 10616
rect 46492 9722 46520 10610
rect 46664 10464 46716 10470
rect 46664 10406 46716 10412
rect 46676 10305 46704 10406
rect 46662 10296 46718 10305
rect 46662 10231 46718 10240
rect 46480 9716 46532 9722
rect 46480 9658 46532 9664
rect 46112 8492 46164 8498
rect 46112 8434 46164 8440
rect 45928 8424 45980 8430
rect 45928 8366 45980 8372
rect 45940 8265 45968 8366
rect 45926 8256 45982 8265
rect 45926 8191 45982 8200
rect 45558 6216 45614 6225
rect 45558 6151 45614 6160
rect 44364 5704 44416 5710
rect 44364 5646 44416 5652
rect 39210 4040 39266 4049
rect 39210 3975 39212 3984
rect 39264 3975 39266 3984
rect 44548 4004 44600 4010
rect 39212 3946 39264 3952
rect 44548 3946 44600 3952
rect 42706 2680 42762 2689
rect 38752 2644 38804 2650
rect 42706 2615 42762 2624
rect 38752 2586 38804 2592
rect 37648 2576 37700 2582
rect 37648 2518 37700 2524
rect 42720 2514 42748 2615
rect 42708 2508 42760 2514
rect 42708 2450 42760 2456
rect 44560 2446 44588 3946
rect 45572 3194 45600 6151
rect 46664 5568 46716 5574
rect 46662 5536 46664 5545
rect 46716 5536 46718 5545
rect 46662 5471 46718 5480
rect 45560 3188 45612 3194
rect 45560 3130 45612 3136
rect 46572 3052 46624 3058
rect 46572 2994 46624 3000
rect 46584 2825 46612 2994
rect 46570 2816 46626 2825
rect 46570 2751 46626 2760
rect 46202 2544 46258 2553
rect 45468 2508 45520 2514
rect 46202 2479 46204 2488
rect 45468 2450 45520 2456
rect 46256 2479 46258 2488
rect 46204 2450 46256 2456
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 34888 2440 34940 2446
rect 34888 2382 34940 2388
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 39304 2440 39356 2446
rect 39304 2382 39356 2388
rect 41880 2440 41932 2446
rect 41880 2382 41932 2388
rect 44548 2440 44600 2446
rect 44548 2382 44600 2388
rect 34612 2372 34664 2378
rect 34612 2314 34664 2320
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 29184 2304 29236 2310
rect 29184 2246 29236 2252
rect 30380 2304 30432 2310
rect 30380 2246 30432 2252
rect 32220 2304 32272 2310
rect 32220 2246 32272 2252
rect 33416 2304 33468 2310
rect 33416 2246 33468 2252
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 27724 800 27752 2246
rect 30392 1442 30420 2246
rect 30300 1414 30420 1442
rect 30300 800 30328 1414
rect 32232 800 32260 2246
rect 34808 800 34836 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 37384 800 37412 2246
rect 39316 800 39344 2382
rect 41892 800 41920 2382
rect 44456 2304 44508 2310
rect 44456 2246 44508 2252
rect 44468 800 44496 2246
rect 18 0 74 800
rect 1950 0 2006 800
rect 4526 0 4582 800
rect 6458 0 6514 800
rect 9034 0 9090 800
rect 11610 0 11666 800
rect 13542 0 13598 800
rect 16118 0 16174 800
rect 18694 0 18750 800
rect 20626 0 20682 800
rect 23202 0 23258 800
rect 25134 0 25190 800
rect 27710 0 27766 800
rect 30286 0 30342 800
rect 32218 0 32274 800
rect 34794 0 34850 800
rect 37370 0 37426 800
rect 39302 0 39358 800
rect 41878 0 41934 800
rect 44454 0 44510 800
rect 45480 785 45508 2450
rect 45650 2408 45706 2417
rect 45650 2343 45706 2352
rect 46388 2372 46440 2378
rect 45664 2310 45692 2343
rect 46388 2314 46440 2320
rect 45652 2304 45704 2310
rect 45652 2246 45704 2252
rect 46400 800 46428 2314
rect 45466 776 45522 785
rect 45466 711 45522 720
rect 46386 0 46442 800
<< via2 >>
rect 1122 46960 1178 47016
rect 1766 49000 1822 49056
rect 4880 47898 4936 47900
rect 4960 47898 5016 47900
rect 5040 47898 5096 47900
rect 5120 47898 5176 47900
rect 4880 47846 4926 47898
rect 4926 47846 4936 47898
rect 4960 47846 4990 47898
rect 4990 47846 5002 47898
rect 5002 47846 5016 47898
rect 5040 47846 5054 47898
rect 5054 47846 5066 47898
rect 5066 47846 5096 47898
rect 5120 47846 5130 47898
rect 5130 47846 5176 47898
rect 4880 47844 4936 47846
rect 4960 47844 5016 47846
rect 5040 47844 5096 47846
rect 5120 47844 5176 47846
rect 938 44260 994 44296
rect 938 44240 940 44260
rect 940 44240 992 44260
rect 992 44240 994 44260
rect 938 41520 994 41576
rect 938 39480 994 39536
rect 938 36760 994 36816
rect 938 32000 994 32056
rect 938 29280 994 29336
rect 938 26560 994 26616
rect 1582 34040 1638 34096
rect 1674 31884 1730 31920
rect 1674 31864 1676 31884
rect 1676 31864 1728 31884
rect 1728 31864 1730 31884
rect 1674 29708 1730 29744
rect 1674 29688 1676 29708
rect 1676 29688 1728 29708
rect 1728 29688 1730 29708
rect 1398 24656 1454 24712
rect 938 24520 994 24576
rect 938 21800 994 21856
rect 1306 19760 1362 19816
rect 938 17040 994 17096
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 1582 17176 1638 17232
rect 938 14320 994 14376
rect 1674 12724 1676 12744
rect 1676 12724 1728 12744
rect 1728 12724 1730 12744
rect 1674 12688 1730 12724
rect 1490 12280 1546 12336
rect 2226 9988 2282 10024
rect 2226 9968 2228 9988
rect 2228 9968 2280 9988
rect 2280 9968 2282 9988
rect 1582 9560 1638 9616
rect 1582 6840 1638 6896
rect 938 4800 994 4856
rect 2226 2916 2282 2952
rect 2226 2896 2228 2916
rect 2228 2896 2280 2916
rect 2280 2896 2282 2916
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 3238 25200 3294 25256
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 6090 35148 6146 35184
rect 6090 35128 6092 35148
rect 6092 35128 6144 35148
rect 6144 35128 6146 35148
rect 10230 41112 10286 41168
rect 5446 31728 5502 31784
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4710 26560 4766 26616
rect 4710 26444 4766 26480
rect 4710 26424 4712 26444
rect 4712 26424 4764 26444
rect 4764 26424 4766 26444
rect 4526 25880 4582 25936
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 3790 23568 3846 23624
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4526 22616 4582 22672
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 3054 18128 3110 18184
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4894 25900 4950 25936
rect 4894 25880 4896 25900
rect 4896 25880 4948 25900
rect 4948 25880 4950 25900
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 5262 23604 5264 23624
rect 5264 23604 5316 23624
rect 5316 23604 5318 23624
rect 5262 23568 5318 23604
rect 5170 23432 5226 23488
rect 5446 23296 5502 23352
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 5446 22888 5502 22944
rect 5262 22616 5318 22672
rect 5722 23160 5778 23216
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 5170 20032 5226 20088
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4250 17584 4306 17640
rect 5170 17584 5226 17640
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 6826 26308 6882 26344
rect 6826 26288 6828 26308
rect 6828 26288 6880 26308
rect 6880 26288 6882 26308
rect 6182 23604 6184 23624
rect 6184 23604 6236 23624
rect 6236 23604 6238 23624
rect 6182 23568 6238 23604
rect 6090 23296 6146 23352
rect 9586 37576 9642 37632
rect 9402 28484 9458 28520
rect 9402 28464 9404 28484
rect 9404 28464 9456 28484
rect 9456 28464 9458 28484
rect 11058 37612 11060 37632
rect 11060 37612 11112 37632
rect 11112 37612 11114 37632
rect 11058 37576 11114 37612
rect 10782 33904 10838 33960
rect 9678 26560 9734 26616
rect 9586 26424 9642 26480
rect 10874 31728 10930 31784
rect 11058 28364 11060 28384
rect 11060 28364 11112 28384
rect 11112 28364 11114 28384
rect 11058 28328 11114 28364
rect 8206 12588 8208 12608
rect 8208 12588 8260 12608
rect 8260 12588 8262 12608
rect 8206 12552 8262 12588
rect 9402 23432 9458 23488
rect 10138 21936 10194 21992
rect 10506 21664 10562 21720
rect 10690 21972 10692 21992
rect 10692 21972 10744 21992
rect 10744 21972 10746 21992
rect 10690 21936 10746 21972
rect 10506 19896 10562 19952
rect 11150 23296 11206 23352
rect 12254 26188 12256 26208
rect 12256 26188 12308 26208
rect 12308 26188 12310 26208
rect 12254 26152 12310 26188
rect 11794 21936 11850 21992
rect 12530 31184 12586 31240
rect 12714 26152 12770 26208
rect 14462 36796 14464 36816
rect 14464 36796 14516 36816
rect 14516 36796 14518 36816
rect 14462 36760 14518 36796
rect 12714 25472 12770 25528
rect 11058 17856 11114 17912
rect 12070 16088 12126 16144
rect 14094 35012 14150 35048
rect 14094 34992 14096 35012
rect 14096 34992 14148 35012
rect 14148 34992 14150 35012
rect 15290 35400 15346 35456
rect 13542 30368 13598 30424
rect 13266 29280 13322 29336
rect 13174 23160 13230 23216
rect 9402 2624 9458 2680
rect 13358 9696 13414 9752
rect 14278 28600 14334 28656
rect 13818 26560 13874 26616
rect 14554 27240 14610 27296
rect 14094 17720 14150 17776
rect 15382 32272 15438 32328
rect 16210 37848 16266 37904
rect 15474 29008 15530 29064
rect 14922 27240 14978 27296
rect 16762 36796 16764 36816
rect 16764 36796 16816 36816
rect 16816 36796 16818 36816
rect 16762 36760 16818 36796
rect 16394 32272 16450 32328
rect 15474 27956 15476 27976
rect 15476 27956 15528 27976
rect 15528 27956 15530 27976
rect 15474 27920 15530 27956
rect 15106 26424 15162 26480
rect 15750 26968 15806 27024
rect 14462 16108 14518 16144
rect 14462 16088 14464 16108
rect 14464 16088 14516 16108
rect 14516 16088 14518 16108
rect 15750 21428 15752 21448
rect 15752 21428 15804 21448
rect 15804 21428 15806 21448
rect 15750 21392 15806 21428
rect 16118 17992 16174 18048
rect 15474 17620 15476 17640
rect 15476 17620 15528 17640
rect 15528 17620 15530 17640
rect 15474 17584 15530 17620
rect 15198 9016 15254 9072
rect 15750 8880 15806 8936
rect 16946 32972 17002 33008
rect 16946 32952 16948 32972
rect 16948 32952 17000 32972
rect 17000 32952 17002 32972
rect 17682 37984 17738 38040
rect 17866 38256 17922 38312
rect 19062 43732 19064 43752
rect 19064 43732 19116 43752
rect 19116 43732 19118 43752
rect 19062 43696 19118 43732
rect 17866 32816 17922 32872
rect 18142 32272 18198 32328
rect 17958 30932 18014 30968
rect 17958 30912 17960 30932
rect 17960 30912 18012 30932
rect 18012 30912 18014 30932
rect 18234 31728 18290 31784
rect 18970 37984 19026 38040
rect 18510 32952 18566 33008
rect 19154 35808 19210 35864
rect 19154 35572 19156 35592
rect 19156 35572 19208 35592
rect 19208 35572 19210 35592
rect 19154 35536 19210 35572
rect 18878 32544 18934 32600
rect 18694 32000 18750 32056
rect 18326 29280 18382 29336
rect 17314 25472 17370 25528
rect 17498 24248 17554 24304
rect 18050 23160 18106 23216
rect 17130 19896 17186 19952
rect 17038 17856 17094 17912
rect 17038 17604 17094 17640
rect 17038 17584 17040 17604
rect 17040 17584 17092 17604
rect 17092 17584 17094 17604
rect 19246 32000 19302 32056
rect 18234 26832 18290 26888
rect 18326 21548 18382 21584
rect 18326 21528 18328 21548
rect 18328 21528 18380 21548
rect 18380 21528 18382 21548
rect 18234 17720 18290 17776
rect 17866 8200 17922 8256
rect 18786 27104 18842 27160
rect 19522 35944 19578 36000
rect 20626 40024 20682 40080
rect 20166 35128 20222 35184
rect 20442 35148 20498 35184
rect 20442 35128 20444 35148
rect 20444 35128 20496 35148
rect 20496 35128 20498 35148
rect 19798 32852 19800 32872
rect 19800 32852 19852 32872
rect 19852 32852 19854 32872
rect 19798 32816 19854 32852
rect 19706 32408 19762 32464
rect 19430 30096 19486 30152
rect 19338 29996 19340 30016
rect 19340 29996 19392 30016
rect 19392 29996 19394 30016
rect 19338 29960 19394 29996
rect 19338 29824 19394 29880
rect 19154 27240 19210 27296
rect 18786 24112 18842 24168
rect 18786 23316 18842 23352
rect 18786 23296 18788 23316
rect 18788 23296 18840 23316
rect 18840 23296 18842 23316
rect 19154 26968 19210 27024
rect 19062 24248 19118 24304
rect 19062 21548 19118 21584
rect 19062 21528 19064 21548
rect 19064 21528 19116 21548
rect 19116 21528 19118 21548
rect 20166 32136 20222 32192
rect 20166 31592 20222 31648
rect 20258 31456 20314 31512
rect 19890 29960 19946 30016
rect 20442 31456 20498 31512
rect 20442 31356 20444 31376
rect 20444 31356 20496 31376
rect 20496 31356 20498 31376
rect 20442 31320 20498 31356
rect 20902 32272 20958 32328
rect 20534 30096 20590 30152
rect 19982 28056 20038 28112
rect 19890 27820 19892 27840
rect 19892 27820 19944 27840
rect 19944 27820 19946 27840
rect 19890 27784 19946 27820
rect 19706 23976 19762 24032
rect 19706 23704 19762 23760
rect 19614 21800 19670 21856
rect 19614 20712 19670 20768
rect 20350 26460 20352 26480
rect 20352 26460 20404 26480
rect 20404 26460 20406 26480
rect 20350 26424 20406 26460
rect 22466 40432 22522 40488
rect 22466 38256 22522 38312
rect 21546 33924 21602 33960
rect 21546 33904 21548 33924
rect 21548 33904 21600 33924
rect 21600 33904 21602 33924
rect 21546 32564 21602 32600
rect 21546 32544 21548 32564
rect 21548 32544 21600 32564
rect 21600 32544 21602 32564
rect 21914 35264 21970 35320
rect 21178 31628 21180 31648
rect 21180 31628 21232 31648
rect 21232 31628 21234 31648
rect 21178 31592 21234 31628
rect 20718 28192 20774 28248
rect 20166 24268 20222 24304
rect 20166 24248 20168 24268
rect 20168 24248 20220 24268
rect 20220 24248 20222 24268
rect 20810 26460 20812 26480
rect 20812 26460 20864 26480
rect 20864 26460 20866 26480
rect 20810 26424 20866 26460
rect 20718 26152 20774 26208
rect 20626 23704 20682 23760
rect 20810 23740 20812 23760
rect 20812 23740 20864 23760
rect 20864 23740 20866 23760
rect 20810 23704 20866 23740
rect 20626 23296 20682 23352
rect 21454 26288 21510 26344
rect 22282 32136 22338 32192
rect 23018 34892 23020 34912
rect 23020 34892 23072 34912
rect 23072 34892 23074 34912
rect 23018 34856 23074 34892
rect 23846 35808 23902 35864
rect 21270 25356 21326 25392
rect 21270 25336 21272 25356
rect 21272 25336 21324 25356
rect 21324 25336 21326 25356
rect 20534 20712 20590 20768
rect 20350 16496 20406 16552
rect 20534 14320 20590 14376
rect 21270 23976 21326 24032
rect 21270 23568 21326 23624
rect 21454 23740 21456 23760
rect 21456 23740 21508 23760
rect 21508 23740 21510 23760
rect 21454 23704 21510 23740
rect 21178 19760 21234 19816
rect 20994 18944 21050 19000
rect 20902 16496 20958 16552
rect 20074 9832 20130 9888
rect 19706 8356 19762 8392
rect 19706 8336 19708 8356
rect 19708 8336 19760 8356
rect 19760 8336 19762 8356
rect 18602 3576 18658 3632
rect 22282 24520 22338 24576
rect 22190 21428 22192 21448
rect 22192 21428 22244 21448
rect 22244 21428 22246 21448
rect 22190 21392 22246 21428
rect 22006 18128 22062 18184
rect 21086 12552 21142 12608
rect 20718 12144 20774 12200
rect 20810 11192 20866 11248
rect 938 2080 994 2136
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 20626 3596 20682 3632
rect 20626 3576 20628 3596
rect 20628 3576 20680 3596
rect 20680 3576 20682 3596
rect 21638 10104 21694 10160
rect 21546 9868 21548 9888
rect 21548 9868 21600 9888
rect 21600 9868 21602 9888
rect 21178 9696 21234 9752
rect 21546 9832 21602 9868
rect 22190 10104 22246 10160
rect 22466 18148 22522 18184
rect 22466 18128 22468 18148
rect 22468 18128 22520 18148
rect 22520 18128 22522 18148
rect 23202 31728 23258 31784
rect 23110 27396 23166 27432
rect 23110 27376 23112 27396
rect 23112 27376 23164 27396
rect 23164 27376 23166 27396
rect 23110 24656 23166 24712
rect 23202 24148 23204 24168
rect 23204 24148 23256 24168
rect 23256 24148 23258 24168
rect 23202 24112 23258 24148
rect 23202 23296 23258 23352
rect 24214 32408 24270 32464
rect 24122 29824 24178 29880
rect 24214 27412 24216 27432
rect 24216 27412 24268 27432
rect 24268 27412 24270 27432
rect 24214 27376 24270 27412
rect 24122 25372 24124 25392
rect 24124 25372 24176 25392
rect 24176 25372 24178 25392
rect 24122 25336 24178 25372
rect 22834 15952 22890 16008
rect 23294 20324 23350 20360
rect 23294 20304 23296 20324
rect 23296 20304 23348 20324
rect 23348 20304 23350 20324
rect 25410 44396 25466 44432
rect 25410 44376 25412 44396
rect 25412 44376 25464 44396
rect 25464 44376 25466 44396
rect 25686 44784 25742 44840
rect 26054 44376 26110 44432
rect 26790 44240 26846 44296
rect 27434 46960 27490 47016
rect 27158 43732 27160 43752
rect 27160 43732 27212 43752
rect 27212 43732 27214 43752
rect 27158 43696 27214 43732
rect 27250 43308 27306 43344
rect 27250 43288 27252 43308
rect 27252 43288 27304 43308
rect 27304 43288 27306 43308
rect 27710 44512 27766 44568
rect 27342 43152 27398 43208
rect 27066 42880 27122 42936
rect 28446 44940 28502 44976
rect 28446 44920 28448 44940
rect 28448 44920 28500 44940
rect 28500 44920 28502 44940
rect 28354 43732 28356 43752
rect 28356 43732 28408 43752
rect 28408 43732 28410 43752
rect 28354 43696 28410 43732
rect 35600 47898 35656 47900
rect 35680 47898 35736 47900
rect 35760 47898 35816 47900
rect 35840 47898 35896 47900
rect 35600 47846 35646 47898
rect 35646 47846 35656 47898
rect 35680 47846 35710 47898
rect 35710 47846 35722 47898
rect 35722 47846 35736 47898
rect 35760 47846 35774 47898
rect 35774 47846 35786 47898
rect 35786 47846 35816 47898
rect 35840 47846 35850 47898
rect 35850 47846 35896 47898
rect 35600 47844 35656 47846
rect 35680 47844 35736 47846
rect 35760 47844 35816 47846
rect 35840 47844 35896 47846
rect 28630 44956 28632 44976
rect 28632 44956 28684 44976
rect 28684 44956 28686 44976
rect 28630 44920 28686 44956
rect 28630 44820 28632 44840
rect 28632 44820 28684 44840
rect 28684 44820 28686 44840
rect 28630 44784 28686 44820
rect 28630 44684 28632 44704
rect 28632 44684 28684 44704
rect 28684 44684 28686 44704
rect 28630 44648 28686 44684
rect 28630 44512 28686 44568
rect 28998 43696 29054 43752
rect 30654 44648 30710 44704
rect 29734 43424 29790 43480
rect 27526 40432 27582 40488
rect 25226 35264 25282 35320
rect 25410 35264 25466 35320
rect 25594 32136 25650 32192
rect 24858 27376 24914 27432
rect 25134 26560 25190 26616
rect 25226 22072 25282 22128
rect 23570 13640 23626 13696
rect 23662 12824 23718 12880
rect 22466 8064 22522 8120
rect 20902 5616 20958 5672
rect 23754 9968 23810 10024
rect 24950 12824 25006 12880
rect 25410 21800 25466 21856
rect 25962 26988 26018 27024
rect 25962 26968 25964 26988
rect 25964 26968 26016 26988
rect 26016 26968 26018 26988
rect 25962 26424 26018 26480
rect 27526 35944 27582 36000
rect 26974 35672 27030 35728
rect 26790 35128 26846 35184
rect 27342 35400 27398 35456
rect 28538 35944 28594 36000
rect 27986 35400 28042 35456
rect 27618 32000 27674 32056
rect 26146 26560 26202 26616
rect 25686 21664 25742 21720
rect 25962 21800 26018 21856
rect 26054 21664 26110 21720
rect 26330 18672 26386 18728
rect 26606 18708 26608 18728
rect 26608 18708 26660 18728
rect 26660 18708 26662 18728
rect 26606 18672 26662 18708
rect 27986 31184 28042 31240
rect 28262 28056 28318 28112
rect 27986 23604 27988 23624
rect 27988 23604 28040 23624
rect 28040 23604 28042 23624
rect 27342 18944 27398 19000
rect 27986 23568 28042 23604
rect 28538 23432 28594 23488
rect 22650 5616 22706 5672
rect 24122 3596 24178 3632
rect 24122 3576 24124 3596
rect 24124 3576 24176 3596
rect 24176 3576 24178 3596
rect 25042 9036 25098 9072
rect 25042 9016 25044 9036
rect 25044 9016 25096 9036
rect 25096 9016 25098 9036
rect 26606 14476 26662 14512
rect 26606 14456 26608 14476
rect 26608 14456 26660 14476
rect 26660 14456 26662 14476
rect 27158 14356 27160 14376
rect 27160 14356 27212 14376
rect 27212 14356 27214 14376
rect 27158 14320 27214 14356
rect 27710 12844 27766 12880
rect 27710 12824 27712 12844
rect 27712 12824 27764 12844
rect 27764 12824 27766 12844
rect 25410 11076 25466 11112
rect 25410 11056 25412 11076
rect 25412 11056 25464 11076
rect 25464 11056 25466 11076
rect 25594 8916 25596 8936
rect 25596 8916 25648 8936
rect 25648 8916 25650 8936
rect 25594 8880 25650 8916
rect 22834 2896 22890 2952
rect 26330 2932 26332 2952
rect 26332 2932 26384 2952
rect 26384 2932 26386 2952
rect 26330 2896 26386 2932
rect 20994 2624 21050 2680
rect 30838 43424 30894 43480
rect 28906 35128 28962 35184
rect 28998 32000 29054 32056
rect 29734 33904 29790 33960
rect 29366 29008 29422 29064
rect 28998 28328 29054 28384
rect 28998 27920 29054 27976
rect 29182 27240 29238 27296
rect 29090 24520 29146 24576
rect 31482 40024 31538 40080
rect 30378 32000 30434 32056
rect 30562 30796 30618 30832
rect 30562 30776 30564 30796
rect 30564 30776 30616 30796
rect 30616 30776 30618 30796
rect 29550 23704 29606 23760
rect 29550 23432 29606 23488
rect 29274 21800 29330 21856
rect 29182 18264 29238 18320
rect 29642 20984 29698 21040
rect 28998 16108 29054 16144
rect 28998 16088 29000 16108
rect 29000 16088 29052 16108
rect 29052 16088 29054 16108
rect 30010 20340 30012 20360
rect 30012 20340 30064 20360
rect 30064 20340 30066 20360
rect 30010 20304 30066 20340
rect 30010 18708 30012 18728
rect 30012 18708 30064 18728
rect 30064 18708 30066 18728
rect 30010 18672 30066 18708
rect 29918 12280 29974 12336
rect 29826 10920 29882 10976
rect 30378 23568 30434 23624
rect 30654 23840 30710 23896
rect 31022 31320 31078 31376
rect 30286 18264 30342 18320
rect 30378 13796 30434 13832
rect 30378 13776 30380 13796
rect 30380 13776 30432 13796
rect 30432 13776 30434 13796
rect 30378 12844 30434 12880
rect 30378 12824 30380 12844
rect 30380 12824 30432 12844
rect 30432 12824 30434 12844
rect 30286 12688 30342 12744
rect 31482 31456 31538 31512
rect 31482 30096 31538 30152
rect 31850 31320 31906 31376
rect 33138 45892 33194 45928
rect 33138 45872 33140 45892
rect 33140 45872 33192 45892
rect 33192 45872 33194 45892
rect 32402 45464 32458 45520
rect 32678 43424 32734 43480
rect 32586 41420 32588 41440
rect 32588 41420 32640 41440
rect 32640 41420 32642 41440
rect 32586 41384 32642 41420
rect 33690 45908 33692 45928
rect 33692 45908 33744 45928
rect 33744 45908 33746 45928
rect 33690 45872 33746 45908
rect 33046 34856 33102 34912
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 35600 46810 35656 46812
rect 35680 46810 35736 46812
rect 35760 46810 35816 46812
rect 35840 46810 35896 46812
rect 35600 46758 35646 46810
rect 35646 46758 35656 46810
rect 35680 46758 35710 46810
rect 35710 46758 35722 46810
rect 35722 46758 35736 46810
rect 35760 46758 35774 46810
rect 35774 46758 35786 46810
rect 35786 46758 35816 46810
rect 35840 46758 35850 46810
rect 35850 46758 35896 46810
rect 35600 46756 35656 46758
rect 35680 46756 35736 46758
rect 35760 46756 35816 46758
rect 35840 46756 35896 46758
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34426 44376 34482 44432
rect 35600 45722 35656 45724
rect 35680 45722 35736 45724
rect 35760 45722 35816 45724
rect 35840 45722 35896 45724
rect 35600 45670 35646 45722
rect 35646 45670 35656 45722
rect 35680 45670 35710 45722
rect 35710 45670 35722 45722
rect 35722 45670 35736 45722
rect 35760 45670 35774 45722
rect 35774 45670 35786 45722
rect 35786 45670 35816 45722
rect 35840 45670 35850 45722
rect 35850 45670 35896 45722
rect 35600 45668 35656 45670
rect 35680 45668 35736 45670
rect 35760 45668 35816 45670
rect 35840 45668 35896 45670
rect 35600 44634 35656 44636
rect 35680 44634 35736 44636
rect 35760 44634 35816 44636
rect 35840 44634 35896 44636
rect 35600 44582 35646 44634
rect 35646 44582 35656 44634
rect 35680 44582 35710 44634
rect 35710 44582 35722 44634
rect 35722 44582 35736 44634
rect 35760 44582 35774 44634
rect 35774 44582 35786 44634
rect 35786 44582 35816 44634
rect 35840 44582 35850 44634
rect 35850 44582 35896 44634
rect 35600 44580 35656 44582
rect 35680 44580 35736 44582
rect 35760 44580 35816 44582
rect 35840 44580 35896 44582
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34702 43152 34758 43208
rect 34518 40704 34574 40760
rect 35600 43546 35656 43548
rect 35680 43546 35736 43548
rect 35760 43546 35816 43548
rect 35840 43546 35896 43548
rect 35600 43494 35646 43546
rect 35646 43494 35656 43546
rect 35680 43494 35710 43546
rect 35710 43494 35722 43546
rect 35722 43494 35736 43546
rect 35760 43494 35774 43546
rect 35774 43494 35786 43546
rect 35786 43494 35816 43546
rect 35840 43494 35850 43546
rect 35850 43494 35896 43546
rect 35600 43492 35656 43494
rect 35680 43492 35736 43494
rect 35760 43492 35816 43494
rect 35840 43492 35896 43494
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 35600 42458 35656 42460
rect 35680 42458 35736 42460
rect 35760 42458 35816 42460
rect 35840 42458 35896 42460
rect 35600 42406 35646 42458
rect 35646 42406 35656 42458
rect 35680 42406 35710 42458
rect 35710 42406 35722 42458
rect 35722 42406 35736 42458
rect 35760 42406 35774 42458
rect 35774 42406 35786 42458
rect 35786 42406 35816 42458
rect 35840 42406 35850 42458
rect 35850 42406 35896 42458
rect 35600 42404 35656 42406
rect 35680 42404 35736 42406
rect 35760 42404 35816 42406
rect 35840 42404 35896 42406
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34886 41656 34942 41712
rect 35162 41520 35218 41576
rect 35714 41656 35770 41712
rect 36266 41520 36322 41576
rect 35600 41370 35656 41372
rect 35680 41370 35736 41372
rect 35760 41370 35816 41372
rect 35840 41370 35896 41372
rect 35600 41318 35646 41370
rect 35646 41318 35656 41370
rect 35680 41318 35710 41370
rect 35710 41318 35722 41370
rect 35722 41318 35736 41370
rect 35760 41318 35774 41370
rect 35774 41318 35786 41370
rect 35786 41318 35816 41370
rect 35840 41318 35850 41370
rect 35850 41318 35896 41370
rect 35600 41316 35656 41318
rect 35680 41316 35736 41318
rect 35760 41316 35816 41318
rect 35840 41316 35896 41318
rect 34702 40704 34758 40760
rect 33414 30776 33470 30832
rect 32862 30640 32918 30696
rect 31298 26832 31354 26888
rect 31574 22072 31630 22128
rect 31850 19896 31906 19952
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 35600 40282 35656 40284
rect 35680 40282 35736 40284
rect 35760 40282 35816 40284
rect 35840 40282 35896 40284
rect 35600 40230 35646 40282
rect 35646 40230 35656 40282
rect 35680 40230 35710 40282
rect 35710 40230 35722 40282
rect 35722 40230 35736 40282
rect 35760 40230 35774 40282
rect 35774 40230 35786 40282
rect 35786 40230 35816 40282
rect 35840 40230 35850 40282
rect 35850 40230 35896 40282
rect 35600 40228 35656 40230
rect 35680 40228 35736 40230
rect 35760 40228 35816 40230
rect 35840 40228 35896 40230
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 35600 39194 35656 39196
rect 35680 39194 35736 39196
rect 35760 39194 35816 39196
rect 35840 39194 35896 39196
rect 35600 39142 35646 39194
rect 35646 39142 35656 39194
rect 35680 39142 35710 39194
rect 35710 39142 35722 39194
rect 35722 39142 35736 39194
rect 35760 39142 35774 39194
rect 35774 39142 35786 39194
rect 35786 39142 35816 39194
rect 35840 39142 35850 39194
rect 35850 39142 35896 39194
rect 35600 39140 35656 39142
rect 35680 39140 35736 39142
rect 35760 39140 35816 39142
rect 35840 39140 35896 39142
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34886 37304 34942 37360
rect 35600 38106 35656 38108
rect 35680 38106 35736 38108
rect 35760 38106 35816 38108
rect 35840 38106 35896 38108
rect 35600 38054 35646 38106
rect 35646 38054 35656 38106
rect 35680 38054 35710 38106
rect 35710 38054 35722 38106
rect 35722 38054 35736 38106
rect 35760 38054 35774 38106
rect 35774 38054 35786 38106
rect 35786 38054 35816 38106
rect 35840 38054 35850 38106
rect 35850 38054 35896 38106
rect 35600 38052 35656 38054
rect 35680 38052 35736 38054
rect 35760 38052 35816 38054
rect 35840 38052 35896 38054
rect 35806 37848 35862 37904
rect 35806 37340 35808 37360
rect 35808 37340 35860 37360
rect 35860 37340 35862 37360
rect 35806 37304 35862 37340
rect 36082 37068 36084 37088
rect 36084 37068 36136 37088
rect 36136 37068 36138 37088
rect 36082 37032 36138 37068
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 37646 43696 37702 43752
rect 37738 42880 37794 42936
rect 36818 39344 36874 39400
rect 36542 39208 36598 39264
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34978 35028 34980 35048
rect 34980 35028 35032 35048
rect 35032 35028 35034 35048
rect 34978 34992 35034 35028
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34886 31864 34942 31920
rect 35990 32272 36046 32328
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 35438 31476 35494 31512
rect 35438 31456 35440 31476
rect 35440 31456 35492 31476
rect 35492 31456 35494 31476
rect 35346 31320 35402 31376
rect 35254 31184 35310 31240
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 33874 25608 33930 25664
rect 30194 7948 30250 7984
rect 30194 7928 30196 7948
rect 30196 7928 30248 7948
rect 30248 7928 30250 7948
rect 33506 20848 33562 20904
rect 33874 21528 33930 21584
rect 34150 20984 34206 21040
rect 35162 30776 35218 30832
rect 34702 28192 34758 28248
rect 34610 24812 34666 24848
rect 34610 24792 34612 24812
rect 34612 24792 34664 24812
rect 34664 24792 34666 24812
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35714 31320 35770 31376
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 35438 29688 35494 29744
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 35806 29008 35862 29064
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34242 20848 34298 20904
rect 33782 19216 33838 19272
rect 33782 18708 33784 18728
rect 33784 18708 33836 18728
rect 33836 18708 33838 18728
rect 33782 18672 33838 18708
rect 31482 12588 31484 12608
rect 31484 12588 31536 12608
rect 31536 12588 31538 12608
rect 31482 12552 31538 12588
rect 31666 3440 31722 3496
rect 32678 4684 32734 4720
rect 32678 4664 32680 4684
rect 32680 4664 32732 4684
rect 32732 4664 32734 4684
rect 33138 8064 33194 8120
rect 34702 20460 34758 20496
rect 34702 20440 34704 20460
rect 34704 20440 34756 20460
rect 34756 20440 34758 20460
rect 33782 13776 33838 13832
rect 34058 12552 34114 12608
rect 34242 7384 34298 7440
rect 33322 4664 33378 4720
rect 33046 3576 33102 3632
rect 33874 3596 33930 3632
rect 33874 3576 33876 3596
rect 33876 3576 33928 3596
rect 33928 3576 33930 3596
rect 35254 23860 35310 23896
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 35254 23840 35256 23860
rect 35256 23840 35308 23860
rect 35308 23840 35310 23860
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 34978 21936 35034 21992
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34886 19252 34888 19272
rect 34888 19252 34940 19272
rect 34940 19252 34942 19272
rect 34886 19216 34942 19252
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 36542 31084 36544 31104
rect 36544 31084 36596 31104
rect 36596 31084 36598 31104
rect 36542 31048 36598 31084
rect 36450 30676 36452 30696
rect 36452 30676 36504 30696
rect 36504 30676 36506 30696
rect 36450 30640 36506 30676
rect 45926 47660 45982 47696
rect 45926 47640 45928 47660
rect 45928 47640 45980 47660
rect 45980 47640 45982 47660
rect 37278 40024 37334 40080
rect 37462 39208 37518 39264
rect 36266 28600 36322 28656
rect 36358 25880 36414 25936
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 36818 29280 36874 29336
rect 37002 25200 37058 25256
rect 36174 18672 36230 18728
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35990 11056 36046 11112
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34794 9560 34850 9616
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35254 3440 35310 3496
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37094 24656 37150 24712
rect 34886 2488 34942 2544
rect 37278 29008 37334 29064
rect 37278 25356 37334 25392
rect 37278 25336 37280 25356
rect 37280 25336 37332 25356
rect 37332 25336 37334 25356
rect 37278 17176 37334 17232
rect 37646 30096 37702 30152
rect 37830 23160 37886 23216
rect 38382 41132 38438 41168
rect 38382 41112 38384 41132
rect 38384 41112 38436 41132
rect 38436 41112 38438 41132
rect 38106 29164 38162 29200
rect 38106 29144 38108 29164
rect 38108 29144 38160 29164
rect 38160 29144 38162 29164
rect 38290 29300 38346 29336
rect 38290 29280 38292 29300
rect 38292 29280 38344 29300
rect 38344 29280 38346 29300
rect 40406 43288 40462 43344
rect 39578 40024 39634 40080
rect 39854 35672 39910 35728
rect 38290 23724 38346 23760
rect 38290 23704 38292 23724
rect 38292 23704 38344 23724
rect 38344 23704 38346 23724
rect 38474 23432 38530 23488
rect 37554 15952 37610 16008
rect 38106 16632 38162 16688
rect 37738 11192 37794 11248
rect 38750 22636 38806 22672
rect 38750 22616 38752 22636
rect 38752 22616 38804 22636
rect 38804 22616 38806 22636
rect 40038 35536 40094 35592
rect 40130 35128 40186 35184
rect 39946 27648 40002 27704
rect 39210 24656 39266 24712
rect 38934 22208 38990 22264
rect 38658 18808 38714 18864
rect 39118 22344 39174 22400
rect 39118 22208 39174 22264
rect 39486 23160 39542 23216
rect 41142 29008 41198 29064
rect 42154 34312 42210 34368
rect 42154 32952 42210 33008
rect 41694 32716 41696 32736
rect 41696 32716 41748 32736
rect 41748 32716 41750 32736
rect 41694 32680 41750 32716
rect 41602 32544 41658 32600
rect 42522 32988 42524 33008
rect 42524 32988 42576 33008
rect 42576 32988 42578 33008
rect 42522 32952 42578 32988
rect 42798 32716 42800 32736
rect 42800 32716 42852 32736
rect 42852 32716 42854 32736
rect 42798 32680 42854 32716
rect 41510 29008 41566 29064
rect 39486 20576 39542 20632
rect 40130 21392 40186 21448
rect 38566 12144 38622 12200
rect 38382 11192 38438 11248
rect 41234 23976 41290 24032
rect 40590 19760 40646 19816
rect 41418 27784 41474 27840
rect 41602 24148 41604 24168
rect 41604 24148 41656 24168
rect 41656 24148 41658 24168
rect 41602 24112 41658 24148
rect 41694 23724 41750 23760
rect 41694 23704 41696 23724
rect 41696 23704 41748 23724
rect 41748 23704 41750 23724
rect 41878 24248 41934 24304
rect 43166 32544 43222 32600
rect 42614 27820 42616 27840
rect 42616 27820 42668 27840
rect 42668 27820 42670 27840
rect 42614 27784 42670 27820
rect 42522 24268 42578 24304
rect 42522 24248 42524 24268
rect 42524 24248 42576 24268
rect 42576 24248 42578 24268
rect 42430 24112 42486 24168
rect 42982 24112 43038 24168
rect 43258 24148 43260 24168
rect 43260 24148 43312 24168
rect 43312 24148 43314 24168
rect 42982 23976 43038 24032
rect 43258 24112 43314 24148
rect 38750 11736 38806 11792
rect 39210 12144 39266 12200
rect 39854 10512 39910 10568
rect 37462 2624 37518 2680
rect 40774 11600 40830 11656
rect 41326 11600 41382 11656
rect 43718 23724 43774 23760
rect 43718 23704 43720 23724
rect 43720 23704 43772 23724
rect 43772 23704 43774 23724
rect 43626 23160 43682 23216
rect 45834 30912 45890 30968
rect 45650 27668 45706 27704
rect 45650 27648 45652 27668
rect 45652 27648 45704 27668
rect 45704 27648 45706 27668
rect 46754 44920 46810 44976
rect 45926 25236 45928 25256
rect 45928 25236 45980 25256
rect 45980 25236 45982 25256
rect 45926 25200 45982 25236
rect 44914 24148 44916 24168
rect 44916 24148 44968 24168
rect 44968 24148 44970 24168
rect 44914 24112 44970 24148
rect 44178 23704 44234 23760
rect 46018 24148 46020 24168
rect 46020 24148 46072 24168
rect 46072 24148 46074 24168
rect 46018 24112 46074 24148
rect 42706 12180 42708 12200
rect 42708 12180 42760 12200
rect 42760 12180 42762 12200
rect 42706 12144 42762 12180
rect 46662 42880 46718 42936
rect 46662 40160 46718 40216
rect 46662 37440 46718 37496
rect 46662 35436 46664 35456
rect 46664 35436 46716 35456
rect 46716 35436 46718 35456
rect 46662 35400 46718 35436
rect 46662 32716 46664 32736
rect 46664 32716 46716 32736
rect 46716 32716 46718 32736
rect 46662 32680 46718 32716
rect 46662 29960 46718 30016
rect 46662 28464 46718 28520
rect 46570 27920 46626 27976
rect 46570 23160 46626 23216
rect 46662 20440 46718 20496
rect 43074 11736 43130 11792
rect 42614 11092 42616 11112
rect 42616 11092 42668 11112
rect 42668 11092 42670 11112
rect 42614 11056 42670 11092
rect 42890 11056 42946 11112
rect 43258 11636 43260 11656
rect 43260 11636 43312 11656
rect 43312 11636 43314 11656
rect 43258 11600 43314 11636
rect 43626 12180 43628 12200
rect 43628 12180 43680 12200
rect 43680 12180 43682 12200
rect 43626 12144 43682 12180
rect 43534 11092 43536 11112
rect 43536 11092 43588 11112
rect 43588 11092 43590 11112
rect 43534 11056 43590 11092
rect 46386 17720 46442 17776
rect 46754 17720 46810 17776
rect 46662 15680 46718 15736
rect 46662 12960 46718 13016
rect 46662 10240 46718 10296
rect 45926 8200 45982 8256
rect 45558 6160 45614 6216
rect 39210 4004 39266 4040
rect 39210 3984 39212 4004
rect 39212 3984 39264 4004
rect 39264 3984 39266 4004
rect 42706 2624 42762 2680
rect 46662 5516 46664 5536
rect 46664 5516 46716 5536
rect 46716 5516 46718 5536
rect 46662 5480 46718 5516
rect 46570 2760 46626 2816
rect 46202 2508 46258 2544
rect 46202 2488 46204 2508
rect 46204 2488 46256 2508
rect 46256 2488 46258 2508
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 45650 2352 45706 2408
rect 45466 720 45522 776
<< metal3 >>
rect 0 49058 800 49088
rect 1761 49058 1827 49061
rect 0 49056 1827 49058
rect 0 49000 1766 49056
rect 1822 49000 1827 49056
rect 0 48998 1827 49000
rect 0 48968 800 48998
rect 1761 48995 1827 48998
rect 4870 47904 5186 47905
rect 4870 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5186 47904
rect 4870 47839 5186 47840
rect 35590 47904 35906 47905
rect 35590 47840 35596 47904
rect 35660 47840 35676 47904
rect 35740 47840 35756 47904
rect 35820 47840 35836 47904
rect 35900 47840 35906 47904
rect 35590 47839 35906 47840
rect 45921 47698 45987 47701
rect 47480 47698 48280 47728
rect 45921 47696 48280 47698
rect 45921 47640 45926 47696
rect 45982 47640 48280 47696
rect 45921 47638 48280 47640
rect 45921 47635 45987 47638
rect 47480 47608 48280 47638
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 0 47018 800 47048
rect 1117 47018 1183 47021
rect 0 47016 1183 47018
rect 0 46960 1122 47016
rect 1178 46960 1183 47016
rect 0 46958 1183 46960
rect 0 46928 800 46958
rect 1117 46955 1183 46958
rect 27429 47018 27495 47021
rect 32254 47018 32260 47020
rect 27429 47016 32260 47018
rect 27429 46960 27434 47016
rect 27490 46960 32260 47016
rect 27429 46958 32260 46960
rect 27429 46955 27495 46958
rect 32254 46956 32260 46958
rect 32324 46956 32330 47020
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 35590 46816 35906 46817
rect 35590 46752 35596 46816
rect 35660 46752 35676 46816
rect 35740 46752 35756 46816
rect 35820 46752 35836 46816
rect 35900 46752 35906 46816
rect 35590 46751 35906 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 33133 45930 33199 45933
rect 33685 45932 33751 45933
rect 33685 45930 33732 45932
rect 33133 45928 33732 45930
rect 33133 45872 33138 45928
rect 33194 45872 33690 45928
rect 33133 45870 33732 45872
rect 33133 45867 33199 45870
rect 33685 45868 33732 45870
rect 33796 45868 33802 45932
rect 33685 45867 33751 45868
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 35590 45728 35906 45729
rect 35590 45664 35596 45728
rect 35660 45664 35676 45728
rect 35740 45664 35756 45728
rect 35820 45664 35836 45728
rect 35900 45664 35906 45728
rect 35590 45663 35906 45664
rect 32397 45524 32463 45525
rect 32397 45522 32444 45524
rect 32352 45520 32444 45522
rect 32352 45464 32402 45520
rect 32352 45462 32444 45464
rect 32397 45460 32444 45462
rect 32508 45460 32514 45524
rect 32397 45459 32463 45460
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 28441 44978 28507 44981
rect 28625 44978 28691 44981
rect 28441 44976 28691 44978
rect 28441 44920 28446 44976
rect 28502 44920 28630 44976
rect 28686 44920 28691 44976
rect 28441 44918 28691 44920
rect 28441 44915 28507 44918
rect 28625 44915 28691 44918
rect 46749 44978 46815 44981
rect 47480 44978 48280 45008
rect 46749 44976 48280 44978
rect 46749 44920 46754 44976
rect 46810 44920 48280 44976
rect 46749 44918 48280 44920
rect 46749 44915 46815 44918
rect 47480 44888 48280 44918
rect 25681 44842 25747 44845
rect 28625 44842 28691 44845
rect 25681 44840 28691 44842
rect 25681 44784 25686 44840
rect 25742 44784 28630 44840
rect 28686 44784 28691 44840
rect 25681 44782 28691 44784
rect 25681 44779 25747 44782
rect 28625 44779 28691 44782
rect 28625 44706 28691 44709
rect 30649 44706 30715 44709
rect 28625 44704 30715 44706
rect 28625 44648 28630 44704
rect 28686 44648 30654 44704
rect 30710 44648 30715 44704
rect 28625 44646 30715 44648
rect 28625 44643 28691 44646
rect 30649 44643 30715 44646
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 35590 44640 35906 44641
rect 35590 44576 35596 44640
rect 35660 44576 35676 44640
rect 35740 44576 35756 44640
rect 35820 44576 35836 44640
rect 35900 44576 35906 44640
rect 35590 44575 35906 44576
rect 27705 44570 27771 44573
rect 28625 44570 28691 44573
rect 27705 44568 28691 44570
rect 27705 44512 27710 44568
rect 27766 44512 28630 44568
rect 28686 44512 28691 44568
rect 27705 44510 28691 44512
rect 27705 44507 27771 44510
rect 28625 44507 28691 44510
rect 25405 44434 25471 44437
rect 26049 44434 26115 44437
rect 34421 44434 34487 44437
rect 25405 44432 34487 44434
rect 25405 44376 25410 44432
rect 25466 44376 26054 44432
rect 26110 44376 34426 44432
rect 34482 44376 34487 44432
rect 25405 44374 34487 44376
rect 25405 44371 25471 44374
rect 26049 44371 26115 44374
rect 34421 44371 34487 44374
rect 0 44298 800 44328
rect 933 44298 999 44301
rect 0 44296 999 44298
rect 0 44240 938 44296
rect 994 44240 999 44296
rect 0 44238 999 44240
rect 0 44208 800 44238
rect 933 44235 999 44238
rect 26785 44298 26851 44301
rect 26918 44298 26924 44300
rect 26785 44296 26924 44298
rect 26785 44240 26790 44296
rect 26846 44240 26924 44296
rect 26785 44238 26924 44240
rect 26785 44235 26851 44238
rect 26918 44236 26924 44238
rect 26988 44236 26994 44300
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19057 43754 19123 43757
rect 19190 43754 19196 43756
rect 19057 43752 19196 43754
rect 19057 43696 19062 43752
rect 19118 43696 19196 43752
rect 19057 43694 19196 43696
rect 19057 43691 19123 43694
rect 19190 43692 19196 43694
rect 19260 43692 19266 43756
rect 27153 43754 27219 43757
rect 28349 43754 28415 43757
rect 27153 43752 28415 43754
rect 27153 43696 27158 43752
rect 27214 43696 28354 43752
rect 28410 43696 28415 43752
rect 27153 43694 28415 43696
rect 27153 43691 27219 43694
rect 28349 43691 28415 43694
rect 28993 43754 29059 43757
rect 37641 43754 37707 43757
rect 28993 43752 37707 43754
rect 28993 43696 28998 43752
rect 29054 43696 37646 43752
rect 37702 43696 37707 43752
rect 28993 43694 37707 43696
rect 28993 43691 29059 43694
rect 37641 43691 37707 43694
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 35590 43552 35906 43553
rect 35590 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35906 43552
rect 35590 43487 35906 43488
rect 29729 43482 29795 43485
rect 30833 43482 30899 43485
rect 32673 43482 32739 43485
rect 29729 43480 32739 43482
rect 29729 43424 29734 43480
rect 29790 43424 30838 43480
rect 30894 43424 32678 43480
rect 32734 43424 32739 43480
rect 29729 43422 32739 43424
rect 29729 43419 29795 43422
rect 30833 43419 30899 43422
rect 32673 43419 32739 43422
rect 27245 43346 27311 43349
rect 40401 43346 40467 43349
rect 27245 43344 40467 43346
rect 27245 43288 27250 43344
rect 27306 43288 40406 43344
rect 40462 43288 40467 43344
rect 27245 43286 40467 43288
rect 27245 43283 27311 43286
rect 40401 43283 40467 43286
rect 27337 43210 27403 43213
rect 34697 43210 34763 43213
rect 27337 43208 34763 43210
rect 27337 43152 27342 43208
rect 27398 43152 34702 43208
rect 34758 43152 34763 43208
rect 27337 43150 34763 43152
rect 27337 43147 27403 43150
rect 34697 43147 34763 43150
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 27061 42940 27127 42941
rect 37733 42940 37799 42941
rect 27061 42936 27108 42940
rect 27172 42938 27178 42940
rect 27061 42880 27066 42936
rect 27061 42876 27108 42880
rect 27172 42878 27218 42938
rect 37733 42936 37780 42940
rect 37844 42938 37850 42940
rect 46657 42938 46723 42941
rect 47480 42938 48280 42968
rect 37733 42880 37738 42936
rect 27172 42876 27178 42878
rect 37733 42876 37780 42880
rect 37844 42878 37890 42938
rect 46657 42936 48280 42938
rect 46657 42880 46662 42936
rect 46718 42880 48280 42936
rect 46657 42878 48280 42880
rect 37844 42876 37850 42878
rect 27061 42875 27127 42876
rect 37733 42875 37799 42876
rect 46657 42875 46723 42878
rect 47480 42848 48280 42878
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 35590 42464 35906 42465
rect 35590 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35906 42464
rect 35590 42399 35906 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 34881 41714 34947 41717
rect 35709 41714 35775 41717
rect 34881 41712 35775 41714
rect 34881 41656 34886 41712
rect 34942 41656 35714 41712
rect 35770 41656 35775 41712
rect 34881 41654 35775 41656
rect 34881 41651 34947 41654
rect 35709 41651 35775 41654
rect 0 41578 800 41608
rect 933 41578 999 41581
rect 0 41576 999 41578
rect 0 41520 938 41576
rect 994 41520 999 41576
rect 0 41518 999 41520
rect 0 41488 800 41518
rect 933 41515 999 41518
rect 35157 41578 35223 41581
rect 36261 41578 36327 41581
rect 35157 41576 36327 41578
rect 35157 41520 35162 41576
rect 35218 41520 36266 41576
rect 36322 41520 36327 41576
rect 35157 41518 36327 41520
rect 35157 41515 35223 41518
rect 36261 41515 36327 41518
rect 32581 41444 32647 41445
rect 32581 41440 32628 41444
rect 32692 41442 32698 41444
rect 32581 41384 32586 41440
rect 32581 41380 32628 41384
rect 32692 41382 32738 41442
rect 32692 41380 32698 41382
rect 32581 41379 32647 41380
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 35590 41376 35906 41377
rect 35590 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35906 41376
rect 35590 41311 35906 41312
rect 10225 41170 10291 41173
rect 38377 41170 38443 41173
rect 10225 41168 38443 41170
rect 10225 41112 10230 41168
rect 10286 41112 38382 41168
rect 38438 41112 38443 41168
rect 10225 41110 38443 41112
rect 10225 41107 10291 41110
rect 38377 41107 38443 41110
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 34513 40762 34579 40765
rect 34697 40762 34763 40765
rect 34513 40760 34763 40762
rect 34513 40704 34518 40760
rect 34574 40704 34702 40760
rect 34758 40704 34763 40760
rect 34513 40702 34763 40704
rect 34513 40699 34579 40702
rect 34697 40699 34763 40702
rect 22461 40490 22527 40493
rect 27521 40490 27587 40493
rect 22461 40488 27587 40490
rect 22461 40432 22466 40488
rect 22522 40432 27526 40488
rect 27582 40432 27587 40488
rect 22461 40430 27587 40432
rect 22461 40427 22527 40430
rect 27521 40427 27587 40430
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 35590 40288 35906 40289
rect 35590 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35906 40288
rect 35590 40223 35906 40224
rect 46657 40218 46723 40221
rect 47480 40218 48280 40248
rect 46657 40216 48280 40218
rect 46657 40160 46662 40216
rect 46718 40160 48280 40216
rect 46657 40158 48280 40160
rect 46657 40155 46723 40158
rect 47480 40128 48280 40158
rect 20478 40020 20484 40084
rect 20548 40082 20554 40084
rect 20621 40082 20687 40085
rect 20548 40080 20687 40082
rect 20548 40024 20626 40080
rect 20682 40024 20687 40080
rect 20548 40022 20687 40024
rect 20548 40020 20554 40022
rect 20621 40019 20687 40022
rect 31477 40082 31543 40085
rect 37273 40082 37339 40085
rect 31477 40080 37339 40082
rect 31477 40024 31482 40080
rect 31538 40024 37278 40080
rect 37334 40024 37339 40080
rect 31477 40022 37339 40024
rect 31477 40019 31543 40022
rect 37273 40019 37339 40022
rect 38878 40020 38884 40084
rect 38948 40082 38954 40084
rect 39573 40082 39639 40085
rect 38948 40080 39639 40082
rect 38948 40024 39578 40080
rect 39634 40024 39639 40080
rect 38948 40022 39639 40024
rect 38948 40020 38954 40022
rect 39573 40019 39639 40022
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 0 39538 800 39568
rect 933 39538 999 39541
rect 0 39536 999 39538
rect 0 39480 938 39536
rect 994 39480 999 39536
rect 0 39478 999 39480
rect 0 39448 800 39478
rect 933 39475 999 39478
rect 12934 39340 12940 39404
rect 13004 39402 13010 39404
rect 36813 39402 36879 39405
rect 13004 39400 36879 39402
rect 13004 39344 36818 39400
rect 36874 39344 36879 39400
rect 13004 39342 36879 39344
rect 13004 39340 13010 39342
rect 36813 39339 36879 39342
rect 36537 39266 36603 39269
rect 37457 39266 37523 39269
rect 36537 39264 37523 39266
rect 36537 39208 36542 39264
rect 36598 39208 37462 39264
rect 37518 39208 37523 39264
rect 36537 39206 37523 39208
rect 36537 39203 36603 39206
rect 37457 39203 37523 39206
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 35590 39200 35906 39201
rect 35590 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35906 39200
rect 35590 39135 35906 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 17861 38314 17927 38317
rect 18822 38314 18828 38316
rect 17861 38312 18828 38314
rect 17861 38256 17866 38312
rect 17922 38256 18828 38312
rect 17861 38254 18828 38256
rect 17861 38251 17927 38254
rect 18822 38252 18828 38254
rect 18892 38314 18898 38316
rect 22461 38314 22527 38317
rect 18892 38312 22527 38314
rect 18892 38256 22466 38312
rect 22522 38256 22527 38312
rect 18892 38254 22527 38256
rect 18892 38252 18898 38254
rect 22461 38251 22527 38254
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 35590 38112 35906 38113
rect 35590 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35906 38112
rect 35590 38047 35906 38048
rect 17677 38042 17743 38045
rect 18965 38042 19031 38045
rect 17677 38040 19031 38042
rect 17677 37984 17682 38040
rect 17738 37984 18970 38040
rect 19026 37984 19031 38040
rect 17677 37982 19031 37984
rect 17677 37979 17743 37982
rect 18965 37979 19031 37982
rect 16205 37906 16271 37909
rect 35801 37906 35867 37909
rect 16205 37904 35867 37906
rect 16205 37848 16210 37904
rect 16266 37848 35806 37904
rect 35862 37848 35867 37904
rect 16205 37846 35867 37848
rect 16205 37843 16271 37846
rect 35801 37843 35867 37846
rect 9581 37634 9647 37637
rect 11053 37634 11119 37637
rect 9581 37632 11119 37634
rect 9581 37576 9586 37632
rect 9642 37576 11058 37632
rect 11114 37576 11119 37632
rect 9581 37574 11119 37576
rect 9581 37571 9647 37574
rect 11053 37571 11119 37574
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 46657 37498 46723 37501
rect 47480 37498 48280 37528
rect 46657 37496 48280 37498
rect 46657 37440 46662 37496
rect 46718 37440 48280 37496
rect 46657 37438 48280 37440
rect 46657 37435 46723 37438
rect 47480 37408 48280 37438
rect 34881 37362 34947 37365
rect 35801 37362 35867 37365
rect 34881 37360 35867 37362
rect 34881 37304 34886 37360
rect 34942 37304 35806 37360
rect 35862 37304 35867 37360
rect 34881 37302 35867 37304
rect 34881 37299 34947 37302
rect 35801 37299 35867 37302
rect 36077 37092 36143 37093
rect 36077 37090 36124 37092
rect 36032 37088 36124 37090
rect 36032 37032 36082 37088
rect 36032 37030 36124 37032
rect 36077 37028 36124 37030
rect 36188 37028 36194 37092
rect 36077 37027 36143 37028
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 0 36818 800 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 800 36758
rect 933 36755 999 36758
rect 14457 36818 14523 36821
rect 16757 36818 16823 36821
rect 14457 36816 16823 36818
rect 14457 36760 14462 36816
rect 14518 36760 16762 36816
rect 16818 36760 16823 36816
rect 14457 36758 16823 36760
rect 14457 36755 14523 36758
rect 16757 36755 16823 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19517 36002 19583 36005
rect 27521 36002 27587 36005
rect 28533 36002 28599 36005
rect 19517 36000 28599 36002
rect 19517 35944 19522 36000
rect 19578 35944 27526 36000
rect 27582 35944 28538 36000
rect 28594 35944 28599 36000
rect 19517 35942 28599 35944
rect 19517 35939 19583 35942
rect 27521 35939 27587 35942
rect 28533 35939 28599 35942
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 19149 35866 19215 35869
rect 23841 35866 23907 35869
rect 19149 35864 23907 35866
rect 19149 35808 19154 35864
rect 19210 35808 23846 35864
rect 23902 35808 23907 35864
rect 19149 35806 23907 35808
rect 19149 35803 19215 35806
rect 23841 35803 23907 35806
rect 26969 35730 27035 35733
rect 39849 35730 39915 35733
rect 26969 35728 39915 35730
rect 26969 35672 26974 35728
rect 27030 35672 39854 35728
rect 39910 35672 39915 35728
rect 26969 35670 39915 35672
rect 26969 35667 27035 35670
rect 39849 35667 39915 35670
rect 19149 35594 19215 35597
rect 40033 35594 40099 35597
rect 19149 35592 40099 35594
rect 19149 35536 19154 35592
rect 19210 35536 40038 35592
rect 40094 35536 40099 35592
rect 19149 35534 40099 35536
rect 19149 35531 19215 35534
rect 40033 35531 40099 35534
rect 15285 35458 15351 35461
rect 27337 35458 27403 35461
rect 27981 35458 28047 35461
rect 15285 35456 28047 35458
rect 15285 35400 15290 35456
rect 15346 35400 27342 35456
rect 27398 35400 27986 35456
rect 28042 35400 28047 35456
rect 15285 35398 28047 35400
rect 15285 35395 15351 35398
rect 27337 35395 27403 35398
rect 27981 35395 28047 35398
rect 46657 35458 46723 35461
rect 47480 35458 48280 35488
rect 46657 35456 48280 35458
rect 46657 35400 46662 35456
rect 46718 35400 48280 35456
rect 46657 35398 48280 35400
rect 46657 35395 46723 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 47480 35368 48280 35398
rect 34930 35327 35246 35328
rect 21909 35322 21975 35325
rect 25221 35322 25287 35325
rect 25405 35322 25471 35325
rect 21909 35320 25471 35322
rect 21909 35264 21914 35320
rect 21970 35264 25226 35320
rect 25282 35264 25410 35320
rect 25466 35264 25471 35320
rect 21909 35262 25471 35264
rect 21909 35259 21975 35262
rect 25221 35259 25287 35262
rect 25405 35259 25471 35262
rect 6085 35186 6151 35189
rect 20161 35186 20227 35189
rect 6085 35184 20227 35186
rect 6085 35128 6090 35184
rect 6146 35128 20166 35184
rect 20222 35128 20227 35184
rect 6085 35126 20227 35128
rect 6085 35123 6151 35126
rect 20161 35123 20227 35126
rect 20437 35186 20503 35189
rect 21398 35186 21404 35188
rect 20437 35184 21404 35186
rect 20437 35128 20442 35184
rect 20498 35128 21404 35184
rect 20437 35126 21404 35128
rect 20437 35123 20503 35126
rect 21398 35124 21404 35126
rect 21468 35186 21474 35188
rect 26785 35186 26851 35189
rect 21468 35184 26851 35186
rect 21468 35128 26790 35184
rect 26846 35128 26851 35184
rect 21468 35126 26851 35128
rect 21468 35124 21474 35126
rect 26785 35123 26851 35126
rect 28901 35186 28967 35189
rect 40125 35186 40191 35189
rect 28901 35184 40191 35186
rect 28901 35128 28906 35184
rect 28962 35128 40130 35184
rect 40186 35128 40191 35184
rect 28901 35126 40191 35128
rect 28901 35123 28967 35126
rect 40125 35123 40191 35126
rect 14089 35050 14155 35053
rect 34973 35050 35039 35053
rect 14089 35048 35039 35050
rect 14089 34992 14094 35048
rect 14150 34992 34978 35048
rect 35034 34992 35039 35048
rect 14089 34990 35039 34992
rect 14089 34987 14155 34990
rect 34973 34987 35039 34990
rect 23013 34914 23079 34917
rect 33041 34914 33107 34917
rect 23013 34912 33107 34914
rect 23013 34856 23018 34912
rect 23074 34856 33046 34912
rect 33102 34856 33107 34912
rect 23013 34854 33107 34856
rect 23013 34851 23079 34854
rect 33041 34851 33107 34854
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 42149 34372 42215 34373
rect 42149 34370 42196 34372
rect 42104 34368 42196 34370
rect 42104 34312 42154 34368
rect 42104 34310 42196 34312
rect 42149 34308 42196 34310
rect 42260 34308 42266 34372
rect 42149 34307 42215 34308
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 0 34098 800 34128
rect 1577 34098 1643 34101
rect 0 34096 1643 34098
rect 0 34040 1582 34096
rect 1638 34040 1643 34096
rect 0 34038 1643 34040
rect 0 34008 800 34038
rect 1577 34035 1643 34038
rect 10777 33962 10843 33965
rect 21541 33962 21607 33965
rect 29729 33962 29795 33965
rect 10777 33960 29795 33962
rect 10777 33904 10782 33960
rect 10838 33904 21546 33960
rect 21602 33904 29734 33960
rect 29790 33904 29795 33960
rect 10777 33902 29795 33904
rect 10777 33899 10843 33902
rect 21541 33899 21607 33902
rect 29729 33899 29795 33902
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 16941 33010 17007 33013
rect 18505 33010 18571 33013
rect 16941 33008 18571 33010
rect 16941 32952 16946 33008
rect 17002 32952 18510 33008
rect 18566 32952 18571 33008
rect 16941 32950 18571 32952
rect 16941 32947 17007 32950
rect 18505 32947 18571 32950
rect 42149 33010 42215 33013
rect 42517 33010 42583 33013
rect 42149 33008 42583 33010
rect 42149 32952 42154 33008
rect 42210 32952 42522 33008
rect 42578 32952 42583 33008
rect 42149 32950 42583 32952
rect 42149 32947 42215 32950
rect 42517 32947 42583 32950
rect 17861 32874 17927 32877
rect 19793 32874 19859 32877
rect 17861 32872 19859 32874
rect 17861 32816 17866 32872
rect 17922 32816 19798 32872
rect 19854 32816 19859 32872
rect 17861 32814 19859 32816
rect 17861 32811 17927 32814
rect 19793 32811 19859 32814
rect 41689 32738 41755 32741
rect 42793 32738 42859 32741
rect 41689 32736 42859 32738
rect 41689 32680 41694 32736
rect 41750 32680 42798 32736
rect 42854 32680 42859 32736
rect 41689 32678 42859 32680
rect 41689 32675 41755 32678
rect 42793 32675 42859 32678
rect 46657 32738 46723 32741
rect 47480 32738 48280 32768
rect 46657 32736 48280 32738
rect 46657 32680 46662 32736
rect 46718 32680 48280 32736
rect 46657 32678 48280 32680
rect 46657 32675 46723 32678
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 47480 32648 48280 32678
rect 35590 32607 35906 32608
rect 18873 32602 18939 32605
rect 21541 32602 21607 32605
rect 18873 32600 21607 32602
rect 18873 32544 18878 32600
rect 18934 32544 21546 32600
rect 21602 32544 21607 32600
rect 18873 32542 21607 32544
rect 18873 32539 18939 32542
rect 21541 32539 21607 32542
rect 41597 32602 41663 32605
rect 43161 32602 43227 32605
rect 41597 32600 43227 32602
rect 41597 32544 41602 32600
rect 41658 32544 43166 32600
rect 43222 32544 43227 32600
rect 41597 32542 43227 32544
rect 41597 32539 41663 32542
rect 43161 32539 43227 32542
rect 19701 32466 19767 32469
rect 24209 32466 24275 32469
rect 19701 32464 24275 32466
rect 19701 32408 19706 32464
rect 19762 32408 24214 32464
rect 24270 32408 24275 32464
rect 19701 32406 24275 32408
rect 19701 32403 19767 32406
rect 24209 32403 24275 32406
rect 15377 32330 15443 32333
rect 15510 32330 15516 32332
rect 15377 32328 15516 32330
rect 15377 32272 15382 32328
rect 15438 32272 15516 32328
rect 15377 32270 15516 32272
rect 15377 32267 15443 32270
rect 15510 32268 15516 32270
rect 15580 32268 15586 32332
rect 16389 32330 16455 32333
rect 18137 32330 18203 32333
rect 16389 32328 18203 32330
rect 16389 32272 16394 32328
rect 16450 32272 18142 32328
rect 18198 32272 18203 32328
rect 16389 32270 18203 32272
rect 16389 32267 16455 32270
rect 18137 32267 18203 32270
rect 20897 32330 20963 32333
rect 35985 32330 36051 32333
rect 20897 32328 36051 32330
rect 20897 32272 20902 32328
rect 20958 32272 35990 32328
rect 36046 32272 36051 32328
rect 20897 32270 36051 32272
rect 20897 32267 20963 32270
rect 35985 32267 36051 32270
rect 20161 32194 20227 32197
rect 22277 32194 22343 32197
rect 25589 32194 25655 32197
rect 20161 32192 25655 32194
rect 20161 32136 20166 32192
rect 20222 32136 22282 32192
rect 22338 32136 25594 32192
rect 25650 32136 25655 32192
rect 20161 32134 25655 32136
rect 20161 32131 20227 32134
rect 22277 32131 22343 32134
rect 25589 32131 25655 32134
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 933 32058 999 32061
rect 0 32056 999 32058
rect 0 32000 938 32056
rect 994 32000 999 32056
rect 0 31998 999 32000
rect 0 31968 800 31998
rect 933 31995 999 31998
rect 18689 32058 18755 32061
rect 19241 32058 19307 32061
rect 27613 32058 27679 32061
rect 18689 32056 27679 32058
rect 18689 32000 18694 32056
rect 18750 32000 19246 32056
rect 19302 32000 27618 32056
rect 27674 32000 27679 32056
rect 18689 31998 27679 32000
rect 18689 31995 18755 31998
rect 19241 31995 19307 31998
rect 27613 31995 27679 31998
rect 28993 32058 29059 32061
rect 30373 32058 30439 32061
rect 28993 32056 30439 32058
rect 28993 32000 28998 32056
rect 29054 32000 30378 32056
rect 30434 32000 30439 32056
rect 28993 31998 30439 32000
rect 28993 31995 29059 31998
rect 30373 31995 30439 31998
rect 1669 31922 1735 31925
rect 34881 31922 34947 31925
rect 1669 31920 34947 31922
rect 1669 31864 1674 31920
rect 1730 31864 34886 31920
rect 34942 31864 34947 31920
rect 1669 31862 34947 31864
rect 1669 31859 1735 31862
rect 34881 31859 34947 31862
rect 5441 31786 5507 31789
rect 10869 31786 10935 31789
rect 5441 31784 10935 31786
rect 5441 31728 5446 31784
rect 5502 31728 10874 31784
rect 10930 31728 10935 31784
rect 5441 31726 10935 31728
rect 5441 31723 5507 31726
rect 10869 31723 10935 31726
rect 18229 31786 18295 31789
rect 23197 31786 23263 31789
rect 18229 31784 23263 31786
rect 18229 31728 18234 31784
rect 18290 31728 23202 31784
rect 23258 31728 23263 31784
rect 18229 31726 23263 31728
rect 18229 31723 18295 31726
rect 23197 31723 23263 31726
rect 20161 31650 20227 31653
rect 21173 31650 21239 31653
rect 20161 31648 21239 31650
rect 20161 31592 20166 31648
rect 20222 31592 21178 31648
rect 21234 31592 21239 31648
rect 20161 31590 21239 31592
rect 20161 31587 20227 31590
rect 21173 31587 21239 31590
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 20253 31514 20319 31517
rect 20437 31514 20503 31517
rect 20253 31512 20503 31514
rect 20253 31456 20258 31512
rect 20314 31456 20442 31512
rect 20498 31456 20503 31512
rect 20253 31454 20503 31456
rect 20253 31451 20319 31454
rect 20437 31451 20503 31454
rect 31477 31514 31543 31517
rect 35433 31514 35499 31517
rect 31477 31512 35499 31514
rect 31477 31456 31482 31512
rect 31538 31456 35438 31512
rect 35494 31456 35499 31512
rect 31477 31454 35499 31456
rect 31477 31451 31543 31454
rect 35433 31451 35499 31454
rect 20437 31378 20503 31381
rect 31017 31378 31083 31381
rect 20437 31376 31083 31378
rect 20437 31320 20442 31376
rect 20498 31320 31022 31376
rect 31078 31320 31083 31376
rect 20437 31318 31083 31320
rect 20437 31315 20503 31318
rect 31017 31315 31083 31318
rect 31845 31378 31911 31381
rect 35341 31378 35407 31381
rect 35709 31378 35775 31381
rect 31845 31376 35775 31378
rect 31845 31320 31850 31376
rect 31906 31320 35346 31376
rect 35402 31320 35714 31376
rect 35770 31320 35775 31376
rect 31845 31318 35775 31320
rect 31845 31315 31911 31318
rect 35341 31315 35407 31318
rect 35709 31315 35775 31318
rect 12525 31242 12591 31245
rect 27981 31242 28047 31245
rect 12525 31240 28047 31242
rect 12525 31184 12530 31240
rect 12586 31184 27986 31240
rect 28042 31184 28047 31240
rect 12525 31182 28047 31184
rect 12525 31179 12591 31182
rect 27981 31179 28047 31182
rect 35249 31242 35315 31245
rect 35249 31240 35450 31242
rect 35249 31184 35254 31240
rect 35310 31184 35450 31240
rect 35249 31182 35450 31184
rect 35249 31179 35315 31182
rect 35390 31106 35450 31182
rect 36537 31106 36603 31109
rect 35390 31104 36603 31106
rect 35390 31048 36542 31104
rect 36598 31048 36603 31104
rect 35390 31046 36603 31048
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 17953 30970 18019 30973
rect 18638 30970 18644 30972
rect 17953 30968 18644 30970
rect 17953 30912 17958 30968
rect 18014 30912 18644 30968
rect 17953 30910 18644 30912
rect 17953 30907 18019 30910
rect 18638 30908 18644 30910
rect 18708 30970 18714 30972
rect 18708 30910 29010 30970
rect 18708 30908 18714 30910
rect 28950 30698 29010 30910
rect 30557 30834 30623 30837
rect 33409 30834 33475 30837
rect 30557 30832 33475 30834
rect 30557 30776 30562 30832
rect 30618 30776 33414 30832
rect 33470 30776 33475 30832
rect 30557 30774 33475 30776
rect 30557 30771 30623 30774
rect 33409 30771 33475 30774
rect 35157 30834 35223 30837
rect 35390 30834 35450 31046
rect 36537 31043 36603 31046
rect 37774 30908 37780 30972
rect 37844 30970 37850 30972
rect 45829 30970 45895 30973
rect 37844 30968 45895 30970
rect 37844 30912 45834 30968
rect 45890 30912 45895 30968
rect 37844 30910 45895 30912
rect 37844 30908 37850 30910
rect 45829 30907 45895 30910
rect 35157 30832 35450 30834
rect 35157 30776 35162 30832
rect 35218 30776 35450 30832
rect 35157 30774 35450 30776
rect 35157 30771 35223 30774
rect 32857 30698 32923 30701
rect 36445 30698 36511 30701
rect 28950 30696 36511 30698
rect 28950 30640 32862 30696
rect 32918 30640 36450 30696
rect 36506 30640 36511 30696
rect 28950 30638 36511 30640
rect 32857 30635 32923 30638
rect 36445 30635 36511 30638
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 13537 30426 13603 30429
rect 13670 30426 13676 30428
rect 13537 30424 13676 30426
rect 13537 30368 13542 30424
rect 13598 30368 13676 30424
rect 13537 30366 13676 30368
rect 13537 30363 13603 30366
rect 13670 30364 13676 30366
rect 13740 30364 13746 30428
rect 19425 30154 19491 30157
rect 20529 30154 20595 30157
rect 19425 30152 20595 30154
rect 19425 30096 19430 30152
rect 19486 30096 20534 30152
rect 20590 30096 20595 30152
rect 19425 30094 20595 30096
rect 19425 30091 19491 30094
rect 20529 30091 20595 30094
rect 31477 30154 31543 30157
rect 37641 30154 37707 30157
rect 31477 30152 37707 30154
rect 31477 30096 31482 30152
rect 31538 30096 37646 30152
rect 37702 30096 37707 30152
rect 31477 30094 37707 30096
rect 31477 30091 31543 30094
rect 37641 30091 37707 30094
rect 19333 30018 19399 30021
rect 19885 30018 19951 30021
rect 19333 30016 19951 30018
rect 19333 29960 19338 30016
rect 19394 29960 19890 30016
rect 19946 29960 19951 30016
rect 19333 29958 19951 29960
rect 19333 29955 19399 29958
rect 19885 29955 19951 29958
rect 46657 30018 46723 30021
rect 47480 30018 48280 30048
rect 46657 30016 48280 30018
rect 46657 29960 46662 30016
rect 46718 29960 48280 30016
rect 46657 29958 48280 29960
rect 46657 29955 46723 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 47480 29928 48280 29958
rect 34930 29887 35246 29888
rect 19333 29882 19399 29885
rect 24117 29882 24183 29885
rect 19333 29880 24183 29882
rect 19333 29824 19338 29880
rect 19394 29824 24122 29880
rect 24178 29824 24183 29880
rect 19333 29822 24183 29824
rect 19333 29819 19399 29822
rect 24117 29819 24183 29822
rect 1669 29746 1735 29749
rect 35433 29746 35499 29749
rect 1669 29744 35499 29746
rect 1669 29688 1674 29744
rect 1730 29688 35438 29744
rect 35494 29688 35499 29744
rect 1669 29686 35499 29688
rect 1669 29683 1735 29686
rect 35433 29683 35499 29686
rect 4870 29408 5186 29409
rect 0 29338 800 29368
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 933 29338 999 29341
rect 0 29336 999 29338
rect 0 29280 938 29336
rect 994 29280 999 29336
rect 0 29278 999 29280
rect 0 29248 800 29278
rect 933 29275 999 29278
rect 13261 29338 13327 29341
rect 18321 29338 18387 29341
rect 13261 29336 18387 29338
rect 13261 29280 13266 29336
rect 13322 29280 18326 29336
rect 18382 29280 18387 29336
rect 13261 29278 18387 29280
rect 13261 29275 13327 29278
rect 18321 29275 18387 29278
rect 36813 29338 36879 29341
rect 38285 29338 38351 29341
rect 36813 29336 38351 29338
rect 36813 29280 36818 29336
rect 36874 29280 38290 29336
rect 38346 29280 38351 29336
rect 36813 29278 38351 29280
rect 36813 29275 36879 29278
rect 38285 29275 38351 29278
rect 38101 29202 38167 29205
rect 22050 29200 38167 29202
rect 22050 29144 38106 29200
rect 38162 29144 38167 29200
rect 22050 29142 38167 29144
rect 15469 29066 15535 29069
rect 22050 29066 22110 29142
rect 38101 29139 38167 29142
rect 15469 29064 22110 29066
rect 15469 29008 15474 29064
rect 15530 29008 22110 29064
rect 15469 29006 22110 29008
rect 29361 29066 29427 29069
rect 35801 29066 35867 29069
rect 29361 29064 35867 29066
rect 29361 29008 29366 29064
rect 29422 29008 35806 29064
rect 35862 29008 35867 29064
rect 29361 29006 35867 29008
rect 15469 29003 15535 29006
rect 29361 29003 29427 29006
rect 35801 29003 35867 29006
rect 37273 29066 37339 29069
rect 37590 29066 37596 29068
rect 37273 29064 37596 29066
rect 37273 29008 37278 29064
rect 37334 29008 37596 29064
rect 37273 29006 37596 29008
rect 37273 29003 37339 29006
rect 37590 29004 37596 29006
rect 37660 29004 37666 29068
rect 41137 29066 41203 29069
rect 41505 29066 41571 29069
rect 41137 29064 41571 29066
rect 41137 29008 41142 29064
rect 41198 29008 41510 29064
rect 41566 29008 41571 29064
rect 41137 29006 41571 29008
rect 41137 29003 41203 29006
rect 41505 29003 41571 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 14273 28658 14339 28661
rect 36261 28658 36327 28661
rect 14273 28656 36327 28658
rect 14273 28600 14278 28656
rect 14334 28600 36266 28656
rect 36322 28600 36327 28656
rect 14273 28598 36327 28600
rect 14273 28595 14339 28598
rect 36261 28595 36327 28598
rect 9397 28522 9463 28525
rect 46657 28522 46723 28525
rect 9397 28520 46723 28522
rect 9397 28464 9402 28520
rect 9458 28464 46662 28520
rect 46718 28464 46723 28520
rect 9397 28462 46723 28464
rect 9397 28459 9463 28462
rect 46657 28459 46723 28462
rect 11053 28386 11119 28389
rect 28993 28386 29059 28389
rect 29862 28386 29868 28388
rect 11053 28384 22110 28386
rect 11053 28328 11058 28384
rect 11114 28328 22110 28384
rect 11053 28326 22110 28328
rect 11053 28323 11119 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 20713 28250 20779 28253
rect 21030 28250 21036 28252
rect 20713 28248 21036 28250
rect 20713 28192 20718 28248
rect 20774 28192 21036 28248
rect 20713 28190 21036 28192
rect 20713 28187 20779 28190
rect 21030 28188 21036 28190
rect 21100 28188 21106 28252
rect 22050 28250 22110 28326
rect 28993 28384 29868 28386
rect 28993 28328 28998 28384
rect 29054 28328 29868 28384
rect 28993 28326 29868 28328
rect 28993 28323 29059 28326
rect 29862 28324 29868 28326
rect 29932 28324 29938 28388
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 34697 28250 34763 28253
rect 22050 28248 34763 28250
rect 22050 28192 34702 28248
rect 34758 28192 34763 28248
rect 22050 28190 34763 28192
rect 34697 28187 34763 28190
rect 19977 28114 20043 28117
rect 28257 28114 28323 28117
rect 19977 28112 28323 28114
rect 19977 28056 19982 28112
rect 20038 28056 28262 28112
rect 28318 28056 28323 28112
rect 19977 28054 28323 28056
rect 19977 28051 20043 28054
rect 28257 28051 28323 28054
rect 15469 27978 15535 27981
rect 28993 27978 29059 27981
rect 15469 27976 29059 27978
rect 15469 27920 15474 27976
rect 15530 27920 28998 27976
rect 29054 27920 29059 27976
rect 15469 27918 29059 27920
rect 15469 27915 15535 27918
rect 28993 27915 29059 27918
rect 46565 27978 46631 27981
rect 47480 27978 48280 28008
rect 46565 27976 48280 27978
rect 46565 27920 46570 27976
rect 46626 27920 48280 27976
rect 46565 27918 48280 27920
rect 46565 27915 46631 27918
rect 47480 27888 48280 27918
rect 19885 27844 19951 27845
rect 19885 27842 19932 27844
rect 19840 27840 19932 27842
rect 19840 27784 19890 27840
rect 19840 27782 19932 27784
rect 19885 27780 19932 27782
rect 19996 27780 20002 27844
rect 41413 27842 41479 27845
rect 42609 27842 42675 27845
rect 41413 27840 42675 27842
rect 41413 27784 41418 27840
rect 41474 27784 42614 27840
rect 42670 27784 42675 27840
rect 41413 27782 42675 27784
rect 19885 27779 19951 27780
rect 41413 27779 41479 27782
rect 42609 27779 42675 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 39941 27706 40007 27709
rect 45645 27706 45711 27709
rect 39941 27704 45711 27706
rect 39941 27648 39946 27704
rect 40002 27648 45650 27704
rect 45706 27648 45711 27704
rect 39941 27646 45711 27648
rect 39941 27643 40007 27646
rect 45645 27643 45711 27646
rect 23105 27434 23171 27437
rect 24209 27434 24275 27437
rect 24853 27434 24919 27437
rect 23105 27432 24919 27434
rect 23105 27376 23110 27432
rect 23166 27376 24214 27432
rect 24270 27376 24858 27432
rect 24914 27376 24919 27432
rect 23105 27374 24919 27376
rect 23105 27371 23171 27374
rect 24209 27371 24275 27374
rect 24853 27371 24919 27374
rect 14549 27298 14615 27301
rect 14917 27298 14983 27301
rect 19149 27298 19215 27301
rect 29177 27300 29243 27301
rect 29126 27298 29132 27300
rect 14549 27296 19215 27298
rect 14549 27240 14554 27296
rect 14610 27240 14922 27296
rect 14978 27240 19154 27296
rect 19210 27240 19215 27296
rect 14549 27238 19215 27240
rect 14549 27235 14615 27238
rect 14917 27235 14983 27238
rect 19149 27235 19215 27238
rect 22050 27238 29132 27298
rect 29196 27298 29243 27300
rect 29196 27296 29288 27298
rect 29238 27240 29288 27296
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 18781 27164 18847 27165
rect 18781 27162 18828 27164
rect 18736 27160 18828 27162
rect 18736 27104 18786 27160
rect 18736 27102 18828 27104
rect 18781 27100 18828 27102
rect 18892 27100 18898 27164
rect 22050 27162 22110 27238
rect 29126 27236 29132 27238
rect 29196 27238 29288 27240
rect 29196 27236 29243 27238
rect 29177 27235 29243 27236
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 35590 27167 35906 27168
rect 19014 27102 22110 27162
rect 18781 27099 18847 27100
rect 15745 27026 15811 27029
rect 19014 27026 19074 27102
rect 15745 27024 19074 27026
rect 15745 26968 15750 27024
rect 15806 26968 19074 27024
rect 15745 26966 19074 26968
rect 19149 27026 19215 27029
rect 25446 27026 25452 27028
rect 19149 27024 25452 27026
rect 19149 26968 19154 27024
rect 19210 26968 25452 27024
rect 19149 26966 25452 26968
rect 15745 26963 15811 26966
rect 19149 26963 19215 26966
rect 25446 26964 25452 26966
rect 25516 27026 25522 27028
rect 25957 27026 26023 27029
rect 25516 27024 26023 27026
rect 25516 26968 25962 27024
rect 26018 26968 26023 27024
rect 25516 26966 26023 26968
rect 25516 26964 25522 26966
rect 25957 26963 26023 26966
rect 18229 26890 18295 26893
rect 31293 26890 31359 26893
rect 18229 26888 31359 26890
rect 18229 26832 18234 26888
rect 18290 26832 31298 26888
rect 31354 26832 31359 26888
rect 18229 26830 31359 26832
rect 18229 26827 18295 26830
rect 31293 26827 31359 26830
rect 4210 26688 4526 26689
rect 0 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 933 26618 999 26621
rect 4705 26620 4771 26621
rect 0 26616 999 26618
rect 0 26560 938 26616
rect 994 26560 999 26616
rect 0 26558 999 26560
rect 0 26528 800 26558
rect 933 26555 999 26558
rect 4654 26556 4660 26620
rect 4724 26618 4771 26620
rect 9673 26618 9739 26621
rect 13813 26618 13879 26621
rect 25129 26618 25195 26621
rect 26141 26618 26207 26621
rect 4724 26616 4816 26618
rect 4766 26560 4816 26616
rect 4724 26558 4816 26560
rect 9673 26616 13879 26618
rect 9673 26560 9678 26616
rect 9734 26560 13818 26616
rect 13874 26560 13879 26616
rect 9673 26558 13879 26560
rect 4724 26556 4771 26558
rect 4705 26555 4771 26556
rect 9673 26555 9739 26558
rect 13813 26555 13879 26558
rect 20670 26616 26207 26618
rect 20670 26560 25134 26616
rect 25190 26560 26146 26616
rect 26202 26560 26207 26616
rect 20670 26558 26207 26560
rect 4705 26482 4771 26485
rect 9581 26482 9647 26485
rect 15101 26482 15167 26485
rect 20345 26484 20411 26485
rect 4705 26480 15167 26482
rect 4705 26424 4710 26480
rect 4766 26424 9586 26480
rect 9642 26424 15106 26480
rect 15162 26424 15167 26480
rect 4705 26422 15167 26424
rect 4705 26419 4771 26422
rect 9581 26419 9647 26422
rect 15101 26419 15167 26422
rect 20294 26420 20300 26484
rect 20364 26482 20411 26484
rect 20670 26482 20730 26558
rect 25129 26555 25195 26558
rect 26141 26555 26207 26558
rect 20364 26480 20730 26482
rect 20406 26424 20730 26480
rect 20364 26422 20730 26424
rect 20805 26482 20871 26485
rect 25957 26482 26023 26485
rect 20805 26480 26023 26482
rect 20805 26424 20810 26480
rect 20866 26424 25962 26480
rect 26018 26424 26023 26480
rect 20805 26422 26023 26424
rect 20364 26420 20411 26422
rect 20345 26419 20411 26420
rect 20805 26419 20871 26422
rect 25957 26419 26023 26422
rect 6821 26346 6887 26349
rect 21449 26346 21515 26349
rect 6821 26344 21515 26346
rect 6821 26288 6826 26344
rect 6882 26288 21454 26344
rect 21510 26288 21515 26344
rect 6821 26286 21515 26288
rect 6821 26283 6887 26286
rect 21449 26283 21515 26286
rect 12249 26210 12315 26213
rect 12709 26210 12775 26213
rect 12249 26208 12775 26210
rect 12249 26152 12254 26208
rect 12310 26152 12714 26208
rect 12770 26152 12775 26208
rect 12249 26150 12775 26152
rect 12249 26147 12315 26150
rect 12709 26147 12775 26150
rect 20713 26210 20779 26213
rect 32438 26210 32444 26212
rect 20713 26208 32444 26210
rect 20713 26152 20718 26208
rect 20774 26152 32444 26208
rect 20713 26150 32444 26152
rect 20713 26147 20779 26150
rect 32438 26148 32444 26150
rect 32508 26148 32514 26212
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 4521 25938 4587 25941
rect 4889 25938 4955 25941
rect 4521 25936 4955 25938
rect 4521 25880 4526 25936
rect 4582 25880 4894 25936
rect 4950 25880 4955 25936
rect 4521 25878 4955 25880
rect 32446 25938 32506 26148
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 36353 25938 36419 25941
rect 32446 25936 36419 25938
rect 32446 25880 36358 25936
rect 36414 25880 36419 25936
rect 32446 25878 36419 25880
rect 4521 25875 4587 25878
rect 4889 25875 4955 25878
rect 36353 25875 36419 25878
rect 33869 25666 33935 25669
rect 34462 25666 34468 25668
rect 33869 25664 34468 25666
rect 33869 25608 33874 25664
rect 33930 25608 34468 25664
rect 33869 25606 34468 25608
rect 33869 25603 33935 25606
rect 34462 25604 34468 25606
rect 34532 25604 34538 25668
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 12709 25530 12775 25533
rect 17309 25530 17375 25533
rect 12709 25528 17375 25530
rect 12709 25472 12714 25528
rect 12770 25472 17314 25528
rect 17370 25472 17375 25528
rect 12709 25470 17375 25472
rect 12709 25467 12775 25470
rect 17309 25467 17375 25470
rect 21265 25394 21331 25397
rect 21398 25394 21404 25396
rect 21265 25392 21404 25394
rect 21265 25336 21270 25392
rect 21326 25336 21404 25392
rect 21265 25334 21404 25336
rect 21265 25331 21331 25334
rect 21398 25332 21404 25334
rect 21468 25332 21474 25396
rect 24117 25394 24183 25397
rect 37273 25394 37339 25397
rect 24117 25392 37339 25394
rect 24117 25336 24122 25392
rect 24178 25336 37278 25392
rect 37334 25336 37339 25392
rect 24117 25334 37339 25336
rect 24117 25331 24183 25334
rect 37273 25331 37339 25334
rect 3233 25258 3299 25261
rect 36997 25258 37063 25261
rect 3233 25256 37063 25258
rect 3233 25200 3238 25256
rect 3294 25200 37002 25256
rect 37058 25200 37063 25256
rect 3233 25198 37063 25200
rect 3233 25195 3299 25198
rect 36997 25195 37063 25198
rect 45921 25258 45987 25261
rect 47480 25258 48280 25288
rect 45921 25256 48280 25258
rect 45921 25200 45926 25256
rect 45982 25200 48280 25256
rect 45921 25198 48280 25200
rect 45921 25195 45987 25198
rect 47480 25168 48280 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 34605 24852 34671 24853
rect 34605 24850 34652 24852
rect 34560 24848 34652 24850
rect 34560 24792 34610 24848
rect 34560 24790 34652 24792
rect 34605 24788 34652 24790
rect 34716 24788 34722 24852
rect 34605 24787 34671 24788
rect 1393 24714 1459 24717
rect 23105 24714 23171 24717
rect 37089 24714 37155 24717
rect 39205 24714 39271 24717
rect 1393 24712 39271 24714
rect 1393 24656 1398 24712
rect 1454 24656 23110 24712
rect 23166 24656 37094 24712
rect 37150 24656 39210 24712
rect 39266 24656 39271 24712
rect 1393 24654 39271 24656
rect 1393 24651 1459 24654
rect 23105 24651 23171 24654
rect 37089 24651 37155 24654
rect 39205 24651 39271 24654
rect 0 24578 800 24608
rect 933 24578 999 24581
rect 0 24576 999 24578
rect 0 24520 938 24576
rect 994 24520 999 24576
rect 0 24518 999 24520
rect 0 24488 800 24518
rect 933 24515 999 24518
rect 22277 24578 22343 24581
rect 29085 24578 29151 24581
rect 22277 24576 29151 24578
rect 22277 24520 22282 24576
rect 22338 24520 29090 24576
rect 29146 24520 29151 24576
rect 22277 24518 29151 24520
rect 22277 24515 22343 24518
rect 29085 24515 29151 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 17493 24306 17559 24309
rect 19057 24306 19123 24309
rect 20161 24306 20227 24309
rect 17493 24304 20227 24306
rect 17493 24248 17498 24304
rect 17554 24248 19062 24304
rect 19118 24248 20166 24304
rect 20222 24248 20227 24304
rect 17493 24246 20227 24248
rect 17493 24243 17559 24246
rect 19057 24243 19123 24246
rect 20161 24243 20227 24246
rect 41873 24306 41939 24309
rect 42517 24306 42583 24309
rect 41873 24304 42583 24306
rect 41873 24248 41878 24304
rect 41934 24248 42522 24304
rect 42578 24248 42583 24304
rect 41873 24246 42583 24248
rect 41873 24243 41939 24246
rect 42517 24243 42583 24246
rect 18781 24170 18847 24173
rect 23197 24170 23263 24173
rect 18781 24168 23263 24170
rect 18781 24112 18786 24168
rect 18842 24112 23202 24168
rect 23258 24112 23263 24168
rect 18781 24110 23263 24112
rect 18781 24107 18847 24110
rect 23197 24107 23263 24110
rect 41597 24170 41663 24173
rect 42425 24170 42491 24173
rect 42977 24170 43043 24173
rect 43253 24170 43319 24173
rect 41597 24168 43319 24170
rect 41597 24112 41602 24168
rect 41658 24112 42430 24168
rect 42486 24112 42982 24168
rect 43038 24112 43258 24168
rect 43314 24112 43319 24168
rect 41597 24110 43319 24112
rect 41597 24107 41663 24110
rect 42425 24107 42491 24110
rect 42977 24107 43043 24110
rect 43253 24107 43319 24110
rect 44909 24170 44975 24173
rect 46013 24170 46079 24173
rect 44909 24168 46079 24170
rect 44909 24112 44914 24168
rect 44970 24112 46018 24168
rect 46074 24112 46079 24168
rect 44909 24110 46079 24112
rect 44909 24107 44975 24110
rect 46013 24107 46079 24110
rect 19701 24034 19767 24037
rect 21265 24034 21331 24037
rect 19701 24032 21331 24034
rect 19701 23976 19706 24032
rect 19762 23976 21270 24032
rect 21326 23976 21331 24032
rect 19701 23974 21331 23976
rect 19701 23971 19767 23974
rect 21265 23971 21331 23974
rect 41229 24034 41295 24037
rect 42977 24034 43043 24037
rect 41229 24032 43043 24034
rect 41229 23976 41234 24032
rect 41290 23976 42982 24032
rect 43038 23976 43043 24032
rect 41229 23974 43043 23976
rect 41229 23971 41295 23974
rect 42977 23971 43043 23974
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 30649 23898 30715 23901
rect 35249 23898 35315 23901
rect 30649 23896 35315 23898
rect 30649 23840 30654 23896
rect 30710 23840 35254 23896
rect 35310 23840 35315 23896
rect 30649 23838 35315 23840
rect 30649 23835 30715 23838
rect 35249 23835 35315 23838
rect 19701 23762 19767 23765
rect 20621 23762 20687 23765
rect 19701 23760 20687 23762
rect 19701 23704 19706 23760
rect 19762 23704 20626 23760
rect 20682 23704 20687 23760
rect 19701 23702 20687 23704
rect 19701 23699 19767 23702
rect 20621 23699 20687 23702
rect 20805 23762 20871 23765
rect 21449 23762 21515 23765
rect 20805 23760 21515 23762
rect 20805 23704 20810 23760
rect 20866 23704 21454 23760
rect 21510 23704 21515 23760
rect 20805 23702 21515 23704
rect 20805 23699 20871 23702
rect 21449 23699 21515 23702
rect 29545 23762 29611 23765
rect 38285 23762 38351 23765
rect 29545 23760 38351 23762
rect 29545 23704 29550 23760
rect 29606 23704 38290 23760
rect 38346 23704 38351 23760
rect 29545 23702 38351 23704
rect 29545 23699 29611 23702
rect 38285 23699 38351 23702
rect 41689 23762 41755 23765
rect 43713 23762 43779 23765
rect 44173 23762 44239 23765
rect 41689 23760 44239 23762
rect 41689 23704 41694 23760
rect 41750 23704 43718 23760
rect 43774 23704 44178 23760
rect 44234 23704 44239 23760
rect 41689 23702 44239 23704
rect 41689 23699 41755 23702
rect 43713 23699 43779 23702
rect 44173 23699 44239 23702
rect 3785 23626 3851 23629
rect 5257 23626 5323 23629
rect 3785 23624 5323 23626
rect 3785 23568 3790 23624
rect 3846 23568 5262 23624
rect 5318 23568 5323 23624
rect 3785 23566 5323 23568
rect 3785 23563 3851 23566
rect 5257 23563 5323 23566
rect 6177 23626 6243 23629
rect 21265 23626 21331 23629
rect 6177 23624 21331 23626
rect 6177 23568 6182 23624
rect 6238 23568 21270 23624
rect 21326 23568 21331 23624
rect 6177 23566 21331 23568
rect 6177 23563 6243 23566
rect 21265 23563 21331 23566
rect 27981 23626 28047 23629
rect 30373 23626 30439 23629
rect 27981 23624 30439 23626
rect 27981 23568 27986 23624
rect 28042 23568 30378 23624
rect 30434 23568 30439 23624
rect 27981 23566 30439 23568
rect 27981 23563 28047 23566
rect 30373 23563 30439 23566
rect 5165 23490 5231 23493
rect 9397 23490 9463 23493
rect 5165 23488 9463 23490
rect 5165 23432 5170 23488
rect 5226 23432 9402 23488
rect 9458 23432 9463 23488
rect 5165 23430 9463 23432
rect 5165 23427 5231 23430
rect 9397 23427 9463 23430
rect 28533 23490 28599 23493
rect 29545 23490 29611 23493
rect 28533 23488 29611 23490
rect 28533 23432 28538 23488
rect 28594 23432 29550 23488
rect 29606 23432 29611 23488
rect 28533 23430 29611 23432
rect 28533 23427 28599 23430
rect 29545 23427 29611 23430
rect 38469 23492 38535 23493
rect 38469 23488 38516 23492
rect 38580 23490 38586 23492
rect 38469 23432 38474 23488
rect 38469 23428 38516 23432
rect 38580 23430 38626 23490
rect 38580 23428 38586 23430
rect 38469 23427 38535 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 5441 23354 5507 23357
rect 6085 23354 6151 23357
rect 5398 23352 5507 23354
rect 5398 23296 5446 23352
rect 5502 23296 5507 23352
rect 5398 23291 5507 23296
rect 5766 23352 6151 23354
rect 5766 23296 6090 23352
rect 6146 23296 6151 23352
rect 5766 23294 6151 23296
rect 5398 22949 5458 23291
rect 5766 23221 5826 23294
rect 6085 23291 6151 23294
rect 11145 23354 11211 23357
rect 18781 23354 18847 23357
rect 11145 23352 18847 23354
rect 11145 23296 11150 23352
rect 11206 23296 18786 23352
rect 18842 23296 18847 23352
rect 11145 23294 18847 23296
rect 11145 23291 11211 23294
rect 18781 23291 18847 23294
rect 20621 23354 20687 23357
rect 23197 23354 23263 23357
rect 20621 23352 23263 23354
rect 20621 23296 20626 23352
rect 20682 23296 23202 23352
rect 23258 23296 23263 23352
rect 20621 23294 23263 23296
rect 20621 23291 20687 23294
rect 23197 23291 23263 23294
rect 5717 23216 5826 23221
rect 5717 23160 5722 23216
rect 5778 23160 5826 23216
rect 5717 23158 5826 23160
rect 13169 23218 13235 23221
rect 18045 23218 18111 23221
rect 13169 23216 18111 23218
rect 13169 23160 13174 23216
rect 13230 23160 18050 23216
rect 18106 23160 18111 23216
rect 13169 23158 18111 23160
rect 5717 23155 5783 23158
rect 13169 23155 13235 23158
rect 18045 23155 18111 23158
rect 32254 23156 32260 23220
rect 32324 23218 32330 23220
rect 37825 23218 37891 23221
rect 32324 23216 37891 23218
rect 32324 23160 37830 23216
rect 37886 23160 37891 23216
rect 32324 23158 37891 23160
rect 32324 23156 32330 23158
rect 37825 23155 37891 23158
rect 39481 23218 39547 23221
rect 43621 23218 43687 23221
rect 39481 23216 43687 23218
rect 39481 23160 39486 23216
rect 39542 23160 43626 23216
rect 43682 23160 43687 23216
rect 39481 23158 43687 23160
rect 39481 23155 39547 23158
rect 43621 23155 43687 23158
rect 46565 23218 46631 23221
rect 47480 23218 48280 23248
rect 46565 23216 48280 23218
rect 46565 23160 46570 23216
rect 46626 23160 48280 23216
rect 46565 23158 48280 23160
rect 46565 23155 46631 23158
rect 47480 23128 48280 23158
rect 5398 22944 5507 22949
rect 5398 22888 5446 22944
rect 5502 22888 5507 22944
rect 5398 22886 5507 22888
rect 5441 22883 5507 22886
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 4521 22674 4587 22677
rect 5257 22674 5323 22677
rect 4521 22672 5323 22674
rect 4521 22616 4526 22672
rect 4582 22616 5262 22672
rect 5318 22616 5323 22672
rect 4521 22614 5323 22616
rect 4521 22611 4587 22614
rect 5257 22611 5323 22614
rect 38745 22674 38811 22677
rect 38878 22674 38884 22676
rect 38745 22672 38884 22674
rect 38745 22616 38750 22672
rect 38806 22616 38884 22672
rect 38745 22614 38884 22616
rect 38745 22611 38811 22614
rect 38878 22612 38884 22614
rect 38948 22612 38954 22676
rect 39113 22404 39179 22405
rect 39062 22402 39068 22404
rect 39022 22342 39068 22402
rect 39132 22400 39179 22404
rect 39174 22344 39179 22400
rect 39062 22340 39068 22342
rect 39132 22340 39179 22344
rect 39113 22339 39179 22340
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 38929 22266 38995 22269
rect 39113 22266 39179 22269
rect 38929 22264 39179 22266
rect 38929 22208 38934 22264
rect 38990 22208 39118 22264
rect 39174 22208 39179 22264
rect 38929 22206 39179 22208
rect 38929 22203 38995 22206
rect 39113 22203 39179 22206
rect 25221 22130 25287 22133
rect 31569 22130 31635 22133
rect 10550 22070 10978 22130
rect 10133 21994 10199 21997
rect 10550 21994 10610 22070
rect 10133 21992 10610 21994
rect 10133 21936 10138 21992
rect 10194 21936 10610 21992
rect 10133 21934 10610 21936
rect 10685 21994 10751 21997
rect 10685 21992 10794 21994
rect 10685 21936 10690 21992
rect 10746 21936 10794 21992
rect 10133 21931 10199 21934
rect 10685 21931 10794 21936
rect 0 21858 800 21888
rect 933 21858 999 21861
rect 0 21856 999 21858
rect 0 21800 938 21856
rect 994 21800 999 21856
rect 0 21798 999 21800
rect 0 21768 800 21798
rect 933 21795 999 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 10501 21722 10567 21725
rect 10734 21722 10794 21931
rect 10918 21858 10978 22070
rect 25221 22128 31635 22130
rect 25221 22072 25226 22128
rect 25282 22072 31574 22128
rect 31630 22072 31635 22128
rect 25221 22070 31635 22072
rect 25221 22067 25287 22070
rect 31569 22067 31635 22070
rect 11789 21994 11855 21997
rect 34646 21994 34652 21996
rect 11789 21992 34652 21994
rect 11789 21936 11794 21992
rect 11850 21936 34652 21992
rect 11789 21934 34652 21936
rect 11789 21931 11855 21934
rect 34646 21932 34652 21934
rect 34716 21994 34722 21996
rect 34973 21994 35039 21997
rect 34716 21992 35039 21994
rect 34716 21936 34978 21992
rect 35034 21936 35039 21992
rect 34716 21934 35039 21936
rect 34716 21932 34722 21934
rect 34973 21931 35039 21934
rect 19609 21858 19675 21861
rect 25405 21860 25471 21861
rect 25405 21858 25452 21860
rect 10918 21856 19675 21858
rect 10918 21800 19614 21856
rect 19670 21800 19675 21856
rect 10918 21798 19675 21800
rect 25360 21856 25452 21858
rect 25360 21800 25410 21856
rect 25360 21798 25452 21800
rect 19609 21795 19675 21798
rect 25405 21796 25452 21798
rect 25516 21796 25522 21860
rect 25957 21858 26023 21861
rect 29269 21858 29335 21861
rect 30230 21858 30236 21860
rect 25957 21856 30236 21858
rect 25957 21800 25962 21856
rect 26018 21800 29274 21856
rect 29330 21800 30236 21856
rect 25957 21798 30236 21800
rect 25405 21795 25471 21796
rect 25957 21795 26023 21798
rect 29269 21795 29335 21798
rect 30230 21796 30236 21798
rect 30300 21796 30306 21860
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 19926 21722 19932 21724
rect 10501 21720 19932 21722
rect 10501 21664 10506 21720
rect 10562 21664 19932 21720
rect 10501 21662 19932 21664
rect 10501 21659 10567 21662
rect 19926 21660 19932 21662
rect 19996 21660 20002 21724
rect 25681 21722 25747 21725
rect 26049 21722 26115 21725
rect 25681 21720 26115 21722
rect 25681 21664 25686 21720
rect 25742 21664 26054 21720
rect 26110 21664 26115 21720
rect 25681 21662 26115 21664
rect 25681 21659 25747 21662
rect 26049 21659 26115 21662
rect 18321 21586 18387 21589
rect 19057 21586 19123 21589
rect 33869 21586 33935 21589
rect 18321 21584 19123 21586
rect 18321 21528 18326 21584
rect 18382 21528 19062 21584
rect 19118 21528 19123 21584
rect 18321 21526 19123 21528
rect 18321 21523 18387 21526
rect 19057 21523 19123 21526
rect 22050 21584 33935 21586
rect 22050 21528 33874 21584
rect 33930 21528 33935 21584
rect 22050 21526 33935 21528
rect 15745 21450 15811 21453
rect 22050 21450 22110 21526
rect 33869 21523 33935 21526
rect 15745 21448 22110 21450
rect 15745 21392 15750 21448
rect 15806 21392 22110 21448
rect 15745 21390 22110 21392
rect 22185 21450 22251 21453
rect 40125 21450 40191 21453
rect 22185 21448 40191 21450
rect 22185 21392 22190 21448
rect 22246 21392 40130 21448
rect 40186 21392 40191 21448
rect 22185 21390 40191 21392
rect 15745 21387 15811 21390
rect 22185 21387 22251 21390
rect 40125 21387 40191 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 29637 21042 29703 21045
rect 34145 21042 34211 21045
rect 29637 21040 34211 21042
rect 29637 20984 29642 21040
rect 29698 20984 34150 21040
rect 34206 20984 34211 21040
rect 29637 20982 34211 20984
rect 29637 20979 29703 20982
rect 34145 20979 34211 20982
rect 33501 20906 33567 20909
rect 34237 20906 34303 20909
rect 33501 20904 34303 20906
rect 33501 20848 33506 20904
rect 33562 20848 34242 20904
rect 34298 20848 34303 20904
rect 33501 20846 34303 20848
rect 33501 20843 33567 20846
rect 34237 20843 34303 20846
rect 19609 20770 19675 20773
rect 20529 20770 20595 20773
rect 19609 20768 20595 20770
rect 19609 20712 19614 20768
rect 19670 20712 20534 20768
rect 20590 20712 20595 20768
rect 19609 20710 20595 20712
rect 19609 20707 19675 20710
rect 20529 20707 20595 20710
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 39481 20636 39547 20637
rect 39430 20634 39436 20636
rect 39390 20574 39436 20634
rect 39500 20632 39547 20636
rect 39542 20576 39547 20632
rect 39430 20572 39436 20574
rect 39500 20572 39547 20576
rect 39481 20571 39547 20572
rect 34462 20436 34468 20500
rect 34532 20498 34538 20500
rect 34697 20498 34763 20501
rect 34532 20496 34763 20498
rect 34532 20440 34702 20496
rect 34758 20440 34763 20496
rect 34532 20438 34763 20440
rect 34532 20436 34538 20438
rect 34697 20435 34763 20438
rect 46657 20498 46723 20501
rect 47480 20498 48280 20528
rect 46657 20496 48280 20498
rect 46657 20440 46662 20496
rect 46718 20440 48280 20496
rect 46657 20438 48280 20440
rect 46657 20435 46723 20438
rect 47480 20408 48280 20438
rect 23289 20362 23355 20365
rect 30005 20362 30071 20365
rect 23289 20360 30071 20362
rect 23289 20304 23294 20360
rect 23350 20304 30010 20360
rect 30066 20304 30071 20360
rect 23289 20302 30071 20304
rect 23289 20299 23355 20302
rect 30005 20299 30071 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 4654 20028 4660 20092
rect 4724 20090 4730 20092
rect 5165 20090 5231 20093
rect 4724 20088 9690 20090
rect 4724 20032 5170 20088
rect 5226 20032 9690 20088
rect 4724 20030 9690 20032
rect 4724 20028 4730 20030
rect 5165 20027 5231 20030
rect 9630 19954 9690 20030
rect 10501 19954 10567 19957
rect 9630 19952 10567 19954
rect 9630 19896 10506 19952
rect 10562 19896 10567 19952
rect 9630 19894 10567 19896
rect 10501 19891 10567 19894
rect 17125 19954 17191 19957
rect 31845 19954 31911 19957
rect 17125 19952 31911 19954
rect 17125 19896 17130 19952
rect 17186 19896 31850 19952
rect 31906 19896 31911 19952
rect 17125 19894 31911 19896
rect 17125 19891 17191 19894
rect 31845 19891 31911 19894
rect 0 19818 800 19848
rect 1301 19818 1367 19821
rect 0 19816 1367 19818
rect 0 19760 1306 19816
rect 1362 19760 1367 19816
rect 0 19758 1367 19760
rect 0 19728 800 19758
rect 1301 19755 1367 19758
rect 21173 19818 21239 19821
rect 39062 19818 39068 19820
rect 21173 19816 39068 19818
rect 21173 19760 21178 19816
rect 21234 19760 39068 19816
rect 21173 19758 39068 19760
rect 21173 19755 21239 19758
rect 39062 19756 39068 19758
rect 39132 19818 39138 19820
rect 40585 19818 40651 19821
rect 39132 19816 40651 19818
rect 39132 19760 40590 19816
rect 40646 19760 40651 19816
rect 39132 19758 40651 19760
rect 39132 19756 39138 19758
rect 40585 19755 40651 19758
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 15510 19212 15516 19276
rect 15580 19274 15586 19276
rect 33777 19274 33843 19277
rect 34881 19274 34947 19277
rect 15580 19272 34947 19274
rect 15580 19216 33782 19272
rect 33838 19216 34886 19272
rect 34942 19216 34947 19272
rect 15580 19214 34947 19216
rect 15580 19212 15586 19214
rect 33777 19211 33843 19214
rect 34881 19211 34947 19214
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 20989 19002 21055 19005
rect 27337 19002 27403 19005
rect 20989 19000 27403 19002
rect 20989 18944 20994 19000
rect 21050 18944 27342 19000
rect 27398 18944 27403 19000
rect 20989 18942 27403 18944
rect 20989 18939 21055 18942
rect 27337 18939 27403 18942
rect 38653 18866 38719 18869
rect 39430 18866 39436 18868
rect 38653 18864 39436 18866
rect 38653 18808 38658 18864
rect 38714 18808 39436 18864
rect 38653 18806 39436 18808
rect 38653 18803 38719 18806
rect 39430 18804 39436 18806
rect 39500 18804 39506 18868
rect 26325 18730 26391 18733
rect 26601 18730 26667 18733
rect 26325 18728 26667 18730
rect 26325 18672 26330 18728
rect 26386 18672 26606 18728
rect 26662 18672 26667 18728
rect 26325 18670 26667 18672
rect 26325 18667 26391 18670
rect 26601 18667 26667 18670
rect 30005 18730 30071 18733
rect 33777 18730 33843 18733
rect 36169 18730 36235 18733
rect 30005 18728 36235 18730
rect 30005 18672 30010 18728
rect 30066 18672 33782 18728
rect 33838 18672 36174 18728
rect 36230 18672 36235 18728
rect 30005 18670 36235 18672
rect 30005 18667 30071 18670
rect 33777 18667 33843 18670
rect 36169 18667 36235 18670
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 29177 18322 29243 18325
rect 30046 18322 30052 18324
rect 29177 18320 30052 18322
rect 29177 18264 29182 18320
rect 29238 18264 30052 18320
rect 29177 18262 30052 18264
rect 29177 18259 29243 18262
rect 30046 18260 30052 18262
rect 30116 18322 30122 18324
rect 30281 18322 30347 18325
rect 30116 18320 30347 18322
rect 30116 18264 30286 18320
rect 30342 18264 30347 18320
rect 30116 18262 30347 18264
rect 30116 18260 30122 18262
rect 30281 18259 30347 18262
rect 3049 18186 3115 18189
rect 12934 18186 12940 18188
rect 3049 18184 12940 18186
rect 3049 18128 3054 18184
rect 3110 18128 12940 18184
rect 3049 18126 12940 18128
rect 3049 18123 3115 18126
rect 12934 18124 12940 18126
rect 13004 18124 13010 18188
rect 22001 18186 22067 18189
rect 22461 18186 22527 18189
rect 22001 18184 22527 18186
rect 22001 18128 22006 18184
rect 22062 18128 22466 18184
rect 22522 18128 22527 18184
rect 22001 18126 22527 18128
rect 22001 18123 22067 18126
rect 22461 18123 22527 18126
rect 15510 17988 15516 18052
rect 15580 18050 15586 18052
rect 16113 18050 16179 18053
rect 15580 18048 16179 18050
rect 15580 17992 16118 18048
rect 16174 17992 16179 18048
rect 15580 17990 16179 17992
rect 15580 17988 15586 17990
rect 16113 17987 16179 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 11053 17914 11119 17917
rect 17033 17914 17099 17917
rect 11053 17912 17099 17914
rect 11053 17856 11058 17912
rect 11114 17856 17038 17912
rect 17094 17856 17099 17912
rect 11053 17854 17099 17856
rect 11053 17851 11119 17854
rect 17033 17851 17099 17854
rect 14089 17778 14155 17781
rect 18229 17778 18295 17781
rect 14089 17776 18295 17778
rect 14089 17720 14094 17776
rect 14150 17720 18234 17776
rect 18290 17720 18295 17776
rect 14089 17718 18295 17720
rect 14089 17715 14155 17718
rect 18229 17715 18295 17718
rect 42190 17716 42196 17780
rect 42260 17778 42266 17780
rect 46381 17778 46447 17781
rect 42260 17776 46447 17778
rect 42260 17720 46386 17776
rect 46442 17720 46447 17776
rect 42260 17718 46447 17720
rect 42260 17716 42266 17718
rect 46381 17715 46447 17718
rect 46749 17778 46815 17781
rect 47480 17778 48280 17808
rect 46749 17776 48280 17778
rect 46749 17720 46754 17776
rect 46810 17720 48280 17776
rect 46749 17718 48280 17720
rect 46749 17715 46815 17718
rect 47480 17688 48280 17718
rect 4245 17642 4311 17645
rect 5165 17642 5231 17645
rect 4245 17640 5231 17642
rect 4245 17584 4250 17640
rect 4306 17584 5170 17640
rect 5226 17584 5231 17640
rect 4245 17582 5231 17584
rect 4245 17579 4311 17582
rect 5165 17579 5231 17582
rect 15469 17642 15535 17645
rect 17033 17642 17099 17645
rect 15469 17640 17099 17642
rect 15469 17584 15474 17640
rect 15530 17584 17038 17640
rect 17094 17584 17099 17640
rect 15469 17582 17099 17584
rect 15469 17579 15535 17582
rect 17033 17579 17099 17582
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 1577 17234 1643 17237
rect 37273 17234 37339 17237
rect 1577 17232 37339 17234
rect 1577 17176 1582 17232
rect 1638 17176 37278 17232
rect 37334 17176 37339 17232
rect 1577 17174 37339 17176
rect 1577 17171 1643 17174
rect 37273 17171 37339 17174
rect 0 17098 800 17128
rect 933 17098 999 17101
rect 0 17096 999 17098
rect 0 17040 938 17096
rect 994 17040 999 17096
rect 0 17038 999 17040
rect 0 17008 800 17038
rect 933 17035 999 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 38101 16692 38167 16693
rect 38101 16688 38148 16692
rect 38212 16690 38218 16692
rect 38101 16632 38106 16688
rect 38101 16628 38148 16632
rect 38212 16630 38258 16690
rect 38212 16628 38218 16630
rect 38101 16627 38167 16628
rect 20345 16556 20411 16557
rect 20294 16554 20300 16556
rect 20254 16494 20300 16554
rect 20364 16552 20411 16556
rect 20406 16496 20411 16552
rect 20294 16492 20300 16494
rect 20364 16492 20411 16496
rect 20345 16491 20411 16492
rect 20897 16554 20963 16557
rect 21030 16554 21036 16556
rect 20897 16552 21036 16554
rect 20897 16496 20902 16552
rect 20958 16496 21036 16552
rect 20897 16494 21036 16496
rect 20897 16491 20963 16494
rect 21030 16492 21036 16494
rect 21100 16492 21106 16556
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 12065 16146 12131 16149
rect 14457 16146 14523 16149
rect 12065 16144 14523 16146
rect 12065 16088 12070 16144
rect 12126 16088 14462 16144
rect 14518 16088 14523 16144
rect 12065 16086 14523 16088
rect 12065 16083 12131 16086
rect 14457 16083 14523 16086
rect 28993 16146 29059 16149
rect 29126 16146 29132 16148
rect 28993 16144 29132 16146
rect 28993 16088 28998 16144
rect 29054 16088 29132 16144
rect 28993 16086 29132 16088
rect 28993 16083 29059 16086
rect 29126 16084 29132 16086
rect 29196 16084 29202 16148
rect 22829 16010 22895 16013
rect 37549 16010 37615 16013
rect 22829 16008 37615 16010
rect 22829 15952 22834 16008
rect 22890 15952 37554 16008
rect 37610 15952 37615 16008
rect 22829 15950 37615 15952
rect 22829 15947 22895 15950
rect 37549 15947 37615 15950
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 46657 15738 46723 15741
rect 47480 15738 48280 15768
rect 46657 15736 48280 15738
rect 46657 15680 46662 15736
rect 46718 15680 48280 15736
rect 46657 15678 48280 15680
rect 46657 15675 46723 15678
rect 47480 15648 48280 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 18822 15132 18828 15196
rect 18892 15194 18898 15196
rect 19742 15194 19748 15196
rect 18892 15134 19748 15194
rect 18892 15132 18898 15134
rect 19742 15132 19748 15134
rect 19812 15132 19818 15196
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19742 14452 19748 14516
rect 19812 14514 19818 14516
rect 26601 14514 26667 14517
rect 19812 14512 26667 14514
rect 19812 14456 26606 14512
rect 26662 14456 26667 14512
rect 19812 14454 26667 14456
rect 19812 14452 19818 14454
rect 26601 14451 26667 14454
rect 0 14378 800 14408
rect 933 14378 999 14381
rect 0 14376 999 14378
rect 0 14320 938 14376
rect 994 14320 999 14376
rect 0 14318 999 14320
rect 0 14288 800 14318
rect 933 14315 999 14318
rect 20529 14378 20595 14381
rect 27153 14378 27219 14381
rect 20529 14376 27219 14378
rect 20529 14320 20534 14376
rect 20590 14320 27158 14376
rect 27214 14320 27219 14376
rect 20529 14318 27219 14320
rect 20529 14315 20595 14318
rect 27153 14315 27219 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 29494 13772 29500 13836
rect 29564 13834 29570 13836
rect 30230 13834 30236 13836
rect 29564 13774 30236 13834
rect 29564 13772 29570 13774
rect 30230 13772 30236 13774
rect 30300 13834 30306 13836
rect 30373 13834 30439 13837
rect 30300 13832 30439 13834
rect 30300 13776 30378 13832
rect 30434 13776 30439 13832
rect 30300 13774 30439 13776
rect 30300 13772 30306 13774
rect 30373 13771 30439 13774
rect 33777 13834 33843 13837
rect 34094 13834 34100 13836
rect 33777 13832 34100 13834
rect 33777 13776 33782 13832
rect 33838 13776 34100 13832
rect 33777 13774 34100 13776
rect 33777 13771 33843 13774
rect 34094 13772 34100 13774
rect 34164 13772 34170 13836
rect 19926 13636 19932 13700
rect 19996 13698 20002 13700
rect 23565 13698 23631 13701
rect 19996 13696 23631 13698
rect 19996 13640 23570 13696
rect 23626 13640 23631 13696
rect 19996 13638 23631 13640
rect 19996 13636 20002 13638
rect 23565 13635 23631 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 46657 13018 46723 13021
rect 47480 13018 48280 13048
rect 46657 13016 48280 13018
rect 46657 12960 46662 13016
rect 46718 12960 48280 13016
rect 46657 12958 48280 12960
rect 46657 12955 46723 12958
rect 47480 12928 48280 12958
rect 23657 12882 23723 12885
rect 24945 12882 25011 12885
rect 23657 12880 25011 12882
rect 23657 12824 23662 12880
rect 23718 12824 24950 12880
rect 25006 12824 25011 12880
rect 23657 12822 25011 12824
rect 23657 12819 23723 12822
rect 24945 12819 25011 12822
rect 27705 12882 27771 12885
rect 30373 12882 30439 12885
rect 27705 12880 30439 12882
rect 27705 12824 27710 12880
rect 27766 12824 30378 12880
rect 30434 12824 30439 12880
rect 27705 12822 30439 12824
rect 27705 12819 27771 12822
rect 30373 12819 30439 12822
rect 1669 12746 1735 12749
rect 30281 12746 30347 12749
rect 1669 12744 30347 12746
rect 1669 12688 1674 12744
rect 1730 12688 30286 12744
rect 30342 12688 30347 12744
rect 1669 12686 30347 12688
rect 1669 12683 1735 12686
rect 30281 12683 30347 12686
rect 8201 12610 8267 12613
rect 21081 12610 21147 12613
rect 8201 12608 21147 12610
rect 8201 12552 8206 12608
rect 8262 12552 21086 12608
rect 21142 12552 21147 12608
rect 8201 12550 21147 12552
rect 8201 12547 8267 12550
rect 21081 12547 21147 12550
rect 31477 12610 31543 12613
rect 34053 12610 34119 12613
rect 31477 12608 34119 12610
rect 31477 12552 31482 12608
rect 31538 12552 34058 12608
rect 34114 12552 34119 12608
rect 31477 12550 34119 12552
rect 31477 12547 31543 12550
rect 34053 12547 34119 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 29913 12340 29979 12341
rect 29862 12338 29868 12340
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 29822 12278 29868 12338
rect 29932 12336 29979 12340
rect 29974 12280 29979 12336
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 29862 12276 29868 12278
rect 29932 12276 29979 12280
rect 29913 12275 29979 12276
rect 20713 12202 20779 12205
rect 38561 12202 38627 12205
rect 39205 12202 39271 12205
rect 20713 12200 39271 12202
rect 20713 12144 20718 12200
rect 20774 12144 38566 12200
rect 38622 12144 39210 12200
rect 39266 12144 39271 12200
rect 20713 12142 39271 12144
rect 20713 12139 20779 12142
rect 38561 12139 38627 12142
rect 39205 12139 39271 12142
rect 42701 12202 42767 12205
rect 43621 12202 43687 12205
rect 42701 12200 43687 12202
rect 42701 12144 42706 12200
rect 42762 12144 43626 12200
rect 43682 12144 43687 12200
rect 42701 12142 43687 12144
rect 42701 12139 42767 12142
rect 43621 12139 43687 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 38745 11794 38811 11797
rect 43069 11794 43135 11797
rect 38745 11792 43135 11794
rect 38745 11736 38750 11792
rect 38806 11736 43074 11792
rect 43130 11736 43135 11792
rect 38745 11734 43135 11736
rect 38745 11731 38811 11734
rect 43069 11731 43135 11734
rect 40769 11658 40835 11661
rect 41321 11658 41387 11661
rect 43253 11658 43319 11661
rect 40769 11656 43319 11658
rect 40769 11600 40774 11656
rect 40830 11600 41326 11656
rect 41382 11600 43258 11656
rect 43314 11600 43319 11656
rect 40769 11598 43319 11600
rect 40769 11595 40835 11598
rect 41321 11595 41387 11598
rect 43253 11595 43319 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 20805 11250 20871 11253
rect 37733 11250 37799 11253
rect 38377 11250 38443 11253
rect 20805 11248 38443 11250
rect 20805 11192 20810 11248
rect 20866 11192 37738 11248
rect 37794 11192 38382 11248
rect 38438 11192 38443 11248
rect 20805 11190 38443 11192
rect 20805 11187 20871 11190
rect 37733 11187 37799 11190
rect 38377 11187 38443 11190
rect 25405 11114 25471 11117
rect 35985 11114 36051 11117
rect 25405 11112 36051 11114
rect 25405 11056 25410 11112
rect 25466 11056 35990 11112
rect 36046 11056 36051 11112
rect 25405 11054 36051 11056
rect 25405 11051 25471 11054
rect 35985 11051 36051 11054
rect 42609 11114 42675 11117
rect 42885 11114 42951 11117
rect 43529 11114 43595 11117
rect 42609 11112 43595 11114
rect 42609 11056 42614 11112
rect 42670 11056 42890 11112
rect 42946 11056 43534 11112
rect 43590 11056 43595 11112
rect 42609 11054 43595 11056
rect 42609 11051 42675 11054
rect 42885 11051 42951 11054
rect 43529 11051 43595 11054
rect 29821 10978 29887 10981
rect 30046 10978 30052 10980
rect 29821 10976 30052 10978
rect 29821 10920 29826 10976
rect 29882 10920 30052 10976
rect 29821 10918 30052 10920
rect 29821 10915 29887 10918
rect 30046 10916 30052 10918
rect 30116 10916 30122 10980
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 26918 10508 26924 10572
rect 26988 10570 26994 10572
rect 39849 10570 39915 10573
rect 26988 10568 39915 10570
rect 26988 10512 39854 10568
rect 39910 10512 39915 10568
rect 26988 10510 39915 10512
rect 26988 10508 26994 10510
rect 39849 10507 39915 10510
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 46657 10298 46723 10301
rect 47480 10298 48280 10328
rect 46657 10296 48280 10298
rect 46657 10240 46662 10296
rect 46718 10240 48280 10296
rect 46657 10238 48280 10240
rect 46657 10235 46723 10238
rect 47480 10208 48280 10238
rect 21633 10162 21699 10165
rect 22185 10162 22251 10165
rect 21633 10160 22251 10162
rect 21633 10104 21638 10160
rect 21694 10104 22190 10160
rect 22246 10104 22251 10160
rect 21633 10102 22251 10104
rect 21633 10099 21699 10102
rect 22185 10099 22251 10102
rect 2221 10026 2287 10029
rect 23749 10026 23815 10029
rect 2221 10024 23815 10026
rect 2221 9968 2226 10024
rect 2282 9968 23754 10024
rect 23810 9968 23815 10024
rect 2221 9966 23815 9968
rect 2221 9963 2287 9966
rect 23749 9963 23815 9966
rect 20069 9890 20135 9893
rect 21541 9890 21607 9893
rect 20069 9888 21607 9890
rect 20069 9832 20074 9888
rect 20130 9832 21546 9888
rect 21602 9832 21607 9888
rect 20069 9830 21607 9832
rect 20069 9827 20135 9830
rect 21541 9827 21607 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 13353 9754 13419 9757
rect 21173 9754 21239 9757
rect 13353 9752 21239 9754
rect 13353 9696 13358 9752
rect 13414 9696 21178 9752
rect 21234 9696 21239 9752
rect 13353 9694 21239 9696
rect 13353 9691 13419 9694
rect 21173 9691 21239 9694
rect 0 9618 800 9648
rect 1577 9618 1643 9621
rect 0 9616 1643 9618
rect 0 9560 1582 9616
rect 1638 9560 1643 9616
rect 0 9558 1643 9560
rect 0 9528 800 9558
rect 1577 9555 1643 9558
rect 34646 9556 34652 9620
rect 34716 9618 34722 9620
rect 34789 9618 34855 9621
rect 34716 9616 34855 9618
rect 34716 9560 34794 9616
rect 34850 9560 34855 9616
rect 34716 9558 34855 9560
rect 34716 9556 34722 9558
rect 34789 9555 34855 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 15193 9074 15259 9077
rect 25037 9074 25103 9077
rect 15193 9072 25103 9074
rect 15193 9016 15198 9072
rect 15254 9016 25042 9072
rect 25098 9016 25103 9072
rect 15193 9014 25103 9016
rect 15193 9011 15259 9014
rect 25037 9011 25103 9014
rect 15745 8938 15811 8941
rect 25589 8938 25655 8941
rect 15745 8936 25655 8938
rect 15745 8880 15750 8936
rect 15806 8880 25594 8936
rect 25650 8880 25655 8936
rect 15745 8878 25655 8880
rect 15745 8875 15811 8878
rect 25589 8875 25655 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 19701 8396 19767 8397
rect 19701 8394 19748 8396
rect 19382 8392 19748 8394
rect 19382 8336 19706 8392
rect 19382 8334 19748 8336
rect 17861 8258 17927 8261
rect 19382 8258 19442 8334
rect 19701 8332 19748 8334
rect 19812 8332 19818 8396
rect 19701 8331 19767 8332
rect 17861 8256 19442 8258
rect 17861 8200 17866 8256
rect 17922 8200 19442 8256
rect 17861 8198 19442 8200
rect 45921 8258 45987 8261
rect 47480 8258 48280 8288
rect 45921 8256 48280 8258
rect 45921 8200 45926 8256
rect 45982 8200 48280 8256
rect 45921 8198 48280 8200
rect 17861 8195 17927 8198
rect 45921 8195 45987 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 47480 8168 48280 8198
rect 34930 8127 35246 8128
rect 22461 8122 22527 8125
rect 33133 8122 33199 8125
rect 22461 8120 33199 8122
rect 22461 8064 22466 8120
rect 22522 8064 33138 8120
rect 33194 8064 33199 8120
rect 22461 8062 33199 8064
rect 22461 8059 22527 8062
rect 33133 8059 33199 8062
rect 29494 7924 29500 7988
rect 29564 7986 29570 7988
rect 30189 7986 30255 7989
rect 29564 7984 30255 7986
rect 29564 7928 30194 7984
rect 30250 7928 30255 7984
rect 29564 7926 30255 7928
rect 29564 7924 29570 7926
rect 30189 7923 30255 7926
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 34094 7380 34100 7444
rect 34164 7442 34170 7444
rect 34237 7442 34303 7445
rect 34164 7440 34303 7442
rect 34164 7384 34242 7440
rect 34298 7384 34303 7440
rect 34164 7382 34303 7384
rect 34164 7380 34170 7382
rect 34237 7379 34303 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 800 6838
rect 1577 6835 1643 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 32622 6156 32628 6220
rect 32692 6218 32698 6220
rect 45553 6218 45619 6221
rect 32692 6216 45619 6218
rect 32692 6160 45558 6216
rect 45614 6160 45619 6216
rect 32692 6158 45619 6160
rect 32692 6156 32698 6158
rect 45553 6155 45619 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 20897 5674 20963 5677
rect 22645 5674 22711 5677
rect 20897 5672 22711 5674
rect 20897 5616 20902 5672
rect 20958 5616 22650 5672
rect 22706 5616 22711 5672
rect 20897 5614 22711 5616
rect 20897 5611 20963 5614
rect 22645 5611 22711 5614
rect 46657 5538 46723 5541
rect 47480 5538 48280 5568
rect 46657 5536 48280 5538
rect 46657 5480 46662 5536
rect 46718 5480 48280 5536
rect 46657 5478 48280 5480
rect 46657 5475 46723 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 47480 5448 48280 5478
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 32673 4722 32739 4725
rect 33317 4722 33383 4725
rect 32673 4720 33383 4722
rect 32673 4664 32678 4720
rect 32734 4664 33322 4720
rect 33378 4664 33383 4720
rect 32673 4662 33383 4664
rect 32673 4659 32739 4662
rect 33317 4659 33383 4662
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 27102 3980 27108 4044
rect 27172 4042 27178 4044
rect 39205 4042 39271 4045
rect 27172 4040 39271 4042
rect 27172 3984 39210 4040
rect 39266 3984 39271 4040
rect 27172 3982 39271 3984
rect 27172 3980 27178 3982
rect 39205 3979 39271 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 18597 3636 18663 3637
rect 18597 3634 18644 3636
rect 18552 3632 18644 3634
rect 18552 3576 18602 3632
rect 18552 3574 18644 3576
rect 18597 3572 18644 3574
rect 18708 3572 18714 3636
rect 20621 3634 20687 3637
rect 24117 3634 24183 3637
rect 20621 3632 24183 3634
rect 20621 3576 20626 3632
rect 20682 3576 24122 3632
rect 24178 3576 24183 3632
rect 20621 3574 24183 3576
rect 18597 3571 18663 3572
rect 20621 3571 20687 3574
rect 24117 3571 24183 3574
rect 33041 3634 33107 3637
rect 33869 3634 33935 3637
rect 33041 3632 33935 3634
rect 33041 3576 33046 3632
rect 33102 3576 33874 3632
rect 33930 3576 33935 3632
rect 33041 3574 33935 3576
rect 33041 3571 33107 3574
rect 33869 3571 33935 3574
rect 31661 3498 31727 3501
rect 34646 3498 34652 3500
rect 31661 3496 34652 3498
rect 31661 3440 31666 3496
rect 31722 3440 34652 3496
rect 31661 3438 34652 3440
rect 31661 3435 31727 3438
rect 34646 3436 34652 3438
rect 34716 3498 34722 3500
rect 35249 3498 35315 3501
rect 34716 3496 35315 3498
rect 34716 3440 35254 3496
rect 35310 3440 35315 3496
rect 34716 3438 35315 3440
rect 34716 3436 34722 3438
rect 35249 3435 35315 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 2221 2954 2287 2957
rect 19190 2954 19196 2956
rect 2221 2952 19196 2954
rect 2221 2896 2226 2952
rect 2282 2896 19196 2952
rect 2221 2894 19196 2896
rect 2221 2891 2287 2894
rect 19190 2892 19196 2894
rect 19260 2892 19266 2956
rect 22829 2954 22895 2957
rect 26325 2954 26391 2957
rect 22829 2952 26391 2954
rect 22829 2896 22834 2952
rect 22890 2896 26330 2952
rect 26386 2896 26391 2952
rect 22829 2894 26391 2896
rect 22829 2891 22895 2894
rect 26325 2891 26391 2894
rect 46565 2818 46631 2821
rect 47480 2818 48280 2848
rect 46565 2816 48280 2818
rect 46565 2760 46570 2816
rect 46626 2760 48280 2816
rect 46565 2758 48280 2760
rect 46565 2755 46631 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 47480 2728 48280 2758
rect 34930 2687 35246 2688
rect 9397 2682 9463 2685
rect 13670 2682 13676 2684
rect 9397 2680 13676 2682
rect 9397 2624 9402 2680
rect 9458 2624 13676 2680
rect 9397 2622 13676 2624
rect 9397 2619 9463 2622
rect 13670 2620 13676 2622
rect 13740 2620 13746 2684
rect 20478 2620 20484 2684
rect 20548 2682 20554 2684
rect 20989 2682 21055 2685
rect 20548 2680 21055 2682
rect 20548 2624 20994 2680
rect 21050 2624 21055 2680
rect 20548 2622 21055 2624
rect 20548 2620 20554 2622
rect 20989 2619 21055 2622
rect 36118 2620 36124 2684
rect 36188 2682 36194 2684
rect 37457 2682 37523 2685
rect 36188 2680 37523 2682
rect 36188 2624 37462 2680
rect 37518 2624 37523 2680
rect 36188 2622 37523 2624
rect 36188 2620 36194 2622
rect 37457 2619 37523 2622
rect 37590 2620 37596 2684
rect 37660 2682 37666 2684
rect 42701 2682 42767 2685
rect 37660 2680 42767 2682
rect 37660 2624 42706 2680
rect 42762 2624 42767 2680
rect 37660 2622 42767 2624
rect 37660 2620 37666 2622
rect 42701 2619 42767 2622
rect 33726 2484 33732 2548
rect 33796 2546 33802 2548
rect 34881 2546 34947 2549
rect 33796 2544 34947 2546
rect 33796 2488 34886 2544
rect 34942 2488 34947 2544
rect 33796 2486 34947 2488
rect 33796 2484 33802 2486
rect 34881 2483 34947 2486
rect 38510 2484 38516 2548
rect 38580 2546 38586 2548
rect 46197 2546 46263 2549
rect 38580 2544 46263 2546
rect 38580 2488 46202 2544
rect 46258 2488 46263 2544
rect 38580 2486 46263 2488
rect 38580 2484 38586 2486
rect 46197 2483 46263 2486
rect 38142 2348 38148 2412
rect 38212 2410 38218 2412
rect 45645 2410 45711 2413
rect 38212 2408 45711 2410
rect 38212 2352 45650 2408
rect 45706 2352 45711 2408
rect 38212 2350 45711 2352
rect 38212 2348 38218 2350
rect 45645 2347 45711 2350
rect 4870 2208 5186 2209
rect 0 2138 800 2168
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 933 2138 999 2141
rect 0 2136 999 2138
rect 0 2080 938 2136
rect 994 2080 999 2136
rect 0 2078 999 2080
rect 0 2048 800 2078
rect 933 2075 999 2078
rect 45461 778 45527 781
rect 47480 778 48280 808
rect 45461 776 48280 778
rect 45461 720 45466 776
rect 45522 720 48280 776
rect 45461 718 48280 720
rect 45461 715 45527 718
rect 47480 688 48280 718
<< via3 >>
rect 4876 47900 4940 47904
rect 4876 47844 4880 47900
rect 4880 47844 4936 47900
rect 4936 47844 4940 47900
rect 4876 47840 4940 47844
rect 4956 47900 5020 47904
rect 4956 47844 4960 47900
rect 4960 47844 5016 47900
rect 5016 47844 5020 47900
rect 4956 47840 5020 47844
rect 5036 47900 5100 47904
rect 5036 47844 5040 47900
rect 5040 47844 5096 47900
rect 5096 47844 5100 47900
rect 5036 47840 5100 47844
rect 5116 47900 5180 47904
rect 5116 47844 5120 47900
rect 5120 47844 5176 47900
rect 5176 47844 5180 47900
rect 5116 47840 5180 47844
rect 35596 47900 35660 47904
rect 35596 47844 35600 47900
rect 35600 47844 35656 47900
rect 35656 47844 35660 47900
rect 35596 47840 35660 47844
rect 35676 47900 35740 47904
rect 35676 47844 35680 47900
rect 35680 47844 35736 47900
rect 35736 47844 35740 47900
rect 35676 47840 35740 47844
rect 35756 47900 35820 47904
rect 35756 47844 35760 47900
rect 35760 47844 35816 47900
rect 35816 47844 35820 47900
rect 35756 47840 35820 47844
rect 35836 47900 35900 47904
rect 35836 47844 35840 47900
rect 35840 47844 35896 47900
rect 35896 47844 35900 47900
rect 35836 47840 35900 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 32260 46956 32324 47020
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 35596 46812 35660 46816
rect 35596 46756 35600 46812
rect 35600 46756 35656 46812
rect 35656 46756 35660 46812
rect 35596 46752 35660 46756
rect 35676 46812 35740 46816
rect 35676 46756 35680 46812
rect 35680 46756 35736 46812
rect 35736 46756 35740 46812
rect 35676 46752 35740 46756
rect 35756 46812 35820 46816
rect 35756 46756 35760 46812
rect 35760 46756 35816 46812
rect 35816 46756 35820 46812
rect 35756 46752 35820 46756
rect 35836 46812 35900 46816
rect 35836 46756 35840 46812
rect 35840 46756 35896 46812
rect 35896 46756 35900 46812
rect 35836 46752 35900 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 33732 45928 33796 45932
rect 33732 45872 33746 45928
rect 33746 45872 33796 45928
rect 33732 45868 33796 45872
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 35596 45724 35660 45728
rect 35596 45668 35600 45724
rect 35600 45668 35656 45724
rect 35656 45668 35660 45724
rect 35596 45664 35660 45668
rect 35676 45724 35740 45728
rect 35676 45668 35680 45724
rect 35680 45668 35736 45724
rect 35736 45668 35740 45724
rect 35676 45664 35740 45668
rect 35756 45724 35820 45728
rect 35756 45668 35760 45724
rect 35760 45668 35816 45724
rect 35816 45668 35820 45724
rect 35756 45664 35820 45668
rect 35836 45724 35900 45728
rect 35836 45668 35840 45724
rect 35840 45668 35896 45724
rect 35896 45668 35900 45724
rect 35836 45664 35900 45668
rect 32444 45520 32508 45524
rect 32444 45464 32458 45520
rect 32458 45464 32508 45520
rect 32444 45460 32508 45464
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 35596 44636 35660 44640
rect 35596 44580 35600 44636
rect 35600 44580 35656 44636
rect 35656 44580 35660 44636
rect 35596 44576 35660 44580
rect 35676 44636 35740 44640
rect 35676 44580 35680 44636
rect 35680 44580 35736 44636
rect 35736 44580 35740 44636
rect 35676 44576 35740 44580
rect 35756 44636 35820 44640
rect 35756 44580 35760 44636
rect 35760 44580 35816 44636
rect 35816 44580 35820 44636
rect 35756 44576 35820 44580
rect 35836 44636 35900 44640
rect 35836 44580 35840 44636
rect 35840 44580 35896 44636
rect 35896 44580 35900 44636
rect 35836 44576 35900 44580
rect 26924 44236 26988 44300
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19196 43692 19260 43756
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 35596 43548 35660 43552
rect 35596 43492 35600 43548
rect 35600 43492 35656 43548
rect 35656 43492 35660 43548
rect 35596 43488 35660 43492
rect 35676 43548 35740 43552
rect 35676 43492 35680 43548
rect 35680 43492 35736 43548
rect 35736 43492 35740 43548
rect 35676 43488 35740 43492
rect 35756 43548 35820 43552
rect 35756 43492 35760 43548
rect 35760 43492 35816 43548
rect 35816 43492 35820 43548
rect 35756 43488 35820 43492
rect 35836 43548 35900 43552
rect 35836 43492 35840 43548
rect 35840 43492 35896 43548
rect 35896 43492 35900 43548
rect 35836 43488 35900 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 27108 42936 27172 42940
rect 27108 42880 27122 42936
rect 27122 42880 27172 42936
rect 27108 42876 27172 42880
rect 37780 42936 37844 42940
rect 37780 42880 37794 42936
rect 37794 42880 37844 42936
rect 37780 42876 37844 42880
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 35596 42460 35660 42464
rect 35596 42404 35600 42460
rect 35600 42404 35656 42460
rect 35656 42404 35660 42460
rect 35596 42400 35660 42404
rect 35676 42460 35740 42464
rect 35676 42404 35680 42460
rect 35680 42404 35736 42460
rect 35736 42404 35740 42460
rect 35676 42400 35740 42404
rect 35756 42460 35820 42464
rect 35756 42404 35760 42460
rect 35760 42404 35816 42460
rect 35816 42404 35820 42460
rect 35756 42400 35820 42404
rect 35836 42460 35900 42464
rect 35836 42404 35840 42460
rect 35840 42404 35896 42460
rect 35896 42404 35900 42460
rect 35836 42400 35900 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 32628 41440 32692 41444
rect 32628 41384 32642 41440
rect 32642 41384 32692 41440
rect 32628 41380 32692 41384
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 35596 41372 35660 41376
rect 35596 41316 35600 41372
rect 35600 41316 35656 41372
rect 35656 41316 35660 41372
rect 35596 41312 35660 41316
rect 35676 41372 35740 41376
rect 35676 41316 35680 41372
rect 35680 41316 35736 41372
rect 35736 41316 35740 41372
rect 35676 41312 35740 41316
rect 35756 41372 35820 41376
rect 35756 41316 35760 41372
rect 35760 41316 35816 41372
rect 35816 41316 35820 41372
rect 35756 41312 35820 41316
rect 35836 41372 35900 41376
rect 35836 41316 35840 41372
rect 35840 41316 35896 41372
rect 35896 41316 35900 41372
rect 35836 41312 35900 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 35596 40284 35660 40288
rect 35596 40228 35600 40284
rect 35600 40228 35656 40284
rect 35656 40228 35660 40284
rect 35596 40224 35660 40228
rect 35676 40284 35740 40288
rect 35676 40228 35680 40284
rect 35680 40228 35736 40284
rect 35736 40228 35740 40284
rect 35676 40224 35740 40228
rect 35756 40284 35820 40288
rect 35756 40228 35760 40284
rect 35760 40228 35816 40284
rect 35816 40228 35820 40284
rect 35756 40224 35820 40228
rect 35836 40284 35900 40288
rect 35836 40228 35840 40284
rect 35840 40228 35896 40284
rect 35896 40228 35900 40284
rect 35836 40224 35900 40228
rect 20484 40020 20548 40084
rect 38884 40020 38948 40084
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 12940 39340 13004 39404
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 35596 39196 35660 39200
rect 35596 39140 35600 39196
rect 35600 39140 35656 39196
rect 35656 39140 35660 39196
rect 35596 39136 35660 39140
rect 35676 39196 35740 39200
rect 35676 39140 35680 39196
rect 35680 39140 35736 39196
rect 35736 39140 35740 39196
rect 35676 39136 35740 39140
rect 35756 39196 35820 39200
rect 35756 39140 35760 39196
rect 35760 39140 35816 39196
rect 35816 39140 35820 39196
rect 35756 39136 35820 39140
rect 35836 39196 35900 39200
rect 35836 39140 35840 39196
rect 35840 39140 35896 39196
rect 35896 39140 35900 39196
rect 35836 39136 35900 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 18828 38252 18892 38316
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 35596 38108 35660 38112
rect 35596 38052 35600 38108
rect 35600 38052 35656 38108
rect 35656 38052 35660 38108
rect 35596 38048 35660 38052
rect 35676 38108 35740 38112
rect 35676 38052 35680 38108
rect 35680 38052 35736 38108
rect 35736 38052 35740 38108
rect 35676 38048 35740 38052
rect 35756 38108 35820 38112
rect 35756 38052 35760 38108
rect 35760 38052 35816 38108
rect 35816 38052 35820 38108
rect 35756 38048 35820 38052
rect 35836 38108 35900 38112
rect 35836 38052 35840 38108
rect 35840 38052 35896 38108
rect 35896 38052 35900 38108
rect 35836 38048 35900 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 36124 37088 36188 37092
rect 36124 37032 36138 37088
rect 36138 37032 36188 37088
rect 36124 37028 36188 37032
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 21404 35124 21468 35188
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 42196 34368 42260 34372
rect 42196 34312 42210 34368
rect 42210 34312 42260 34368
rect 42196 34308 42260 34312
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 15516 32268 15580 32332
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 18644 30908 18708 30972
rect 37780 30908 37844 30972
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 13676 30364 13740 30428
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 37596 29004 37660 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 21036 28188 21100 28252
rect 29868 28324 29932 28388
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 19932 27840 19996 27844
rect 19932 27784 19946 27840
rect 19946 27784 19996 27840
rect 19932 27780 19996 27784
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 29132 27296 29196 27300
rect 29132 27240 29182 27296
rect 29182 27240 29196 27296
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 18828 27160 18892 27164
rect 18828 27104 18842 27160
rect 18842 27104 18892 27160
rect 18828 27100 18892 27104
rect 29132 27236 29196 27240
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 25452 26964 25516 27028
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4660 26616 4724 26620
rect 4660 26560 4710 26616
rect 4710 26560 4724 26616
rect 4660 26556 4724 26560
rect 20300 26480 20364 26484
rect 20300 26424 20350 26480
rect 20350 26424 20364 26480
rect 20300 26420 20364 26424
rect 32444 26148 32508 26212
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 34468 25604 34532 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 21404 25332 21468 25396
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 34652 24848 34716 24852
rect 34652 24792 34666 24848
rect 34666 24792 34716 24848
rect 34652 24788 34716 24792
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 38516 23488 38580 23492
rect 38516 23432 38530 23488
rect 38530 23432 38580 23488
rect 38516 23428 38580 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 32260 23156 32324 23220
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 38884 22612 38948 22676
rect 39068 22400 39132 22404
rect 39068 22344 39118 22400
rect 39118 22344 39132 22400
rect 39068 22340 39132 22344
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 34652 21932 34716 21996
rect 25452 21856 25516 21860
rect 25452 21800 25466 21856
rect 25466 21800 25516 21856
rect 25452 21796 25516 21800
rect 30236 21796 30300 21860
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 19932 21660 19996 21724
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 39436 20632 39500 20636
rect 39436 20576 39486 20632
rect 39486 20576 39500 20632
rect 39436 20572 39500 20576
rect 34468 20436 34532 20500
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4660 20028 4724 20092
rect 39068 19756 39132 19820
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 15516 19212 15580 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 39436 18804 39500 18868
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 30052 18260 30116 18324
rect 12940 18124 13004 18188
rect 15516 17988 15580 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 42196 17716 42260 17780
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 38148 16688 38212 16692
rect 38148 16632 38162 16688
rect 38162 16632 38212 16688
rect 38148 16628 38212 16632
rect 20300 16552 20364 16556
rect 20300 16496 20350 16552
rect 20350 16496 20364 16552
rect 20300 16492 20364 16496
rect 21036 16492 21100 16556
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 29132 16084 29196 16148
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 18828 15132 18892 15196
rect 19748 15132 19812 15196
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19748 14452 19812 14516
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 29500 13772 29564 13836
rect 30236 13772 30300 13836
rect 34100 13772 34164 13836
rect 19932 13636 19996 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 29868 12336 29932 12340
rect 29868 12280 29918 12336
rect 29918 12280 29932 12336
rect 29868 12276 29932 12280
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 30052 10916 30116 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 26924 10508 26988 10572
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 34652 9556 34716 9620
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 19748 8392 19812 8396
rect 19748 8336 19762 8392
rect 19762 8336 19812 8392
rect 19748 8332 19812 8336
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 29500 7924 29564 7988
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 34100 7380 34164 7444
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 32628 6156 32692 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 27108 3980 27172 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 18644 3632 18708 3636
rect 18644 3576 18658 3632
rect 18658 3576 18708 3632
rect 18644 3572 18708 3576
rect 34652 3436 34716 3500
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 19196 2892 19260 2956
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 13676 2620 13740 2684
rect 20484 2620 20548 2684
rect 36124 2620 36188 2684
rect 37596 2620 37660 2684
rect 33732 2484 33796 2548
rect 38516 2484 38580 2548
rect 38148 2348 38212 2412
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 47360 4528 47920
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4868 47904 5188 47920
rect 4868 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5188 47904
rect 4868 46816 5188 47840
rect 34928 47360 35248 47920
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 32259 47020 32325 47021
rect 32259 46956 32260 47020
rect 32324 46956 32325 47020
rect 32259 46955 32325 46956
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 26923 44300 26989 44301
rect 26923 44236 26924 44300
rect 26988 44236 26989 44300
rect 26923 44235 26989 44236
rect 19195 43756 19261 43757
rect 19195 43692 19196 43756
rect 19260 43692 19261 43756
rect 19195 43691 19261 43692
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 12939 39404 13005 39405
rect 12939 39340 12940 39404
rect 13004 39340 13005 39404
rect 12939 39339 13005 39340
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4659 26620 4725 26621
rect 4659 26556 4660 26620
rect 4724 26556 4725 26620
rect 4659 26555 4725 26556
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4662 20093 4722 26555
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4659 20092 4725 20093
rect 4659 20028 4660 20092
rect 4724 20028 4725 20092
rect 4659 20027 4725 20028
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 12942 18189 13002 39339
rect 18827 38316 18893 38317
rect 18827 38252 18828 38316
rect 18892 38252 18893 38316
rect 18827 38251 18893 38252
rect 15515 32332 15581 32333
rect 15515 32268 15516 32332
rect 15580 32268 15581 32332
rect 15515 32267 15581 32268
rect 13675 30428 13741 30429
rect 13675 30364 13676 30428
rect 13740 30364 13741 30428
rect 13675 30363 13741 30364
rect 12939 18188 13005 18189
rect 12939 18124 12940 18188
rect 13004 18124 13005 18188
rect 12939 18123 13005 18124
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 13678 2685 13738 30363
rect 15518 19277 15578 32267
rect 18643 30972 18709 30973
rect 18643 30908 18644 30972
rect 18708 30908 18709 30972
rect 18643 30907 18709 30908
rect 15515 19276 15581 19277
rect 15515 19212 15516 19276
rect 15580 19212 15581 19276
rect 15515 19211 15581 19212
rect 15518 18053 15578 19211
rect 15515 18052 15581 18053
rect 15515 17988 15516 18052
rect 15580 17988 15581 18052
rect 15515 17987 15581 17988
rect 18646 3637 18706 30907
rect 18830 27165 18890 38251
rect 18827 27164 18893 27165
rect 18827 27100 18828 27164
rect 18892 27100 18893 27164
rect 18827 27099 18893 27100
rect 18830 15197 18890 27099
rect 18827 15196 18893 15197
rect 18827 15132 18828 15196
rect 18892 15132 18893 15196
rect 18827 15131 18893 15132
rect 18643 3636 18709 3637
rect 18643 3572 18644 3636
rect 18708 3572 18709 3636
rect 18643 3571 18709 3572
rect 19198 2957 19258 43691
rect 20483 40084 20549 40085
rect 20483 40020 20484 40084
rect 20548 40020 20549 40084
rect 20483 40019 20549 40020
rect 19931 27844 19997 27845
rect 19931 27780 19932 27844
rect 19996 27780 19997 27844
rect 19931 27779 19997 27780
rect 19934 21725 19994 27779
rect 20299 26484 20365 26485
rect 20299 26420 20300 26484
rect 20364 26420 20365 26484
rect 20299 26419 20365 26420
rect 19931 21724 19997 21725
rect 19931 21660 19932 21724
rect 19996 21660 19997 21724
rect 19931 21659 19997 21660
rect 19747 15196 19813 15197
rect 19747 15132 19748 15196
rect 19812 15132 19813 15196
rect 19747 15131 19813 15132
rect 19750 14517 19810 15131
rect 19747 14516 19813 14517
rect 19747 14452 19748 14516
rect 19812 14452 19813 14516
rect 19747 14451 19813 14452
rect 19750 8397 19810 14451
rect 19934 13701 19994 21659
rect 20302 16557 20362 26419
rect 20299 16556 20365 16557
rect 20299 16492 20300 16556
rect 20364 16492 20365 16556
rect 20299 16491 20365 16492
rect 19931 13700 19997 13701
rect 19931 13636 19932 13700
rect 19996 13636 19997 13700
rect 19931 13635 19997 13636
rect 19747 8396 19813 8397
rect 19747 8332 19748 8396
rect 19812 8332 19813 8396
rect 19747 8331 19813 8332
rect 19195 2956 19261 2957
rect 19195 2892 19196 2956
rect 19260 2892 19261 2956
rect 19195 2891 19261 2892
rect 20486 2685 20546 40019
rect 21403 35188 21469 35189
rect 21403 35124 21404 35188
rect 21468 35124 21469 35188
rect 21403 35123 21469 35124
rect 21035 28252 21101 28253
rect 21035 28188 21036 28252
rect 21100 28188 21101 28252
rect 21035 28187 21101 28188
rect 21038 16557 21098 28187
rect 21406 25397 21466 35123
rect 25451 27028 25517 27029
rect 25451 26964 25452 27028
rect 25516 26964 25517 27028
rect 25451 26963 25517 26964
rect 21403 25396 21469 25397
rect 21403 25332 21404 25396
rect 21468 25332 21469 25396
rect 21403 25331 21469 25332
rect 25454 21861 25514 26963
rect 25451 21860 25517 21861
rect 25451 21796 25452 21860
rect 25516 21796 25517 21860
rect 25451 21795 25517 21796
rect 21035 16556 21101 16557
rect 21035 16492 21036 16556
rect 21100 16492 21101 16556
rect 21035 16491 21101 16492
rect 26926 10573 26986 44235
rect 27107 42940 27173 42941
rect 27107 42876 27108 42940
rect 27172 42876 27173 42940
rect 27107 42875 27173 42876
rect 26923 10572 26989 10573
rect 26923 10508 26924 10572
rect 26988 10508 26989 10572
rect 26923 10507 26989 10508
rect 27110 4045 27170 42875
rect 29867 28388 29933 28389
rect 29867 28324 29868 28388
rect 29932 28324 29933 28388
rect 29867 28323 29933 28324
rect 29131 27300 29197 27301
rect 29131 27236 29132 27300
rect 29196 27236 29197 27300
rect 29131 27235 29197 27236
rect 29134 16149 29194 27235
rect 29131 16148 29197 16149
rect 29131 16084 29132 16148
rect 29196 16084 29197 16148
rect 29131 16083 29197 16084
rect 29499 13836 29565 13837
rect 29499 13772 29500 13836
rect 29564 13772 29565 13836
rect 29499 13771 29565 13772
rect 29502 7989 29562 13771
rect 29870 12341 29930 28323
rect 32262 23221 32322 46955
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 33731 45932 33797 45933
rect 33731 45868 33732 45932
rect 33796 45868 33797 45932
rect 33731 45867 33797 45868
rect 32443 45524 32509 45525
rect 32443 45460 32444 45524
rect 32508 45460 32509 45524
rect 32443 45459 32509 45460
rect 32446 26213 32506 45459
rect 32627 41444 32693 41445
rect 32627 41380 32628 41444
rect 32692 41380 32693 41444
rect 32627 41379 32693 41380
rect 32443 26212 32509 26213
rect 32443 26148 32444 26212
rect 32508 26148 32509 26212
rect 32443 26147 32509 26148
rect 32259 23220 32325 23221
rect 32259 23156 32260 23220
rect 32324 23156 32325 23220
rect 32259 23155 32325 23156
rect 30235 21860 30301 21861
rect 30235 21796 30236 21860
rect 30300 21796 30301 21860
rect 30235 21795 30301 21796
rect 30051 18324 30117 18325
rect 30051 18260 30052 18324
rect 30116 18260 30117 18324
rect 30051 18259 30117 18260
rect 29867 12340 29933 12341
rect 29867 12276 29868 12340
rect 29932 12276 29933 12340
rect 29867 12275 29933 12276
rect 30054 10981 30114 18259
rect 30238 13837 30298 21795
rect 30235 13836 30301 13837
rect 30235 13772 30236 13836
rect 30300 13772 30301 13836
rect 30235 13771 30301 13772
rect 30051 10980 30117 10981
rect 30051 10916 30052 10980
rect 30116 10916 30117 10980
rect 30051 10915 30117 10916
rect 29499 7988 29565 7989
rect 29499 7924 29500 7988
rect 29564 7924 29565 7988
rect 29499 7923 29565 7924
rect 32630 6221 32690 41379
rect 32627 6220 32693 6221
rect 32627 6156 32628 6220
rect 32692 6156 32693 6220
rect 32627 6155 32693 6156
rect 27107 4044 27173 4045
rect 27107 3980 27108 4044
rect 27172 3980 27173 4044
rect 27107 3979 27173 3980
rect 13675 2684 13741 2685
rect 13675 2620 13676 2684
rect 13740 2620 13741 2684
rect 13675 2619 13741 2620
rect 20483 2684 20549 2685
rect 20483 2620 20484 2684
rect 20548 2620 20549 2684
rect 20483 2619 20549 2620
rect 33734 2549 33794 45867
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36260 35248 36416
rect 34928 36024 34970 36260
rect 35206 36024 35248 36260
rect 34928 35392 35248 36024
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34467 25668 34533 25669
rect 34467 25604 34468 25668
rect 34532 25604 34533 25668
rect 34467 25603 34533 25604
rect 34470 20501 34530 25603
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34651 24852 34717 24853
rect 34651 24788 34652 24852
rect 34716 24788 34717 24852
rect 34651 24787 34717 24788
rect 34654 21997 34714 24787
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34651 21996 34717 21997
rect 34651 21932 34652 21996
rect 34716 21932 34717 21996
rect 34651 21931 34717 21932
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34467 20500 34533 20501
rect 34467 20436 34468 20500
rect 34532 20436 34533 20500
rect 34467 20435 34533 20436
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34099 13836 34165 13837
rect 34099 13772 34100 13836
rect 34164 13772 34165 13836
rect 34099 13771 34165 13772
rect 34102 7445 34162 13771
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34651 9620 34717 9621
rect 34651 9556 34652 9620
rect 34716 9556 34717 9620
rect 34651 9555 34717 9556
rect 34099 7444 34165 7445
rect 34099 7380 34100 7444
rect 34164 7380 34165 7444
rect 34099 7379 34165 7380
rect 34654 3501 34714 9555
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34651 3500 34717 3501
rect 34651 3436 34652 3500
rect 34716 3436 34717 3500
rect 34651 3435 34717 3436
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 33731 2548 33797 2549
rect 33731 2484 33732 2548
rect 33796 2484 33797 2548
rect 33731 2483 33797 2484
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 2128 35248 2688
rect 35588 47904 35908 47920
rect 35588 47840 35596 47904
rect 35660 47840 35676 47904
rect 35740 47840 35756 47904
rect 35820 47840 35836 47904
rect 35900 47840 35908 47904
rect 35588 46816 35908 47840
rect 35588 46752 35596 46816
rect 35660 46752 35676 46816
rect 35740 46752 35756 46816
rect 35820 46752 35836 46816
rect 35900 46752 35908 46816
rect 35588 45728 35908 46752
rect 35588 45664 35596 45728
rect 35660 45664 35676 45728
rect 35740 45664 35756 45728
rect 35820 45664 35836 45728
rect 35900 45664 35908 45728
rect 35588 44640 35908 45664
rect 35588 44576 35596 44640
rect 35660 44576 35676 44640
rect 35740 44576 35756 44640
rect 35820 44576 35836 44640
rect 35900 44576 35908 44640
rect 35588 43552 35908 44576
rect 35588 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35908 43552
rect 35588 42464 35908 43488
rect 37779 42940 37845 42941
rect 37779 42876 37780 42940
rect 37844 42876 37845 42940
rect 37779 42875 37845 42876
rect 35588 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35908 42464
rect 35588 41376 35908 42400
rect 35588 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35908 41376
rect 35588 40288 35908 41312
rect 35588 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35908 40288
rect 35588 39200 35908 40224
rect 35588 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35908 39200
rect 35588 38112 35908 39136
rect 35588 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35908 38112
rect 35588 37024 35908 38048
rect 36123 37092 36189 37093
rect 36123 37028 36124 37092
rect 36188 37028 36189 37092
rect 36123 37027 36189 37028
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 36920 35908 36960
rect 35588 36684 35630 36920
rect 35866 36684 35908 36920
rect 35588 35936 35908 36684
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 36126 2685 36186 37027
rect 37782 30973 37842 42875
rect 38883 40084 38949 40085
rect 38883 40020 38884 40084
rect 38948 40020 38949 40084
rect 38883 40019 38949 40020
rect 37779 30972 37845 30973
rect 37779 30908 37780 30972
rect 37844 30908 37845 30972
rect 37779 30907 37845 30908
rect 37595 29068 37661 29069
rect 37595 29004 37596 29068
rect 37660 29004 37661 29068
rect 37595 29003 37661 29004
rect 37598 2685 37658 29003
rect 38515 23492 38581 23493
rect 38515 23428 38516 23492
rect 38580 23428 38581 23492
rect 38515 23427 38581 23428
rect 38147 16692 38213 16693
rect 38147 16628 38148 16692
rect 38212 16628 38213 16692
rect 38147 16627 38213 16628
rect 36123 2684 36189 2685
rect 36123 2620 36124 2684
rect 36188 2620 36189 2684
rect 36123 2619 36189 2620
rect 37595 2684 37661 2685
rect 37595 2620 37596 2684
rect 37660 2620 37661 2684
rect 37595 2619 37661 2620
rect 38150 2413 38210 16627
rect 38518 2549 38578 23427
rect 38886 22677 38946 40019
rect 42195 34372 42261 34373
rect 42195 34308 42196 34372
rect 42260 34308 42261 34372
rect 42195 34307 42261 34308
rect 38883 22676 38949 22677
rect 38883 22612 38884 22676
rect 38948 22612 38949 22676
rect 38883 22611 38949 22612
rect 39067 22404 39133 22405
rect 39067 22340 39068 22404
rect 39132 22340 39133 22404
rect 39067 22339 39133 22340
rect 39070 19821 39130 22339
rect 39435 20636 39501 20637
rect 39435 20572 39436 20636
rect 39500 20572 39501 20636
rect 39435 20571 39501 20572
rect 39067 19820 39133 19821
rect 39067 19756 39068 19820
rect 39132 19756 39133 19820
rect 39067 19755 39133 19756
rect 39438 18869 39498 20571
rect 39435 18868 39501 18869
rect 39435 18804 39436 18868
rect 39500 18804 39501 18868
rect 39435 18803 39501 18804
rect 42198 17781 42258 34307
rect 42195 17780 42261 17781
rect 42195 17716 42196 17780
rect 42260 17716 42261 17780
rect 42195 17715 42261 17716
rect 38515 2548 38581 2549
rect 38515 2484 38516 2548
rect 38580 2484 38581 2548
rect 38515 2483 38581 2484
rect 38147 2412 38213 2413
rect 38147 2348 38148 2412
rect 38212 2348 38213 2412
rect 38147 2347 38213 2348
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
<< via4 >>
rect 4250 36024 4486 36260
rect 4910 36684 5146 36920
rect 4250 5388 4486 5624
rect 4910 6048 5146 6284
rect 34970 36024 35206 36260
rect 34970 5388 35206 5624
rect 35630 36684 35866 36920
rect 35630 6048 35866 6284
<< metal5 >>
rect 1056 36920 47152 36962
rect 1056 36684 4910 36920
rect 5146 36684 35630 36920
rect 35866 36684 47152 36920
rect 1056 36642 47152 36684
rect 1056 36260 47152 36302
rect 1056 36024 4250 36260
rect 4486 36024 34970 36260
rect 35206 36024 47152 36260
rect 1056 35982 47152 36024
rect 1056 6284 47152 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 47152 6284
rect 1056 6006 47152 6048
rect 1056 5624 47152 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 47152 5624
rect 1056 5346 47152 5388
use sky130_fd_sc_hd__clkbuf_2  _1484_
timestamp 0
transform 1 0 39284 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1485_
timestamp 0
transform 1 0 39284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1486_
timestamp 0
transform 1 0 38548 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1487_
timestamp 0
transform 1 0 39560 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1488_
timestamp 0
transform 1 0 38824 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1489_
timestamp 0
transform 1 0 39560 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1490_
timestamp 0
transform 1 0 38548 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _1491_
timestamp 0
transform 1 0 38180 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 0
transform 1 0 39836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1493_
timestamp 0
transform 1 0 38732 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1494_
timestamp 0
transform 1 0 39468 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1495_
timestamp 0
transform 1 0 37352 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 0
transform 1 0 38088 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1497_
timestamp 0
transform 1 0 38272 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 0
transform 1 0 39008 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1499_
timestamp 0
transform 1 0 38456 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 0
transform 1 0 39100 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1501_
timestamp 0
transform 1 0 40020 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1502_
timestamp 0
transform 1 0 45448 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1503_
timestamp 0
transform 1 0 42504 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1504_
timestamp 0
transform 1 0 45264 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _1505_
timestamp 0
transform 1 0 45724 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1506_
timestamp 0
transform 1 0 46184 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1507_
timestamp 0
transform 1 0 45724 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1508_
timestamp 0
transform 1 0 45356 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1509_
timestamp 0
transform 1 0 46276 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1510_
timestamp 0
transform 1 0 46368 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1511_
timestamp 0
transform 1 0 46276 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1512_
timestamp 0
transform 1 0 45908 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1513_
timestamp 0
transform 1 0 45724 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1514_
timestamp 0
transform 1 0 46000 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1515_
timestamp 0
transform 1 0 45724 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1516_
timestamp 0
transform 1 0 45908 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1517_
timestamp 0
transform 1 0 45172 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1518_
timestamp 0
transform 1 0 46184 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1519_
timestamp 0
transform 1 0 44988 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1520_
timestamp 0
transform 1 0 45264 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1521_
timestamp 0
transform 1 0 43516 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1522_
timestamp 0
transform 1 0 43976 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1523_
timestamp 0
transform 1 0 41676 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1524_
timestamp 0
transform 1 0 41124 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1525_
timestamp 0
transform 1 0 41124 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1526_
timestamp 0
transform 1 0 40112 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1527_
timestamp 0
transform 1 0 37996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1528_
timestamp 0
transform 1 0 43700 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1529_
timestamp 0
transform 1 0 44988 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1530_
timestamp 0
transform 1 0 44988 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1531_
timestamp 0
transform 1 0 45448 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1532_
timestamp 0
transform 1 0 38364 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1533_
timestamp 0
transform 1 0 38548 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1534_
timestamp 0
transform 1 0 36064 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1535_
timestamp 0
transform 1 0 38824 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _1536_
timestamp 0
transform 1 0 38732 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_1  _1537_
timestamp 0
transform 1 0 37996 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1538_
timestamp 0
transform 1 0 38640 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1539_
timestamp 0
transform 1 0 38456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1540_
timestamp 0
transform 1 0 37352 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1541_
timestamp 0
transform 1 0 37168 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_4  _1542_
timestamp 0
transform 1 0 37628 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1543_
timestamp 0
transform 1 0 35696 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1544_
timestamp 0
transform 1 0 35512 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1545_
timestamp 0
transform 1 0 36156 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1546_
timestamp 0
transform 1 0 35880 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1547_
timestamp 0
transform 1 0 38916 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1548_
timestamp 0
transform 1 0 38180 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1549_
timestamp 0
transform 1 0 37444 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1550_
timestamp 0
transform 1 0 37260 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1551_
timestamp 0
transform 1 0 35052 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1552_
timestamp 0
transform 1 0 39836 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a311oi_4  _1553_
timestamp 0
transform 1 0 38640 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _1554_
timestamp 0
transform 1 0 37536 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1555_
timestamp 0
transform 1 0 37444 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1556_
timestamp 0
transform 1 0 36800 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1557_
timestamp 0
transform 1 0 36524 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1558_
timestamp 0
transform 1 0 37260 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1559_
timestamp 0
transform 1 0 34776 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_4  _1560_
timestamp 0
transform 1 0 35420 0 -1 39168
box -38 -48 1602 592
use sky130_fd_sc_hd__nor3b_2  _1561_
timestamp 0
transform 1 0 37260 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1562_
timestamp 0
transform 1 0 37812 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1563_
timestamp 0
transform 1 0 36892 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _1564_
timestamp 0
transform 1 0 33396 0 1 38080
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _1565_
timestamp 0
transform 1 0 7544 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1566_
timestamp 0
transform 1 0 7728 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1567_
timestamp 0
transform 1 0 8372 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1568_
timestamp 0
transform 1 0 7268 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1569_
timestamp 0
transform 1 0 7728 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1570_
timestamp 0
transform 1 0 6624 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1571_
timestamp 0
transform 1 0 7176 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1572_
timestamp 0
transform 1 0 6808 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1573_
timestamp 0
transform 1 0 7452 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1574_
timestamp 0
transform 1 0 20056 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1575_
timestamp 0
transform 1 0 19964 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _1576_
timestamp 0
transform 1 0 18308 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1577_
timestamp 0
transform 1 0 20056 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _1578_
timestamp 0
transform 1 0 18952 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1579_
timestamp 0
transform 1 0 21804 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1580_
timestamp 0
transform 1 0 23276 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1581_
timestamp 0
transform 1 0 20976 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1582_
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1583_
timestamp 0
transform 1 0 20608 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1584_
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1585_
timestamp 0
transform 1 0 8924 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1586_
timestamp 0
transform 1 0 21804 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1587_
timestamp 0
transform 1 0 20792 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1588_
timestamp 0
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1589_
timestamp 0
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1590_
timestamp 0
transform 1 0 19688 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1591_
timestamp 0
transform 1 0 22448 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1592_
timestamp 0
transform 1 0 20056 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1593_
timestamp 0
transform 1 0 20056 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1594_
timestamp 0
transform 1 0 24380 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1595_
timestamp 0
transform 1 0 26128 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1596_
timestamp 0
transform 1 0 25944 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1597_
timestamp 0
transform 1 0 25852 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1598_
timestamp 0
transform 1 0 32108 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _1599_
timestamp 0
transform 1 0 23000 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1600_
timestamp 0
transform 1 0 24104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1601_
timestamp 0
transform 1 0 27508 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1602_
timestamp 0
transform 1 0 26956 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1603_
timestamp 0
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1604_
timestamp 0
transform 1 0 18032 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1605_
timestamp 0
transform 1 0 13892 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _1606_
timestamp 0
transform 1 0 21988 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1607_
timestamp 0
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1608_
timestamp 0
transform 1 0 21620 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1609_
timestamp 0
transform 1 0 19412 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1610_
timestamp 0
transform 1 0 19504 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1611_
timestamp 0
transform 1 0 19228 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1612_
timestamp 0
transform 1 0 20608 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1613_
timestamp 0
transform 1 0 4048 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1614_
timestamp 0
transform 1 0 21160 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1615_
timestamp 0
transform 1 0 20792 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1616_
timestamp 0
transform 1 0 19412 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1617_
timestamp 0
transform 1 0 19504 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1618_
timestamp 0
transform 1 0 17204 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1619_
timestamp 0
transform 1 0 20240 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1620_
timestamp 0
transform 1 0 20424 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1621_
timestamp 0
transform 1 0 17204 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1622_
timestamp 0
transform 1 0 19228 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1623_
timestamp 0
transform 1 0 11500 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1624_
timestamp 0
transform 1 0 20240 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1625_
timestamp 0
transform 1 0 18860 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1626_
timestamp 0
transform 1 0 18584 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1627_
timestamp 0
transform 1 0 15548 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_4  _1628_
timestamp 0
transform 1 0 21252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1629_
timestamp 0
transform 1 0 20700 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1630_
timestamp 0
transform 1 0 10028 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _1631_
timestamp 0
transform 1 0 19412 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1632_
timestamp 0
transform 1 0 17480 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1633_
timestamp 0
transform 1 0 19136 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1634_
timestamp 0
transform 1 0 9200 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _1635_
timestamp 0
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1636_
timestamp 0
transform 1 0 21160 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1637_
timestamp 0
transform 1 0 23460 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1638_
timestamp 0
transform 1 0 25208 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1639_
timestamp 0
transform 1 0 23552 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1640_
timestamp 0
transform 1 0 26956 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_4  _1641_
timestamp 0
transform 1 0 21160 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1642_
timestamp 0
transform 1 0 21160 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1643_
timestamp 0
transform 1 0 32108 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_4  _1644_
timestamp 0
transform 1 0 21804 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1645_
timestamp 0
transform 1 0 27232 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1646_
timestamp 0
transform 1 0 25576 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1647_
timestamp 0
transform 1 0 24104 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1648_
timestamp 0
transform 1 0 26864 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1649_
timestamp 0
transform 1 0 4232 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1650_
timestamp 0
transform 1 0 19780 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1651_
timestamp 0
transform 1 0 27600 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1652_
timestamp 0
transform 1 0 28428 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1653_
timestamp 0
transform 1 0 29900 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1654_
timestamp 0
transform 1 0 29348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1655_
timestamp 0
transform 1 0 28796 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1656_
timestamp 0
transform 1 0 4048 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1657_
timestamp 0
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1658_
timestamp 0
transform 1 0 23184 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1659_
timestamp 0
transform 1 0 25116 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1660_
timestamp 0
transform 1 0 29532 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1661_
timestamp 0
transform 1 0 32660 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1662_
timestamp 0
transform 1 0 30176 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1663_
timestamp 0
transform 1 0 25208 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1664_
timestamp 0
transform 1 0 17020 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1665_
timestamp 0
transform 1 0 18952 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1666_
timestamp 0
transform 1 0 4508 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1667_
timestamp 0
transform 1 0 19964 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1668_
timestamp 0
transform 1 0 29256 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1669_
timestamp 0
transform 1 0 30452 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1670_
timestamp 0
transform 1 0 33488 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1671_
timestamp 0
transform 1 0 30452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1672_
timestamp 0
transform 1 0 29532 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1673_
timestamp 0
transform 1 0 19504 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1674_
timestamp 0
transform 1 0 21252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1675_
timestamp 0
transform 1 0 4324 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1676_
timestamp 0
transform 1 0 20884 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1677_
timestamp 0
transform 1 0 27876 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1678_
timestamp 0
transform 1 0 29072 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1679_
timestamp 0
transform 1 0 33396 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1680_
timestamp 0
transform 1 0 29992 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1681_
timestamp 0
transform 1 0 29532 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1682_
timestamp 0
transform 1 0 14812 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1683_
timestamp 0
transform 1 0 25484 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1684_
timestamp 0
transform 1 0 10488 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1685_
timestamp 0
transform 1 0 23000 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1686_
timestamp 0
transform 1 0 20700 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _1687_
timestamp 0
transform 1 0 37628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1688_
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1689_
timestamp 0
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1690_
timestamp 0
transform 1 0 18308 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1691_
timestamp 0
transform 1 0 24104 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1692_
timestamp 0
transform 1 0 29716 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1693_
timestamp 0
transform 1 0 33396 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1694_
timestamp 0
transform 1 0 30636 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1695_
timestamp 0
transform 1 0 24656 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1696_
timestamp 0
transform 1 0 9476 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1697_
timestamp 0
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1698_
timestamp 0
transform 1 0 19688 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1699_
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1700_
timestamp 0
transform 1 0 25300 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1701_
timestamp 0
transform 1 0 33488 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1702_
timestamp 0
transform 1 0 26956 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1703_
timestamp 0
transform 1 0 22172 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1704_
timestamp 0
transform 1 0 22356 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1705_
timestamp 0
transform 1 0 23460 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1706_
timestamp 0
transform 1 0 25944 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1707_
timestamp 0
transform 1 0 22632 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1708_
timestamp 0
transform 1 0 4140 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1709_
timestamp 0
transform 1 0 20056 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1710_
timestamp 0
transform 1 0 19688 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1711_
timestamp 0
transform 1 0 21620 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1712_
timestamp 0
transform 1 0 22172 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1713_
timestamp 0
transform 1 0 16928 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1714_
timestamp 0
transform 1 0 25852 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1715_
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1716_
timestamp 0
transform 1 0 20700 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1717_
timestamp 0
transform 1 0 28612 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1718_
timestamp 0
transform 1 0 29532 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1719_
timestamp 0
transform 1 0 32108 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1720_
timestamp 0
transform 1 0 29992 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1721_
timestamp 0
transform 1 0 29164 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1722_
timestamp 0
transform 1 0 7912 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1723_
timestamp 0
transform 1 0 21988 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1724_
timestamp 0
transform 1 0 19044 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1725_
timestamp 0
transform 1 0 21160 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1726_
timestamp 0
transform 1 0 29532 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1727_
timestamp 0
transform 1 0 32660 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1728_
timestamp 0
transform 1 0 30360 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1729_
timestamp 0
transform 1 0 22356 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1730_
timestamp 0
transform 1 0 11224 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1731_
timestamp 0
transform 1 0 21436 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1732_
timestamp 0
transform 1 0 17204 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1733_
timestamp 0
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1734_
timestamp 0
transform 1 0 14444 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1735_
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1736_
timestamp 0
transform 1 0 21988 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1737_
timestamp 0
transform 1 0 21712 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1738_
timestamp 0
transform 1 0 17848 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1739_
timestamp 0
transform 1 0 24840 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1740_
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1741_
timestamp 0
transform 1 0 20700 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1742_
timestamp 0
transform 1 0 24012 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1743_
timestamp 0
transform 1 0 26036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1744_
timestamp 0
transform 1 0 25576 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1745_
timestamp 0
transform 1 0 26588 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1746_
timestamp 0
transform 1 0 25392 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1747_
timestamp 0
transform 1 0 11592 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1748_
timestamp 0
transform 1 0 11040 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1749_
timestamp 0
transform 1 0 10304 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1750_
timestamp 0
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1751_
timestamp 0
transform 1 0 8556 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _1752_
timestamp 0
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1753_
timestamp 0
transform 1 0 13432 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1754_
timestamp 0
transform 1 0 12144 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1755_
timestamp 0
transform 1 0 11684 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1756_
timestamp 0
transform 1 0 14904 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1757_
timestamp 0
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1758_
timestamp 0
transform 1 0 17664 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1759_
timestamp 0
transform 1 0 16376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1760_
timestamp 0
transform 1 0 21160 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1761_
timestamp 0
transform 1 0 22724 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1762_
timestamp 0
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1763_
timestamp 0
transform 1 0 21896 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1764_
timestamp 0
transform 1 0 15916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1765_
timestamp 0
transform 1 0 23736 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1766_
timestamp 0
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1767_
timestamp 0
transform 1 0 20976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1768_
timestamp 0
transform 1 0 24380 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_4  _1769_
timestamp 0
transform 1 0 15824 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1770_
timestamp 0
transform 1 0 15824 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1771_
timestamp 0
transform 1 0 31740 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _1772_
timestamp 0
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1773_
timestamp 0
transform 1 0 25208 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1774_
timestamp 0
transform 1 0 23000 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1775_
timestamp 0
transform 1 0 4048 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _1776_
timestamp 0
transform 1 0 13156 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1777_
timestamp 0
transform 1 0 11776 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1778_
timestamp 0
transform 1 0 17388 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1779_
timestamp 0
transform 1 0 19320 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1780_
timestamp 0
transform 1 0 18952 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1781_
timestamp 0
transform 1 0 14168 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1782_
timestamp 0
transform 1 0 20700 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1783_
timestamp 0
transform 1 0 20884 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1784_
timestamp 0
transform 1 0 11224 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1785_
timestamp 0
transform 1 0 13064 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1786_
timestamp 0
transform 1 0 16928 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1787_
timestamp 0
transform 1 0 18308 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1788_
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1789_
timestamp 0
transform 1 0 11408 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1790_
timestamp 0
transform 1 0 9476 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _1791_
timestamp 0
transform 1 0 13340 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1792_
timestamp 0
transform 1 0 13156 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _1793_
timestamp 0
transform 1 0 11960 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1794_
timestamp 0
transform 1 0 12420 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1795_
timestamp 0
transform 1 0 14628 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1796_
timestamp 0
transform 1 0 13708 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1797_
timestamp 0
transform 1 0 14076 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1798_
timestamp 0
transform 1 0 23552 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1799_
timestamp 0
transform 1 0 25668 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1800_
timestamp 0
transform 1 0 9476 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1801_
timestamp 0
transform 1 0 11868 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1802_
timestamp 0
transform 1 0 14444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1803_
timestamp 0
transform 1 0 26588 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1804_
timestamp 0
transform 1 0 28520 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1805_
timestamp 0
transform 1 0 32108 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _1806_
timestamp 0
transform 1 0 19044 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1807_
timestamp 0
transform 1 0 28152 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1808_
timestamp 0
transform 1 0 27508 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1809_
timestamp 0
transform 1 0 24380 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1810_
timestamp 0
transform 1 0 26312 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1811_
timestamp 0
transform 1 0 4232 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1812_
timestamp 0
transform 1 0 11960 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1813_
timestamp 0
transform 1 0 27324 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1814_
timestamp 0
transform 1 0 28060 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1815_
timestamp 0
transform 1 0 29900 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1816_
timestamp 0
transform 1 0 28612 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1817_
timestamp 0
transform 1 0 27416 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1818_
timestamp 0
transform 1 0 10212 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1819_
timestamp 0
transform 1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1820_
timestamp 0
transform 1 0 3956 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _1821_
timestamp 0
transform 1 0 12144 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1822_
timestamp 0
transform 1 0 12052 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1823_
timestamp 0
transform 1 0 22908 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1824_
timestamp 0
transform 1 0 23368 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1825_
timestamp 0
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1826_
timestamp 0
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1827_
timestamp 0
transform 1 0 28888 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1828_
timestamp 0
transform 1 0 33028 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_4  _1829_
timestamp 0
transform 1 0 24656 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1830_
timestamp 0
transform 1 0 30176 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1831_
timestamp 0
transform 1 0 23092 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1832_
timestamp 0
transform 1 0 4324 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1833_
timestamp 0
transform 1 0 12144 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1834_
timestamp 0
transform 1 0 17112 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1835_
timestamp 0
transform 1 0 19228 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1836_
timestamp 0
transform 1 0 29808 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1837_
timestamp 0
transform 1 0 33488 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1838_
timestamp 0
transform 1 0 31004 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1839_
timestamp 0
transform 1 0 20332 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1840_
timestamp 0
transform 1 0 19504 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1841_
timestamp 0
transform 1 0 21620 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1842_
timestamp 0
transform 1 0 4508 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1843_
timestamp 0
transform 1 0 11776 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1844_
timestamp 0
transform 1 0 27416 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1845_
timestamp 0
transform 1 0 23184 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1846_
timestamp 0
transform 1 0 33396 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1847_
timestamp 0
transform 1 0 22816 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1848_
timestamp 0
transform 1 0 22172 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1849_
timestamp 0
transform 1 0 25576 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1850_
timestamp 0
transform 1 0 23092 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1851_
timestamp 0
transform 1 0 24380 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1852_
timestamp 0
transform 1 0 14536 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1853_
timestamp 0
transform 1 0 10304 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1854_
timestamp 0
transform 1 0 15364 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1855_
timestamp 0
transform 1 0 20148 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1856_
timestamp 0
transform 1 0 19872 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1857_
timestamp 0
transform 1 0 8740 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1858_
timestamp 0
transform 1 0 12696 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1859_
timestamp 0
transform 1 0 19964 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1860_
timestamp 0
transform 1 0 17204 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1861_
timestamp 0
transform 1 0 17204 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1862_
timestamp 0
transform 1 0 18032 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1863_
timestamp 0
transform 1 0 19780 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1864_
timestamp 0
transform 1 0 29900 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_4  _1865_
timestamp 0
transform 1 0 23184 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1866_
timestamp 0
transform 1 0 23368 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1867_
timestamp 0
transform 1 0 33212 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1868_
timestamp 0
transform 1 0 31464 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1869_
timestamp 0
transform 1 0 20332 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1870_
timestamp 0
transform 1 0 19688 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1871_
timestamp 0
transform 1 0 21804 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1872_
timestamp 0
transform 1 0 9476 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1873_
timestamp 0
transform 1 0 12512 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1874_
timestamp 0
transform 1 0 24748 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1875_
timestamp 0
transform 1 0 22908 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1876_
timestamp 0
transform 1 0 33396 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1877_
timestamp 0
transform 1 0 23184 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1878_
timestamp 0
transform 1 0 22540 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1879_
timestamp 0
transform 1 0 4140 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1880_
timestamp 0
transform 1 0 11960 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1881_
timestamp 0
transform 1 0 19136 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1882_
timestamp 0
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1883_
timestamp 0
transform 1 0 26956 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1884_
timestamp 0
transform 1 0 23000 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1885_
timestamp 0
transform 1 0 24380 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1886_
timestamp 0
transform 1 0 22816 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1887_
timestamp 0
transform 1 0 5796 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1888_
timestamp 0
transform 1 0 12144 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1889_
timestamp 0
transform 1 0 17112 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1890_
timestamp 0
transform 1 0 19872 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1891_
timestamp 0
transform 1 0 29532 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1892_
timestamp 0
transform 1 0 32108 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1893_
timestamp 0
transform 1 0 31464 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1894_
timestamp 0
transform 1 0 19228 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1895_
timestamp 0
transform 1 0 7636 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1896_
timestamp 0
transform 1 0 12880 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1897_
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1898_
timestamp 0
transform 1 0 20792 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1899_
timestamp 0
transform 1 0 29440 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1900_
timestamp 0
transform 1 0 32936 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1901_
timestamp 0
transform 1 0 30728 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1902_
timestamp 0
transform 1 0 22632 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1903_
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1904_
timestamp 0
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1905_
timestamp 0
transform 1 0 17112 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1906_
timestamp 0
transform 1 0 19780 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1907_
timestamp 0
transform 1 0 14536 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1908_
timestamp 0
transform 1 0 21620 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1909_
timestamp 0
transform 1 0 20884 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1910_
timestamp 0
transform 1 0 20700 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1911_
timestamp 0
transform 1 0 11592 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1912_
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1913_
timestamp 0
transform 1 0 17848 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1914_
timestamp 0
transform 1 0 19780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1915_
timestamp 0
transform 1 0 24380 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1916_
timestamp 0
transform 1 0 24932 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1917_
timestamp 0
transform 1 0 24932 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1918_
timestamp 0
transform 1 0 20056 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1919_
timestamp 0
transform 1 0 24380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1920_
timestamp 0
transform 1 0 33120 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1921_
timestamp 0
transform 1 0 32936 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1922_
timestamp 0
transform 1 0 19228 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1923_
timestamp 0
transform 1 0 19412 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1924_
timestamp 0
transform 1 0 15640 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1925_
timestamp 0
transform 1 0 18584 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1926_
timestamp 0
transform 1 0 18860 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1927_
timestamp 0
transform 1 0 15088 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1928_
timestamp 0
transform 1 0 17388 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1929_
timestamp 0
transform 1 0 16468 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1930_
timestamp 0
transform 1 0 16836 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1931_
timestamp 0
transform 1 0 3772 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1932_
timestamp 0
transform 1 0 17388 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1933_
timestamp 0
transform 1 0 17848 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1934_
timestamp 0
transform 1 0 44712 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1935_
timestamp 0
transform 1 0 44896 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1936_
timestamp 0
transform 1 0 44528 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1937_
timestamp 0
transform 1 0 45448 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1938_
timestamp 0
transform 1 0 44988 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1939_
timestamp 0
transform 1 0 46000 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1940_
timestamp 0
transform 1 0 45264 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1941_
timestamp 0
transform 1 0 44252 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1942_
timestamp 0
transform 1 0 42412 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_2  _1943_
timestamp 0
transform 1 0 41124 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1944_
timestamp 0
transform 1 0 43332 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1945_
timestamp 0
transform 1 0 44988 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1946_
timestamp 0
transform 1 0 44528 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_2  _1947_
timestamp 0
transform 1 0 43884 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_1  _1948_
timestamp 0
transform 1 0 45724 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1949_
timestamp 0
transform 1 0 45540 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1950_
timestamp 0
transform 1 0 44988 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1951_
timestamp 0
transform 1 0 46276 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1952_
timestamp 0
transform 1 0 45908 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1953_
timestamp 0
transform 1 0 39836 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1954_
timestamp 0
transform 1 0 40204 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1955_
timestamp 0
transform 1 0 40664 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _1956_
timestamp 0
transform 1 0 40756 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1957_
timestamp 0
transform 1 0 43148 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1958_
timestamp 0
transform 1 0 44988 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1959_
timestamp 0
transform 1 0 40940 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1960_
timestamp 0
transform 1 0 40480 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_1  _1961_
timestamp 0
transform 1 0 41584 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1962_
timestamp 0
transform 1 0 40848 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1963_
timestamp 0
transform 1 0 40112 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1964_
timestamp 0
transform 1 0 41308 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1965_
timestamp 0
transform 1 0 41492 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1966_
timestamp 0
transform 1 0 40480 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2oi_2  _1967_
timestamp 0
transform 1 0 41032 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1968_
timestamp 0
transform 1 0 41768 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1969_
timestamp 0
transform 1 0 40572 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1970_
timestamp 0
transform 1 0 40848 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1971_
timestamp 0
transform 1 0 41400 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1972_
timestamp 0
transform 1 0 38272 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1973_
timestamp 0
transform 1 0 42596 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1974_
timestamp 0
transform 1 0 43148 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1975_
timestamp 0
transform 1 0 43056 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1976_
timestamp 0
transform 1 0 41308 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1977_
timestamp 0
transform 1 0 41860 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1978_
timestamp 0
transform 1 0 40940 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1979_
timestamp 0
transform 1 0 38732 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1980_
timestamp 0
transform 1 0 44160 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1981_
timestamp 0
transform 1 0 43700 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1982_
timestamp 0
transform 1 0 43516 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_2  _1983_
timestamp 0
transform 1 0 42228 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__a2bb2oi_2  _1984_
timestamp 0
transform 1 0 43792 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1985_
timestamp 0
transform 1 0 43884 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1986_
timestamp 0
transform 1 0 44068 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1987_
timestamp 0
transform 1 0 44988 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1988_
timestamp 0
transform 1 0 44528 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1989_
timestamp 0
transform 1 0 39192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1990_
timestamp 0
transform 1 0 44988 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1991_
timestamp 0
transform 1 0 45908 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1992_
timestamp 0
transform 1 0 44620 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_4  _1993_
timestamp 0
transform 1 0 45264 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1994_
timestamp 0
transform 1 0 46460 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _1995_
timestamp 0
transform 1 0 45448 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1996_
timestamp 0
transform 1 0 46368 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1997_
timestamp 0
transform 1 0 43240 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1998_
timestamp 0
transform 1 0 42780 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1999_
timestamp 0
transform 1 0 43332 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2000_
timestamp 0
transform 1 0 44620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2001_
timestamp 0
transform 1 0 44988 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _2002_
timestamp 0
transform 1 0 44252 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2003_
timestamp 0
transform 1 0 38732 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _2004_
timestamp 0
transform 1 0 41124 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _2005_
timestamp 0
transform 1 0 43056 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _2006_
timestamp 0
transform 1 0 44160 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2007_
timestamp 0
transform 1 0 44068 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2008_
timestamp 0
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2009_
timestamp 0
transform 1 0 44068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _2010_
timestamp 0
transform 1 0 44620 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _2011_
timestamp 0
transform 1 0 38548 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _2012_
timestamp 0
transform 1 0 42412 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2013_
timestamp 0
transform 1 0 43792 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_2  _2014_
timestamp 0
transform 1 0 43976 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _2015_
timestamp 0
transform 1 0 44804 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2016_
timestamp 0
transform 1 0 41952 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2017_
timestamp 0
transform 1 0 42504 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2018_
timestamp 0
transform 1 0 43608 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2019_
timestamp 0
transform 1 0 45264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2020_
timestamp 0
transform 1 0 44804 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2021_
timestamp 0
transform 1 0 42780 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _2022_
timestamp 0
transform 1 0 43148 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2023_
timestamp 0
transform 1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2024_
timestamp 0
transform 1 0 43884 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2025_
timestamp 0
transform 1 0 44988 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2026_
timestamp 0
transform 1 0 42964 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _2027_
timestamp 0
transform 1 0 43148 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2028_
timestamp 0
transform 1 0 39836 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _2029_
timestamp 0
transform 1 0 42964 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2030_
timestamp 0
transform 1 0 42964 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2031_
timestamp 0
transform 1 0 43884 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2032_
timestamp 0
transform 1 0 43884 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2033_
timestamp 0
transform 1 0 41032 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _2034_
timestamp 0
transform 1 0 41124 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _2035_
timestamp 0
transform 1 0 41768 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2036_
timestamp 0
transform 1 0 43424 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2037_
timestamp 0
transform 1 0 43792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2038_
timestamp 0
transform 1 0 43148 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2039_
timestamp 0
transform 1 0 42780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2040_
timestamp 0
transform 1 0 42780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_2  _2041_
timestamp 0
transform 1 0 42412 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _2042_
timestamp 0
transform 1 0 42780 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2043_
timestamp 0
transform 1 0 37904 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2044_
timestamp 0
transform 1 0 38088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2045_
timestamp 0
transform 1 0 39100 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2046_
timestamp 0
transform 1 0 41492 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _2047_
timestamp 0
transform 1 0 41492 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__xor2_1  _2048_
timestamp 0
transform 1 0 40204 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2049_
timestamp 0
transform 1 0 37720 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2050_
timestamp 0
transform 1 0 38180 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2051_
timestamp 0
transform 1 0 37536 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2052_
timestamp 0
transform 1 0 39008 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2053_
timestamp 0
transform 1 0 39192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2054_
timestamp 0
transform 1 0 41124 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _2055_
timestamp 0
transform 1 0 38640 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2oi_1  _2056_
timestamp 0
transform 1 0 38364 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2057_
timestamp 0
transform 1 0 39560 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2058_
timestamp 0
transform 1 0 34684 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2059_
timestamp 0
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2060_
timestamp 0
transform 1 0 36340 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _2061_
timestamp 0
transform 1 0 36800 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2062_
timestamp 0
transform 1 0 36708 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2063_
timestamp 0
transform 1 0 39192 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _2064_
timestamp 0
transform 1 0 36892 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2065_
timestamp 0
transform 1 0 39284 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2066_
timestamp 0
transform 1 0 39836 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2067_
timestamp 0
transform 1 0 43884 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2068_
timestamp 0
transform 1 0 39744 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _2069_
timestamp 0
transform 1 0 38456 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _2070_
timestamp 0
transform 1 0 36064 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _2071_
timestamp 0
transform 1 0 31096 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2072_
timestamp 0
transform 1 0 15180 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2073_
timestamp 0
transform 1 0 12604 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2074_
timestamp 0
transform 1 0 11684 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _2075_
timestamp 0
transform 1 0 14996 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2076_
timestamp 0
transform 1 0 11500 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_4  _2077_
timestamp 0
transform 1 0 14996 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _2078_
timestamp 0
transform 1 0 17388 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2079_
timestamp 0
transform 1 0 32384 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2080_
timestamp 0
transform 1 0 30636 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2081_
timestamp 0
transform 1 0 44988 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2082_
timestamp 0
transform 1 0 45080 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2083_
timestamp 0
transform 1 0 45448 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2084_
timestamp 0
transform 1 0 43516 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _2085_
timestamp 0
transform 1 0 46092 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2086_
timestamp 0
transform 1 0 40204 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2087_
timestamp 0
transform 1 0 40388 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2088_
timestamp 0
transform 1 0 44344 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2089_
timestamp 0
transform 1 0 44160 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2090_
timestamp 0
transform 1 0 37628 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2091_
timestamp 0
transform 1 0 37260 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2092_
timestamp 0
transform 1 0 36616 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2093_
timestamp 0
transform 1 0 37260 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2094_
timestamp 0
transform 1 0 37260 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _2095_
timestamp 0
transform 1 0 36892 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2096_
timestamp 0
transform 1 0 16652 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2097_
timestamp 0
transform 1 0 12604 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2098_
timestamp 0
transform 1 0 12236 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2099_
timestamp 0
transform 1 0 39836 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _2100_
timestamp 0
transform 1 0 41768 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2101_
timestamp 0
transform 1 0 41952 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _2102_
timestamp 0
transform 1 0 43884 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _2103_
timestamp 0
transform 1 0 39836 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2104_
timestamp 0
transform 1 0 41032 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2105_
timestamp 0
transform 1 0 42504 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _2106_
timestamp 0
transform 1 0 41676 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2107_
timestamp 0
transform 1 0 41584 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _2108_
timestamp 0
transform 1 0 31096 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2109_
timestamp 0
transform 1 0 36156 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _2110_
timestamp 0
transform 1 0 36064 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2111_
timestamp 0
transform 1 0 14628 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2112_
timestamp 0
transform 1 0 11776 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2113_
timestamp 0
transform 1 0 11132 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2114_
timestamp 0
transform 1 0 41216 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2115_
timestamp 0
transform 1 0 42228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _2116_
timestamp 0
transform 1 0 42412 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2117_
timestamp 0
transform 1 0 41676 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2118_
timestamp 0
transform 1 0 41308 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2119_
timestamp 0
transform 1 0 39836 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _2120_
timestamp 0
transform 1 0 38732 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _2121_
timestamp 0
transform 1 0 34684 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2122_
timestamp 0
transform 1 0 31004 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _2123_
timestamp 0
transform 1 0 32108 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2124_
timestamp 0
transform 1 0 30268 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2125_
timestamp 0
transform 1 0 40204 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2126_
timestamp 0
transform 1 0 42412 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2127_
timestamp 0
transform 1 0 41584 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2128_
timestamp 0
transform 1 0 43148 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2129_
timestamp 0
transform 1 0 44252 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2130_
timestamp 0
transform 1 0 42320 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2131_
timestamp 0
transform 1 0 43884 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _2132_
timestamp 0
transform 1 0 42780 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2133_
timestamp 0
transform 1 0 42136 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2134_
timestamp 0
transform 1 0 38180 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _2135_
timestamp 0
transform 1 0 34684 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _2136_
timestamp 0
transform 1 0 29992 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2137_
timestamp 0
transform 1 0 29808 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2138_
timestamp 0
transform 1 0 29716 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2139_
timestamp 0
transform 1 0 42412 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2140_
timestamp 0
transform 1 0 41768 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2141_
timestamp 0
transform 1 0 41768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2142_
timestamp 0
transform 1 0 42412 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2143_
timestamp 0
transform 1 0 37904 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2144_
timestamp 0
transform 1 0 39744 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2145_
timestamp 0
transform 1 0 35512 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _2146_
timestamp 0
transform 1 0 36708 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2147_
timestamp 0
transform 1 0 33580 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _2148_
timestamp 0
transform 1 0 32016 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2149_
timestamp 0
transform 1 0 31740 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _2150_
timestamp 0
transform 1 0 44528 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_2  _2151_
timestamp 0
transform 1 0 43056 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2152_
timestamp 0
transform 1 0 41584 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2153_
timestamp 0
transform 1 0 42412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _2154_
timestamp 0
transform 1 0 42228 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_2  _2155_
timestamp 0
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _2156_
timestamp 0
transform 1 0 40480 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2157_
timestamp 0
transform 1 0 41124 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2158_
timestamp 0
transform 1 0 35420 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _2159_
timestamp 0
transform 1 0 36248 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2160_
timestamp 0
transform 1 0 33672 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _2161_
timestamp 0
transform 1 0 32476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2162_
timestamp 0
transform 1 0 34684 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2163_
timestamp 0
transform 1 0 34040 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2164_
timestamp 0
transform 1 0 41584 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2165_
timestamp 0
transform 1 0 46184 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2166_
timestamp 0
transform 1 0 41216 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _2167_
timestamp 0
transform 1 0 41492 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _2168_
timestamp 0
transform 1 0 39192 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _2169_
timestamp 0
transform 1 0 39284 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _2170_
timestamp 0
transform 1 0 40204 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2171_
timestamp 0
transform 1 0 38272 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2172_
timestamp 0
transform 1 0 33028 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _2173_
timestamp 0
transform 1 0 33580 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2174_
timestamp 0
transform 1 0 33120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2175_
timestamp 0
transform 1 0 38364 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _2176_
timestamp 0
transform 1 0 42596 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2177_
timestamp 0
transform 1 0 43884 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _2178_
timestamp 0
transform 1 0 42872 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2179_
timestamp 0
transform 1 0 43240 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _2180_
timestamp 0
transform 1 0 42412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _2181_
timestamp 0
transform 1 0 43056 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2182_
timestamp 0
transform 1 0 41952 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2183_
timestamp 0
transform 1 0 42136 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2184_
timestamp 0
transform 1 0 43332 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2185_
timestamp 0
transform 1 0 42412 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _2186_
timestamp 0
transform 1 0 37812 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _2187_
timestamp 0
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2188_
timestamp 0
transform 1 0 23184 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2189_
timestamp 0
transform 1 0 23000 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2190_
timestamp 0
transform 1 0 42412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2191_
timestamp 0
transform 1 0 41676 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2192_
timestamp 0
transform 1 0 41492 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2193_
timestamp 0
transform 1 0 40848 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2194_
timestamp 0
transform 1 0 37904 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _2195_
timestamp 0
transform 1 0 37536 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2196_
timestamp 0
transform 1 0 33580 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _2197_
timestamp 0
transform 1 0 33764 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2198_
timestamp 0
transform 1 0 34224 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _2199_
timestamp 0
transform 1 0 40204 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _2200_
timestamp 0
transform 1 0 41768 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _2201_
timestamp 0
transform 1 0 41124 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _2202_
timestamp 0
transform 1 0 40756 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2203_
timestamp 0
transform 1 0 41492 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _2204_
timestamp 0
transform 1 0 40572 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _2205_
timestamp 0
transform 1 0 40020 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _2206_
timestamp 0
transform 1 0 38364 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _2207_
timestamp 0
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2208_
timestamp 0
transform 1 0 33672 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2209_
timestamp 0
transform 1 0 33396 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2210_
timestamp 0
transform 1 0 38364 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2211_
timestamp 0
transform 1 0 41124 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2212_
timestamp 0
transform 1 0 40480 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2213_
timestamp 0
transform 1 0 39836 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_4  _2214_
timestamp 0
transform 1 0 39928 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__o2bb2ai_4  _2215_
timestamp 0
transform 1 0 36800 0 1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_2  _2216_
timestamp 0
transform 1 0 22448 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2217_
timestamp 0
transform 1 0 23000 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2218_
timestamp 0
transform 1 0 22816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2219_
timestamp 0
transform 1 0 39928 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2220_
timestamp 0
transform 1 0 40572 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _2221_
timestamp 0
transform 1 0 42412 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2222_
timestamp 0
transform 1 0 42780 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_2  _2223_
timestamp 0
transform 1 0 42228 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _2224_
timestamp 0
transform 1 0 43332 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2225_
timestamp 0
transform 1 0 42504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2226_
timestamp 0
transform 1 0 44160 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2227_
timestamp 0
transform 1 0 43056 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _2228_
timestamp 0
transform 1 0 35880 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _2229_
timestamp 0
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2230_
timestamp 0
transform 1 0 33396 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2231_
timestamp 0
transform 1 0 31924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2232_
timestamp 0
transform 1 0 42412 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2233_
timestamp 0
transform 1 0 42688 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2234_
timestamp 0
transform 1 0 43056 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2235_
timestamp 0
transform 1 0 42964 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2236_
timestamp 0
transform 1 0 42596 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2237_
timestamp 0
transform 1 0 39836 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _2238_
timestamp 0
transform 1 0 37444 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _2239_
timestamp 0
transform 1 0 33672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2240_
timestamp 0
transform 1 0 31832 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2241_
timestamp 0
transform 1 0 32292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2242_
timestamp 0
transform 1 0 43424 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2243_
timestamp 0
transform 1 0 42688 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2244_
timestamp 0
transform 1 0 40756 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2245_
timestamp 0
transform 1 0 40388 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2246_
timestamp 0
transform 1 0 40020 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2247_
timestamp 0
transform 1 0 40112 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _2248_
timestamp 0
transform 1 0 40572 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2249_
timestamp 0
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _2250_
timestamp 0
transform 1 0 36156 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2251_
timestamp 0
transform 1 0 15548 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _2252_
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2253_
timestamp 0
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2254_
timestamp 0
transform 1 0 38548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2255_
timestamp 0
transform 1 0 38548 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2256_
timestamp 0
transform 1 0 38732 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _2257_
timestamp 0
transform 1 0 39192 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2258_
timestamp 0
transform 1 0 39376 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _2259_
timestamp 0
transform 1 0 38640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2260_
timestamp 0
transform 1 0 38364 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _2261_
timestamp 0
transform 1 0 38272 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2262_
timestamp 0
transform 1 0 24748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2263_
timestamp 0
transform 1 0 24564 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2264_
timestamp 0
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2265_
timestamp 0
transform 1 0 14720 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _2266_
timestamp 0
transform 1 0 17480 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _2267_
timestamp 0
transform 1 0 12696 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2268_
timestamp 0
transform 1 0 14720 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_4  _2269_
timestamp 0
transform 1 0 16652 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  _2270_
timestamp 0
transform 1 0 18216 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2271_
timestamp 0
transform 1 0 32108 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2272_
timestamp 0
transform 1 0 31372 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2273_
timestamp 0
transform 1 0 14536 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2274_
timestamp 0
transform 1 0 13340 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2275_
timestamp 0
transform 1 0 13156 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2276_
timestamp 0
transform 1 0 12236 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2277_
timestamp 0
transform 1 0 32108 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2278_
timestamp 0
transform 1 0 31924 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2279_
timestamp 0
transform 1 0 30176 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2280_
timestamp 0
transform 1 0 29716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2281_
timestamp 0
transform 1 0 33028 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2282_
timestamp 0
transform 1 0 33856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2283_
timestamp 0
transform 1 0 33764 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2284_
timestamp 0
transform 1 0 34684 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2285_
timestamp 0
transform 1 0 35236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2286_
timestamp 0
transform 1 0 35328 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2287_
timestamp 0
transform 1 0 34776 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2288_
timestamp 0
transform 1 0 24380 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2289_
timestamp 0
transform 1 0 23368 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2290_
timestamp 0
transform 1 0 33764 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2291_
timestamp 0
transform 1 0 33488 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2292_
timestamp 0
transform 1 0 34684 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2293_
timestamp 0
transform 1 0 35512 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2294_
timestamp 0
transform 1 0 24380 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2295_
timestamp 0
transform 1 0 24932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2296_
timestamp 0
transform 1 0 32568 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2297_
timestamp 0
transform 1 0 31832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2298_
timestamp 0
transform 1 0 33580 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2299_
timestamp 0
transform 1 0 34132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2300_
timestamp 0
transform 1 0 22264 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2301_
timestamp 0
transform 1 0 23092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2302_
timestamp 0
transform 1 0 25760 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2303_
timestamp 0
transform 1 0 25944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2304_
timestamp 0
transform 1 0 11960 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_4  _2305_
timestamp 0
transform 1 0 16468 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  _2306_
timestamp 0
transform 1 0 17756 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2307_
timestamp 0
transform 1 0 30820 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2308_
timestamp 0
transform 1 0 30544 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2309_
timestamp 0
transform 1 0 12604 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2310_
timestamp 0
transform 1 0 11500 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2311_
timestamp 0
transform 1 0 12420 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2312_
timestamp 0
transform 1 0 10488 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2313_
timestamp 0
transform 1 0 31096 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2314_
timestamp 0
transform 1 0 30820 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2315_
timestamp 0
transform 1 0 30452 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2316_
timestamp 0
transform 1 0 29532 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2317_
timestamp 0
transform 1 0 31832 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2318_
timestamp 0
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2319_
timestamp 0
transform 1 0 32108 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2320_
timestamp 0
transform 1 0 33028 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2321_
timestamp 0
transform 1 0 32660 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2322_
timestamp 0
transform 1 0 32384 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2323_
timestamp 0
transform 1 0 32200 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2324_
timestamp 0
transform 1 0 22264 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2325_
timestamp 0
transform 1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2326_
timestamp 0
transform 1 0 32936 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2327_
timestamp 0
transform 1 0 32476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2328_
timestamp 0
transform 1 0 32476 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2329_
timestamp 0
transform 1 0 32200 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2330_
timestamp 0
transform 1 0 23092 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2331_
timestamp 0
transform 1 0 21988 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2332_
timestamp 0
transform 1 0 31004 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2333_
timestamp 0
transform 1 0 30820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2334_
timestamp 0
transform 1 0 32016 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2335_
timestamp 0
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2336_
timestamp 0
transform 1 0 19964 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2337_
timestamp 0
transform 1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2338_
timestamp 0
transform 1 0 23460 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2339_
timestamp 0
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2340_
timestamp 0
transform 1 0 12420 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_4  _2341_
timestamp 0
transform 1 0 16376 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  _2342_
timestamp 0
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2343_
timestamp 0
transform 1 0 21804 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2344_
timestamp 0
transform 1 0 21896 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2345_
timestamp 0
transform 1 0 16284 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2346_
timestamp 0
transform 1 0 16100 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2347_
timestamp 0
transform 1 0 15180 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2348_
timestamp 0
transform 1 0 14628 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2349_
timestamp 0
transform 1 0 27140 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2350_
timestamp 0
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2351_
timestamp 0
transform 1 0 26956 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2352_
timestamp 0
transform 1 0 26220 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2353_
timestamp 0
transform 1 0 27600 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2354_
timestamp 0
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2355_
timestamp 0
transform 1 0 19872 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2356_
timestamp 0
transform 1 0 31372 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2357_
timestamp 0
transform 1 0 32108 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2358_
timestamp 0
transform 1 0 30820 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2359_
timestamp 0
transform 1 0 30820 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2360_
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2361_
timestamp 0
transform 1 0 18676 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2362_
timestamp 0
transform 1 0 31556 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2363_
timestamp 0
transform 1 0 32384 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2364_
timestamp 0
transform 1 0 23460 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2365_
timestamp 0
transform 1 0 22448 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2366_
timestamp 0
transform 1 0 21712 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2367_
timestamp 0
transform 1 0 20240 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2368_
timestamp 0
transform 1 0 17664 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2369_
timestamp 0
transform 1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2370_
timestamp 0
transform 1 0 20424 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2371_
timestamp 0
transform 1 0 18676 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2372_
timestamp 0
transform 1 0 17112 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2373_
timestamp 0
transform 1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2374_
timestamp 0
transform 1 0 19228 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2375_
timestamp 0
transform 1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2376_
timestamp 0
transform 1 0 13708 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _2377_
timestamp 0
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _2378_
timestamp 0
transform 1 0 14628 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _2379_
timestamp 0
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2380_
timestamp 0
transform 1 0 24012 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2381_
timestamp 0
transform 1 0 23920 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2382_
timestamp 0
transform 1 0 19044 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2383_
timestamp 0
transform 1 0 18308 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2384_
timestamp 0
transform 1 0 17296 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2385_
timestamp 0
transform 1 0 16744 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2386_
timestamp 0
transform 1 0 30360 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2387_
timestamp 0
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2388_
timestamp 0
transform 1 0 27876 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2389_
timestamp 0
transform 1 0 27140 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2390_
timestamp 0
transform 1 0 29164 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2391_
timestamp 0
transform 1 0 29992 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2392_
timestamp 0
transform 1 0 29808 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2393_
timestamp 0
transform 1 0 31188 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2394_
timestamp 0
transform 1 0 31096 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2395_
timestamp 0
transform 1 0 31188 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2396_
timestamp 0
transform 1 0 30084 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2397_
timestamp 0
transform 1 0 27416 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2398_
timestamp 0
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2399_
timestamp 0
transform 1 0 31188 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2400_
timestamp 0
transform 1 0 31188 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2401_
timestamp 0
transform 1 0 27232 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2402_
timestamp 0
transform 1 0 27784 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2403_
timestamp 0
transform 1 0 27048 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2404_
timestamp 0
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2405_
timestamp 0
transform 1 0 29532 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2406_
timestamp 0
transform 1 0 28980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2407_
timestamp 0
transform 1 0 29716 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2408_
timestamp 0
transform 1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2409_
timestamp 0
transform 1 0 14720 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2410_
timestamp 0
transform 1 0 14536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2411_
timestamp 0
transform 1 0 25668 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2412_
timestamp 0
transform 1 0 24472 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2413_
timestamp 0
transform 1 0 20792 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2414_
timestamp 0
transform 1 0 12144 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _2415_
timestamp 0
transform 1 0 13340 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2416_
timestamp 0
transform 1 0 6164 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2417_
timestamp 0
transform 1 0 6624 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2418_
timestamp 0
transform 1 0 6256 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2419_
timestamp 0
transform 1 0 15824 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2420_
timestamp 0
transform 1 0 3128 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2421_
timestamp 0
transform 1 0 1472 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2422_
timestamp 0
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2423_
timestamp 0
transform 1 0 8004 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2424_
timestamp 0
transform 1 0 6256 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2425_
timestamp 0
transform 1 0 23460 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2426_
timestamp 0
transform 1 0 7820 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2427_
timestamp 0
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2428_
timestamp 0
transform 1 0 23000 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2429_
timestamp 0
transform 1 0 3036 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2430_
timestamp 0
transform 1 0 3588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2431_
timestamp 0
transform 1 0 23092 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2432_
timestamp 0
transform 1 0 2392 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2433_
timestamp 0
transform 1 0 2024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2434_
timestamp 0
transform 1 0 15824 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2435_
timestamp 0
transform 1 0 6532 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2436_
timestamp 0
transform 1 0 2576 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2437_
timestamp 0
transform 1 0 2116 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2438_
timestamp 0
transform 1 0 17480 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2439_
timestamp 0
transform 1 0 3220 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2440_
timestamp 0
transform 1 0 2208 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2441_
timestamp 0
transform 1 0 15364 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _2442_
timestamp 0
transform 1 0 7452 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2443_
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2444_
timestamp 0
transform 1 0 16836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2445_
timestamp 0
transform 1 0 6624 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2446_
timestamp 0
transform 1 0 5520 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2447_
timestamp 0
transform 1 0 17296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2448_
timestamp 0
transform 1 0 8464 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2449_
timestamp 0
transform 1 0 7452 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2450_
timestamp 0
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2451_
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2452_
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2453_
timestamp 0
transform 1 0 16560 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2454_
timestamp 0
transform 1 0 5152 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2455_
timestamp 0
transform 1 0 4232 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2456_
timestamp 0
transform 1 0 17848 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2457_
timestamp 0
transform 1 0 7636 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2458_
timestamp 0
transform 1 0 5888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2459_
timestamp 0
transform 1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2460_
timestamp 0
transform 1 0 10580 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2461_
timestamp 0
transform 1 0 9476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2462_
timestamp 0
transform 1 0 17204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2463_
timestamp 0
transform 1 0 9660 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2464_
timestamp 0
transform 1 0 9292 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _2465_
timestamp 0
transform 1 0 11592 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2466_
timestamp 0
transform 1 0 6256 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2467_
timestamp 0
transform 1 0 6624 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2468_
timestamp 0
transform 1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2469_
timestamp 0
transform 1 0 2576 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2470_
timestamp 0
transform 1 0 2208 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2471_
timestamp 0
transform 1 0 7084 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2472_
timestamp 0
transform 1 0 6808 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2473_
timestamp 0
transform 1 0 6992 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2474_
timestamp 0
transform 1 0 6716 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2475_
timestamp 0
transform 1 0 3772 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2476_
timestamp 0
transform 1 0 1840 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2477_
timestamp 0
transform 1 0 2576 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2478_
timestamp 0
transform 1 0 2116 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2479_
timestamp 0
transform 1 0 6992 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2480_
timestamp 0
transform 1 0 2576 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2481_
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2482_
timestamp 0
transform 1 0 2576 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2483_
timestamp 0
transform 1 0 2116 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2484_
timestamp 0
transform 1 0 7544 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2485_
timestamp 0
transform 1 0 6624 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2486_
timestamp 0
transform 1 0 6532 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2487_
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2488_
timestamp 0
transform 1 0 7636 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2489_
timestamp 0
transform 1 0 6900 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2490_
timestamp 0
transform 1 0 3772 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2491_
timestamp 0
transform 1 0 2760 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2492_
timestamp 0
transform 1 0 4784 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2493_
timestamp 0
transform 1 0 4140 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2494_
timestamp 0
transform 1 0 6716 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2495_
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2496_
timestamp 0
transform 1 0 10396 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2497_
timestamp 0
transform 1 0 9200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2498_
timestamp 0
transform 1 0 10488 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2499_
timestamp 0
transform 1 0 9384 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _2500_
timestamp 0
transform 1 0 12328 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2501_
timestamp 0
transform 1 0 8188 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2502_
timestamp 0
transform 1 0 7636 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2503_
timestamp 0
transform 1 0 7360 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2504_
timestamp 0
transform 1 0 4416 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2505_
timestamp 0
transform 1 0 3680 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2506_
timestamp 0
transform 1 0 8924 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2507_
timestamp 0
transform 1 0 8188 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2508_
timestamp 0
transform 1 0 8004 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2509_
timestamp 0
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2510_
timestamp 0
transform 1 0 4048 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2511_
timestamp 0
transform 1 0 3496 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2512_
timestamp 0
transform 1 0 3772 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2513_
timestamp 0
transform 1 0 3128 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2514_
timestamp 0
transform 1 0 7636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2515_
timestamp 0
transform 1 0 3496 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2516_
timestamp 0
transform 1 0 3956 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2517_
timestamp 0
transform 1 0 4508 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2518_
timestamp 0
transform 1 0 4232 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2519_
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2520_
timestamp 0
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2521_
timestamp 0
transform 1 0 8004 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2522_
timestamp 0
transform 1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2523_
timestamp 0
transform 1 0 8740 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2524_
timestamp 0
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2525_
timestamp 0
transform 1 0 4140 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2526_
timestamp 0
transform 1 0 3864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2527_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2528_
timestamp 0
transform 1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2529_
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2530_
timestamp 0
transform 1 0 7728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2531_
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2532_
timestamp 0
transform 1 0 10396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2533_
timestamp 0
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2534_
timestamp 0
transform 1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2535_
timestamp 0
transform 1 0 13432 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _2536_
timestamp 0
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2537_
timestamp 0
transform 1 0 9660 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2538_
timestamp 0
transform 1 0 10488 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2539_
timestamp 0
transform 1 0 9292 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2540_
timestamp 0
transform 1 0 4048 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2541_
timestamp 0
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2542_
timestamp 0
transform 1 0 10672 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2543_
timestamp 0
transform 1 0 9384 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2544_
timestamp 0
transform 1 0 9660 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2545_
timestamp 0
transform 1 0 9016 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2546_
timestamp 0
transform 1 0 5244 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2547_
timestamp 0
transform 1 0 4140 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2548_
timestamp 0
transform 1 0 4324 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2549_
timestamp 0
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2550_
timestamp 0
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2551_
timestamp 0
transform 1 0 6440 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2552_
timestamp 0
transform 1 0 5336 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2553_
timestamp 0
transform 1 0 5336 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2554_
timestamp 0
transform 1 0 4508 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2555_
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2556_
timestamp 0
transform 1 0 9660 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2557_
timestamp 0
transform 1 0 9752 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2558_
timestamp 0
transform 1 0 10672 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2559_
timestamp 0
transform 1 0 10304 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2560_
timestamp 0
transform 1 0 10028 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2561_
timestamp 0
transform 1 0 5060 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2562_
timestamp 0
transform 1 0 3864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2563_
timestamp 0
transform 1 0 7728 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2564_
timestamp 0
transform 1 0 6900 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2565_
timestamp 0
transform 1 0 8004 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2566_
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2567_
timestamp 0
transform 1 0 11684 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2568_
timestamp 0
transform 1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2569_
timestamp 0
transform 1 0 13432 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2570_
timestamp 0
transform 1 0 11500 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _2571_
timestamp 0
transform 1 0 12604 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _2572_
timestamp 0
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2573_
timestamp 0
transform 1 0 14168 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2574_
timestamp 0
transform 1 0 19688 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2575_
timestamp 0
transform 1 0 20700 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2576_
timestamp 0
transform 1 0 16652 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2577_
timestamp 0
transform 1 0 15456 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2578_
timestamp 0
transform 1 0 14996 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2579_
timestamp 0
transform 1 0 13432 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2580_
timestamp 0
transform 1 0 22356 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2581_
timestamp 0
transform 1 0 23184 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2582_
timestamp 0
transform 1 0 21896 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2583_
timestamp 0
transform 1 0 21620 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2584_
timestamp 0
transform 1 0 21804 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2585_
timestamp 0
transform 1 0 21528 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2586_
timestamp 0
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2587_
timestamp 0
transform 1 0 13248 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2588_
timestamp 0
transform 1 0 12972 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2589_
timestamp 0
transform 1 0 14076 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2590_
timestamp 0
transform 1 0 15180 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2591_
timestamp 0
transform 1 0 13064 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2592_
timestamp 0
transform 1 0 12880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2593_
timestamp 0
transform 1 0 13524 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2594_
timestamp 0
transform 1 0 11776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2595_
timestamp 0
transform 1 0 14352 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2596_
timestamp 0
transform 1 0 13248 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2597_
timestamp 0
transform 1 0 12788 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2598_
timestamp 0
transform 1 0 12512 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2599_
timestamp 0
transform 1 0 14536 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2600_
timestamp 0
transform 1 0 14444 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2601_
timestamp 0
transform 1 0 13524 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2602_
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2603_
timestamp 0
transform 1 0 13156 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2604_
timestamp 0
transform 1 0 14352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2605_
timestamp 0
transform 1 0 14076 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2606_
timestamp 0
transform 1 0 13800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _2607_
timestamp 0
transform 1 0 15548 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _2608_
timestamp 0
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2609_
timestamp 0
transform 1 0 19504 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2610_
timestamp 0
transform 1 0 19320 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2611_
timestamp 0
transform 1 0 15548 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2612_
timestamp 0
transform 1 0 15180 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2613_
timestamp 0
transform 1 0 14260 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2614_
timestamp 0
transform 1 0 13708 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2615_
timestamp 0
transform 1 0 21988 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2616_
timestamp 0
transform 1 0 21988 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2617_
timestamp 0
transform 1 0 20884 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2618_
timestamp 0
transform 1 0 20608 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2619_
timestamp 0
transform 1 0 21804 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2620_
timestamp 0
transform 1 0 21068 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2621_
timestamp 0
transform 1 0 16008 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2622_
timestamp 0
transform 1 0 14996 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2623_
timestamp 0
transform 1 0 14720 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2624_
timestamp 0
transform 1 0 16652 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2625_
timestamp 0
transform 1 0 15732 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2626_
timestamp 0
transform 1 0 14168 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2627_
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2628_
timestamp 0
transform 1 0 14904 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2629_
timestamp 0
transform 1 0 14628 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2630_
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2631_
timestamp 0
transform 1 0 15364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2632_
timestamp 0
transform 1 0 15272 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2633_
timestamp 0
transform 1 0 14536 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2634_
timestamp 0
transform 1 0 15732 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2635_
timestamp 0
transform 1 0 15088 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2636_
timestamp 0
transform 1 0 16008 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2637_
timestamp 0
transform 1 0 15916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2638_
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2639_
timestamp 0
transform 1 0 14628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2640_
timestamp 0
transform 1 0 15456 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2641_
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_4  _2642_
timestamp 0
transform 1 0 14720 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _2643_
timestamp 0
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2644_
timestamp 0
transform 1 0 24840 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2645_
timestamp 0
transform 1 0 24196 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2646_
timestamp 0
transform 1 0 18308 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2647_
timestamp 0
transform 1 0 18032 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2648_
timestamp 0
transform 1 0 17756 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2649_
timestamp 0
transform 1 0 18584 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2650_
timestamp 0
transform 1 0 29532 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2651_
timestamp 0
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2652_
timestamp 0
transform 1 0 29348 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2653_
timestamp 0
transform 1 0 28888 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2654_
timestamp 0
transform 1 0 29348 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2655_
timestamp 0
transform 1 0 28796 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2656_
timestamp 0
transform 1 0 28980 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2657_
timestamp 0
transform 1 0 32108 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2658_
timestamp 0
transform 1 0 31556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2659_
timestamp 0
transform 1 0 30452 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2660_
timestamp 0
transform 1 0 30268 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2661_
timestamp 0
transform 1 0 27508 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2662_
timestamp 0
transform 1 0 28704 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2663_
timestamp 0
transform 1 0 32108 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2664_
timestamp 0
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2665_
timestamp 0
transform 1 0 28980 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2666_
timestamp 0
transform 1 0 28704 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2667_
timestamp 0
transform 1 0 28888 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2668_
timestamp 0
transform 1 0 27692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2669_
timestamp 0
transform 1 0 29532 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2670_
timestamp 0
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2671_
timestamp 0
transform 1 0 29624 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2672_
timestamp 0
transform 1 0 31280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2673_
timestamp 0
transform 1 0 14996 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2674_
timestamp 0
transform 1 0 14260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2675_
timestamp 0
transform 1 0 25668 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2676_
timestamp 0
transform 1 0 26496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_4  _2677_
timestamp 0
transform 1 0 15640 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  _2678_
timestamp 0
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2679_
timestamp 0
transform 1 0 23092 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2680_
timestamp 0
transform 1 0 21436 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2681_
timestamp 0
transform 1 0 18308 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2682_
timestamp 0
transform 1 0 18216 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2683_
timestamp 0
transform 1 0 16652 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2684_
timestamp 0
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2685_
timestamp 0
transform 1 0 24380 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2686_
timestamp 0
transform 1 0 25208 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2687_
timestamp 0
transform 1 0 23276 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2688_
timestamp 0
transform 1 0 23828 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2689_
timestamp 0
transform 1 0 23460 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2690_
timestamp 0
transform 1 0 22816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2691_
timestamp 0
transform 1 0 18124 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2692_
timestamp 0
transform 1 0 17572 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2693_
timestamp 0
transform 1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2694_
timestamp 0
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2695_
timestamp 0
transform 1 0 19228 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2696_
timestamp 0
transform 1 0 16560 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2697_
timestamp 0
transform 1 0 16284 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2698_
timestamp 0
transform 1 0 17480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2699_
timestamp 0
transform 1 0 17204 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2700_
timestamp 0
transform 1 0 18308 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2701_
timestamp 0
transform 1 0 17388 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2702_
timestamp 0
transform 1 0 17480 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2703_
timestamp 0
transform 1 0 17204 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2704_
timestamp 0
transform 1 0 19044 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2705_
timestamp 0
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2706_
timestamp 0
transform 1 0 19136 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2707_
timestamp 0
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2708_
timestamp 0
transform 1 0 17296 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2709_
timestamp 0
transform 1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2710_
timestamp 0
transform 1 0 17480 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2711_
timestamp 0
transform 1 0 17572 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2712_
timestamp 0
transform 1 0 37260 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2713_
timestamp 0
transform 1 0 35420 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2714_
timestamp 0
transform 1 0 34776 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2715_
timestamp 0
transform 1 0 37260 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2716_
timestamp 0
transform 1 0 36524 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2717_
timestamp 0
transform 1 0 32108 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2718_
timestamp 0
transform 1 0 31464 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2719_
timestamp 0
transform 1 0 31096 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2720_
timestamp 0
transform 1 0 32108 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2721_
timestamp 0
transform 1 0 37260 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2722_
timestamp 0
transform 1 0 36524 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2723_
timestamp 0
transform 1 0 37536 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2724_
timestamp 0
transform 1 0 2944 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2725_
timestamp 0
transform 1 0 13064 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2726_
timestamp 0
transform 1 0 13432 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2727_
timestamp 0
transform 1 0 13248 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2728_
timestamp 0
transform 1 0 13248 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2729_
timestamp 0
transform 1 0 1932 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2730_
timestamp 0
transform 1 0 2760 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2731_
timestamp 0
transform 1 0 8924 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2732_
timestamp 0
transform 1 0 8004 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2733_
timestamp 0
transform 1 0 12696 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2734_
timestamp 0
transform 1 0 10948 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2735_
timestamp 0
transform 1 0 1932 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2736_
timestamp 0
transform 1 0 2024 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2737_
timestamp 0
transform 1 0 5428 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2738_
timestamp 0
transform 1 0 4232 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2739_
timestamp 0
transform 1 0 2208 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2740_
timestamp 0
transform 1 0 1840 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2741_
timestamp 0
transform 1 0 39836 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2742_
timestamp 0
transform 1 0 38732 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2743_
timestamp 0
transform 1 0 1748 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2744_
timestamp 0
transform 1 0 3128 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2745_
timestamp 0
transform 1 0 20148 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2746_
timestamp 0
transform 1 0 20700 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2747_
timestamp 0
transform 1 0 33488 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _2748_
timestamp 0
transform 1 0 27968 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2749_
timestamp 0
transform 1 0 29164 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2750_
timestamp 0
transform 1 0 25668 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2751_
timestamp 0
transform 1 0 28152 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2752_
timestamp 0
transform 1 0 26036 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2753_
timestamp 0
transform 1 0 25392 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2754_
timestamp 0
transform 1 0 33120 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2755_
timestamp 0
transform 1 0 27600 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2756_
timestamp 0
transform 1 0 26220 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2757_
timestamp 0
transform 1 0 21804 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2758_
timestamp 0
transform 1 0 25484 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2759_
timestamp 0
transform 1 0 26956 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2760_
timestamp 0
transform 1 0 29072 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _2761_
timestamp 0
transform 1 0 28520 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  _2762_
timestamp 0
transform 1 0 26404 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2763_
timestamp 0
transform 1 0 26864 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2764_
timestamp 0
transform 1 0 25484 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2765_
timestamp 0
transform 1 0 30360 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2766_
timestamp 0
transform 1 0 31096 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2767_
timestamp 0
transform 1 0 30636 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2768_
timestamp 0
transform 1 0 30360 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2769_
timestamp 0
transform 1 0 33028 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2770_
timestamp 0
transform 1 0 33488 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2771_
timestamp 0
transform 1 0 33396 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2772_
timestamp 0
transform 1 0 32752 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _2773_
timestamp 0
transform 1 0 32292 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _2774_
timestamp 0
transform 1 0 31280 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _2775_
timestamp 0
transform 1 0 30084 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2776_
timestamp 0
transform 1 0 30452 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2777_
timestamp 0
transform 1 0 29900 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2778_
timestamp 0
transform 1 0 29348 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _2779_
timestamp 0
transform 1 0 29532 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2780_
timestamp 0
transform 1 0 30176 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2781_
timestamp 0
transform 1 0 29716 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _2782_
timestamp 0
transform 1 0 29532 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2783_
timestamp 0
transform 1 0 30176 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2784_
timestamp 0
transform 1 0 29532 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2785_
timestamp 0
transform 1 0 28796 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _2786_
timestamp 0
transform 1 0 27876 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2787_
timestamp 0
transform 1 0 29164 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2788_
timestamp 0
transform 1 0 29532 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2789_
timestamp 0
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2790_
timestamp 0
transform 1 0 29348 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2791_
timestamp 0
transform 1 0 29992 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2792_
timestamp 0
transform 1 0 28980 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2793_
timestamp 0
transform 1 0 29624 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _2794_
timestamp 0
transform 1 0 28428 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _2795_
timestamp 0
transform 1 0 27324 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2796_
timestamp 0
transform 1 0 22908 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2797_
timestamp 0
transform 1 0 23000 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _2798_
timestamp 0
transform 1 0 28428 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2799_
timestamp 0
transform 1 0 23092 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2800_
timestamp 0
transform 1 0 25300 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _2801_
timestamp 0
transform 1 0 22356 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2802_
timestamp 0
transform 1 0 21436 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2803_
timestamp 0
transform 1 0 20332 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2804_
timestamp 0
transform 1 0 22540 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2805_
timestamp 0
transform 1 0 23276 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2806_
timestamp 0
transform 1 0 21896 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_2  _2807_
timestamp 0
transform 1 0 22080 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _2808_
timestamp 0
transform 1 0 23000 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2809_
timestamp 0
transform 1 0 22540 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2810_
timestamp 0
transform 1 0 19320 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2811_
timestamp 0
transform 1 0 18860 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2812_
timestamp 0
transform 1 0 19780 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2813_
timestamp 0
transform 1 0 21068 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_1  _2814_
timestamp 0
transform 1 0 26956 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2815_
timestamp 0
transform 1 0 21804 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2816_
timestamp 0
transform 1 0 20608 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2817_
timestamp 0
transform 1 0 19964 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2818_
timestamp 0
transform 1 0 19688 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2819_
timestamp 0
transform 1 0 20884 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2820_
timestamp 0
transform 1 0 20148 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _2821_
timestamp 0
transform 1 0 20792 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2822_
timestamp 0
transform 1 0 20884 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2823_
timestamp 0
transform 1 0 20148 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _2824_
timestamp 0
transform 1 0 25300 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2825_
timestamp 0
transform 1 0 35512 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _2826_
timestamp 0
transform 1 0 34960 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _2827_
timestamp 0
transform 1 0 35236 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2828_
timestamp 0
transform 1 0 34316 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2829_
timestamp 0
transform 1 0 33948 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2830_
timestamp 0
transform 1 0 32568 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_4  _2831_
timestamp 0
transform 1 0 16652 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  _2832_
timestamp 0
transform 1 0 35420 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2833_
timestamp 0
transform 1 0 33672 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2834_
timestamp 0
transform 1 0 34684 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2835_
timestamp 0
transform 1 0 14904 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2836_
timestamp 0
transform 1 0 13616 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2837_
timestamp 0
transform 1 0 13156 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2838_
timestamp 0
transform 1 0 12604 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2839_
timestamp 0
transform 1 0 35144 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2840_
timestamp 0
transform 1 0 33948 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2841_
timestamp 0
transform 1 0 32108 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2842_
timestamp 0
transform 1 0 31464 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2843_
timestamp 0
transform 1 0 35236 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2844_
timestamp 0
transform 1 0 34960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2845_
timestamp 0
transform 1 0 36156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2846_
timestamp 0
transform 1 0 35696 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2847_
timestamp 0
transform 1 0 35696 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2848_
timestamp 0
transform 1 0 36340 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2849_
timestamp 0
transform 1 0 35880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2850_
timestamp 0
transform 1 0 37260 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2851_
timestamp 0
transform 1 0 36616 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2852_
timestamp 0
transform 1 0 37260 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2853_
timestamp 0
transform 1 0 36064 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2854_
timestamp 0
transform 1 0 36340 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2855_
timestamp 0
transform 1 0 36800 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2856_
timestamp 0
transform 1 0 36156 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2857_
timestamp 0
transform 1 0 35420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2858_
timestamp 0
transform 1 0 35052 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2859_
timestamp 0
transform 1 0 35052 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2860_
timestamp 0
transform 1 0 35880 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2861_
timestamp 0
transform 1 0 34960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2862_
timestamp 0
transform 1 0 22448 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2863_
timestamp 0
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2864_
timestamp 0
transform 1 0 27324 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2865_
timestamp 0
transform 1 0 27324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _2866_
timestamp 0
transform 1 0 13800 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _2867_
timestamp 0
transform 1 0 25852 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2868_
timestamp 0
transform 1 0 24104 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2869_
timestamp 0
transform 1 0 23920 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2870_
timestamp 0
transform 1 0 17204 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2871_
timestamp 0
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2872_
timestamp 0
transform 1 0 16376 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2873_
timestamp 0
transform 1 0 17480 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2874_
timestamp 0
transform 1 0 26312 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2875_
timestamp 0
transform 1 0 26036 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2876_
timestamp 0
transform 1 0 27784 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2877_
timestamp 0
transform 1 0 27048 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2878_
timestamp 0
transform 1 0 27324 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2879_
timestamp 0
transform 1 0 28520 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2880_
timestamp 0
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2881_
timestamp 0
transform 1 0 29532 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2882_
timestamp 0
transform 1 0 29164 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2883_
timestamp 0
transform 1 0 27048 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2884_
timestamp 0
transform 1 0 27140 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2885_
timestamp 0
transform 1 0 26404 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2886_
timestamp 0
transform 1 0 26404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2887_
timestamp 0
transform 1 0 29256 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2888_
timestamp 0
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2889_
timestamp 0
transform 1 0 25208 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2890_
timestamp 0
transform 1 0 24748 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2891_
timestamp 0
transform 1 0 26956 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2892_
timestamp 0
transform 1 0 26312 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2893_
timestamp 0
transform 1 0 28428 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2894_
timestamp 0
transform 1 0 27508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2895_
timestamp 0
transform 1 0 28704 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2896_
timestamp 0
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2897_
timestamp 0
transform 1 0 13616 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2898_
timestamp 0
transform 1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2899_
timestamp 0
transform 1 0 26312 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2900_
timestamp 0
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _2901_
timestamp 0
transform 1 0 14076 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _2902_
timestamp 0
transform 1 0 26128 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2903_
timestamp 0
transform 1 0 23184 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2904_
timestamp 0
transform 1 0 23000 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2905_
timestamp 0
transform 1 0 18124 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2906_
timestamp 0
transform 1 0 16008 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2907_
timestamp 0
transform 1 0 16652 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2908_
timestamp 0
transform 1 0 16008 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2909_
timestamp 0
transform 1 0 25024 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2910_
timestamp 0
transform 1 0 24748 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2911_
timestamp 0
transform 1 0 26496 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2912_
timestamp 0
transform 1 0 26496 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2913_
timestamp 0
transform 1 0 26220 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2914_
timestamp 0
transform 1 0 25944 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2915_
timestamp 0
transform 1 0 27876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2916_
timestamp 0
transform 1 0 28612 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2917_
timestamp 0
transform 1 0 29532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2918_
timestamp 0
transform 1 0 26312 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2919_
timestamp 0
transform 1 0 26036 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2920_
timestamp 0
transform 1 0 25944 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2921_
timestamp 0
transform 1 0 24840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2922_
timestamp 0
transform 1 0 28612 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2923_
timestamp 0
transform 1 0 28980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2924_
timestamp 0
transform 1 0 24472 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2925_
timestamp 0
transform 1 0 24472 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2926_
timestamp 0
transform 1 0 25484 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2927_
timestamp 0
transform 1 0 25392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2928_
timestamp 0
transform 1 0 27232 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2929_
timestamp 0
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2930_
timestamp 0
transform 1 0 27508 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2931_
timestamp 0
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2932_
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2933_
timestamp 0
transform 1 0 12972 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2934_
timestamp 0
transform 1 0 23092 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2935_
timestamp 0
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2936_
timestamp 0
transform 1 0 36432 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2937_
timestamp 0
transform 1 0 37352 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2938_
timestamp 0
transform 1 0 37168 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2939_
timestamp 0
transform 1 0 34040 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2940_
timestamp 0
transform 1 0 33396 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _2941_
timestamp 0
transform 1 0 36156 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2942_
timestamp 0
transform 1 0 37260 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _2943_
timestamp 0
transform 1 0 36064 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2944_
timestamp 0
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2945_
timestamp 0
transform 1 0 18124 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2946_
timestamp 0
transform 1 0 16652 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2947_
timestamp 0
transform 1 0 16560 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2948_
timestamp 0
transform 1 0 16284 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2949_
timestamp 0
transform 1 0 16652 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2950_
timestamp 0
transform 1 0 15364 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2951_
timestamp 0
transform 1 0 17112 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2952_
timestamp 0
transform 1 0 16928 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2953_
timestamp 0
transform 1 0 7360 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2954_
timestamp 0
transform 1 0 6992 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2955_
timestamp 0
transform 1 0 6992 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2956_
timestamp 0
transform 1 0 6624 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2957_
timestamp 0
transform 1 0 6348 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2958_
timestamp 0
transform 1 0 5428 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2959_
timestamp 0
transform 1 0 6348 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2960_
timestamp 0
transform 1 0 5428 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2961_
timestamp 0
transform 1 0 9108 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2962_
timestamp 0
transform 1 0 9752 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2963_
timestamp 0
transform 1 0 11500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2964_
timestamp 0
transform 1 0 12696 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2965_
timestamp 0
transform 1 0 11868 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2966_
timestamp 0
transform 1 0 11776 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2967_
timestamp 0
transform 1 0 10396 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2968_
timestamp 0
transform 1 0 9660 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2969_
timestamp 0
transform 1 0 10028 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2970_
timestamp 0
transform 1 0 10580 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2971_
timestamp 0
transform 1 0 10488 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2972_
timestamp 0
transform 1 0 10580 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2973_
timestamp 0
transform 1 0 36432 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2974_
timestamp 0
transform 1 0 36892 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2975_
timestamp 0
transform 1 0 35788 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2976_
timestamp 0
transform 1 0 36340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2977_
timestamp 0
transform 1 0 34500 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2978_
timestamp 0
transform 1 0 36340 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2979_
timestamp 0
transform 1 0 35328 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _2980_
timestamp 0
transform 1 0 34500 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2981_
timestamp 0
transform 1 0 9660 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2982_
timestamp 0
transform 1 0 8832 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2983_
timestamp 0
transform 1 0 26036 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2984_
timestamp 0
transform 1 0 26128 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _2985_
timestamp 0
transform 1 0 35880 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _2986_
timestamp 0
transform 1 0 18216 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2987_
timestamp 0
transform 1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2988_
timestamp 0
transform 1 0 34684 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2989_
timestamp 0
transform 1 0 33396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2990_
timestamp 0
transform 1 0 38364 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2991_
timestamp 0
transform 1 0 39192 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2992_
timestamp 0
transform 1 0 15548 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2993_
timestamp 0
transform 1 0 13432 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2994_
timestamp 0
transform 1 0 9384 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2995_
timestamp 0
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2996_
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2997_
timestamp 0
transform 1 0 10672 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2998_
timestamp 0
transform 1 0 34684 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _2999_
timestamp 0
transform 1 0 35052 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _3000_
timestamp 0
transform 1 0 35696 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _3001_
timestamp 0
transform 1 0 35144 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _3002_
timestamp 0
transform 1 0 34868 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _3003_
timestamp 0
transform 1 0 35328 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _3004_
timestamp 0
transform 1 0 33580 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _3005_
timestamp 0
transform 1 0 30912 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3006_
timestamp 0
transform 1 0 11868 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3007_
timestamp 0
transform 1 0 11500 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3008_
timestamp 0
transform 1 0 30544 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3009_
timestamp 0
transform 1 0 29532 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3010_
timestamp 0
transform 1 0 32108 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3011_
timestamp 0
transform 1 0 34684 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3012_
timestamp 0
transform 1 0 33120 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3013_
timestamp 0
transform 1 0 22632 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3014_
timestamp 0
transform 1 0 33212 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3015_
timestamp 0
transform 1 0 33120 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3016_
timestamp 0
transform 1 0 22448 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3017_
timestamp 0
transform 1 0 32108 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3018_
timestamp 0
transform 1 0 32108 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3019_
timestamp 0
transform 1 0 20792 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3020_
timestamp 0
transform 1 0 24380 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3021_
timestamp 0
transform 1 0 31648 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3022_
timestamp 0
transform 1 0 13064 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3023_
timestamp 0
transform 1 0 12512 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3024_
timestamp 0
transform 1 0 32200 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3025_
timestamp 0
transform 1 0 29992 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3026_
timestamp 0
transform 1 0 33580 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3027_
timestamp 0
transform 1 0 34316 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3028_
timestamp 0
transform 1 0 35328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3029_
timestamp 0
transform 1 0 22816 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3030_
timestamp 0
transform 1 0 34684 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3031_
timestamp 0
transform 1 0 35328 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3032_
timestamp 0
transform 1 0 24380 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3033_
timestamp 0
transform 1 0 32752 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3034_
timestamp 0
transform 1 0 34408 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3035_
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3036_
timestamp 0
transform 1 0 25944 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtp_1  _3037_
timestamp 0
transform 1 0 39560 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3038_
timestamp 0
transform 1 0 37628 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3039_
timestamp 0
transform 1 0 39744 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3040_
timestamp 0
transform 1 0 37352 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3041_
timestamp 0
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3042_
timestamp 0
transform 1 0 36064 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3043_
timestamp 0
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3044_
timestamp 0
transform 1 0 38088 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3045_
timestamp 0
transform 1 0 38548 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3046_
timestamp 0
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3047_
timestamp 0
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3048_
timestamp 0
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3049_
timestamp 0
transform 1 0 35604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3050_
timestamp 0
transform 1 0 37444 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3051_
timestamp 0
transform 1 0 35880 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3052_
timestamp 0
transform 1 0 35696 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3053_
timestamp 0
transform 1 0 34408 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3054_
timestamp 0
transform 1 0 35696 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3055_
timestamp 0
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3056_
timestamp 0
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3057_
timestamp 0
transform 1 0 34408 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3058_
timestamp 0
transform 1 0 23092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3059_
timestamp 0
transform 1 0 37076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3060_
timestamp 0
transform 1 0 22080 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3061_
timestamp 0
transform 1 0 20148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3062_
timestamp 0
transform 1 0 20240 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3063_
timestamp 0
transform 1 0 37168 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3064_
timestamp 0
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3065_
timestamp 0
transform 1 0 19872 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3066_
timestamp 0
transform 1 0 35144 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3067_
timestamp 0
transform 1 0 36248 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _3068_
timestamp 0
transform 1 0 20148 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _3069_
timestamp 0
transform 1 0 30176 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3070_
timestamp 0
transform 1 0 11776 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3071_
timestamp 0
transform 1 0 10764 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3072_
timestamp 0
transform 1 0 30544 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3073_
timestamp 0
transform 1 0 28980 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3074_
timestamp 0
transform 1 0 31740 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3075_
timestamp 0
transform 1 0 32936 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3076_
timestamp 0
transform 1 0 31924 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3077_
timestamp 0
transform 1 0 22632 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3078_
timestamp 0
transform 1 0 32752 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3079_
timestamp 0
transform 1 0 31924 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3080_
timestamp 0
transform 1 0 21620 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3081_
timestamp 0
transform 1 0 30452 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3082_
timestamp 0
transform 1 0 32108 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3083_
timestamp 0
transform 1 0 19504 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3084_
timestamp 0
transform 1 0 23460 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3085_
timestamp 0
transform 1 0 9016 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3086_
timestamp 0
transform 1 0 8004 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3087_
timestamp 0
transform 1 0 7544 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _3088_
timestamp 0
transform 1 0 8096 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _3089_
timestamp 0
transform 1 0 21804 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3090_
timestamp 0
transform 1 0 16652 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3091_
timestamp 0
transform 1 0 14168 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3092_
timestamp 0
transform 1 0 26956 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3093_
timestamp 0
transform 1 0 25668 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3094_
timestamp 0
transform 1 0 26128 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3095_
timestamp 0
transform 1 0 30544 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3096_
timestamp 0
transform 1 0 30544 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3097_
timestamp 0
transform 1 0 17664 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3098_
timestamp 0
transform 1 0 32108 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3099_
timestamp 0
transform 1 0 21988 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3100_
timestamp 0
transform 1 0 19688 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3101_
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3102_
timestamp 0
transform 1 0 18952 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3103_
timestamp 0
transform 1 0 16744 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3104_
timestamp 0
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3105_
timestamp 0
transform 1 0 24380 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3106_
timestamp 0
transform 1 0 17664 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3107_
timestamp 0
transform 1 0 16284 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3108_
timestamp 0
transform 1 0 29532 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3109_
timestamp 0
transform 1 0 27416 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3110_
timestamp 0
transform 1 0 29532 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3111_
timestamp 0
transform 1 0 30728 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3112_
timestamp 0
transform 1 0 29716 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3113_
timestamp 0
transform 1 0 25392 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3114_
timestamp 0
transform 1 0 30820 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3115_
timestamp 0
transform 1 0 27232 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3116_
timestamp 0
transform 1 0 26956 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3117_
timestamp 0
transform 1 0 28612 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3118_
timestamp 0
transform 1 0 29808 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3119_
timestamp 0
transform 1 0 14076 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3120_
timestamp 0
transform 1 0 24196 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3121_
timestamp 0
transform 1 0 6348 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3122_
timestamp 0
transform 1 0 1656 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3123_
timestamp 0
transform 1 0 6532 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3124_
timestamp 0
transform 1 0 6348 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3125_
timestamp 0
transform 1 0 2116 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3126_
timestamp 0
transform 1 0 1564 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3127_
timestamp 0
transform 1 0 1656 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3128_
timestamp 0
transform 1 0 1748 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3129_
timestamp 0
transform 1 0 6900 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3130_
timestamp 0
transform 1 0 5796 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3131_
timestamp 0
transform 1 0 7176 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3132_
timestamp 0
transform 1 0 2024 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3133_
timestamp 0
transform 1 0 3680 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3134_
timestamp 0
transform 1 0 6164 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3135_
timestamp 0
transform 1 0 9752 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3136_
timestamp 0
transform 1 0 8924 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3137_
timestamp 0
transform 1 0 5612 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3138_
timestamp 0
transform 1 0 1748 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3139_
timestamp 0
transform 1 0 6532 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3140_
timestamp 0
transform 1 0 6348 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3141_
timestamp 0
transform 1 0 2116 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3142_
timestamp 0
transform 1 0 1656 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3143_
timestamp 0
transform 1 0 1656 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3144_
timestamp 0
transform 1 0 1748 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3145_
timestamp 0
transform 1 0 6900 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3146_
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3147_
timestamp 0
transform 1 0 7176 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3148_
timestamp 0
transform 1 0 2300 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3149_
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3150_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3151_
timestamp 0
transform 1 0 9568 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3152_
timestamp 0
transform 1 0 9016 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3153_
timestamp 0
transform 1 0 7084 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3154_
timestamp 0
transform 1 0 3956 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3155_
timestamp 0
transform 1 0 8004 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3156_
timestamp 0
transform 1 0 7912 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3157_
timestamp 0
transform 1 0 3772 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3158_
timestamp 0
transform 1 0 2576 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3159_
timestamp 0
transform 1 0 3496 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3160_
timestamp 0
transform 1 0 3864 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3161_
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3162_
timestamp 0
transform 1 0 7912 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3163_
timestamp 0
transform 1 0 8924 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3164_
timestamp 0
transform 1 0 3404 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3165_
timestamp 0
transform 1 0 5336 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3166_
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3167_
timestamp 0
transform 1 0 9936 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3168_
timestamp 0
transform 1 0 9292 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3169_
timestamp 0
transform 1 0 9016 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3170_
timestamp 0
transform 1 0 3312 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3171_
timestamp 0
transform 1 0 9660 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3172_
timestamp 0
transform 1 0 9292 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3173_
timestamp 0
transform 1 0 3772 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3174_
timestamp 0
transform 1 0 3772 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3175_
timestamp 0
transform 1 0 4968 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3176_
timestamp 0
transform 1 0 4784 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3177_
timestamp 0
transform 1 0 9936 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3178_
timestamp 0
transform 1 0 9384 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3179_
timestamp 0
transform 1 0 10028 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3180_
timestamp 0
transform 1 0 4416 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3181_
timestamp 0
transform 1 0 6440 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3182_
timestamp 0
transform 1 0 7360 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3183_
timestamp 0
transform 1 0 10212 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3184_
timestamp 0
transform 1 0 11776 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3185_
timestamp 0
transform 1 0 19228 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3186_
timestamp 0
transform 1 0 15732 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3187_
timestamp 0
transform 1 0 14076 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3188_
timestamp 0
transform 1 0 22264 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3189_
timestamp 0
transform 1 0 21804 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3190_
timestamp 0
transform 1 0 21252 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3191_
timestamp 0
transform 1 0 12512 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3192_
timestamp 0
transform 1 0 13708 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3193_
timestamp 0
transform 1 0 12512 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3194_
timestamp 0
transform 1 0 12052 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3195_
timestamp 0
transform 1 0 12880 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3196_
timestamp 0
transform 1 0 12144 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3197_
timestamp 0
transform 1 0 14260 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3198_
timestamp 0
transform 1 0 12512 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3199_
timestamp 0
transform 1 0 12420 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3200_
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3201_
timestamp 0
transform 1 0 19044 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3202_
timestamp 0
transform 1 0 15088 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3203_
timestamp 0
transform 1 0 13524 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3204_
timestamp 0
transform 1 0 21804 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3205_
timestamp 0
transform 1 0 20792 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3206_
timestamp 0
transform 1 0 19780 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3207_
timestamp 0
transform 1 0 14444 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3208_
timestamp 0
transform 1 0 16008 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3209_
timestamp 0
transform 1 0 13064 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3210_
timestamp 0
transform 1 0 14444 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3211_
timestamp 0
transform 1 0 15640 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3212_
timestamp 0
transform 1 0 14812 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3213_
timestamp 0
transform 1 0 14720 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3214_
timestamp 0
transform 1 0 15732 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3215_
timestamp 0
transform 1 0 14904 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3216_
timestamp 0
transform 1 0 14904 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3217_
timestamp 0
transform 1 0 24472 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3218_
timestamp 0
transform 1 0 19228 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3219_
timestamp 0
transform 1 0 17020 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3220_
timestamp 0
transform 1 0 28888 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3221_
timestamp 0
transform 1 0 27876 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3222_
timestamp 0
transform 1 0 29532 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3223_
timestamp 0
transform 1 0 31832 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3224_
timestamp 0
transform 1 0 29900 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3225_
timestamp 0
transform 1 0 27232 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3226_
timestamp 0
transform 1 0 31832 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3227_
timestamp 0
transform 1 0 28060 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3228_
timestamp 0
transform 1 0 27416 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3229_
timestamp 0
transform 1 0 28888 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3230_
timestamp 0
transform 1 0 29624 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3231_
timestamp 0
transform 1 0 14260 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3232_
timestamp 0
transform 1 0 24656 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3233_
timestamp 0
transform 1 0 21804 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3234_
timestamp 0
transform 1 0 19320 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3235_
timestamp 0
transform 1 0 16652 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3236_
timestamp 0
transform 1 0 22816 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3237_
timestamp 0
transform 1 0 23644 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3238_
timestamp 0
transform 1 0 24380 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3239_
timestamp 0
transform 1 0 17112 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3240_
timestamp 0
transform 1 0 17756 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3241_
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3242_
timestamp 0
transform 1 0 16928 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3243_
timestamp 0
transform 1 0 17664 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3244_
timestamp 0
transform 1 0 16928 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3245_
timestamp 0
transform 1 0 16836 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3246_
timestamp 0
transform 1 0 19228 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3247_
timestamp 0
transform 1 0 16744 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3248_
timestamp 0
transform 1 0 16928 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3249_
timestamp 0
transform 1 0 33948 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3250_
timestamp 0
transform 1 0 36064 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3251_
timestamp 0
transform 1 0 30544 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _3252_
timestamp 0
transform 1 0 31924 0 1 46784
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _3253_
timestamp 0
transform 1 0 22816 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3254_
timestamp 0
transform 1 0 13708 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3255_
timestamp 0
transform 1 0 14076 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _3256_
timestamp 0
transform 1 0 1840 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _3257_
timestamp 0
transform 1 0 7544 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3258_
timestamp 0
transform 1 0 11224 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3259_
timestamp 0
transform 1 0 1748 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3260_
timestamp 0
transform 1 0 4508 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _3261_
timestamp 0
transform 1 0 2116 0 1 40256
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _3262_
timestamp 0
transform 1 0 38180 0 1 43520
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _3263_
timestamp 0
transform 1 0 1564 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _3264_
timestamp 0
transform 1 0 20240 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3265_
timestamp 0
transform 1 0 19228 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3266_
timestamp 0
transform 1 0 18768 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3267_
timestamp 0
transform 1 0 17388 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _3268_
timestamp 0
transform 1 0 18216 0 -1 46784
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _3269_
timestamp 0
transform 1 0 24748 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3270_
timestamp 0
transform 1 0 30176 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _3271_
timestamp 0
transform 1 0 26956 0 1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _3272_
timestamp 0
transform 1 0 26956 0 -1 46784
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _3273_
timestamp 0
transform 1 0 21712 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _3274_
timestamp 0
transform 1 0 22724 0 -1 43520
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _3275_
timestamp 0
transform 1 0 20240 0 1 43520
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _3276_
timestamp 0
transform 1 0 20148 0 -1 46784
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _3277_
timestamp 0
transform 1 0 23460 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3278_
timestamp 0
transform 1 0 24380 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _3278__182
timestamp 0
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _3279__181
timestamp 0
transform 1 0 27416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _3279_
timestamp 0
transform 1 0 27048 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3280_
timestamp 0
transform 1 0 4600 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _3280__180
timestamp 0
transform 1 0 4876 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _3281__179
timestamp 0
transform 1 0 38088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _3281_
timestamp 0
transform 1 0 37812 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _3282__178
timestamp 0
transform 1 0 17940 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _3282_
timestamp 0
transform 1 0 19228 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _3283__177
timestamp 0
transform 1 0 39468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _3283_
timestamp 0
transform 1 0 38456 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _3284_
timestamp 0
transform 1 0 39008 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _3284__176
timestamp 0
transform 1 0 39376 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _3285_
timestamp 0
transform 1 0 32108 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3286_
timestamp 0
transform 1 0 32568 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3287_
timestamp 0
transform 1 0 14168 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3288_
timestamp 0
transform 1 0 11132 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3289_
timestamp 0
transform 1 0 33672 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3290_
timestamp 0
transform 1 0 31740 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3291_
timestamp 0
transform 1 0 35236 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3292_
timestamp 0
transform 1 0 35420 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3293_
timestamp 0
transform 1 0 36800 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3294_
timestamp 0
transform 1 0 36892 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3295_
timestamp 0
transform 1 0 35788 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3296_
timestamp 0
transform 1 0 37260 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3297_
timestamp 0
transform 1 0 35696 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3298_
timestamp 0
transform 1 0 34776 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3299_
timestamp 0
transform 1 0 35236 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3300_
timestamp 0
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3301_
timestamp 0
transform 1 0 27508 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3302_
timestamp 0
transform 1 0 24380 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3303_
timestamp 0
transform 1 0 16652 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3304_
timestamp 0
transform 1 0 15364 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3305_
timestamp 0
transform 1 0 25392 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3306_
timestamp 0
transform 1 0 26956 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3307_
timestamp 0
transform 1 0 27048 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3308_
timestamp 0
transform 1 0 28980 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3309_
timestamp 0
transform 1 0 26956 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3310_
timestamp 0
transform 1 0 26956 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3311_
timestamp 0
transform 1 0 29532 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3312_
timestamp 0
transform 1 0 24380 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3313_
timestamp 0
transform 1 0 26036 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3314_
timestamp 0
transform 1 0 27784 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3315_
timestamp 0
transform 1 0 27232 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3316_
timestamp 0
transform 1 0 12512 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3317_
timestamp 0
transform 1 0 24656 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3318_
timestamp 0
transform 1 0 22632 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3319_
timestamp 0
transform 1 0 16376 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3320_
timestamp 0
transform 1 0 15088 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3321_
timestamp 0
transform 1 0 24472 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3322_
timestamp 0
transform 1 0 26312 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3323_
timestamp 0
transform 1 0 26956 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3324_
timestamp 0
transform 1 0 28520 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3325_
timestamp 0
transform 1 0 25392 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3326_
timestamp 0
transform 1 0 24472 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3327_
timestamp 0
transform 1 0 28796 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3328_
timestamp 0
transform 1 0 24288 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3329_
timestamp 0
transform 1 0 25116 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3330_
timestamp 0
transform 1 0 26956 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3331_
timestamp 0
transform 1 0 27140 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3332_
timestamp 0
transform 1 0 12420 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3333_
timestamp 0
transform 1 0 22540 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3334_
timestamp 0
transform 1 0 38088 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3335_
timestamp 0
transform 1 0 37536 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3336_
timestamp 0
transform 1 0 34684 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3337_
timestamp 0
transform 1 0 32936 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3338_
timestamp 0
transform 1 0 13524 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3339_
timestamp 0
transform 1 0 16928 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3340_
timestamp 0
transform 1 0 16652 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3341_
timestamp 0
transform 1 0 14996 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3342_
timestamp 0
transform 1 0 16652 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3343_
timestamp 0
transform 1 0 6532 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3344_
timestamp 0
transform 1 0 6256 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3345_
timestamp 0
transform 1 0 4968 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3346_
timestamp 0
transform 1 0 4784 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3347_
timestamp 0
transform 1 0 9936 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3348_
timestamp 0
transform 1 0 11316 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3349_
timestamp 0
transform 1 0 9200 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3350_
timestamp 0
transform 1 0 10672 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3351_
timestamp 0
transform 1 0 35972 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3352_
timestamp 0
transform 1 0 35696 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3353_
timestamp 0
transform 1 0 33028 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3354_
timestamp 0
transform 1 0 34684 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3355_
timestamp 0
transform 1 0 8924 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3356_
timestamp 0
transform 1 0 25852 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3357_
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3358_
timestamp 0
transform 1 0 33580 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3359_
timestamp 0
transform 1 0 38824 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3360_
timestamp 0
transform 1 0 13708 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3361_
timestamp 0
transform 1 0 7912 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3362_
timestamp 0
transform 1 0 9936 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3363_
timestamp 0
transform 1 0 34960 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3364_
timestamp 0
transform 1 0 36064 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3365_
timestamp 0
transform 1 0 33396 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3366_
timestamp 0
transform 1 0 32384 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3367_
timestamp 0
transform 1 0 37904 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3368_
timestamp 0
transform 1 0 37444 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3369_
timestamp 0
transform 1 0 38180 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _3370_
timestamp 0
transform 1 0 38272 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _3378_
timestamp 0
transform 1 0 3036 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _3379_
timestamp 0
transform 1 0 45448 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3380_
timestamp 0
transform 1 0 45632 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3381_
timestamp 0
transform 1 0 45632 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3382_
timestamp 0
transform 1 0 39376 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3383_
timestamp 0
transform 1 0 39468 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3384_
timestamp 0
transform 1 0 38180 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3385_
timestamp 0
transform 1 0 40112 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3386_
timestamp 0
transform 1 0 39836 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3387_
timestamp 0
transform 1 0 45540 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3388_
timestamp 0
transform 1 0 45264 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3389_
timestamp 0
transform 1 0 45632 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _3390_
timestamp 0
transform 1 0 45540 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _3391_
timestamp 0
transform 1 0 44896 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3392_
timestamp 0
transform 1 0 43240 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3393_
timestamp 0
transform 1 0 40940 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _3394_
timestamp 0
transform 1 0 39836 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 0
transform 1 0 9292 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 0
transform 1 0 17940 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 0
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 0
transform 1 0 1932 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 0
transform 1 0 25116 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 0
transform 1 0 22540 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 0
transform 1 0 36616 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 0
transform 1 0 1564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 0
transform 1 0 1932 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 0
transform 1 0 17756 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 0
transform 1 0 36432 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 0
transform 1 0 6808 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 0
transform 1 0 38088 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 0
transform 1 0 12328 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 0
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 0
transform 1 0 2300 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 0
transform 1 0 17848 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 0
transform 1 0 7176 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 0
transform 1 0 2668 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 0
transform 1 0 7544 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 0
transform 1 0 1932 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 0
transform 1 0 5704 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 0
transform 1 0 6072 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 0
transform 1 0 6440 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 0
transform 1 0 6808 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 0
transform 1 0 6808 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 0
transform 1 0 7176 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 0
transform 1 0 7544 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 0
transform 1 0 7912 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 0
transform 1 0 8280 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 0
transform 1 0 8648 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 0
transform 1 0 9292 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 0
transform 1 0 39008 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout84
timestamp 0
transform 1 0 39284 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout85
timestamp 0
transform 1 0 23736 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout86
timestamp 0
transform 1 0 37260 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout87
timestamp 0
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout88
timestamp 0
transform 1 0 38548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout89
timestamp 0
transform 1 0 39468 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout90
timestamp 0
transform 1 0 37444 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout91
timestamp 0
transform 1 0 35512 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp 0
transform 1 0 30820 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout93
timestamp 0
transform 1 0 25760 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout94
timestamp 0
transform 1 0 36984 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout95
timestamp 0
transform 1 0 2576 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout96
timestamp 0
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout97
timestamp 0
transform 1 0 9016 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout98
timestamp 0
transform 1 0 10120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout99
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout100
timestamp 0
transform 1 0 19228 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout101
timestamp 0
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout102
timestamp 0
transform 1 0 19964 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout103
timestamp 0
transform 1 0 20792 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout104
timestamp 0
transform 1 0 19872 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout105
timestamp 0
transform 1 0 18216 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout106
timestamp 0
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout107
timestamp 0
transform 1 0 8556 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout108
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout109
timestamp 0
transform 1 0 9016 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout110
timestamp 0
transform 1 0 9108 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout111
timestamp 0
transform 1 0 9936 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout112
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout113
timestamp 0
transform 1 0 18124 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout114
timestamp 0
transform 1 0 16652 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout115
timestamp 0
transform 1 0 17756 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout116
timestamp 0
transform 1 0 18032 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout117
timestamp 0
transform 1 0 18124 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout118
timestamp 0
transform 1 0 24288 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout119
timestamp 0
transform 1 0 28888 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout120
timestamp 0
transform 1 0 29716 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout121
timestamp 0
transform 1 0 28244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout122
timestamp 0
transform 1 0 29532 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout123
timestamp 0
transform 1 0 29072 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout124
timestamp 0
transform 1 0 32200 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout125
timestamp 0
transform 1 0 35880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout126
timestamp 0
transform 1 0 38548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout127
timestamp 0
transform 1 0 35512 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout128
timestamp 0
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout129
timestamp 0
transform 1 0 29532 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout130
timestamp 0
transform 1 0 28060 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout131
timestamp 0
transform 1 0 26956 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout132
timestamp 0
transform 1 0 34316 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout133
timestamp 0
transform 1 0 33488 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout134
timestamp 0
transform 1 0 36156 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout135
timestamp 0
transform 1 0 36248 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout136
timestamp 0
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout137
timestamp 0
transform 1 0 4600 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout138
timestamp 0
transform 1 0 10028 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout139
timestamp 0
transform 1 0 10396 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout140
timestamp 0
transform 1 0 2208 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout141
timestamp 0
transform 1 0 9384 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout142
timestamp 0
transform 1 0 9752 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout143
timestamp 0
transform 1 0 18124 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout144
timestamp 0
transform 1 0 18584 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout145
timestamp 0
transform 1 0 18860 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout146
timestamp 0
transform 1 0 18216 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout147
timestamp 0
transform 1 0 11500 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout148
timestamp 0
transform 1 0 10856 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout149
timestamp 0
transform 1 0 11040 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout150
timestamp 0
transform 1 0 14260 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout151
timestamp 0
transform 1 0 17112 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout152
timestamp 0
transform 1 0 18216 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout153
timestamp 0
transform 1 0 19228 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout154
timestamp 0
transform 1 0 18216 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout155
timestamp 0
transform 1 0 18216 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout156
timestamp 0
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout157
timestamp 0
transform 1 0 28520 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout158
timestamp 0
transform 1 0 24472 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout159
timestamp 0
transform 1 0 29532 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout160
timestamp 0
transform 1 0 29072 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout161
timestamp 0
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout162
timestamp 0
transform 1 0 36064 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout163
timestamp 0
transform 1 0 39100 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout164
timestamp 0
transform 1 0 24472 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout165
timestamp 0
transform 1 0 27876 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout166
timestamp 0
transform 1 0 24380 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout167
timestamp 0
transform 1 0 27324 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout168
timestamp 0
transform 1 0 28244 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout169
timestamp 0
transform 1 0 33672 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout170
timestamp 0
transform 1 0 38272 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout171
timestamp 0
transform 1 0 33028 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout172
timestamp 0
transform 1 0 38548 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout173
timestamp 0
transform 1 0 39468 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout174
timestamp 0
transform 1 0 38180 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout175
timestamp 0
transform 1 0 38824 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7
timestamp 0
transform 1 0 1748 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp 0
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42
timestamp 0
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 0
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62
timestamp 0
transform 1 0 6808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74
timestamp 0
transform 1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 0
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119
timestamp 0
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 0
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 0
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151
timestamp 0
transform 1 0 14996 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 0
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 0
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_179
timestamp 0
transform 1 0 17572 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_191
timestamp 0
transform 1 0 18676 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 0
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 0
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 0
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 0
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244
timestamp 0
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 0
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 0
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 0
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_281
timestamp 0
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_289
timestamp 0
transform 1 0 27692 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_294
timestamp 0
transform 1 0 28152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_302
timestamp 0
transform 1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309
timestamp 0
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_315
timestamp 0
transform 1 0 30084 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_322
timestamp 0
transform 1 0 30728 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 0
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 0
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_343
timestamp 0
transform 1 0 32660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_354
timestamp 0
transform 1 0 33672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 0
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 0
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_371
timestamp 0
transform 1 0 35236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 0
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 0
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 0
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_399
timestamp 0
transform 1 0 37812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_411
timestamp 0
transform 1 0 38916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_415
timestamp 0
transform 1 0 39284 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 0
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 0
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 0
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 0
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_459
timestamp 0
transform 1 0 43332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_471
timestamp 0
transform 1 0 44436 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_477
timestamp 0
transform 1 0 44988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_483
timestamp 0
transform 1 0 45540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 0
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_13
timestamp 0
transform 1 0 2300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_25
timestamp 0
transform 1 0 3404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_37
timestamp 0
transform 1 0 4508 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 0
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 0
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_185
timestamp 0
transform 1 0 18124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_197
timestamp 0
transform 1 0 19228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 0
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_241
timestamp 0
transform 1 0 23276 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_262
timestamp 0
transform 1 0 25208 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 0
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_281
timestamp 0
transform 1 0 26956 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_298
timestamp 0
transform 1 0 28520 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_318
timestamp 0
transform 1 0 30360 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_324
timestamp 0
transform 1 0 30912 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 0
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_369
timestamp 0
transform 1 0 35052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_381
timestamp 0
transform 1 0 36156 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_389
timestamp 0
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 0
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 0
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 0
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 0
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 0
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 0
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 0
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 0
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 0
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_485
timestamp 0
transform 1 0 45724 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 0
transform 1 0 14812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_160
timestamp 0
transform 1 0 15824 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_166
timestamp 0
transform 1 0 16376 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 0
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 0
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_201
timestamp 0
transform 1 0 19596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_242
timestamp 0
transform 1 0 23368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_269
timestamp 0
transform 1 0 25852 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 0
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 0
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 0
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_318
timestamp 0
transform 1 0 30360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_338
timestamp 0
transform 1 0 32200 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 0
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_374
timestamp 0
transform 1 0 35512 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_386
timestamp 0
transform 1 0 36616 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_398
timestamp 0
transform 1 0 37720 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_410
timestamp 0
transform 1 0 38824 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 0
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 0
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 0
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 0
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 0
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 0
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 0
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 0
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_489
timestamp 0
transform 1 0 46092 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_137
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_157
timestamp 0
transform 1 0 15548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 0
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_183
timestamp 0
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_187
timestamp 0
transform 1 0 18308 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_207
timestamp 0
transform 1 0 20148 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_215
timestamp 0
transform 1 0 20884 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 0
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_234
timestamp 0
transform 1 0 22632 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_249
timestamp 0
transform 1 0 24012 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_264
timestamp 0
transform 1 0 25392 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 0
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 0
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_281
timestamp 0
transform 1 0 26956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_288
timestamp 0
transform 1 0 27600 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_296
timestamp 0
transform 1 0 28336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_315
timestamp 0
transform 1 0 30084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_326
timestamp 0
transform 1 0 31096 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 0
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_337
timestamp 0
transform 1 0 32108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_343
timestamp 0
transform 1 0 32660 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_360
timestamp 0
transform 1 0 34224 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_372
timestamp 0
transform 1 0 35328 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_384
timestamp 0
transform 1 0 36432 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_393
timestamp 0
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_416
timestamp 0
transform 1 0 39376 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_428
timestamp 0
transform 1 0 40480 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_440
timestamp 0
transform 1 0 41584 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 0
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 0
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 0
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 0
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 0
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 0
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_103
timestamp 0
transform 1 0 10580 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_107
timestamp 0
transform 1 0 10948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_119
timestamp 0
transform 1 0 12052 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_131
timestamp 0
transform 1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_147
timestamp 0
transform 1 0 14628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_167
timestamp 0
transform 1 0 16468 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_178
timestamp 0
transform 1 0 17480 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 0
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 0
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_206
timestamp 0
transform 1 0 20056 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_218
timestamp 0
transform 1 0 21160 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_230
timestamp 0
transform 1 0 22264 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 0
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 0
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 0
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 0
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 0
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_318
timestamp 0
transform 1 0 30360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_330
timestamp 0
transform 1 0 31464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_358
timestamp 0
transform 1 0 34040 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp 0
transform 1 0 34684 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_378
timestamp 0
transform 1 0 35880 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_390
timestamp 0
transform 1 0 36984 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_405
timestamp 0
transform 1 0 38364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_417
timestamp 0
transform 1 0 39468 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 0
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 0
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 0
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 0
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 0
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 0
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 0
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_489
timestamp 0
transform 1 0 46092 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7
timestamp 0
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_19
timestamp 0
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_31
timestamp 0
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_43
timestamp 0
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_122
timestamp 0
transform 1 0 12328 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_142
timestamp 0
transform 1 0 14168 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_154
timestamp 0
transform 1 0 15272 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 0
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_185
timestamp 0
transform 1 0 18124 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 0
transform 1 0 18860 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_199
timestamp 0
transform 1 0 19412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_211
timestamp 0
transform 1 0 20516 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_219
timestamp 0
transform 1 0 21252 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_243
timestamp 0
transform 1 0 23460 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_255
timestamp 0
transform 1 0 24564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_281
timestamp 0
transform 1 0 26956 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_294
timestamp 0
transform 1 0 28152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_306
timestamp 0
transform 1 0 29256 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_319
timestamp 0
transform 1 0 30452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 0
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 0
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_358
timestamp 0
transform 1 0 34040 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_382
timestamp 0
transform 1 0 36248 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 0
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 0
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 0
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 0
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 0
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 0
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 0
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 0
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 0
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 0
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 0
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_121
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_150
timestamp 0
transform 1 0 14904 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_162
timestamp 0
transform 1 0 16008 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 0
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 0
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 0
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_207
timestamp 0
transform 1 0 20148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 0
transform 1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_244
timestamp 0
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_253
timestamp 0
transform 1 0 24380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_261
timestamp 0
transform 1 0 25116 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_276
timestamp 0
transform 1 0 26496 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_288
timestamp 0
transform 1 0 27600 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_300
timestamp 0
transform 1 0 28704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_309
timestamp 0
transform 1 0 29532 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_326
timestamp 0
transform 1 0 31096 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_338
timestamp 0
transform 1 0 32200 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_350
timestamp 0
transform 1 0 33304 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 0
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_365
timestamp 0
transform 1 0 34684 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_372
timestamp 0
transform 1 0 35328 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_384
timestamp 0
transform 1 0 36432 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_396
timestamp 0
transform 1 0 37536 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_408
timestamp 0
transform 1 0 38640 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 0
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 0
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 0
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 0
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 0
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 0
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 0
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_489
timestamp 0
transform 1 0 46092 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 0
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 0
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 0
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_190
timestamp 0
transform 1 0 18584 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 0
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 0
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_246
timestamp 0
transform 1 0 23736 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_250
timestamp 0
transform 1 0 24104 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 0
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 0
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_293
timestamp 0
transform 1 0 28060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_301
timestamp 0
transform 1 0 28796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_331
timestamp 0
transform 1 0 31556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 0
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 0
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 0
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 0
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 0
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 0
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 0
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 0
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 0
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 0
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 0
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 0
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 0
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 0
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 0
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 0
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 0
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_104
timestamp 0
transform 1 0 10672 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_116
timestamp 0
transform 1 0 11776 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_128
timestamp 0
transform 1 0 12880 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_145
timestamp 0
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_167
timestamp 0
transform 1 0 16468 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_175
timestamp 0
transform 1 0 17204 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_185
timestamp 0
transform 1 0 18124 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_213
timestamp 0
transform 1 0 20700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_225
timestamp 0
transform 1 0 21804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_237
timestamp 0
transform 1 0 22908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 0
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp 0
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_272
timestamp 0
transform 1 0 26128 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_280
timestamp 0
transform 1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_299
timestamp 0
transform 1 0 28612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 0
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 0
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_324
timestamp 0
transform 1 0 30912 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_345
timestamp 0
transform 1 0 32844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_353
timestamp 0
transform 1 0 33580 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_358
timestamp 0
transform 1 0 34040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 0
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 0
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 0
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 0
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 0
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 0
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 0
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 0
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 0
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 0
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 0
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 0
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 0
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 0
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_489
timestamp 0
transform 1 0 46092 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 0
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 0
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 0
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 0
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 0
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_85
timestamp 0
transform 1 0 8924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_122
timestamp 0
transform 1 0 12328 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_139
timestamp 0
transform 1 0 13892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_151
timestamp 0
transform 1 0 14996 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_159
timestamp 0
transform 1 0 15732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 0
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_186
timestamp 0
transform 1 0 18216 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_192
timestamp 0
transform 1 0 18768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 0
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_236
timestamp 0
transform 1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_248
timestamp 0
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_262
timestamp 0
transform 1 0 25208 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_274
timestamp 0
transform 1 0 26312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_309
timestamp 0
transform 1 0 29532 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_320
timestamp 0
transform 1 0 30544 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_332
timestamp 0
transform 1 0 31648 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp 0
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 0
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 0
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 0
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 0
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 0
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 0
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 0
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 0
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 0
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 0
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 0
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_94
timestamp 0
transform 1 0 9752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_98
timestamp 0
transform 1 0 10120 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_147
timestamp 0
transform 1 0 14628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_152
timestamp 0
transform 1 0 15088 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 0
transform 1 0 15640 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_218
timestamp 0
transform 1 0 21160 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_230
timestamp 0
transform 1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp 0
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_253
timestamp 0
transform 1 0 24380 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_268
timestamp 0
transform 1 0 25760 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_280
timestamp 0
transform 1 0 26864 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_286
timestamp 0
transform 1 0 27416 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_296
timestamp 0
transform 1 0 28336 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_330
timestamp 0
transform 1 0 31464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_365
timestamp 0
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_387
timestamp 0
transform 1 0 36708 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_399
timestamp 0
transform 1 0 37812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_410
timestamp 0
transform 1 0 38824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp 0
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 0
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 0
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 0
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 0
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 0
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 0
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 0
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_489
timestamp 0
transform 1 0 46092 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_84
timestamp 0
transform 1 0 8832 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_96
timestamp 0
transform 1 0 9936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_144
timestamp 0
transform 1 0 14352 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 0
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_173
timestamp 0
transform 1 0 17020 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 0
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_231
timestamp 0
transform 1 0 22356 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_240
timestamp 0
transform 1 0 23184 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_252
timestamp 0
transform 1 0 24288 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_272
timestamp 0
transform 1 0 26128 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 0
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 0
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_305
timestamp 0
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 0
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 0
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 0
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_342
timestamp 0
transform 1 0 32568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_367
timestamp 0
transform 1 0 34868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_375
timestamp 0
transform 1 0 35604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_382
timestamp 0
transform 1 0 36248 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 0
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 0
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_404
timestamp 0
transform 1 0 38272 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_423
timestamp 0
transform 1 0 40020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_435
timestamp 0
transform 1 0 41124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 0
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 0
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 0
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 0
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_485
timestamp 0
transform 1 0 45724 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_112
timestamp 0
transform 1 0 11408 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_124
timestamp 0
transform 1 0 12512 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_130
timestamp 0
transform 1 0 13064 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_171
timestamp 0
transform 1 0 16836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_183
timestamp 0
transform 1 0 17940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 0
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_209
timestamp 0
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_217
timestamp 0
transform 1 0 21068 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_238
timestamp 0
transform 1 0 23000 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_246
timestamp 0
transform 1 0 23736 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_283
timestamp 0
transform 1 0 27140 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_293
timestamp 0
transform 1 0 28060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_305
timestamp 0
transform 1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_309
timestamp 0
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_317
timestamp 0
transform 1 0 30268 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_327
timestamp 0
transform 1 0 31188 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_335
timestamp 0
transform 1 0 31924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_353
timestamp 0
transform 1 0 33580 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_361
timestamp 0
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 0
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_377
timestamp 0
transform 1 0 35788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_389
timestamp 0
transform 1 0 36892 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_411
timestamp 0
transform 1 0 38916 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 0
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 0
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_445
timestamp 0
transform 1 0 42044 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_451
timestamp 0
transform 1 0 42596 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_456
timestamp 0
transform 1 0 43056 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_468
timestamp 0
transform 1 0 44160 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 0
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_489
timestamp 0
transform 1 0 46092 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 0
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 0
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_73
timestamp 0
transform 1 0 7820 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_95
timestamp 0
transform 1 0 9844 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_100
timestamp 0
transform 1 0 10304 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 0
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 0
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 0
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 0
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 0
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_209
timestamp 0
transform 1 0 20332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_213
timestamp 0
transform 1 0 20700 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 0
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 0
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 0
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_270
timestamp 0
transform 1 0 25944 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_276
timestamp 0
transform 1 0 26496 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_306
timestamp 0
transform 1 0 29256 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_318
timestamp 0
transform 1 0 30360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_331
timestamp 0
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 0
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_337
timestamp 0
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_348
timestamp 0
transform 1 0 33120 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_360
timestamp 0
transform 1 0 34224 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_372
timestamp 0
transform 1 0 35328 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 0
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_393
timestamp 0
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_401
timestamp 0
transform 1 0 37996 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_409
timestamp 0
transform 1 0 38732 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_421
timestamp 0
transform 1 0 39836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_431
timestamp 0
transform 1 0 40756 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_463
timestamp 0
transform 1 0 43700 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_475
timestamp 0
transform 1 0 44804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_487
timestamp 0
transform 1 0 45908 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_495
timestamp 0
transform 1 0 46644 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_9
timestamp 0
transform 1 0 1932 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_13
timestamp 0
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 0
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_49
timestamp 0
transform 1 0 5612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 0
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_131
timestamp 0
transform 1 0 13156 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_157
timestamp 0
transform 1 0 15548 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_169
timestamp 0
transform 1 0 16652 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_188
timestamp 0
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_197
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_205
timestamp 0
transform 1 0 19964 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_220
timestamp 0
transform 1 0 21344 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_233
timestamp 0
transform 1 0 22540 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_241
timestamp 0
transform 1 0 23276 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 0
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 0
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 0
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_277
timestamp 0
transform 1 0 26588 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_285
timestamp 0
transform 1 0 27324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 0
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_339
timestamp 0
transform 1 0 32292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_351
timestamp 0
transform 1 0 33396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 0
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_365
timestamp 0
transform 1 0 34684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_369
timestamp 0
transform 1 0 35052 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_394
timestamp 0
transform 1 0 37352 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_406
timestamp 0
transform 1 0 38456 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_414
timestamp 0
transform 1 0 39192 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_439
timestamp 0
transform 1 0 41492 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_458
timestamp 0
transform 1 0 43240 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_470
timestamp 0
transform 1 0 44344 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 0
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_489
timestamp 0
transform 1 0 46092 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 0
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 0
transform 1 0 6624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_70
timestamp 0
transform 1 0 7544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 0
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_134
timestamp 0
transform 1 0 13432 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 0
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_203
timestamp 0
transform 1 0 19780 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 0
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 0
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 0
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_233
timestamp 0
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_239
timestamp 0
transform 1 0 23092 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_251
timestamp 0
transform 1 0 24196 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_263
timestamp 0
transform 1 0 25300 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 0
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 0
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 0
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 0
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_320
timestamp 0
transform 1 0 30544 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_326
timestamp 0
transform 1 0 31096 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_330
timestamp 0
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 0
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_365
timestamp 0
transform 1 0 34684 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_373
timestamp 0
transform 1 0 35420 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 0
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_393
timestamp 0
transform 1 0 37260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_399
timestamp 0
transform 1 0 37812 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_414
timestamp 0
transform 1 0 39192 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_422
timestamp 0
transform 1 0 39928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_431
timestamp 0
transform 1 0 40756 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_438
timestamp 0
transform 1 0 41400 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_446
timestamp 0
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_449
timestamp 0
transform 1 0 42412 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_465
timestamp 0
transform 1 0 43884 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_477
timestamp 0
transform 1 0 44988 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_489
timestamp 0
transform 1 0 46092 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_45
timestamp 0
transform 1 0 5244 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_62
timestamp 0
transform 1 0 6808 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_74
timestamp 0
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 0
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp 0
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 0
transform 1 0 9660 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_110
timestamp 0
transform 1 0 11224 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_122
timestamp 0
transform 1 0 12328 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 0
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 0
transform 1 0 14812 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_177
timestamp 0
transform 1 0 17388 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 0
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 0
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 0
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 0
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_221
timestamp 0
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_229
timestamp 0
transform 1 0 22172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 0
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 0
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_257
timestamp 0
transform 1 0 24748 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_283
timestamp 0
transform 1 0 27140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_295
timestamp 0
transform 1 0 28244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 0
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_315
timestamp 0
transform 1 0 30084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_339
timestamp 0
transform 1 0 32292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 0
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_365
timestamp 0
transform 1 0 34684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_373
timestamp 0
transform 1 0 35420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_387
timestamp 0
transform 1 0 36708 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_395
timestamp 0
transform 1 0 37444 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_406
timestamp 0
transform 1 0 38456 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 0
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 0
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_445
timestamp 0
transform 1 0 42044 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_449
timestamp 0
transform 1 0 42412 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_470
timestamp 0
transform 1 0 44344 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 0
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_489
timestamp 0
transform 1 0 46092 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_27
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_36
timestamp 0
transform 1 0 4416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_49
timestamp 0
transform 1 0 5612 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 0
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_66
timestamp 0
transform 1 0 7176 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_78
timestamp 0
transform 1 0 8280 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 0
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 0
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 0
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 0
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 0
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 0
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 0
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 0
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_230
timestamp 0
transform 1 0 22264 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_247
timestamp 0
transform 1 0 23828 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_259
timestamp 0
transform 1 0 24932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_271
timestamp 0
transform 1 0 26036 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_297
timestamp 0
transform 1 0 28428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_312
timestamp 0
transform 1 0 29808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_320
timestamp 0
transform 1 0 30544 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_326
timestamp 0
transform 1 0 31096 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_343
timestamp 0
transform 1 0 32660 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_364
timestamp 0
transform 1 0 34592 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_376
timestamp 0
transform 1 0 35696 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_388
timestamp 0
transform 1 0 36800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_393
timestamp 0
transform 1 0 37260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_405
timestamp 0
transform 1 0 38364 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_418
timestamp 0
transform 1 0 39560 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_430
timestamp 0
transform 1 0 40664 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_438
timestamp 0
transform 1 0 41400 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_463
timestamp 0
transform 1 0 43700 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_472
timestamp 0
transform 1 0 44528 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_484
timestamp 0
transform 1 0 45632 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_496
timestamp 0
transform 1 0 46736 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_45
timestamp 0
transform 1 0 5244 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 0
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_102
timestamp 0
transform 1 0 10488 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 0
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 0
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_155
timestamp 0
transform 1 0 15364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_167
timestamp 0
transform 1 0 16468 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 0
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_216
timestamp 0
transform 1 0 20976 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_222
timestamp 0
transform 1 0 21528 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 0
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_275
timestamp 0
transform 1 0 26404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_281
timestamp 0
transform 1 0 26956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_291
timestamp 0
transform 1 0 27876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 0
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 0
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_309
timestamp 0
transform 1 0 29532 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_316
timestamp 0
transform 1 0 30176 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_328
timestamp 0
transform 1 0 31280 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_340
timestamp 0
transform 1 0 32384 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 0
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 0
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 0
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 0
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_377
timestamp 0
transform 1 0 35788 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_386
timestamp 0
transform 1 0 36616 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_398
timestamp 0
transform 1 0 37720 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_404
timestamp 0
transform 1 0 38272 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 0
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_426
timestamp 0
transform 1 0 40296 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_434
timestamp 0
transform 1 0 41032 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 0
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 0
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_489
timestamp 0
transform 1 0 46092 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_7
timestamp 0
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_19
timestamp 0
transform 1 0 2852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_27
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 0
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_78
timestamp 0
transform 1 0 8280 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_84
timestamp 0
transform 1 0 8832 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 0
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_210
timestamp 0
transform 1 0 20424 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 0
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 0
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 0
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_237
timestamp 0
transform 1 0 22908 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_262
timestamp 0
transform 1 0 25208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 0
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_281
timestamp 0
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_292
timestamp 0
transform 1 0 27968 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_300
timestamp 0
transform 1 0 28704 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 0
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 0
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 0
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 0
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_370
timestamp 0
transform 1 0 35144 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_378
timestamp 0
transform 1 0 35880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_383
timestamp 0
transform 1 0 36340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 0
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 0
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_405
timestamp 0
transform 1 0 38364 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_413
timestamp 0
transform 1 0 39100 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_421
timestamp 0
transform 1 0 39836 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_432
timestamp 0
transform 1 0 40848 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_444
timestamp 0
transform 1 0 41952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_449
timestamp 0
transform 1 0 42412 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_459
timestamp 0
transform 1 0 43332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_471
timestamp 0
transform 1 0 44436 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_475
timestamp 0
transform 1 0 44804 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_484
timestamp 0
transform 1 0 45632 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_496
timestamp 0
transform 1 0 46736 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_33
timestamp 0
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_37
timestamp 0
transform 1 0 4508 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_49
timestamp 0
transform 1 0 5612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_57
timestamp 0
transform 1 0 6348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_74
timestamp 0
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 0
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_108
timestamp 0
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_112
timestamp 0
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 0
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_164
timestamp 0
transform 1 0 16192 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_170
timestamp 0
transform 1 0 16744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 0
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 0
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 0
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_205
timestamp 0
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_211
timestamp 0
transform 1 0 20516 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_223
timestamp 0
transform 1 0 21620 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_262
timestamp 0
transform 1 0 25208 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_274
timestamp 0
transform 1 0 26312 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_302
timestamp 0
transform 1 0 28888 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 0
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_309
timestamp 0
transform 1 0 29532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_350
timestamp 0
transform 1 0 33304 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_390
timestamp 0
transform 1 0 36984 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_397
timestamp 0
transform 1 0 37628 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_409
timestamp 0
transform 1 0 38732 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_417
timestamp 0
transform 1 0 39468 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 0
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 0
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_445
timestamp 0
transform 1 0 42044 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_453
timestamp 0
transform 1 0 42780 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_459
timestamp 0
transform 1 0 43332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_471
timestamp 0
transform 1 0 44436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 0
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_477
timestamp 0
transform 1 0 44988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_483
timestamp 0
transform 1 0 45540 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_491
timestamp 0
transform 1 0 46276 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 0
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 0
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 0
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 0
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_66
timestamp 0
transform 1 0 7176 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_78
timestamp 0
transform 1 0 8280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_86
timestamp 0
transform 1 0 9016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_92
timestamp 0
transform 1 0 9568 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 0
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 0
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 0
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_128
timestamp 0
transform 1 0 12880 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_135
timestamp 0
transform 1 0 13524 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_147
timestamp 0
transform 1 0 14628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_151
timestamp 0
transform 1 0 14996 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_155
timestamp 0
transform 1 0 15364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 0
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_193
timestamp 0
transform 1 0 18860 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_201
timestamp 0
transform 1 0 19596 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 0
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_225
timestamp 0
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_231
timestamp 0
transform 1 0 22356 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_236
timestamp 0
transform 1 0 22816 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_246
timestamp 0
transform 1 0 23736 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_258
timestamp 0
transform 1 0 24840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 0
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_332
timestamp 0
transform 1 0 31648 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_346
timestamp 0
transform 1 0 32936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_350
timestamp 0
transform 1 0 33304 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_372
timestamp 0
transform 1 0 35328 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_402
timestamp 0
transform 1 0 38088 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_414
timestamp 0
transform 1 0 39192 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_422
timestamp 0
transform 1 0 39928 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_427
timestamp 0
transform 1 0 40388 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 0
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 0
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_449
timestamp 0
transform 1 0 42412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_457
timestamp 0
transform 1 0 43148 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_469
timestamp 0
transform 1 0 44252 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_483
timestamp 0
transform 1 0 45540 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_495
timestamp 0
transform 1 0 46644 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_7
timestamp 0
transform 1 0 1748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 0
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_33
timestamp 0
transform 1 0 4140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_45
timestamp 0
transform 1 0 5244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_57
timestamp 0
transform 1 0 6348 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_68
timestamp 0
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 0
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_117
timestamp 0
transform 1 0 11868 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_124
timestamp 0
transform 1 0 12512 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 0
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_153
timestamp 0
transform 1 0 15180 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_159
timestamp 0
transform 1 0 15732 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_166
timestamp 0
transform 1 0 16376 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_178
timestamp 0
transform 1 0 17480 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_197
timestamp 0
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_203
timestamp 0
transform 1 0 19780 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_218
timestamp 0
transform 1 0 21160 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_233
timestamp 0
transform 1 0 22540 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_239
timestamp 0
transform 1 0 23092 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 0
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_262
timestamp 0
transform 1 0 25208 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_267
timestamp 0
transform 1 0 25668 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 0
transform 1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_319
timestamp 0
transform 1 0 30452 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_339
timestamp 0
transform 1 0 32292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_351
timestamp 0
transform 1 0 33396 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 0
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 0
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_393
timestamp 0
transform 1 0 37260 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_406
timestamp 0
transform 1 0 38456 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 0
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_447
timestamp 0
transform 1 0 42228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_455
timestamp 0
transform 1 0 42964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_460
timestamp 0
transform 1 0 43424 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_467
timestamp 0
transform 1 0 44068 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 0
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 0
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_489
timestamp 0
transform 1 0 46092 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 0
transform 1 0 3220 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_41
timestamp 0
transform 1 0 4876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 0
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_73
timestamp 0
transform 1 0 7820 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_90
timestamp 0
transform 1 0 9384 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_103
timestamp 0
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_121
timestamp 0
transform 1 0 12236 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_136
timestamp 0
transform 1 0 13616 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_148
timestamp 0
transform 1 0 14720 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 0
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_188
timestamp 0
transform 1 0 18400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 0
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 0
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_233
timestamp 0
transform 1 0 22540 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_240
timestamp 0
transform 1 0 23184 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_252
timestamp 0
transform 1 0 24288 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_264
timestamp 0
transform 1 0 25392 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_272
timestamp 0
transform 1 0 26128 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 0
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_290
timestamp 0
transform 1 0 27784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_302
timestamp 0
transform 1 0 28888 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_315
timestamp 0
transform 1 0 30084 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_327
timestamp 0
transform 1 0 31188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 0
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 0
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_349
timestamp 0
transform 1 0 33212 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_359
timestamp 0
transform 1 0 34132 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_371
timestamp 0
transform 1 0 35236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_384
timestamp 0
transform 1 0 36432 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 0
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_405
timestamp 0
transform 1 0 38364 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_422
timestamp 0
transform 1 0 39928 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_434
timestamp 0
transform 1 0 41032 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_438
timestamp 0
transform 1 0 41400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 0
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_449
timestamp 0
transform 1 0 42412 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_453
timestamp 0
transform 1 0 42780 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_467
timestamp 0
transform 1 0 44068 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 0
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 0
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_42
timestamp 0
transform 1 0 4968 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_67
timestamp 0
transform 1 0 7268 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_71
timestamp 0
transform 1 0 7636 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_106
timestamp 0
transform 1 0 10856 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_118
timestamp 0
transform 1 0 11960 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 0
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 0
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_165
timestamp 0
transform 1 0 16284 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_187
timestamp 0
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 0
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 0
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_201
timestamp 0
transform 1 0 19596 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_229
timestamp 0
transform 1 0 22172 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_241
timestamp 0
transform 1 0 23276 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 0
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 0
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_265
timestamp 0
transform 1 0 25484 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_287
timestamp 0
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_299
timestamp 0
transform 1 0 28612 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_325
timestamp 0
transform 1 0 31004 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_343
timestamp 0
transform 1 0 32660 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_355
timestamp 0
transform 1 0 33764 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 0
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_374
timestamp 0
transform 1 0 35512 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_380
timestamp 0
transform 1 0 36064 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_385
timestamp 0
transform 1 0 36524 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 0
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_413
timestamp 0
transform 1 0 39100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 0
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 0
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 0
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 0
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 0
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 0
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 0
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_477
timestamp 0
transform 1 0 44988 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_493
timestamp 0
transform 1 0 46460 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 0
transform 1 0 2116 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_38
timestamp 0
transform 1 0 4600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 0
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 0
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_144
timestamp 0
transform 1 0 14352 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_161
timestamp 0
transform 1 0 15916 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 0
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_208
timestamp 0
transform 1 0 20240 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_216
timestamp 0
transform 1 0 20976 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_249
timestamp 0
transform 1 0 24012 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_263
timestamp 0
transform 1 0 25300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_275
timestamp 0
transform 1 0 26404 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_287
timestamp 0
transform 1 0 27508 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_299
timestamp 0
transform 1 0 28612 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_307
timestamp 0
transform 1 0 29348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_319
timestamp 0
transform 1 0 30452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_325
timestamp 0
transform 1 0 31004 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 0
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 0
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_353
timestamp 0
transform 1 0 33580 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_357
timestamp 0
transform 1 0 33948 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_377
timestamp 0
transform 1 0 35788 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 0
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 0
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_417
timestamp 0
transform 1 0 39468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_443
timestamp 0
transform 1 0 41860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 0
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_449
timestamp 0
transform 1 0 42412 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_459
timestamp 0
transform 1 0 43332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_471
timestamp 0
transform 1 0 44436 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_492
timestamp 0
transform 1 0 46368 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 0
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 0
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_38
timestamp 0
transform 1 0 4600 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_42
timestamp 0
transform 1 0 4968 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_52
timestamp 0
transform 1 0 5888 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_64
timestamp 0
transform 1 0 6992 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_76
timestamp 0
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_89
timestamp 0
transform 1 0 9292 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_106
timestamp 0
transform 1 0 10856 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_134
timestamp 0
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_159
timestamp 0
transform 1 0 15732 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_171
timestamp 0
transform 1 0 16836 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 0
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_216
timestamp 0
transform 1 0 20976 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_228
timestamp 0
transform 1 0 22080 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 0
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 0
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 0
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_261
timestamp 0
transform 1 0 25116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_273
timestamp 0
transform 1 0 26220 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_284
timestamp 0
transform 1 0 27232 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_296
timestamp 0
transform 1 0 28336 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 0
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_321
timestamp 0
transform 1 0 30636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_338
timestamp 0
transform 1 0 32200 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_342
timestamp 0
transform 1 0 32568 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 0
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_381
timestamp 0
transform 1 0 36156 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_387
timestamp 0
transform 1 0 36708 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 0
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 0
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_440
timestamp 0
transform 1 0 41584 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_467
timestamp 0
transform 1 0 44068 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 0
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_482
timestamp 0
transform 1 0 45448 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_492
timestamp 0
transform 1 0 46368 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_496
timestamp 0
transform 1 0 46736 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_6
timestamp 0
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_26
timestamp 0
transform 1 0 3496 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_32
timestamp 0
transform 1 0 4048 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 0
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_63
timestamp 0
transform 1 0 6900 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_78
timestamp 0
transform 1 0 8280 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_90
timestamp 0
transform 1 0 9384 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_102
timestamp 0
transform 1 0 10488 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 0
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_137
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 0
transform 1 0 14076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_151
timestamp 0
transform 1 0 14996 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 0
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 0
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_205
timestamp 0
transform 1 0 19964 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_233
timestamp 0
transform 1 0 22540 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_250
timestamp 0
transform 1 0 24104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 0
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_297
timestamp 0
transform 1 0 28428 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_314
timestamp 0
transform 1 0 29992 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_326
timestamp 0
transform 1 0 31096 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_337
timestamp 0
transform 1 0 32108 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_345
timestamp 0
transform 1 0 32844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_356
timestamp 0
transform 1 0 33856 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_360
timestamp 0
transform 1 0 34224 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_374
timestamp 0
transform 1 0 35512 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_386
timestamp 0
transform 1 0 36616 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_412
timestamp 0
transform 1 0 39008 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_420
timestamp 0
transform 1 0 39744 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_426
timestamp 0
transform 1 0 40296 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_435
timestamp 0
transform 1 0 41124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 0
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_454
timestamp 0
transform 1 0 42872 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_466
timestamp 0
transform 1 0 43976 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_484
timestamp 0
transform 1 0 45632 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_496
timestamp 0
transform 1 0 46736 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp 0
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_58
timestamp 0
transform 1 0 6440 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_68
timestamp 0
transform 1 0 7360 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_79
timestamp 0
transform 1 0 8372 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_94
timestamp 0
transform 1 0 9752 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_121
timestamp 0
transform 1 0 12236 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_129
timestamp 0
transform 1 0 12972 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_151
timestamp 0
transform 1 0 14996 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 0
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 0
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 0
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 0
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_213
timestamp 0
transform 1 0 20700 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_225
timestamp 0
transform 1 0 21804 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_237
timestamp 0
transform 1 0 22908 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_241
timestamp 0
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 0
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 0
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_265
timestamp 0
transform 1 0 25484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_273
timestamp 0
transform 1 0 26220 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_278
timestamp 0
transform 1 0 26680 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_290
timestamp 0
transform 1 0 27784 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_298
timestamp 0
transform 1 0 28520 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 0
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 0
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 0
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 0
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_374
timestamp 0
transform 1 0 35512 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_386
timestamp 0
transform 1 0 36616 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_398
timestamp 0
transform 1 0 37720 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 0
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 0
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 0
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_457
timestamp 0
transform 1 0 43148 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_473
timestamp 0
transform 1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_477
timestamp 0
transform 1 0 44988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_22
timestamp 0
transform 1 0 3128 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_34
timestamp 0
transform 1 0 4232 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 0
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_79
timestamp 0
transform 1 0 8372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 0
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_122
timestamp 0
transform 1 0 12328 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 0
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_189
timestamp 0
transform 1 0 18492 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_194
timestamp 0
transform 1 0 18952 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_202
timestamp 0
transform 1 0 19688 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_215
timestamp 0
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 0
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_229
timestamp 0
transform 1 0 22172 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_237
timestamp 0
transform 1 0 22908 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_259
timestamp 0
transform 1 0 24932 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_271
timestamp 0
transform 1 0 26036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 0
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 0
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 0
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_305
timestamp 0
transform 1 0 29164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_327
timestamp 0
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 0
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_346
timestamp 0
transform 1 0 32936 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_373
timestamp 0
transform 1 0 35420 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_385
timestamp 0
transform 1 0 36524 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_389
timestamp 0
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_402
timestamp 0
transform 1 0 38088 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_414
timestamp 0
transform 1 0 39192 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_426
timestamp 0
transform 1 0 40296 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 0
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_455
timestamp 0
transform 1 0 42964 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_463
timestamp 0
transform 1 0 43700 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_468
timestamp 0
transform 1 0 44160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_474
timestamp 0
transform 1 0 44712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_482
timestamp 0
transform 1 0 45448 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_492
timestamp 0
transform 1 0 46368 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_496
timestamp 0
transform 1 0 46736 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 0
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 0
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 0
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_53
timestamp 0
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_61
timestamp 0
transform 1 0 6716 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 0
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 0
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_101
timestamp 0
transform 1 0 10396 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_123
timestamp 0
transform 1 0 12420 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_144
timestamp 0
transform 1 0 14352 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_148
timestamp 0
transform 1 0 14720 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_170
timestamp 0
transform 1 0 16744 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_174
timestamp 0
transform 1 0 17112 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_179
timestamp 0
transform 1 0 17572 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_212
timestamp 0
transform 1 0 20608 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 0
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_262
timestamp 0
transform 1 0 25208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_295
timestamp 0
transform 1 0 28244 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_303
timestamp 0
transform 1 0 28980 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_318
timestamp 0
transform 1 0 30360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_330
timestamp 0
transform 1 0 31464 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_350
timestamp 0
transform 1 0 33304 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_365
timestamp 0
transform 1 0 34684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 0
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 0
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 0
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_429
timestamp 0
transform 1 0 40572 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_442
timestamp 0
transform 1 0 41768 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_454
timestamp 0
transform 1 0 42872 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_477
timestamp 0
transform 1 0 44988 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_485
timestamp 0
transform 1 0 45724 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_490
timestamp 0
transform 1 0 46184 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_496
timestamp 0
transform 1 0 46736 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_7
timestamp 0
transform 1 0 1748 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_15
timestamp 0
transform 1 0 2484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_25
timestamp 0
transform 1 0 3404 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_42
timestamp 0
transform 1 0 4968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 0
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 0
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 0
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 0
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_93
timestamp 0
transform 1 0 9660 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_99
timestamp 0
transform 1 0 10212 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 0
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_117
timestamp 0
transform 1 0 11868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_125
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_131
timestamp 0
transform 1 0 13156 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_143
timestamp 0
transform 1 0 14260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 0
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 0
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_188
timestamp 0
transform 1 0 18400 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_200
timestamp 0
transform 1 0 19504 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_206
timestamp 0
transform 1 0 20056 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 0
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 0
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_229
timestamp 0
transform 1 0 22172 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_260
timestamp 0
transform 1 0 25024 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 0
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 0
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_349
timestamp 0
transform 1 0 33212 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_373
timestamp 0
transform 1 0 35420 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_379
timestamp 0
transform 1 0 35972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 0
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_393
timestamp 0
transform 1 0 37260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_419
timestamp 0
transform 1 0 39652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_449
timestamp 0
transform 1 0 42412 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_455
timestamp 0
transform 1 0 42964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_462
timestamp 0
transform 1 0 43608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_466
timestamp 0
transform 1 0 43976 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_474
timestamp 0
transform 1 0 44712 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_486
timestamp 0
transform 1 0 45816 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_494
timestamp 0
transform 1 0 46552 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_22
timestamp 0
transform 1 0 3128 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_34
timestamp 0
transform 1 0 4232 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_67
timestamp 0
transform 1 0 7268 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_79
timestamp 0
transform 1 0 8372 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 0
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 0
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_121
timestamp 0
transform 1 0 12236 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_129
timestamp 0
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 0
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_153
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_158
timestamp 0
transform 1 0 15640 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 0
transform 1 0 16744 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_174
timestamp 0
transform 1 0 17112 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_188
timestamp 0
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 0
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_203
timestamp 0
transform 1 0 19780 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_219
timestamp 0
transform 1 0 21252 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_231
timestamp 0
transform 1 0 22356 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_235
timestamp 0
transform 1 0 22724 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_262
timestamp 0
transform 1 0 25208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_296
timestamp 0
transform 1 0 28336 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_325
timestamp 0
transform 1 0 31004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_338
timestamp 0
transform 1 0 32200 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_346
timestamp 0
transform 1 0 32936 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 0
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 0
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_389
timestamp 0
transform 1 0 36892 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_395
timestamp 0
transform 1 0 37444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_404
timestamp 0
transform 1 0 38272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_411
timestamp 0
transform 1 0 38916 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 0
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 0
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_433
timestamp 0
transform 1 0 40940 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_442
timestamp 0
transform 1 0 41768 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_450
timestamp 0
transform 1 0 42504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_461
timestamp 0
transform 1 0 43516 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_467
timestamp 0
transform 1 0 44068 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_477
timestamp 0
transform 1 0 44988 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_491
timestamp 0
transform 1 0 46276 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_22
timestamp 0
transform 1 0 3128 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_67
timestamp 0
transform 1 0 7268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_91
timestamp 0
transform 1 0 9476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_98
timestamp 0
transform 1 0 10120 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 0
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 0
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 0
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_128
timestamp 0
transform 1 0 12880 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_141
timestamp 0
transform 1 0 14076 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_147
timestamp 0
transform 1 0 14628 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 0
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_190
timestamp 0
transform 1 0 18584 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_200
timestamp 0
transform 1 0 19504 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_204
timestamp 0
transform 1 0 19872 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_211
timestamp 0
transform 1 0 20516 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 0
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 0
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_237
timestamp 0
transform 1 0 22908 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_241
timestamp 0
transform 1 0 23276 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_245
timestamp 0
transform 1 0 23644 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_257
timestamp 0
transform 1 0 24748 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 0
transform 1 0 25852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 0
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 0
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 0
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_305
timestamp 0
transform 1 0 29164 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 0
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_340
timestamp 0
transform 1 0 32384 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 0
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 0
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 0
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 0
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_413
timestamp 0
transform 1 0 39100 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_425
timestamp 0
transform 1 0 40204 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_431
timestamp 0
transform 1 0 40756 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_439
timestamp 0
transform 1 0 41492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_458
timestamp 0
transform 1 0 43240 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_462
timestamp 0
transform 1 0 43608 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_474
timestamp 0
transform 1 0 44712 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_491
timestamp 0
transform 1 0 46276 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_3
timestamp 0
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_14
timestamp 0
transform 1 0 2392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_25
timestamp 0
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_41
timestamp 0
transform 1 0 4876 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_58
timestamp 0
transform 1 0 6440 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_66
timestamp 0
transform 1 0 7176 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_72
timestamp 0
transform 1 0 7728 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_113
timestamp 0
transform 1 0 11500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_165
timestamp 0
transform 1 0 16284 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 0
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_220
timestamp 0
transform 1 0 21344 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_232
timestamp 0
transform 1 0 22448 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 0
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 0
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 0
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 0
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 0
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 0
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 0
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 0
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 0
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_333
timestamp 0
transform 1 0 31740 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 0
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_369
timestamp 0
transform 1 0 35052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_381
timestamp 0
transform 1 0 36156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_389
timestamp 0
transform 1 0 36892 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_403
timestamp 0
transform 1 0 38180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_415
timestamp 0
transform 1 0 39284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 0
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 0
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 0
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_457
timestamp 0
transform 1 0 43148 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_466
timestamp 0
transform 1 0 43976 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_477
timestamp 0
transform 1 0 44988 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 0
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 0
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 0
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 0
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 0
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_65
timestamp 0
transform 1 0 7084 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_82
timestamp 0
transform 1 0 8648 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_94
timestamp 0
transform 1 0 9752 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 0
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 0
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 0
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_149
timestamp 0
transform 1 0 14812 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_157
timestamp 0
transform 1 0 15548 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 0
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 0
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_195
timestamp 0
transform 1 0 19044 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_203
timestamp 0
transform 1 0 19780 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_215
timestamp 0
transform 1 0 20884 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 0
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_236
timestamp 0
transform 1 0 22816 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_244
timestamp 0
transform 1 0 23552 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_252
timestamp 0
transform 1 0 24288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 0
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_309
timestamp 0
transform 1 0 29532 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_321
timestamp 0
transform 1 0 30636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 0
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_337
timestamp 0
transform 1 0 32108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_350
timestamp 0
transform 1 0 33304 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 0
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_409
timestamp 0
transform 1 0 38732 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_427
timestamp 0
transform 1 0 40388 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_433
timestamp 0
transform 1 0 40940 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_438
timestamp 0
transform 1 0 41400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 0
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 0
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 0
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_485
timestamp 0
transform 1 0 45724 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_490
timestamp 0
transform 1 0 46184 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_496
timestamp 0
transform 1 0 46736 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_6
timestamp 0
transform 1 0 1656 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_10
timestamp 0
transform 1 0 2024 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_14
timestamp 0
transform 1 0 2392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_25
timestamp 0
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_29
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_55
timestamp 0
transform 1 0 6164 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 0
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_118
timestamp 0
transform 1 0 11960 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_130
timestamp 0
transform 1 0 13064 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_135
timestamp 0
transform 1 0 13524 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 0
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_145
timestamp 0
transform 1 0 14444 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_157
timestamp 0
transform 1 0 15548 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_165
timestamp 0
transform 1 0 16284 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_170
timestamp 0
transform 1 0 16744 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_186
timestamp 0
transform 1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 0
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 0
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_223
timestamp 0
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_253
timestamp 0
transform 1 0 24380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_303
timestamp 0
transform 1 0 28980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 0
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 0
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_336
timestamp 0
transform 1 0 32016 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_348
timestamp 0
transform 1 0 33120 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 0
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_377
timestamp 0
transform 1 0 35788 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_404
timestamp 0
transform 1 0 38272 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_413
timestamp 0
transform 1 0 39100 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 0
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_445
timestamp 0
transform 1 0 42044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 0
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 0
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 0
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 0
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_489
timestamp 0
transform 1 0 46092 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_32
timestamp 0
transform 1 0 4048 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_36
timestamp 0
transform 1 0 4416 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_69
timestamp 0
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_89
timestamp 0
transform 1 0 9292 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_123
timestamp 0
transform 1 0 12420 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_127
timestamp 0
transform 1 0 12788 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_153
timestamp 0
transform 1 0 15180 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_161
timestamp 0
transform 1 0 15916 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 0
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_178
timestamp 0
transform 1 0 17480 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_186
timestamp 0
transform 1 0 18216 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_196
timestamp 0
transform 1 0 19136 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 0
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_231
timestamp 0
transform 1 0 22356 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_235
timestamp 0
transform 1 0 22724 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_243
timestamp 0
transform 1 0 23460 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_251
timestamp 0
transform 1 0 24196 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_268
timestamp 0
transform 1 0 25760 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_281
timestamp 0
transform 1 0 26956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_312
timestamp 0
transform 1 0 29808 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_318
timestamp 0
transform 1 0 30360 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_328
timestamp 0
transform 1 0 31280 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 0
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 0
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 0
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 0
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 0
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 0
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_403
timestamp 0
transform 1 0 38180 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_410
timestamp 0
transform 1 0 38824 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_418
timestamp 0
transform 1 0 39560 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_430
timestamp 0
transform 1 0 40664 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_442
timestamp 0
transform 1 0 41768 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_455
timestamp 0
transform 1 0 42964 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_467
timestamp 0
transform 1 0 44068 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_479
timestamp 0
transform 1 0 45172 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_491
timestamp 0
transform 1 0 46276 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 0
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 0
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_33
timestamp 0
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_58
timestamp 0
transform 1 0 6440 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_70
timestamp 0
transform 1 0 7544 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_78
timestamp 0
transform 1 0 8280 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_101
timestamp 0
transform 1 0 10396 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_107
timestamp 0
transform 1 0 10948 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_114
timestamp 0
transform 1 0 11592 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_126
timestamp 0
transform 1 0 12696 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 0
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 0
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_154
timestamp 0
transform 1 0 15272 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_174
timestamp 0
transform 1 0 17112 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 0
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 0
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_221
timestamp 0
transform 1 0 21436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_231
timestamp 0
transform 1 0 22356 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 0
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 0
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 0
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 0
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 0
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 0
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 0
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_309
timestamp 0
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_329
timestamp 0
transform 1 0 31372 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_341
timestamp 0
transform 1 0 32476 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 0
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 0
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 0
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_377
timestamp 0
transform 1 0 35788 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_381
timestamp 0
transform 1 0 36156 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_392
timestamp 0
transform 1 0 37168 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_404
timestamp 0
transform 1 0 38272 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_414
timestamp 0
transform 1 0 39192 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 0
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_433
timestamp 0
transform 1 0 40940 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_441
timestamp 0
transform 1 0 41676 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_456
timestamp 0
transform 1 0 43056 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_472
timestamp 0
transform 1 0 44528 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_3
timestamp 0
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_11
timestamp 0
transform 1 0 2116 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 0
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_27
timestamp 0
transform 1 0 3588 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 0
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 0
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_81
timestamp 0
transform 1 0 8556 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_92
timestamp 0
transform 1 0 9568 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_104
timestamp 0
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 0
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_119
timestamp 0
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_132
timestamp 0
transform 1 0 13248 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_156
timestamp 0
transform 1 0 15456 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_182
timestamp 0
transform 1 0 17848 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_192
timestamp 0
transform 1 0 18768 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_210
timestamp 0
transform 1 0 20424 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_214
timestamp 0
transform 1 0 20792 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 0
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 0
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 0
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_249
timestamp 0
transform 1 0 24012 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_255
timestamp 0
transform 1 0 24564 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_271
timestamp 0
transform 1 0 26036 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 0
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_281
timestamp 0
transform 1 0 26956 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_312
timestamp 0
transform 1 0 29808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_316
timestamp 0
transform 1 0 30176 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_320
timestamp 0
transform 1 0 30544 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 0
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_337
timestamp 0
transform 1 0 32108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_349
timestamp 0
transform 1 0 33212 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 0
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_393
timestamp 0
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_401
timestamp 0
transform 1 0 37996 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_414
timestamp 0
transform 1 0 39192 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_423
timestamp 0
transform 1 0 40020 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_432
timestamp 0
transform 1 0 40848 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_443
timestamp 0
transform 1 0 41860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 0
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_453
timestamp 0
transform 1 0 42780 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_461
timestamp 0
transform 1 0 43516 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_479
timestamp 0
transform 1 0 45172 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_496
timestamp 0
transform 1 0 46736 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 0
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 0
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 0
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_29
timestamp 0
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_46
timestamp 0
transform 1 0 5336 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 0
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_75
timestamp 0
transform 1 0 8004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 0
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 0
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_97
timestamp 0
transform 1 0 10028 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_105
timestamp 0
transform 1 0 10764 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 0
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 0
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_149
timestamp 0
transform 1 0 14812 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_154
timestamp 0
transform 1 0 15272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_158
timestamp 0
transform 1 0 15640 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_178
timestamp 0
transform 1 0 17480 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_184
timestamp 0
transform 1 0 18032 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 0
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 0
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_221
timestamp 0
transform 1 0 21436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_242
timestamp 0
transform 1 0 23368 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_269
timestamp 0
transform 1 0 25852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 0
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_316
timestamp 0
transform 1 0 30176 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_322
timestamp 0
transform 1 0 30728 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_332
timestamp 0
transform 1 0 31648 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_351
timestamp 0
transform 1 0 33396 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 0
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_365
timestamp 0
transform 1 0 34684 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_371
timestamp 0
transform 1 0 35236 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_413
timestamp 0
transform 1 0 39100 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_429
timestamp 0
transform 1 0 40572 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_437
timestamp 0
transform 1 0 41308 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_452
timestamp 0
transform 1 0 42688 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_461
timestamp 0
transform 1 0 43516 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_473
timestamp 0
transform 1 0 44620 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_495
timestamp 0
transform 1 0 46644 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 0
transform 1 0 1748 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_21
timestamp 0
transform 1 0 3036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_33
timestamp 0
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 0
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 0
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 0
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_69
timestamp 0
transform 1 0 7452 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_102
timestamp 0
transform 1 0 10488 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 0
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_113
timestamp 0
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_124
timestamp 0
transform 1 0 12512 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_136
timestamp 0
transform 1 0 13616 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_148
timestamp 0
transform 1 0 14720 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_160
timestamp 0
transform 1 0 15824 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_179
timestamp 0
transform 1 0 17572 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 0
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 0
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_246
timestamp 0
transform 1 0 23736 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_254
timestamp 0
transform 1 0 24472 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_260
timestamp 0
transform 1 0 25024 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_297
timestamp 0
transform 1 0 28428 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_303
timestamp 0
transform 1 0 28980 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_310
timestamp 0
transform 1 0 29624 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_337
timestamp 0
transform 1 0 32108 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_341
timestamp 0
transform 1 0 32476 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_347
timestamp 0
transform 1 0 33028 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_372
timestamp 0
transform 1 0 35328 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_386
timestamp 0
transform 1 0 36616 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 0
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_401
timestamp 0
transform 1 0 37996 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_408
timestamp 0
transform 1 0 38640 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_442
timestamp 0
transform 1 0 41768 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 0
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_461
timestamp 0
transform 1 0 43516 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_468
timestamp 0
transform 1 0 44160 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_475
timestamp 0
transform 1 0 44804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_487
timestamp 0
transform 1 0 45908 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_496
timestamp 0
transform 1 0 46736 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 0
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_7
timestamp 0
transform 1 0 1748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 0
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_45
timestamp 0
transform 1 0 5244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_57
timestamp 0
transform 1 0 6348 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_63
timestamp 0
transform 1 0 6900 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_76
timestamp 0
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 0
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 0
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 0
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_117
timestamp 0
transform 1 0 11868 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_127
timestamp 0
transform 1 0 12788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 0
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_144
timestamp 0
transform 1 0 14352 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_180
timestamp 0
transform 1 0 17664 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 0
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 0
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_209
timestamp 0
transform 1 0 20332 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_217
timestamp 0
transform 1 0 21068 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_225
timestamp 0
transform 1 0 21804 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_237
timestamp 0
transform 1 0 22908 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 0
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 0
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_265
timestamp 0
transform 1 0 25484 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_269
timestamp 0
transform 1 0 25852 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_276
timestamp 0
transform 1 0 26496 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_280
timestamp 0
transform 1 0 26864 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_284
timestamp 0
transform 1 0 27232 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_296
timestamp 0
transform 1 0 28336 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 0
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_321
timestamp 0
transform 1 0 30636 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_326
timestamp 0
transform 1 0 31096 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_338
timestamp 0
transform 1 0 32200 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_346
timestamp 0
transform 1 0 32936 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_365
timestamp 0
transform 1 0 34684 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_369
timestamp 0
transform 1 0 35052 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_381
timestamp 0
transform 1 0 36156 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_418
timestamp 0
transform 1 0 39560 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_432
timestamp 0
transform 1 0 40848 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_444
timestamp 0
transform 1 0 41952 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_456
timestamp 0
transform 1 0 43056 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_483
timestamp 0
transform 1 0 45540 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_3
timestamp 0
transform 1 0 1380 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_9
timestamp 0
transform 1 0 1932 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_13
timestamp 0
transform 1 0 2300 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_23
timestamp 0
transform 1 0 3220 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 0
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_57
timestamp 0
transform 1 0 6348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_63
timestamp 0
transform 1 0 6900 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_73
timestamp 0
transform 1 0 7820 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_82
timestamp 0
transform 1 0 8648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_106
timestamp 0
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_139
timestamp 0
transform 1 0 13892 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_150
timestamp 0
transform 1 0 14904 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_163
timestamp 0
transform 1 0 16100 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 0
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 0
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_179
timestamp 0
transform 1 0 17572 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_183
timestamp 0
transform 1 0 17940 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_199
timestamp 0
transform 1 0 19412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_211
timestamp 0
transform 1 0 20516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 0
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 0
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_237
timestamp 0
transform 1 0 22908 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_250
timestamp 0
transform 1 0 24104 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_262
timestamp 0
transform 1 0 25208 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_268
timestamp 0
transform 1 0 25760 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 0
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 0
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 0
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 0
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 0
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 0
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 0
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 0
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 0
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_349
timestamp 0
transform 1 0 33212 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_362
timestamp 0
transform 1 0 34408 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_374
timestamp 0
transform 1 0 35512 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_389
timestamp 0
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 0
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 0
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_420
timestamp 0
transform 1 0 39744 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_432
timestamp 0
transform 1 0 40848 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_444
timestamp 0
transform 1 0 41952 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_471
timestamp 0
transform 1 0 44436 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_483
timestamp 0
transform 1 0 45540 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_491
timestamp 0
transform 1 0 46276 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 0
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 0
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 0
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_53
timestamp 0
transform 1 0 5980 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_59
timestamp 0
transform 1 0 6532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_63
timestamp 0
transform 1 0 6900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_67
timestamp 0
transform 1 0 7268 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_71
timestamp 0
transform 1 0 7636 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 0
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_85
timestamp 0
transform 1 0 8924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_147
timestamp 0
transform 1 0 14628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_160
timestamp 0
transform 1 0 15824 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_166
timestamp 0
transform 1 0 16376 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_182
timestamp 0
transform 1 0 17848 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_188
timestamp 0
transform 1 0 18400 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 0
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 0
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_205
timestamp 0
transform 1 0 19964 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_220
timestamp 0
transform 1 0 21344 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_232
timestamp 0
transform 1 0 22448 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_240
timestamp 0
transform 1 0 23184 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 0
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 0
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_265
timestamp 0
transform 1 0 25484 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_271
timestamp 0
transform 1 0 26036 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_278
timestamp 0
transform 1 0 26680 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_290
timestamp 0
transform 1 0 27784 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_302
timestamp 0
transform 1 0 28888 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_309
timestamp 0
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_315
timestamp 0
transform 1 0 30084 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_325
timestamp 0
transform 1 0 31004 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_349
timestamp 0
transform 1 0 33212 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_361
timestamp 0
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_365
timestamp 0
transform 1 0 34684 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_379
timestamp 0
transform 1 0 35972 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_391
timestamp 0
transform 1 0 37076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_415
timestamp 0
transform 1 0 39284 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 0
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 0
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_433
timestamp 0
transform 1 0 40940 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_439
timestamp 0
transform 1 0 41492 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_462
timestamp 0
transform 1 0 43608 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_474
timestamp 0
transform 1 0 44712 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_477
timestamp 0
transform 1 0 44988 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_7
timestamp 0
transform 1 0 1748 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_19
timestamp 0
transform 1 0 2852 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_31
timestamp 0
transform 1 0 3956 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_44
timestamp 0
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 0
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_75
timestamp 0
transform 1 0 8004 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_100
timestamp 0
transform 1 0 10304 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_106
timestamp 0
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_113
timestamp 0
transform 1 0 11500 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_130
timestamp 0
transform 1 0 13064 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_147
timestamp 0
transform 1 0 14628 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 0
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 0
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_180
timestamp 0
transform 1 0 17664 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_215
timestamp 0
transform 1 0 20884 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 0
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_234
timestamp 0
transform 1 0 22632 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_258
timestamp 0
transform 1 0 24840 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_275
timestamp 0
transform 1 0 26404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 0
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_297
timestamp 0
transform 1 0 28428 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_301
timestamp 0
transform 1 0 28796 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_323
timestamp 0
transform 1 0 30820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 0
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_340
timestamp 0
transform 1 0 32384 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_346
timestamp 0
transform 1 0 32936 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_368
timestamp 0
transform 1 0 34960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_393
timestamp 0
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_401
timestamp 0
transform 1 0 37996 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_405
timestamp 0
transform 1 0 38364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_412
timestamp 0
transform 1 0 39008 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_429
timestamp 0
transform 1 0 40572 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 0
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_449
timestamp 0
transform 1 0 42412 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 0
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_473
timestamp 0
transform 1 0 44620 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_495
timestamp 0
transform 1 0 46644 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_3
timestamp 0
transform 1 0 1380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_25
timestamp 0
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_38
timestamp 0
transform 1 0 4600 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_46
timestamp 0
transform 1 0 5336 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_60
timestamp 0
transform 1 0 6624 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 0
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 0
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_111
timestamp 0
transform 1 0 11316 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_117
timestamp 0
transform 1 0 11868 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_124
timestamp 0
transform 1 0 12512 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 0
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_141
timestamp 0
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_158
timestamp 0
transform 1 0 15640 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_183
timestamp 0
transform 1 0 17940 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_235
timestamp 0
transform 1 0 22724 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_269
timestamp 0
transform 1 0 25852 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_301
timestamp 0
transform 1 0 28796 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_330
timestamp 0
transform 1 0 31464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_365
timestamp 0
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_417
timestamp 0
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_431
timestamp 0
transform 1 0 40756 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_444
timestamp 0
transform 1 0 41952 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_456
timestamp 0
transform 1 0 43056 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_468
timestamp 0
transform 1 0 44160 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_477
timestamp 0
transform 1 0 44988 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_481
timestamp 0
transform 1 0 45356 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_493
timestamp 0
transform 1 0 46460 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_3
timestamp 0
transform 1 0 1380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_14
timestamp 0
transform 1 0 2392 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_32
timestamp 0
transform 1 0 4048 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_48
timestamp 0
transform 1 0 5520 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_57
timestamp 0
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_65
timestamp 0
transform 1 0 7084 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_72
timestamp 0
transform 1 0 7728 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_84
timestamp 0
transform 1 0 8832 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_96
timestamp 0
transform 1 0 9936 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 0
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 0
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_132
timestamp 0
transform 1 0 13248 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_156
timestamp 0
transform 1 0 15456 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 0
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_175
timestamp 0
transform 1 0 17204 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_183
timestamp 0
transform 1 0 17940 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_216
timestamp 0
transform 1 0 20976 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_234
timestamp 0
transform 1 0 22632 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_267
timestamp 0
transform 1 0 25668 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_275
timestamp 0
transform 1 0 26404 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 0
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_294
timestamp 0
transform 1 0 28152 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_300
timestamp 0
transform 1 0 28704 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_304
timestamp 0
transform 1 0 29072 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_325
timestamp 0
transform 1 0 31004 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_363
timestamp 0
transform 1 0 34500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_375
timestamp 0
transform 1 0 35604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_387
timestamp 0
transform 1 0 36708 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 0
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_393
timestamp 0
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_401
timestamp 0
transform 1 0 37996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_411
timestamp 0
transform 1 0 38916 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_419
timestamp 0
transform 1 0 39652 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_427
timestamp 0
transform 1 0 40388 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_435
timestamp 0
transform 1 0 41124 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 0
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_454
timestamp 0
transform 1 0 42872 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_460
timestamp 0
transform 1 0 43424 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_485
timestamp 0
transform 1 0 45724 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 0
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_15
timestamp 0
transform 1 0 2484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_25
timestamp 0
transform 1 0 3404 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_29
timestamp 0
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_33
timestamp 0
transform 1 0 4140 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_53
timestamp 0
transform 1 0 5980 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_61
timestamp 0
transform 1 0 6716 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_71
timestamp 0
transform 1 0 7636 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_78
timestamp 0
transform 1 0 8280 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_48_112
timestamp 0
transform 1 0 11408 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_135
timestamp 0
transform 1 0 13524 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 0
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_147
timestamp 0
transform 1 0 14628 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_156
timestamp 0
transform 1 0 15456 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_168
timestamp 0
transform 1 0 16560 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_180
timestamp 0
transform 1 0 17664 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 0
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 0
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_197
timestamp 0
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_204
timestamp 0
transform 1 0 19872 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_212
timestamp 0
transform 1 0 20608 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_216
timestamp 0
transform 1 0 20976 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_220
timestamp 0
transform 1 0 21344 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_225
timestamp 0
transform 1 0 21804 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_237
timestamp 0
transform 1 0 22908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 0
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 0
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_265
timestamp 0
transform 1 0 25484 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_271
timestamp 0
transform 1 0 26036 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_297
timestamp 0
transform 1 0 28428 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_301
timestamp 0
transform 1 0 28796 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_325
timestamp 0
transform 1 0 31004 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_333
timestamp 0
transform 1 0 31740 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_345
timestamp 0
transform 1 0 32844 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_359
timestamp 0
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 0
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 0
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 0
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_396
timestamp 0
transform 1 0 37536 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_404
timestamp 0
transform 1 0 38272 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_411
timestamp 0
transform 1 0 38916 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 0
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 0
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_433
timestamp 0
transform 1 0 40940 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_441
timestamp 0
transform 1 0 41676 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_446
timestamp 0
transform 1 0 42136 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_458
timestamp 0
transform 1 0 43240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_462
timestamp 0
transform 1 0 43608 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 0
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_480
timestamp 0
transform 1 0 45264 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_492
timestamp 0
transform 1 0 46368 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_496
timestamp 0
transform 1 0 46736 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 0
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 0
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 0
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_39
timestamp 0
transform 1 0 4692 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_66
timestamp 0
transform 1 0 7176 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_86
timestamp 0
transform 1 0 9016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_116
timestamp 0
transform 1 0 11776 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_124
timestamp 0
transform 1 0 12512 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_151
timestamp 0
transform 1 0 14996 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_169
timestamp 0
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_214
timestamp 0
transform 1 0 20792 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 0
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 0
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 0
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 0
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 0
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 0
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 0
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 0
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 0
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 0
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 0
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 0
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 0
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_349
timestamp 0
transform 1 0 33212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_369
timestamp 0
transform 1 0 35052 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_377
timestamp 0
transform 1 0 35788 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_389
timestamp 0
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_400
timestamp 0
transform 1 0 37904 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_404
timestamp 0
transform 1 0 38272 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_414
timestamp 0
transform 1 0 39192 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_426
timestamp 0
transform 1 0 40296 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_435
timestamp 0
transform 1 0 41124 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 0
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_455
timestamp 0
transform 1 0 42964 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_467
timestamp 0
transform 1 0 44068 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_479
timestamp 0
transform 1 0 45172 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_491
timestamp 0
transform 1 0 46276 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_13
timestamp 0
transform 1 0 2300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_25
timestamp 0
transform 1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 0
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_41
timestamp 0
transform 1 0 4876 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_50
timestamp 0
transform 1 0 5704 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_58
timestamp 0
transform 1 0 6440 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_69
timestamp 0
transform 1 0 7452 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_74
timestamp 0
transform 1 0 7912 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_80
timestamp 0
transform 1 0 8464 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 0
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_89
timestamp 0
transform 1 0 9292 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_99
timestamp 0
transform 1 0 10212 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_127
timestamp 0
transform 1 0 12788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 0
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 0
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_197
timestamp 0
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_205
timestamp 0
transform 1 0 19964 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_224
timestamp 0
transform 1 0 21712 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_231
timestamp 0
transform 1 0 22356 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_236
timestamp 0
transform 1 0 22816 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 0
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 0
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_261
timestamp 0
transform 1 0 25116 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_268
timestamp 0
transform 1 0 25760 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_280
timestamp 0
transform 1 0 26864 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_292
timestamp 0
transform 1 0 27968 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_325
timestamp 0
transform 1 0 31004 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_337
timestamp 0
transform 1 0 32108 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_349
timestamp 0
transform 1 0 33212 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_361
timestamp 0
transform 1 0 34316 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_365
timestamp 0
transform 1 0 34684 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_380
timestamp 0
transform 1 0 36064 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_392
timestamp 0
transform 1 0 37168 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_396
timestamp 0
transform 1 0 37536 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_401
timestamp 0
transform 1 0 37996 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_410
timestamp 0
transform 1 0 38824 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 0
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_425
timestamp 0
transform 1 0 40204 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_460
timestamp 0
transform 1 0 43424 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_472
timestamp 0
transform 1 0 44528 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_487
timestamp 0
transform 1 0 45908 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_496
timestamp 0
transform 1 0 46736 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_3
timestamp 0
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_18
timestamp 0
transform 1 0 2760 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_40
timestamp 0
transform 1 0 4784 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_46
timestamp 0
transform 1 0 5336 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_50
timestamp 0
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_66
timestamp 0
transform 1 0 7176 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_90
timestamp 0
transform 1 0 9384 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_96
timestamp 0
transform 1 0 9936 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_107
timestamp 0
transform 1 0 10948 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 0
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 0
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_119
timestamp 0
transform 1 0 12052 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_131
timestamp 0
transform 1 0 13156 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_141
timestamp 0
transform 1 0 14076 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_153
timestamp 0
transform 1 0 15180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 0
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_178
timestamp 0
transform 1 0 17480 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_182
timestamp 0
transform 1 0 17848 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_185
timestamp 0
transform 1 0 18124 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_196
timestamp 0
transform 1 0 19136 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_204
timestamp 0
transform 1 0 19872 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_212
timestamp 0
transform 1 0 20608 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_235
timestamp 0
transform 1 0 22724 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_242
timestamp 0
transform 1 0 23368 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_264
timestamp 0
transform 1 0 25392 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_273
timestamp 0
transform 1 0 26220 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_297
timestamp 0
transform 1 0 28428 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_309
timestamp 0
transform 1 0 29532 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_317
timestamp 0
transform 1 0 30268 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_358
timestamp 0
transform 1 0 34040 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_370
timestamp 0
transform 1 0 35144 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_378
timestamp 0
transform 1 0 35880 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_387
timestamp 0
transform 1 0 36708 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 0
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_397
timestamp 0
transform 1 0 37628 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_432
timestamp 0
transform 1 0 40848 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_449
timestamp 0
transform 1 0 42412 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_455
timestamp 0
transform 1 0 42964 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_492
timestamp 0
transform 1 0 46368 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_496
timestamp 0
transform 1 0 46736 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 0
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_23
timestamp 0
transform 1 0 3220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 0
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_41
timestamp 0
transform 1 0 4876 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_58
timestamp 0
transform 1 0 6440 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_70
timestamp 0
transform 1 0 7544 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 0
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 0
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_97
timestamp 0
transform 1 0 10028 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_110
timestamp 0
transform 1 0 11224 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_122
timestamp 0
transform 1 0 12328 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 0
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 0
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 0
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 0
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 0
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 0
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 0
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 0
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_209
timestamp 0
transform 1 0 20332 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_218
timestamp 0
transform 1 0 21160 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_222
timestamp 0
transform 1 0 21528 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_231
timestamp 0
transform 1 0 22356 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_235
timestamp 0
transform 1 0 22724 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 0
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_277
timestamp 0
transform 1 0 26588 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_283
timestamp 0
transform 1 0 27140 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_293
timestamp 0
transform 1 0 28060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_305
timestamp 0
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_309
timestamp 0
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_336
timestamp 0
transform 1 0 32016 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_358
timestamp 0
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_388
timestamp 0
transform 1 0 36800 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_406
timestamp 0
transform 1 0 38456 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_418
timestamp 0
transform 1 0 39560 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_434
timestamp 0
transform 1 0 41032 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_446
timestamp 0
transform 1 0 42136 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_458
timestamp 0
transform 1 0 43240 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_470
timestamp 0
transform 1 0 44344 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_52_477
timestamp 0
transform 1 0 44988 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_490
timestamp 0
transform 1 0 46184 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_496
timestamp 0
transform 1 0 46736 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 0
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_9
timestamp 0
transform 1 0 1932 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_13
timestamp 0
transform 1 0 2300 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_25
timestamp 0
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_37
timestamp 0
transform 1 0 4508 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_49
timestamp 0
transform 1 0 5612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 0
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 0
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 0
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 0
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_102
timestamp 0
transform 1 0 10488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 0
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_113
timestamp 0
transform 1 0 11500 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_124
timestamp 0
transform 1 0 12512 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_136
timestamp 0
transform 1 0 13616 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_148
timestamp 0
transform 1 0 14720 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_159
timestamp 0
transform 1 0 15732 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 0
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 0
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 0
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 0
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_205
timestamp 0
transform 1 0 19964 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_209
timestamp 0
transform 1 0 20332 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 0
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 0
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_236
timestamp 0
transform 1 0 22816 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_265
timestamp 0
transform 1 0 25484 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 0
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 0
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_281
timestamp 0
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_300
timestamp 0
transform 1 0 28704 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_312
timestamp 0
transform 1 0 29808 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_320
timestamp 0
transform 1 0 30544 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 0
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_346
timestamp 0
transform 1 0 32936 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_379
timestamp 0
transform 1 0 35972 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 0
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_393
timestamp 0
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_399
timestamp 0
transform 1 0 37812 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_411
timestamp 0
transform 1 0 38916 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_423
timestamp 0
transform 1 0 40020 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_435
timestamp 0
transform 1 0 41124 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_445
timestamp 0
transform 1 0 42044 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 0
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 0
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_473
timestamp 0
transform 1 0 44620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_480
timestamp 0
transform 1 0 45264 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_492
timestamp 0
transform 1 0 46368 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_496
timestamp 0
transform 1 0 46736 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_13
timestamp 0
transform 1 0 2300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_25
timestamp 0
transform 1 0 3404 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 0
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 0
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_53
timestamp 0
transform 1 0 5980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_73
timestamp 0
transform 1 0 7820 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_109
timestamp 0
transform 1 0 11132 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_134
timestamp 0
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_141
timestamp 0
transform 1 0 14076 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_158
timestamp 0
transform 1 0 15640 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_164
timestamp 0
transform 1 0 16192 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_182
timestamp 0
transform 1 0 17848 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 0
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_224
timestamp 0
transform 1 0 21712 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_241
timestamp 0
transform 1 0 23276 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_249
timestamp 0
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 0
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 0
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_304
timestamp 0
transform 1 0 29072 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_335
timestamp 0
transform 1 0 31924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_347
timestamp 0
transform 1 0 33028 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_355
timestamp 0
transform 1 0 33764 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 0
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_374
timestamp 0
transform 1 0 35512 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_389
timestamp 0
transform 1 0 36892 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_409
timestamp 0
transform 1 0 38732 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_417
timestamp 0
transform 1 0 39468 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_431
timestamp 0
transform 1 0 40756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_443
timestamp 0
transform 1 0 41860 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_447
timestamp 0
transform 1 0 42228 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_452
timestamp 0
transform 1 0 42688 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_464
timestamp 0
transform 1 0 43792 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_480
timestamp 0
transform 1 0 45264 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_492
timestamp 0
transform 1 0 46368 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_496
timestamp 0
transform 1 0 46736 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_3
timestamp 0
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_31
timestamp 0
transform 1 0 3956 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_73
timestamp 0
transform 1 0 7820 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_90
timestamp 0
transform 1 0 9384 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_132
timestamp 0
transform 1 0 13248 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_160
timestamp 0
transform 1 0 15824 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 0
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 0
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_230
timestamp 0
transform 1 0 22264 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_242
timestamp 0
transform 1 0 23368 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_247
timestamp 0
transform 1 0 23828 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_255
timestamp 0
transform 1 0 24564 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_269
timestamp 0
transform 1 0 25852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 0
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_327
timestamp 0
transform 1 0 31188 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 0
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_346
timestamp 0
transform 1 0 32936 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_358
timestamp 0
transform 1 0 34040 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_370
timestamp 0
transform 1 0 35144 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_382
timestamp 0
transform 1 0 36248 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_393
timestamp 0
transform 1 0 37260 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_401
timestamp 0
transform 1 0 37996 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_413
timestamp 0
transform 1 0 39100 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_433
timestamp 0
transform 1 0 40940 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_439
timestamp 0
transform 1 0 41492 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_461
timestamp 0
transform 1 0 43516 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_480
timestamp 0
transform 1 0 45264 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_491
timestamp 0
transform 1 0 46276 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_3
timestamp 0
transform 1 0 1380 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_23
timestamp 0
transform 1 0 3220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 0
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_29
timestamp 0
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_53
timestamp 0
transform 1 0 5980 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 0
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_85
timestamp 0
transform 1 0 8924 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_105
timestamp 0
transform 1 0 10764 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 0
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 0
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_141
timestamp 0
transform 1 0 14076 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_163
timestamp 0
transform 1 0 16100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_173
timestamp 0
transform 1 0 17020 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_222
timestamp 0
transform 1 0 21528 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_230
timestamp 0
transform 1 0 22264 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_243
timestamp 0
transform 1 0 23460 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 0
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_253
timestamp 0
transform 1 0 24380 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_270
timestamp 0
transform 1 0 25944 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_283
timestamp 0
transform 1 0 27140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_295
timestamp 0
transform 1 0 28244 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_303
timestamp 0
transform 1 0 28980 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_318
timestamp 0
transform 1 0 30360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_330
timestamp 0
transform 1 0 31464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_334
timestamp 0
transform 1 0 31832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_354
timestamp 0
transform 1 0 33672 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 0
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_365
timestamp 0
transform 1 0 34684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_373
timestamp 0
transform 1 0 35420 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_394
timestamp 0
transform 1 0 37352 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_400
timestamp 0
transform 1 0 37904 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_405
timestamp 0
transform 1 0 38364 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_412
timestamp 0
transform 1 0 39008 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_56_421
timestamp 0
transform 1 0 39836 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_427
timestamp 0
transform 1 0 40388 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_436
timestamp 0
transform 1 0 41216 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_454
timestamp 0
transform 1 0 42872 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_466
timestamp 0
transform 1 0 43976 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_489
timestamp 0
transform 1 0 46092 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_3
timestamp 0
transform 1 0 1380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_11
timestamp 0
transform 1 0 2116 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_15
timestamp 0
transform 1 0 2484 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_25
timestamp 0
transform 1 0 3404 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_47
timestamp 0
transform 1 0 5428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 0
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 0
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 0
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_81
timestamp 0
transform 1 0 8556 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_89
timestamp 0
transform 1 0 9292 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_100
timestamp 0
transform 1 0 10304 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 0
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_124
timestamp 0
transform 1 0 12512 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_134
timestamp 0
transform 1 0 13432 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_146
timestamp 0
transform 1 0 14536 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_158
timestamp 0
transform 1 0 15640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 0
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 0
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_181
timestamp 0
transform 1 0 17756 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_189
timestamp 0
transform 1 0 18492 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_197
timestamp 0
transform 1 0 19228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_209
timestamp 0
transform 1 0 20332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 0
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_225
timestamp 0
transform 1 0 21804 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_229
timestamp 0
transform 1 0 22172 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_246
timestamp 0
transform 1 0 23736 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 0
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 0
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 0
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 0
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 0
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 0
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_346
timestamp 0
transform 1 0 32936 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_358
timestamp 0
transform 1 0 34040 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_374
timestamp 0
transform 1 0 35512 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_386
timestamp 0
transform 1 0 36616 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_57_393
timestamp 0
transform 1 0 37260 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_412
timestamp 0
transform 1 0 39008 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_427
timestamp 0
transform 1 0 40388 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_438
timestamp 0
transform 1 0 41400 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 0
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_457
timestamp 0
transform 1 0 43148 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_496
timestamp 0
transform 1 0 46736 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 0
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 0
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 0
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_29
timestamp 0
transform 1 0 3772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_35
timestamp 0
transform 1 0 4324 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_45
timestamp 0
transform 1 0 5244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_57
timestamp 0
transform 1 0 6348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_69
timestamp 0
transform 1 0 7452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_81
timestamp 0
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 0
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 0
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 0
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 0
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 0
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 0
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 0
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_174
timestamp 0
transform 1 0 17112 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_186
timestamp 0
transform 1 0 18216 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_190
timestamp 0
transform 1 0 18584 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 0
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_209
timestamp 0
transform 1 0 20332 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_225
timestamp 0
transform 1 0 21804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_230
timestamp 0
transform 1 0 22264 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_242
timestamp 0
transform 1 0 23368 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 0
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 0
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 0
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 0
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 0
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 0
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 0
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 0
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_321
timestamp 0
transform 1 0 30636 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_329
timestamp 0
transform 1 0 31372 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_349
timestamp 0
transform 1 0 33212 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_357
timestamp 0
transform 1 0 33948 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_381
timestamp 0
transform 1 0 36156 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_389
timestamp 0
transform 1 0 36892 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_400
timestamp 0
transform 1 0 37904 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_412
timestamp 0
transform 1 0 39008 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_421
timestamp 0
transform 1 0 39836 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_429
timestamp 0
transform 1 0 40572 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_437
timestamp 0
transform 1 0 41308 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_443
timestamp 0
transform 1 0 41860 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_450
timestamp 0
transform 1 0 42504 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_456
timestamp 0
transform 1 0 43056 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_460
timestamp 0
transform 1 0 43424 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_472
timestamp 0
transform 1 0 44528 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_481
timestamp 0
transform 1 0 45356 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_493
timestamp 0
transform 1 0 46460 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_9
timestamp 0
transform 1 0 1932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_30
timestamp 0
transform 1 0 3864 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_42
timestamp 0
transform 1 0 4968 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 0
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 0
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 0
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_123
timestamp 0
transform 1 0 12420 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_129
timestamp 0
transform 1 0 12972 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_155
timestamp 0
transform 1 0 15364 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 0
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_189
timestamp 0
transform 1 0 18492 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_204
timestamp 0
transform 1 0 19872 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_216
timestamp 0
transform 1 0 20976 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 0
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_237
timestamp 0
transform 1 0 22908 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_261
timestamp 0
transform 1 0 25116 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_271
timestamp 0
transform 1 0 26036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 0
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_281
timestamp 0
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_285
timestamp 0
transform 1 0 27324 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_305
timestamp 0
transform 1 0 29164 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 0
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 0
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 0
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_361
timestamp 0
transform 1 0 34316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_378
timestamp 0
transform 1 0 35880 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 0
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_393
timestamp 0
transform 1 0 37260 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_400
timestamp 0
transform 1 0 37904 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_430
timestamp 0
transform 1 0 40664 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_434
timestamp 0
transform 1 0 41032 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_453
timestamp 0
transform 1 0 42780 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_465
timestamp 0
transform 1 0 43884 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_477
timestamp 0
transform 1 0 44988 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_489
timestamp 0
transform 1 0 46092 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_3
timestamp 0
transform 1 0 1380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 0
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_29
timestamp 0
transform 1 0 3772 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_33
timestamp 0
transform 1 0 4140 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_55
timestamp 0
transform 1 0 6164 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_94
timestamp 0
transform 1 0 9752 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_126
timestamp 0
transform 1 0 12696 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_130
timestamp 0
transform 1 0 13064 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 0
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_148
timestamp 0
transform 1 0 14720 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_160
timestamp 0
transform 1 0 15824 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_172
timestamp 0
transform 1 0 16928 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 0
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_203
timestamp 0
transform 1 0 19780 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_210
timestamp 0
transform 1 0 20424 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_230
timestamp 0
transform 1 0 22264 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_245
timestamp 0
transform 1 0 23644 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 0
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_286
timestamp 0
transform 1 0 27416 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_293
timestamp 0
transform 1 0 28060 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_312
timestamp 0
transform 1 0 29808 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_334
timestamp 0
transform 1 0 31832 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_346
timestamp 0
transform 1 0 32936 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_358
timestamp 0
transform 1 0 34040 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_377
timestamp 0
transform 1 0 35788 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_395
timestamp 0
transform 1 0 37444 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_60_407
timestamp 0
transform 1 0 38548 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_60_417
timestamp 0
transform 1 0 39468 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 0
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 0
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 0
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 0
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 0
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 0
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_489
timestamp 0
transform 1 0 46092 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 0
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_7
timestamp 0
transform 1 0 1748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_30
timestamp 0
transform 1 0 3864 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 0
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_57
timestamp 0
transform 1 0 6348 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_61
timestamp 0
transform 1 0 6716 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_74
timestamp 0
transform 1 0 7912 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_80
timestamp 0
transform 1 0 8464 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_88
timestamp 0
transform 1 0 9200 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_109
timestamp 0
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 0
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_125
timestamp 0
transform 1 0 12604 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_129
timestamp 0
transform 1 0 12972 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_136
timestamp 0
transform 1 0 13616 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_143
timestamp 0
transform 1 0 14260 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_185
timestamp 0
transform 1 0 18124 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_209
timestamp 0
transform 1 0 20332 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_61_271
timestamp 0
transform 1 0 26036 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 0
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_288
timestamp 0
transform 1 0 27600 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_296
timestamp 0
transform 1 0 28336 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_328
timestamp 0
transform 1 0 31280 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_358
timestamp 0
transform 1 0 34040 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_370
timestamp 0
transform 1 0 35144 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 0
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 0
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_417
timestamp 0
transform 1 0 39468 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_432
timestamp 0
transform 1 0 40848 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_444
timestamp 0
transform 1 0 41952 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 0
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 0
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 0
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_485
timestamp 0
transform 1 0 45724 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 0
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_11
timestamp 0
transform 1 0 2116 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_22
timestamp 0
transform 1 0 3128 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_38
timestamp 0
transform 1 0 4600 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_50
timestamp 0
transform 1 0 5704 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_62
timestamp 0
transform 1 0 6808 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_74
timestamp 0
transform 1 0 7912 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 0
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_85
timestamp 0
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_93
timestamp 0
transform 1 0 9660 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_113
timestamp 0
transform 1 0 11500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_125
timestamp 0
transform 1 0 12604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_137
timestamp 0
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_145
timestamp 0
transform 1 0 14444 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_193
timestamp 0
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_197
timestamp 0
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_201
timestamp 0
transform 1 0 19596 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_214
timestamp 0
transform 1 0 20792 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_222
timestamp 0
transform 1 0 21528 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 0
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 0
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 0
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 0
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 0
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 0
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_301
timestamp 0
transform 1 0 28796 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 0
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_313
timestamp 0
transform 1 0 29900 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_325
timestamp 0
transform 1 0 31004 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 0
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_368
timestamp 0
transform 1 0 34960 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_376
timestamp 0
transform 1 0 35696 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_395
timestamp 0
transform 1 0 37444 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_407
timestamp 0
transform 1 0 38548 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 0
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 0
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 0
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 0
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 0
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 0
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 0
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 0
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_489
timestamp 0
transform 1 0 46092 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 0
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 0
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_27
timestamp 0
transform 1 0 3588 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_31
timestamp 0
transform 1 0 3956 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_41
timestamp 0
transform 1 0 4876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 0
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_57
timestamp 0
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 0
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 0
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 0
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 0
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 0
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 0
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 0
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 0
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 0
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_161
timestamp 0
transform 1 0 15916 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_178
timestamp 0
transform 1 0 17480 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_190
timestamp 0
transform 1 0 18584 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_196
timestamp 0
transform 1 0 19136 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_203
timestamp 0
transform 1 0 19780 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_215
timestamp 0
transform 1 0 20884 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 0
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 0
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_237
timestamp 0
transform 1 0 22908 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_242
timestamp 0
transform 1 0 23368 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_254
timestamp 0
transform 1 0 24472 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_266
timestamp 0
transform 1 0 25576 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 0
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_297
timestamp 0
transform 1 0 28428 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_309
timestamp 0
transform 1 0 29532 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_313
timestamp 0
transform 1 0 29900 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_318
timestamp 0
transform 1 0 30360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 0
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 0
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_341
timestamp 0
transform 1 0 32476 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_358
timestamp 0
transform 1 0 34040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_362
timestamp 0
transform 1 0 34408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_371
timestamp 0
transform 1 0 35236 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_379
timestamp 0
transform 1 0 35972 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_389
timestamp 0
transform 1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 0
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_405
timestamp 0
transform 1 0 38364 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_409
timestamp 0
transform 1 0 38732 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_426
timestamp 0
transform 1 0 40296 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_438
timestamp 0
transform 1 0 41400 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_446
timestamp 0
transform 1 0 42136 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 0
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 0
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 0
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 0
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_6
timestamp 0
transform 1 0 1656 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_18
timestamp 0
transform 1 0 2760 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 0
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 0
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_59
timestamp 0
transform 1 0 6532 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_69
timestamp 0
transform 1 0 7452 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 0
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_106
timestamp 0
transform 1 0 10856 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 0
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_152
timestamp 0
transform 1 0 15088 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_164
timestamp 0
transform 1 0 16192 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_176
timestamp 0
transform 1 0 17296 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 0
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_197
timestamp 0
transform 1 0 19228 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 0
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 0
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 0
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 0
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 0
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_274
timestamp 0
transform 1 0 26312 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 0
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 0
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_330
timestamp 0
transform 1 0 31464 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_342
timestamp 0
transform 1 0 32568 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_358
timestamp 0
transform 1 0 34040 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_64_381
timestamp 0
transform 1 0 36156 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_388
timestamp 0
transform 1 0 36800 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_400
timestamp 0
transform 1 0 37904 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_404
timestamp 0
transform 1 0 38272 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 0
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 0
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 0
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 0
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 0
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 0
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 0
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 0
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_489
timestamp 0
transform 1 0 46092 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 0
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_15
timestamp 0
transform 1 0 2484 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_23
timestamp 0
transform 1 0 3220 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_45
timestamp 0
transform 1 0 5244 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_73
timestamp 0
transform 1 0 7820 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 0
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_134
timestamp 0
transform 1 0 13432 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_160
timestamp 0
transform 1 0 15824 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_169
timestamp 0
transform 1 0 16652 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_193
timestamp 0
transform 1 0 18860 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_211
timestamp 0
transform 1 0 20516 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_218
timestamp 0
transform 1 0 21160 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_246
timestamp 0
transform 1 0 23736 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_252
timestamp 0
transform 1 0 24288 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_274
timestamp 0
transform 1 0 26312 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 0
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_281
timestamp 0
transform 1 0 26956 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_285
timestamp 0
transform 1 0 27324 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_309
timestamp 0
transform 1 0 29532 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_314
timestamp 0
transform 1 0 29992 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_325
timestamp 0
transform 1 0 31004 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_333
timestamp 0
transform 1 0 31740 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_346
timestamp 0
transform 1 0 32936 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_354
timestamp 0
transform 1 0 33672 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_366
timestamp 0
transform 1 0 34776 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_378
timestamp 0
transform 1 0 35880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_389
timestamp 0
transform 1 0 36892 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_398
timestamp 0
transform 1 0 37720 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_402
timestamp 0
transform 1 0 38088 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_419
timestamp 0
transform 1 0 39652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_431
timestamp 0
transform 1 0 40756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_443
timestamp 0
transform 1 0 41860 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 0
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 0
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 0
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 0
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_485
timestamp 0
transform 1 0 45724 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 0
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 0
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 0
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_29
timestamp 0
transform 1 0 3772 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_36
timestamp 0
transform 1 0 4416 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_48
timestamp 0
transform 1 0 5520 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_81
timestamp 0
transform 1 0 8556 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_85
timestamp 0
transform 1 0 8924 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_102
timestamp 0
transform 1 0 10488 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_108
timestamp 0
transform 1 0 11040 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_128
timestamp 0
transform 1 0 12880 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_157
timestamp 0
transform 1 0 15548 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_161
timestamp 0
transform 1 0 15916 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_165
timestamp 0
transform 1 0 16284 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_216
timestamp 0
transform 1 0 20976 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 0
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_269
timestamp 0
transform 1 0 25852 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_273
timestamp 0
transform 1 0 26220 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_299
timestamp 0
transform 1 0 28612 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 0
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_325
timestamp 0
transform 1 0 31004 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_348
timestamp 0
transform 1 0 33120 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_365
timestamp 0
transform 1 0 34684 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_396
timestamp 0
transform 1 0 37536 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_416
timestamp 0
transform 1 0 39376 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 0
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 0
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 0
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 0
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 0
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 0
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 0
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_489
timestamp 0
transform 1 0 46092 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 0
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 0
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 0
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 0
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 0
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 0
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_57
timestamp 0
transform 1 0 6348 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_65
timestamp 0
transform 1 0 7084 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_71
timestamp 0
transform 1 0 7636 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_83
timestamp 0
transform 1 0 8740 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_92
timestamp 0
transform 1 0 9568 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_104
timestamp 0
transform 1 0 10672 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 0
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 0
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 0
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_149
timestamp 0
transform 1 0 14812 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 0
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_193
timestamp 0
transform 1 0 18860 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_197
timestamp 0
transform 1 0 19228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_201
timestamp 0
transform 1 0 19596 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_211
timestamp 0
transform 1 0 20516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 0
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_241
timestamp 0
transform 1 0 23276 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_249
timestamp 0
transform 1 0 24012 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_259
timestamp 0
transform 1 0 24932 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_271
timestamp 0
transform 1 0 26036 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 0
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 0
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 0
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_305
timestamp 0
transform 1 0 29164 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_311
timestamp 0
transform 1 0 29716 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_321
timestamp 0
transform 1 0 30636 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_325
timestamp 0
transform 1 0 31004 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_330
timestamp 0
transform 1 0 31464 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_337
timestamp 0
transform 1 0 32108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_345
timestamp 0
transform 1 0 32844 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_371
timestamp 0
transform 1 0 35236 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_390
timestamp 0
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_399
timestamp 0
transform 1 0 37812 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_403
timestamp 0
transform 1 0 38180 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_408
timestamp 0
transform 1 0 38640 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_420
timestamp 0
transform 1 0 39744 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_432
timestamp 0
transform 1 0 40848 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_444
timestamp 0
transform 1 0 41952 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 0
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 0
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 0
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 0
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_3
timestamp 0
transform 1 0 1380 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_11
timestamp 0
transform 1 0 2116 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_15
timestamp 0
transform 1 0 2484 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_19
timestamp 0
transform 1 0 2852 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 0
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 0
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 0
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_53
timestamp 0
transform 1 0 5980 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_61
timestamp 0
transform 1 0 6716 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_64
timestamp 0
transform 1 0 6992 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_76
timestamp 0
transform 1 0 8096 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_85
timestamp 0
transform 1 0 8924 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_91
timestamp 0
transform 1 0 9476 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_103
timestamp 0
transform 1 0 10580 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_115
timestamp 0
transform 1 0 11684 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_125
timestamp 0
transform 1 0 12604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_137
timestamp 0
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_141
timestamp 0
transform 1 0 14076 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_151
timestamp 0
transform 1 0 14996 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_171
timestamp 0
transform 1 0 16836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_183
timestamp 0
transform 1 0 17940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 0
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 0
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 0
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 0
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_233
timestamp 0
transform 1 0 22540 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_239
timestamp 0
transform 1 0 23092 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_249
timestamp 0
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 0
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 0
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 0
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_289
timestamp 0
transform 1 0 27692 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_300
timestamp 0
transform 1 0 28704 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 0
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_349
timestamp 0
transform 1 0 33212 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_361
timestamp 0
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 0
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_377
timestamp 0
transform 1 0 35788 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_382
timestamp 0
transform 1 0 36248 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_393
timestamp 0
transform 1 0 37260 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 0
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 0
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 0
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 0
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 0
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 0
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 0
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_489
timestamp 0
transform 1 0 46092 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_7
timestamp 0
transform 1 0 1748 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_11
timestamp 0
transform 1 0 2116 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_21
timestamp 0
transform 1 0 3036 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_33
timestamp 0
transform 1 0 4140 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_45
timestamp 0
transform 1 0 5244 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_53
timestamp 0
transform 1 0 5980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_57
timestamp 0
transform 1 0 6348 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_61
timestamp 0
transform 1 0 6716 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_64
timestamp 0
transform 1 0 6992 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_68
timestamp 0
transform 1 0 7360 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_72
timestamp 0
transform 1 0 7728 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_76
timestamp 0
transform 1 0 8096 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_80
timestamp 0
transform 1 0 8464 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_87
timestamp 0
transform 1 0 9108 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_91
timestamp 0
transform 1 0 9476 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_102
timestamp 0
transform 1 0 10488 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_108
timestamp 0
transform 1 0 11040 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_129
timestamp 0
transform 1 0 12972 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_140
timestamp 0
transform 1 0 13984 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_146
timestamp 0
transform 1 0 14536 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_150
timestamp 0
transform 1 0 14904 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_162
timestamp 0
transform 1 0 16008 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_169
timestamp 0
transform 1 0 16652 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_175
timestamp 0
transform 1 0 17204 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_185
timestamp 0
transform 1 0 18124 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_197
timestamp 0
transform 1 0 19228 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_209
timestamp 0
transform 1 0 20332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_221
timestamp 0
transform 1 0 21436 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 0
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_237
timestamp 0
transform 1 0 22908 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_241
timestamp 0
transform 1 0 23276 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_69_267
timestamp 0
transform 1 0 25668 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_276
timestamp 0
transform 1 0 26496 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_290
timestamp 0
transform 1 0 27784 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_316
timestamp 0
transform 1 0 30176 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_332
timestamp 0
transform 1 0 31648 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 0
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_349
timestamp 0
transform 1 0 33212 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_359
timestamp 0
transform 1 0 34132 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_371
timestamp 0
transform 1 0 35236 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_379
timestamp 0
transform 1 0 35972 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_390
timestamp 0
transform 1 0 36984 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_397
timestamp 0
transform 1 0 37628 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 0
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 0
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 0
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 0
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 0
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 0
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 0
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 0
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_7
timestamp 0
transform 1 0 1748 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 0
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_41
timestamp 0
transform 1 0 4876 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_49
timestamp 0
transform 1 0 5612 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_52
timestamp 0
transform 1 0 5888 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_56
timestamp 0
transform 1 0 6256 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_60
timestamp 0
transform 1 0 6624 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_64
timestamp 0
transform 1 0 6992 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_68
timestamp 0
transform 1 0 7360 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_72
timestamp 0
transform 1 0 7728 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_101
timestamp 0
transform 1 0 10396 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_141
timestamp 0
transform 1 0 14076 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_162
timestamp 0
transform 1 0 16008 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_193
timestamp 0
transform 1 0 18860 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_197
timestamp 0
transform 1 0 19228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_205
timestamp 0
transform 1 0 19964 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_216
timestamp 0
transform 1 0 20976 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_224
timestamp 0
transform 1 0 21712 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 0
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_253
timestamp 0
transform 1 0 24380 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_264
timestamp 0
transform 1 0 25392 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_305
timestamp 0
transform 1 0 29164 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_70_309
timestamp 0
transform 1 0 29532 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_315
timestamp 0
transform 1 0 30084 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_332
timestamp 0
transform 1 0 31648 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_344
timestamp 0
transform 1 0 32752 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_362
timestamp 0
transform 1 0 34408 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_365
timestamp 0
transform 1 0 34684 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_373
timestamp 0
transform 1 0 35420 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_384
timestamp 0
transform 1 0 36432 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_392
timestamp 0
transform 1 0 37168 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_70_403
timestamp 0
transform 1 0 38180 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 0
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_428
timestamp 0
transform 1 0 40480 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_440
timestamp 0
transform 1 0 41584 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_452
timestamp 0
transform 1 0 42688 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_464
timestamp 0
transform 1 0 43792 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 0
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_489
timestamp 0
transform 1 0 46092 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 0
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 0
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 0
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 0
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 0
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 0
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 0
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 0
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 0
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 0
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_105
timestamp 0
transform 1 0 10764 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_109
timestamp 0
transform 1 0 11132 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_71_117
timestamp 0
transform 1 0 11868 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_71_132
timestamp 0
transform 1 0 13248 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_140
timestamp 0
transform 1 0 13984 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_158
timestamp 0
transform 1 0 15640 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_166
timestamp 0
transform 1 0 16376 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_169
timestamp 0
transform 1 0 16652 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_189
timestamp 0
transform 1 0 18492 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_71_241
timestamp 0
transform 1 0 23276 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_247
timestamp 0
transform 1 0 23828 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_270
timestamp 0
transform 1 0 25944 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_278
timestamp 0
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_281
timestamp 0
transform 1 0 26956 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_289
timestamp 0
transform 1 0 27692 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_301
timestamp 0
transform 1 0 28796 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_313
timestamp 0
transform 1 0 29900 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_325
timestamp 0
transform 1 0 31004 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_333
timestamp 0
transform 1 0 31740 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 0
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_349
timestamp 0
transform 1 0 33212 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_71_361
timestamp 0
transform 1 0 34316 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_367
timestamp 0
transform 1 0 34868 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_379
timestamp 0
transform 1 0 35972 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_390
timestamp 0
transform 1 0 36984 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_419
timestamp 0
transform 1 0 39652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_431
timestamp 0
transform 1 0 40756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_443
timestamp 0
transform 1 0 41860 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 0
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 0
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 0
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 0
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 0
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_7
timestamp 0
transform 1 0 1748 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_11
timestamp 0
transform 1 0 2116 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_23
timestamp 0
transform 1 0 3220 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 0
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 0
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 0
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 0
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 0
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 0
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 0
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 0
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_97
timestamp 0
transform 1 0 10028 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_105
timestamp 0
transform 1 0 10764 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_118
timestamp 0
transform 1 0 11960 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_130
timestamp 0
transform 1 0 13064 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_137
timestamp 0
transform 1 0 13708 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 0
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 0
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_165
timestamp 0
transform 1 0 16284 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_173
timestamp 0
transform 1 0 17020 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_184
timestamp 0
transform 1 0 18032 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_192
timestamp 0
transform 1 0 18768 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_216
timestamp 0
transform 1 0 20976 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_224
timestamp 0
transform 1 0 21712 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_229
timestamp 0
transform 1 0 22172 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_241
timestamp 0
transform 1 0 23276 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_249
timestamp 0
transform 1 0 24012 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_269
timestamp 0
transform 1 0 25852 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_281
timestamp 0
transform 1 0 26956 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_293
timestamp 0
transform 1 0 28060 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_305
timestamp 0
transform 1 0 29164 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 0
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_321
timestamp 0
transform 1 0 30636 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_325
timestamp 0
transform 1 0 31004 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_332
timestamp 0
transform 1 0 31648 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_336
timestamp 0
transform 1 0 32016 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_350
timestamp 0
transform 1 0 33304 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_358
timestamp 0
transform 1 0 34040 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_72_380
timestamp 0
transform 1 0 36064 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_72_388
timestamp 0
transform 1 0 36800 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_394
timestamp 0
transform 1 0 37352 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_406
timestamp 0
transform 1 0 38456 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_412
timestamp 0
transform 1 0 39008 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 0
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 0
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 0
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 0
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 0
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 0
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 0
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_489
timestamp 0
transform 1 0 46092 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 0
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 0
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 0
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 0
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 0
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 0
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 0
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 0
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 0
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 0
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 0
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 0
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 0
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_125
timestamp 0
transform 1 0 12604 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_131
timestamp 0
transform 1 0 13156 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_135
timestamp 0
transform 1 0 13524 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_153
timestamp 0
transform 1 0 15180 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_157
timestamp 0
transform 1 0 15548 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_162
timestamp 0
transform 1 0 16008 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 0
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_181
timestamp 0
transform 1 0 17756 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_189
timestamp 0
transform 1 0 18492 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_202
timestamp 0
transform 1 0 19688 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_214
timestamp 0
transform 1 0 20792 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 0
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 0
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 0
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 0
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 0
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 0
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 0
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 0
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 0
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_305
timestamp 0
transform 1 0 29164 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_310
timestamp 0
transform 1 0 29624 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_316
timestamp 0
transform 1 0 30176 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_361
timestamp 0
transform 1 0 34316 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_369
timestamp 0
transform 1 0 35052 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_377
timestamp 0
transform 1 0 35788 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_389
timestamp 0
transform 1 0 36892 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 0
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 0
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 0
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 0
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 0
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 0
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 0
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 0
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 0
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 0
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 0
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 0
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 0
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 0
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 0
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 0
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 0
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 0
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 0
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 0
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 0
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 0
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 0
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 0
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 0
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_166
timestamp 0
transform 1 0 16376 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_181
timestamp 0
transform 1 0 17756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_193
timestamp 0
transform 1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_206
timestamp 0
transform 1 0 20056 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_218
timestamp 0
transform 1 0 21160 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_230
timestamp 0
transform 1 0 22264 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_236
timestamp 0
transform 1 0 22816 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_248
timestamp 0
transform 1 0 23920 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 0
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 0
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_277
timestamp 0
transform 1 0 26588 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_298
timestamp 0
transform 1 0 28520 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_74_321
timestamp 0
transform 1 0 30636 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_329
timestamp 0
transform 1 0 31372 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_333
timestamp 0
transform 1 0 31740 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_341
timestamp 0
transform 1 0 32476 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_348
timestamp 0
transform 1 0 33120 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_360
timestamp 0
transform 1 0 34224 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_365
timestamp 0
transform 1 0 34684 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_369
timestamp 0
transform 1 0 35052 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_373
timestamp 0
transform 1 0 35420 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_385
timestamp 0
transform 1 0 36524 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_393
timestamp 0
transform 1 0 37260 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_411
timestamp 0
transform 1 0 38916 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_415
timestamp 0
transform 1 0 39284 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 0
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 0
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 0
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 0
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 0
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 0
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 0
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 0
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_489
timestamp 0
transform 1 0 46092 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 0
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 0
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 0
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 0
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 0
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 0
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 0
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 0
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 0
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 0
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 0
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 0
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 0
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_125
timestamp 0
transform 1 0 12604 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_133
timestamp 0
transform 1 0 13340 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_153
timestamp 0
transform 1 0 15180 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_194
timestamp 0
transform 1 0 18952 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_206
timestamp 0
transform 1 0 20056 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_75_214
timestamp 0
transform 1 0 20792 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_231
timestamp 0
transform 1 0 22356 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_252
timestamp 0
transform 1 0 24288 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_264
timestamp 0
transform 1 0 25392 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_276
timestamp 0
transform 1 0 26496 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_287
timestamp 0
transform 1 0 27508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_299
timestamp 0
transform 1 0 28612 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_323
timestamp 0
transform 1 0 30820 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 0
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 0
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_349
timestamp 0
transform 1 0 33212 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_384
timestamp 0
transform 1 0 36432 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_388
timestamp 0
transform 1 0 36800 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_402
timestamp 0
transform 1 0 38088 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_408
timestamp 0
transform 1 0 38640 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_428
timestamp 0
transform 1 0 40480 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_440
timestamp 0
transform 1 0 41584 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 0
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 0
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 0
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_485
timestamp 0
transform 1 0 45724 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 0
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 0
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 0
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_35
timestamp 0
transform 1 0 4324 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_47
timestamp 0
transform 1 0 5428 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_59
timestamp 0
transform 1 0 6532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_71
timestamp 0
transform 1 0 7636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 0
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 0
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 0
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 0
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 0
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 0
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 0
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_141
timestamp 0
transform 1 0 14076 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_149
timestamp 0
transform 1 0 14812 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_156
timestamp 0
transform 1 0 15456 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_168
timestamp 0
transform 1 0 16560 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_188
timestamp 0
transform 1 0 18400 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_192
timestamp 0
transform 1 0 18768 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_197
timestamp 0
transform 1 0 19228 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_225
timestamp 0
transform 1 0 21804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_234
timestamp 0
transform 1 0 22632 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_284
timestamp 0
transform 1 0 27232 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_290
timestamp 0
transform 1 0 27784 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_299
timestamp 0
transform 1 0 28612 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_322
timestamp 0
transform 1 0 30728 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_334
timestamp 0
transform 1 0 31832 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_76_356
timestamp 0
transform 1 0 33856 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_365
timestamp 0
transform 1 0 34684 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_377
timestamp 0
transform 1 0 35788 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_76_402
timestamp 0
transform 1 0 38088 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_430
timestamp 0
transform 1 0 40664 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_442
timestamp 0
transform 1 0 41768 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_454
timestamp 0
transform 1 0 42872 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_466
timestamp 0
transform 1 0 43976 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_474
timestamp 0
transform 1 0 44712 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 0
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_489
timestamp 0
transform 1 0 46092 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_7
timestamp 0
transform 1 0 1748 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_19
timestamp 0
transform 1 0 2852 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_31
timestamp 0
transform 1 0 3956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_43
timestamp 0
transform 1 0 5060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 0
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 0
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 0
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 0
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 0
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 0
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 0
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 0
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 0
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 0
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_149
timestamp 0
transform 1 0 14812 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_77_158
timestamp 0
transform 1 0 15640 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_166
timestamp 0
transform 1 0 16376 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_169
timestamp 0
transform 1 0 16652 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_77_174
timestamp 0
transform 1 0 17112 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_193
timestamp 0
transform 1 0 18860 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_201
timestamp 0
transform 1 0 19596 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_207
timestamp 0
transform 1 0 20148 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_211
timestamp 0
transform 1 0 20516 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_215
timestamp 0
transform 1 0 20884 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 0
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_225
timestamp 0
transform 1 0 21804 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_243
timestamp 0
transform 1 0 23460 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_255
timestamp 0
transform 1 0 24564 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_263
timestamp 0
transform 1 0 25300 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_271
timestamp 0
transform 1 0 26036 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 0
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_290
timestamp 0
transform 1 0 27784 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_303
timestamp 0
transform 1 0 28980 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_313
timestamp 0
transform 1 0 29900 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_325
timestamp 0
transform 1 0 31004 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_333
timestamp 0
transform 1 0 31740 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_337
timestamp 0
transform 1 0 32108 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_345
timestamp 0
transform 1 0 32844 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_77_362
timestamp 0
transform 1 0 34408 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_77_384
timestamp 0
transform 1 0 36432 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_77_397
timestamp 0
transform 1 0 37628 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_77_411
timestamp 0
transform 1 0 38916 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_427
timestamp 0
transform 1 0 40388 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_439
timestamp 0
transform 1 0 41492 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 0
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 0
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 0
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 0
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 0
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 0
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 0
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 0
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 0
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 0
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 0
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 0
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 0
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 0
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 0
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 0
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 0
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 0
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 0
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 0
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_141
timestamp 0
transform 1 0 14076 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_149
timestamp 0
transform 1 0 14812 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_176
timestamp 0
transform 1 0 17296 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_188
timestamp 0
transform 1 0 18400 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_197
timestamp 0
transform 1 0 19228 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_205
timestamp 0
transform 1 0 19964 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_223
timestamp 0
transform 1 0 21620 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_232
timestamp 0
transform 1 0 22448 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_236
timestamp 0
transform 1 0 22816 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_242
timestamp 0
transform 1 0 23368 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_250
timestamp 0
transform 1 0 24104 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_253
timestamp 0
transform 1 0 24380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_261
timestamp 0
transform 1 0 25116 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_78_272
timestamp 0
transform 1 0 26128 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_78_282
timestamp 0
transform 1 0 27048 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_291
timestamp 0
transform 1 0 27876 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_297
timestamp 0
transform 1 0 28428 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_303
timestamp 0
transform 1 0 28980 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_309
timestamp 0
transform 1 0 29532 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_317
timestamp 0
transform 1 0 30268 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_334
timestamp 0
transform 1 0 31832 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_338
timestamp 0
transform 1 0 32200 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_347
timestamp 0
transform 1 0 33028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_359
timestamp 0
transform 1 0 34132 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 0
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 0
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 0
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 0
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_401
timestamp 0
transform 1 0 37996 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_409
timestamp 0
transform 1 0 38732 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_414
timestamp 0
transform 1 0 39192 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 0
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 0
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 0
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 0
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 0
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 0
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 0
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_489
timestamp 0
transform 1 0 46092 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 0
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 0
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 0
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 0
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 0
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 0
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 0
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 0
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 0
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 0
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 0
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 0
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 0
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 0
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 0
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 0
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 0
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 0
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_178
timestamp 0
transform 1 0 17480 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_185
timestamp 0
transform 1 0 18124 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_197
timestamp 0
transform 1 0 19228 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_208
timestamp 0
transform 1 0 20240 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_220
timestamp 0
transform 1 0 21344 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 0
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 0
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 0
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 0
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 0
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 0
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 0
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_293
timestamp 0
transform 1 0 28060 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_312
timestamp 0
transform 1 0 29808 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_79_334
timestamp 0
transform 1 0 31832 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_337
timestamp 0
transform 1 0 32108 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_343
timestamp 0
transform 1 0 32660 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_358
timestamp 0
transform 1 0 34040 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_370
timestamp 0
transform 1 0 35144 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_382
timestamp 0
transform 1 0 36248 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_402
timestamp 0
transform 1 0 38088 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_414
timestamp 0
transform 1 0 39192 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_426
timestamp 0
transform 1 0 40296 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_438
timestamp 0
transform 1 0 41400 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_446
timestamp 0
transform 1 0 42136 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 0
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 0
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 0
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_485
timestamp 0
transform 1 0 45724 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_493
timestamp 0
transform 1 0 46460 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 0
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 0
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 0
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 0
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 0
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 0
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 0
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 0
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 0
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 0
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 0
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 0
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 0
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 0
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 0
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 0
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 0
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_165
timestamp 0
transform 1 0 16284 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_171
timestamp 0
transform 1 0 16836 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_175
timestamp 0
transform 1 0 17204 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_197
timestamp 0
transform 1 0 19228 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_205
timestamp 0
transform 1 0 19964 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_213
timestamp 0
transform 1 0 20700 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 0
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_244
timestamp 0
transform 1 0 23552 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_80_275
timestamp 0
transform 1 0 26404 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_283
timestamp 0
transform 1 0 27140 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_293
timestamp 0
transform 1 0 28060 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_303
timestamp 0
transform 1 0 28980 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 0
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_309
timestamp 0
transform 1 0 29532 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_327
timestamp 0
transform 1 0 31188 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_339
timestamp 0
transform 1 0 32292 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_80_355
timestamp 0
transform 1 0 33764 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 0
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_371
timestamp 0
transform 1 0 35236 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_379
timestamp 0
transform 1 0 35972 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_396
timestamp 0
transform 1 0 37536 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_408
timestamp 0
transform 1 0 38640 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 0
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 0
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 0
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 0
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 0
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 0
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 0
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_489
timestamp 0
transform 1 0 46092 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_9
timestamp 0
transform 1 0 1932 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_21
timestamp 0
transform 1 0 3036 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_33
timestamp 0
transform 1 0 4140 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_44
timestamp 0
transform 1 0 5152 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 0
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 0
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 0
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 0
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 0
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 0
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 0
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 0
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 0
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 0
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 0
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 0
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_185
timestamp 0
transform 1 0 18124 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_203
timestamp 0
transform 1 0 19780 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_225
timestamp 0
transform 1 0 21804 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_81_259
timestamp 0
transform 1 0 24932 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_263
timestamp 0
transform 1 0 25300 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_298
timestamp 0
transform 1 0 28520 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_302
timestamp 0
transform 1 0 28888 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_313
timestamp 0
transform 1 0 29900 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 0
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_340
timestamp 0
transform 1 0 32384 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_346
timestamp 0
transform 1 0 32936 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_382
timestamp 0
transform 1 0 36248 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_388
timestamp 0
transform 1 0 36800 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 0
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 0
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 0
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 0
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 0
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 0
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 0
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 0
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 0
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 0
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 0
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_7
timestamp 0
transform 1 0 1748 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_13
timestamp 0
transform 1 0 2300 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_24
timestamp 0
transform 1 0 3312 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_29
timestamp 0
transform 1 0 3772 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_37
timestamp 0
transform 1 0 4508 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_54
timestamp 0
transform 1 0 6072 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_66
timestamp 0
transform 1 0 7176 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_78
timestamp 0
transform 1 0 8280 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 0
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 0
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 0
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 0
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 0
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 0
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 0
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 0
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_165
timestamp 0
transform 1 0 16284 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_173
timestamp 0
transform 1 0 17020 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_213
timestamp 0
transform 1 0 20700 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_218
timestamp 0
transform 1 0 21160 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_82_240
timestamp 0
transform 1 0 23184 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_248
timestamp 0
transform 1 0 23920 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_318
timestamp 0
transform 1 0 30360 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_354
timestamp 0
transform 1 0 33672 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_362
timestamp 0
transform 1 0 34408 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_365
timestamp 0
transform 1 0 34684 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_369
timestamp 0
transform 1 0 35052 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_381
timestamp 0
transform 1 0 36156 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_393
timestamp 0
transform 1 0 37260 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_405
timestamp 0
transform 1 0 38364 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_417
timestamp 0
transform 1 0 39468 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 0
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 0
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 0
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 0
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 0
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 0
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 0
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_489
timestamp 0
transform 1 0 46092 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_493
timestamp 0
transform 1 0 46460 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_3
timestamp 0
transform 1 0 1380 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_11
timestamp 0
transform 1 0 2116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_23
timestamp 0
transform 1 0 3220 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_29
timestamp 0
transform 1 0 3772 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_41
timestamp 0
transform 1 0 4876 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_49
timestamp 0
transform 1 0 5612 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 0
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_69
timestamp 0
transform 1 0 7452 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_77
timestamp 0
transform 1 0 8188 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_83_83
timestamp 0
transform 1 0 8740 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_85
timestamp 0
transform 1 0 8924 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_97
timestamp 0
transform 1 0 10028 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 0
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 0
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 0
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_125
timestamp 0
transform 1 0 12604 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_133
timestamp 0
transform 1 0 13340 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_139
timestamp 0
transform 1 0 13892 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_141
timestamp 0
transform 1 0 14076 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_153
timestamp 0
transform 1 0 15180 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 0
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 0
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_169
timestamp 0
transform 1 0 16652 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_175
timestamp 0
transform 1 0 17204 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_180
timestamp 0
transform 1 0 17664 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_184
timestamp 0
transform 1 0 18032 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_83_201
timestamp 0
transform 1 0 19596 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_211
timestamp 0
transform 1 0 20516 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 0
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_225
timestamp 0
transform 1 0 21804 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_233
timestamp 0
transform 1 0 22540 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_238
timestamp 0
transform 1 0 23000 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_250
timestamp 0
transform 1 0 24104 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_253
timestamp 0
transform 1 0 24380 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_265
timestamp 0
transform 1 0 25484 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_277
timestamp 0
transform 1 0 26588 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_83_281
timestamp 0
transform 1 0 26956 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_287
timestamp 0
transform 1 0 27508 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_299
timestamp 0
transform 1 0 28612 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_303
timestamp 0
transform 1 0 28980 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_309
timestamp 0
transform 1 0 29532 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_321
timestamp 0
transform 1 0 30636 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_333
timestamp 0
transform 1 0 31740 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_343
timestamp 0
transform 1 0 32660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_355
timestamp 0
transform 1 0 33764 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_359
timestamp 0
transform 1 0 34132 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_365
timestamp 0
transform 1 0 34684 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_377
timestamp 0
transform 1 0 35788 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 0
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 0
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 0
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_405
timestamp 0
transform 1 0 38364 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_412
timestamp 0
transform 1 0 39008 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_421
timestamp 0
transform 1 0 39836 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_433
timestamp 0
transform 1 0 40940 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_443
timestamp 0
transform 1 0 41860 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 0
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_449
timestamp 0
transform 1 0 42412 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_457
timestamp 0
transform 1 0 43148 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_468
timestamp 0
transform 1 0 44160 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_83_477
timestamp 0
transform 1 0 44988 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_483
timestamp 0
transform 1 0 45540 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 0
transform 1 0 45908 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 0
transform 1 0 43240 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 0
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 0
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform 1 0 39376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 0
transform 1 0 42412 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 0
transform 1 0 45908 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 0
transform 1 0 5888 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 0
transform 1 0 1380 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 0
transform 1 0 24564 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 0
transform 1 0 1380 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 0
transform 1 0 45908 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 0
transform 1 0 45632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 0
transform 1 0 27140 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 0
transform 1 0 45632 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 0
transform 1 0 1380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 0
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 0
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 0
transform 1 0 46552 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 0
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 0
transform 1 0 46552 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 0
transform 1 0 46460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 0
transform 1 0 8464 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 0
transform 1 0 45908 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 0
transform 1 0 9108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 0
transform 1 0 46460 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 0
transform 1 0 25208 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 0
transform 1 0 38732 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 0
transform 1 0 46460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 0
transform 1 0 36156 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 0
transform 1 0 46276 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 0
transform 1 0 46460 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 0
transform 1 0 46460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 0
transform 1 0 46460 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 0
transform 1 0 46460 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 0
transform 1 0 46276 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 0
transform 1 0 46460 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 0
transform 1 0 46460 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output46
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 0
transform 1 0 46460 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 0
transform 1 0 1380 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 0
transform 1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output50
timestamp 0
transform 1 0 1564 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 0
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 0
transform 1 0 29072 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 0
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output54
timestamp 0
transform 1 0 30176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 0
transform 1 0 46460 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 0
transform 1 0 15548 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 0
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 0
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 0
transform 1 0 34224 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 0
transform 1 0 1380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 0
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output63
timestamp 0
transform 1 0 1380 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 0
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 0
transform 1 0 17296 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 0
transform 1 0 46460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 0
transform 1 0 46460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 0
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output69
timestamp 0
transform 1 0 1380 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 0
transform 1 0 12972 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 0
transform 1 0 22632 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 0
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 0
transform 1 0 20148 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 0
transform 1 0 32108 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 0
transform 1 0 41308 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 0
transform 1 0 3312 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 0
transform 1 0 10396 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 0
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 0
transform 1 0 1380 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 47104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 47104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 47104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 47104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 47104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 47104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 47104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 47104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 47104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 47104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 47104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 47104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 47104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 47104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 47104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 47104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 47104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 47104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 47104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 47104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 47104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 47104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 47104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 47104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 47104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 47104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 47104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 0
transform -1 0 47104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 0
transform -1 0 47104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 0
transform -1 0 47104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 0
transform -1 0 47104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 0
transform -1 0 47104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 0
transform -1 0 47104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 0
transform -1 0 47104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 0
transform -1 0 47104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 0
transform -1 0 47104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 0
transform -1 0 47104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 0
transform -1 0 47104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 0
transform -1 0 47104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 0
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 0
transform -1 0 47104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 0
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 0
transform -1 0 47104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 0
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 0
transform -1 0 47104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 0
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 0
transform -1 0 47104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 0
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 0
transform -1 0 47104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 0
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 0
transform -1 0 47104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 0
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 0
transform -1 0 47104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 0
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 0
transform -1 0 47104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 0
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 0
transform -1 0 47104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 0
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 0
transform -1 0 47104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 0
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 0
transform -1 0 47104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 0
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 0
transform -1 0 47104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 0
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 0
transform -1 0 47104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 0
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 0
transform -1 0 47104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 0
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 0
transform -1 0 47104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 0
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 0
transform -1 0 47104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 0
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 0
transform -1 0 47104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 0
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 0
transform -1 0 47104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 0
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 0
transform -1 0 47104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 0
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 0
transform -1 0 47104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 0
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 0
transform -1 0 47104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 0
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 0
transform -1 0 47104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 0
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 0
transform -1 0 47104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 0
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 0
transform -1 0 47104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 0
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 0
transform -1 0 47104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 0
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 0
transform -1 0 47104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 0
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 0
transform -1 0 47104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 0
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 0
transform -1 0 47104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 0
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 0
transform -1 0 47104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 0
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 0
transform -1 0 47104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 0
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 0
transform -1 0 47104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 0
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 0
transform -1 0 47104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 0
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 0
transform -1 0 47104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 0
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 0
transform -1 0 47104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 0
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 0
transform -1 0 47104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 0
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 0
transform -1 0 47104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 0
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 0
transform -1 0 47104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 0
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 0
transform -1 0 47104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 0
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 0
transform -1 0 47104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 0
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 0
transform -1 0 47104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 0
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 0
transform -1 0 47104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 0
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 0
transform -1 0 47104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 0
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 0
transform -1 0 47104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 0
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 0
transform -1 0 47104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 0
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 0
transform -1 0 47104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 0
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 0
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 0
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 0
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 0
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 0
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 0
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 0
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 0
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 0
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 0
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 0
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 0
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 0
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 0
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 0
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 0
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 0
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 0
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 0
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 0
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 0
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 0
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 0
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 0
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 0
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 0
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 0
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 0
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 0
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 0
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 0
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 0
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 0
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 0
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 0
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 0
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 0
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 0
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 0
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 0
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 0
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 0
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 0
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 0
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 0
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 0
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 0
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 0
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 0
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 0
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 0
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 0
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 0
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 0
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 0
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 0
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 0
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 0
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 0
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 0
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 0
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 0
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 0
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 0
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 0
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 0
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 0
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 0
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 0
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 0
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 0
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 0
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 0
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 0
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 0
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 0
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 0
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 0
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 0
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 0
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 0
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 0
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 0
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 0
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 0
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 0
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 0
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 0
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 0
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 0
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 0
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 0
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 0
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 0
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 0
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 0
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 0
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 0
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 0
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 0
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 0
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 0
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 0
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 0
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 0
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 0
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 0
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 0
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 0
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 0
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 0
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 0
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 0
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 0
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 0
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 0
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 0
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 0
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 0
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 0
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 0
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 0
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 0
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 0
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 0
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 0
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 0
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 0
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 0
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 0
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 0
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 0
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 0
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 0
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 0
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 0
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 0
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 0
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 0
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 0
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 0
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 0
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 0
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 0
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 0
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 0
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 0
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 0
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 0
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 0
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 0
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 0
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 0
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 0
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 0
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 0
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 0
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 0
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 0
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 0
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 0
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 0
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 0
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 0
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 0
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 0
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 0
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 0
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 0
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 0
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 0
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 0
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 0
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 0
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 0
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 0
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 0
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 0
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 0
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 0
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 0
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 0
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 0
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 0
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 0
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 0
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 0
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 0
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 0
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 0
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 0
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 0
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 0
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 0
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 0
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 0
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 0
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 0
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 0
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 0
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 0
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 0
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 0
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 0
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 0
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 0
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 0
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 0
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 0
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 0
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 0
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 0
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 0
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 0
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 0
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 0
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 0
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 0
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 0
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 0
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 0
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 0
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 0
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 0
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 0
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 0
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 0
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 0
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 0
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 0
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 0
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 0
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 0
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 0
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 0
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 0
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 0
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 0
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 0
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 0
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 0
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 0
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 0
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 0
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 0
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 0
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 0
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 0
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 0
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 0
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 0
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 0
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 0
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 0
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 0
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 0
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 0
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 0
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 0
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 0
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 0
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 0
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 0
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 0
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 0
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 0
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 0
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 0
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 0
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 0
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 0
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 0
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 0
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 0
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 0
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 0
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 0
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 0
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 0
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 0
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 0
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 0
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 0
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 0
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 0
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 0
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 0
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 0
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 0
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 0
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 0
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 0
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 0
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 0
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 0
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 0
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 0
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 0
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 0
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 0
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 0
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 0
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 0
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 0
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 0
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 0
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 0
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 0
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 0
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 0
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 0
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 0
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 0
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 0
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 0
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 0
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 0
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 0
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 0
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 0
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 0
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 0
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 0
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 0
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 0
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 0
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 0
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 0
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 0
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 0
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 0
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 0
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 0
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 0
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 0
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 0
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 0
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 0
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 0
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 0
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 0
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 0
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 0
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 0
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 0
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 0
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 0
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 0
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 0
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 0
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 0
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 0
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 0
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 0
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 0
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 0
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 0
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 0
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 0
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 0
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 0
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 0
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 0
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 0
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 0
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 0
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 0
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 0
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 0
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 0
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 0
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 0
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 0
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 0
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 0
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 0
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 0
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 0
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 0
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 0
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 0
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 0
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 0
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 0
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 0
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 0
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 0
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 0
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 0
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 0
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 0
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 0
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 0
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 0
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 0
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 0
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 0
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 0
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 0
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 0
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 0
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 0
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 0
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 0
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 0
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 0
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 0
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 0
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 0
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 0
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 0
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 0
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 0
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 0
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 0
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 0
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 0
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 0
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 0
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 0
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 0
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 0
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 0
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 0
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 0
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 0
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 0
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 0
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 0
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 0
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 0
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 0
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 0
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 0
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 0
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 0
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 0
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 0
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 0
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 0
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 0
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 0
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 0
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 0
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 0
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 0
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 0
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 0
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 0
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 0
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 0
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 0
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 0
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 0
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 0
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 0
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 0
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 0
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 0
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 0
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 0
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 0
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 0
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 0
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 0
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 0
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 0
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 0
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 0
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 0
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 0
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 0
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 0
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 0
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 0
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 0
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 0
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 0
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 0
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 0
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 0
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 0
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 0
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 0
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 0
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 0
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 0
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 0
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 0
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 0
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 0
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 0
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 0
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 0
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 0
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 0
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 0
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 0
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 0
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 0
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 0
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 0
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 0
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 0
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 0
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 0
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 0
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 0
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 0
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 0
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 0
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 0
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 0
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 0
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 0
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 0
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 0
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 0
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 0
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 0
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 0
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 0
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 0
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 0
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 0
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 0
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 0
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 0
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 0
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 0
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 0
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 0
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 0
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 0
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 0
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 0
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 0
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 0
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 0
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 0
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 0
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 0
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 0
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 0
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 0
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 0
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 0
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 0
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 0
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 0
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 0
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 0
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 0
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 0
transform 1 0 3680 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 0
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 0
transform 1 0 8832 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 0
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 0
transform 1 0 13984 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 0
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 0
transform 1 0 19136 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 0
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 0
transform 1 0 24288 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 0
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 0
transform 1 0 29440 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 0
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 0
transform 1 0 34592 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 0
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 0
transform 1 0 39744 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 0
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 0
transform 1 0 44896 0 -1 47872
box -38 -48 130 592
<< labels >>
rlabel metal1 s 24104 47872 24104 47872 4 VGND
rlabel metal1 s 24104 47328 24104 47328 4 VPWR
rlabel metal2 s 45954 8313 45954 8313 4 D_R_data[0]
rlabel metal2 s 43286 48671 43286 48671 4 D_R_data[10]
rlabel metal3 s 820 24548 820 24548 4 D_R_data[11]
rlabel metal3 s 1096 12308 1096 12308 4 D_R_data[12]
rlabel metal2 s 13570 1588 13570 1588 4 D_R_data[13]
rlabel metal2 s 23230 1588 23230 1588 4 D_R_data[14]
rlabel metal2 s 39330 1588 39330 1588 4 D_R_data[15]
rlabel metal2 s 41906 1588 41906 1588 4 D_R_data[1]
rlabel metal3 s 45954 47651 45954 47651 4 D_R_data[2]
rlabel metal2 s 6026 48705 6026 48705 4 D_R_data[3]
rlabel metal3 s 820 32028 820 32028 4 D_R_data[4]
rlabel metal2 s 24610 48671 24610 48671 4 D_R_data[5]
rlabel metal3 s 820 29308 820 29308 4 D_R_data[6]
rlabel metal2 s 45494 1615 45494 1615 4 D_R_data[7]
rlabel metal2 s 46414 1554 46414 1554 4 D_R_data[8]
rlabel metal2 s 27278 48705 27278 48705 4 D_R_data[9]
rlabel metal1 s 36248 47770 36248 47770 4 D_W_data[0]
rlabel metal3 s 46690 5525 46690 5525 4 D_W_data[10]
rlabel metal3 s 46690 32725 46690 32725 4 D_W_data[11]
rlabel metal3 s 1142 6868 1142 6868 4 D_W_data[12]
rlabel metal2 s 46690 15793 46690 15793 4 D_W_data[13]
rlabel metal3 s 46690 35445 46690 35445 4 D_W_data[14]
rlabel metal3 s 820 2108 820 2108 4 D_W_data[15]
rlabel metal2 s 46690 42993 46690 42993 4 D_W_data[1]
rlabel metal2 s 46782 17697 46782 17697 4 D_W_data[2]
rlabel metal2 s 46690 29631 46690 29631 4 D_W_data[3]
rlabel metal2 s 46690 13073 46690 13073 4 D_W_data[4]
rlabel metal3 s 1142 9588 1142 9588 4 D_W_data[5]
rlabel metal2 s 46690 40273 46690 40273 4 D_W_data[6]
rlabel metal3 s 820 41548 820 41548 4 D_W_data[7]
rlabel metal3 s 912 46988 912 46988 4 D_W_data[8]
rlabel metal3 s 1234 49028 1234 49028 4 D_W_data[9]
rlabel metal2 s 4554 1520 4554 1520 4 D_addr[0]
rlabel metal1 s 29164 47770 29164 47770 4 D_addr[1]
rlabel metal2 s 18722 1520 18722 1520 4 D_addr[2]
rlabel metal2 s 30314 1095 30314 1095 4 D_addr[3]
rlabel metal2 s 46690 37553 46690 37553 4 D_addr[4]
rlabel metal2 s 15778 48739 15778 48739 4 D_addr[5]
rlabel metal1 s 1472 19482 1472 19482 4 D_addr[6]
rlabel metal2 s 11638 1520 11638 1520 4 D_addr[7]
rlabel metal2 s 37398 1520 37398 1520 4 D_rd
rlabel metal2 s 34454 48739 34454 48739 4 D_wr
rlabel metal3 s 820 39508 820 39508 4 I_addr[0]
rlabel metal2 s 27738 1520 27738 1520 4 I_addr[10]
rlabel metal1 s 1472 46682 1472 46682 4 I_addr[11]
rlabel metal2 s 44482 1520 44482 1520 4 I_addr[12]
rlabel metal1 s 17480 47770 17480 47770 4 I_addr[13]
rlabel metal2 s 46690 10353 46690 10353 4 I_addr[14]
rlabel metal2 s 46690 20519 46690 20519 4 I_addr[15]
rlabel metal2 s 34822 1520 34822 1520 4 I_addr[1]
rlabel metal3 s 1142 34068 1142 34068 4 I_addr[2]
rlabel metal2 s 13202 48739 13202 48739 4 I_addr[3]
rlabel metal1 s 22724 47770 22724 47770 4 I_addr[4]
rlabel metal3 s 820 4828 820 4828 4 I_addr[5]
rlabel metal2 s 46 1792 46 1792 4 I_addr[6]
rlabel metal3 s 820 26588 820 26588 4 I_addr[7]
rlabel metal1 s 20194 47770 20194 47770 4 I_addr[8]
rlabel metal1 s 32062 47770 32062 47770 4 I_addr[9]
rlabel metal2 s 45862 48671 45862 48671 4 I_data[0]
rlabel metal3 s 820 36788 820 36788 4 I_data[10]
rlabel metal2 s 6486 1588 6486 1588 4 I_data[11]
rlabel metal2 s 1978 1588 1978 1588 4 I_data[12]
rlabel metal1 s 47242 47022 47242 47022 4 I_data[13]
rlabel metal3 s 820 17068 820 17068 4 I_data[14]
rlabel metal2 s 20654 1554 20654 1554 4 I_data[15]
rlabel metal2 s 46782 45203 46782 45203 4 I_data[1]
rlabel metal2 s 46598 2907 46598 2907 4 I_data[2]
rlabel metal2 s 8694 48671 8694 48671 4 I_data[3]
rlabel metal3 s 45954 25245 45954 25245 4 I_data[4]
rlabel metal2 s 9062 1588 9062 1588 4 I_data[5]
rlabel metal2 s 16146 1588 16146 1588 4 I_data[6]
rlabel metal3 s 820 21828 820 21828 4 I_data[7]
rlabel metal2 s 46598 27999 46598 27999 4 I_data[8]
rlabel metal2 s 25162 1588 25162 1588 4 I_data[9]
rlabel metal1 s 41492 47770 41492 47770 4 I_rd
rlabel metal1 s 11178 20910 11178 20910 4 _0000_
rlabel metal1 s 9936 19346 9936 19346 4 _0001_
rlabel metal2 s 14122 24412 14122 24412 4 _0002_
rlabel metal1 s 12236 14382 12236 14382 4 _0003_
rlabel metal2 s 21298 32853 21298 32853 4 _0004_
rlabel metal1 s 20608 40902 20608 40902 4 _0005_
rlabel metal1 s 19412 44166 19412 44166 4 _0006_
rlabel metal1 s 21574 17238 21574 17238 4 _0007_
rlabel metal1 s 8862 24854 8862 24854 4 _0008_
rlabel metal2 s 8321 20502 8321 20502 4 _0009_
rlabel metal1 s 7626 24786 7626 24786 4 _0010_
rlabel metal2 s 8413 27030 8413 27030 4 _0011_
rlabel metal2 s 19545 41582 19545 41582 4 _0012_
rlabel metal1 s 18982 41174 18982 41174 4 _0013_
rlabel metal1 s 17280 44438 17280 44438 4 _0014_
rlabel metal1 s 17940 45322 17940 45322 4 _0015_
rlabel metal1 s 30942 39338 30942 39338 4 _0016_
rlabel metal2 s 12185 32878 12185 32878 4 _0017_
rlabel metal1 s 11484 40086 11484 40086 4 _0018_
rlabel metal2 s 30861 30294 30861 30294 4 _0019_
rlabel metal1 s 29808 37978 29808 37978 4 _0020_
rlabel metal1 s 32092 28118 32092 28118 4 _0021_
rlabel metal2 s 34086 16354 34086 16354 4 _0022_
rlabel metal1 s 33212 24922 33212 24922 4 _0023_
rlabel metal1 s 22995 17238 22995 17238 4 _0024_
rlabel metal1 s 33897 10710 33897 10710 4 _0025_
rlabel metal2 s 33437 19822 33437 19822 4 _0026_
rlabel metal2 s 22862 10914 22862 10914 4 _0027_
rlabel metal1 s 32184 3094 32184 3094 4 _0028_
rlabel metal1 s 32384 8602 32384 8602 4 _0029_
rlabel metal2 s 21109 3502 21109 3502 4 _0030_
rlabel metal2 s 24978 3298 24978 3298 4 _0031_
rlabel metal1 s 31839 38250 31839 38250 4 _0032_
rlabel metal2 s 13386 34374 13386 34374 4 _0033_
rlabel metal1 s 12611 40426 12611 40426 4 _0034_
rlabel metal1 s 32466 32810 32466 32810 4 _0035_
rlabel metal1 s 30022 37162 30022 37162 4 _0036_
rlabel metal2 s 33902 28934 33902 28934 4 _0037_
rlabel metal2 s 34633 16150 34633 16150 4 _0038_
rlabel metal1 s 35548 24174 35548 24174 4 _0039_
rlabel metal1 s 23271 19822 23271 19822 4 _0040_
rlabel metal1 s 34904 13294 34904 13294 4 _0041_
rlabel metal1 s 35875 21590 35875 21590 4 _0042_
rlabel metal2 s 24840 12308 24840 12308 4 _0043_
rlabel metal1 s 32460 4182 32460 4182 4 _0044_
rlabel metal1 s 34362 6630 34362 6630 4 _0045_
rlabel metal1 s 22627 3094 22627 3094 4 _0046_
rlabel metal1 s 26164 3502 26164 3502 4 _0047_
rlabel metal2 s 30590 40290 30590 40290 4 _0048_
rlabel metal2 s 12093 32402 12093 32402 4 _0049_
rlabel metal1 s 10794 40426 10794 40426 4 _0050_
rlabel metal2 s 30861 30702 30861 30702 4 _0051_
rlabel metal2 s 29578 35462 29578 35462 4 _0052_
rlabel metal2 s 32057 26350 32057 26350 4 _0053_
rlabel metal1 s 32966 16490 32966 16490 4 _0054_
rlabel metal2 s 32241 24174 32241 24174 4 _0055_
rlabel metal2 s 22494 18530 22494 18530 4 _0056_
rlabel metal1 s 32972 11118 32972 11118 4 _0057_
rlabel metal2 s 32241 20910 32241 20910 4 _0058_
rlabel metal2 s 22034 12002 22034 12002 4 _0059_
rlabel metal2 s 30769 3502 30769 3502 4 _0060_
rlabel metal1 s 32092 7446 32092 7446 4 _0061_
rlabel metal2 s 19821 3026 19821 3026 4 _0062_
rlabel metal2 s 23777 3094 23777 3094 4 _0063_
rlabel metal2 s 22121 41174 22121 41174 4 _0064_
rlabel metal1 s 16544 34646 16544 34646 4 _0065_
rlabel metal1 s 14582 40154 14582 40154 4 _0066_
rlabel metal1 s 27273 30226 27273 30226 4 _0067_
rlabel metal2 s 26266 40290 26266 40290 4 _0068_
rlabel metal2 s 26634 28322 26634 28322 4 _0069_
rlabel metal1 s 32154 20536 32154 20536 4 _0070_
rlabel metal2 s 30861 24854 30861 24854 4 _0071_
rlabel metal2 s 18722 18530 18722 18530 4 _0072_
rlabel metal2 s 32430 15878 32430 15878 4 _0073_
rlabel metal1 s 22397 21930 22397 21930 4 _0074_
rlabel metal2 s 20286 13702 20286 13702 4 _0075_
rlabel metal2 s 17250 4998 17250 4998 4 _0076_
rlabel metal1 s 18982 6358 18982 6358 4 _0077_
rlabel metal1 s 16774 3434 16774 3434 4 _0078_
rlabel metal1 s 18850 4114 18850 4114 4 _0079_
rlabel metal1 s 24318 41514 24318 41514 4 _0080_
rlabel metal2 s 18354 34578 18354 34578 4 _0081_
rlabel metal2 s 16601 40494 16601 40494 4 _0082_
rlabel metal1 s 29752 31790 29752 31790 4 _0083_
rlabel metal1 s 27446 40426 27446 40426 4 _0084_
rlabel metal2 s 30038 29274 30038 29274 4 _0085_
rlabel metal2 s 31142 16354 31142 16354 4 _0086_
rlabel metal2 s 30033 21998 30033 21998 4 _0087_
rlabel metal1 s 26353 19414 26353 19414 4 _0088_
rlabel metal2 s 31234 10914 31234 10914 4 _0089_
rlabel metal2 s 27830 21794 27830 21794 4 _0090_
rlabel metal1 s 26940 11798 26940 11798 4 _0091_
rlabel metal1 s 28975 4114 28975 4114 4 _0092_
rlabel metal1 s 30401 6358 30401 6358 4 _0093_
rlabel metal1 s 14490 3706 14490 3706 4 _0094_
rlabel metal2 s 24518 6086 24518 6086 4 _0095_
rlabel metal1 s 6302 37298 6302 37298 4 _0096_
rlabel metal1 s 1732 32470 1732 32470 4 _0097_
rlabel metal1 s 6562 34646 6562 34646 4 _0098_
rlabel metal2 s 6665 31790 6665 31790 4 _0099_
rlabel metal2 s 3634 35258 3634 35258 4 _0100_
rlabel metal1 s 1973 26282 1973 26282 4 _0101_
rlabel metal1 s 2065 20502 2065 20502 4 _0102_
rlabel metal2 s 2065 23086 2065 23086 4 _0103_
rlabel metal1 s 6394 18360 6394 18360 4 _0104_
rlabel metal1 s 5826 15402 5826 15402 4 _0105_
rlabel metal2 s 7498 21318 7498 21318 4 _0106_
rlabel metal1 s 2438 16762 2438 16762 4 _0107_
rlabel metal1 s 4135 12886 4135 12886 4 _0108_
rlabel metal1 s 6194 9962 6194 9962 4 _0109_
rlabel metal1 s 9782 9962 9782 9962 4 _0110_
rlabel metal1 s 9287 12886 9287 12886 4 _0111_
rlabel metal2 s 6026 38114 6026 38114 4 _0112_
rlabel metal2 s 2065 32878 2065 32878 4 _0113_
rlabel metal2 s 6849 35054 6849 35054 4 _0114_
rlabel metal1 s 6711 32470 6711 32470 4 _0115_
rlabel metal1 s 2146 35734 2146 35734 4 _0116_
rlabel metal2 s 1973 27438 1973 27438 4 _0117_
rlabel metal2 s 1973 19822 1973 19822 4 _0118_
rlabel metal1 s 2116 22202 2116 22202 4 _0119_
rlabel metal2 s 6670 18530 6670 18530 4 _0120_
rlabel metal1 s 6516 15062 6516 15062 4 _0121_
rlabel metal1 s 7206 21930 7206 21930 4 _0122_
rlabel metal1 s 2714 15674 2714 15674 4 _0123_
rlabel metal2 s 4186 12002 4186 12002 4 _0124_
rlabel metal1 s 6516 9622 6516 9622 4 _0125_
rlabel metal1 s 9384 10234 9384 10234 4 _0126_
rlabel metal1 s 9384 11322 9384 11322 4 _0127_
rlabel metal2 s 7401 38318 7401 38318 4 _0128_
rlabel metal1 s 3986 33558 3986 33558 4 _0129_
rlabel metal2 s 8321 34578 8321 34578 4 _0130_
rlabel metal2 s 8970 32198 8970 32198 4 _0131_
rlabel metal2 s 4089 37230 4089 37230 4 _0132_
rlabel metal2 s 3174 27846 3174 27846 4 _0133_
rlabel metal1 s 3905 19414 3905 19414 4 _0134_
rlabel metal1 s 4411 21998 4411 21998 4 _0135_
rlabel metal2 s 8602 18258 8602 18258 4 _0136_
rlabel metal1 s 7988 15062 7988 15062 4 _0137_
rlabel metal1 s 8908 23018 8908 23018 4 _0138_
rlabel metal1 s 3818 14586 3818 14586 4 _0139_
rlabel metal2 s 5653 11118 5653 11118 4 _0140_
rlabel metal2 s 7769 7446 7769 7446 4 _0141_
rlabel metal1 s 10350 6970 10350 6970 4 _0142_
rlabel metal1 s 10207 13226 10207 13226 4 _0143_
rlabel metal2 s 9333 38318 9333 38318 4 _0144_
rlabel metal1 s 3721 30294 3721 30294 4 _0145_
rlabel metal1 s 9690 35734 9690 35734 4 _0146_
rlabel metal1 s 9322 32810 9322 32810 4 _0147_
rlabel metal1 s 4135 37910 4135 37910 4 _0148_
rlabel metal1 s 3992 25262 3992 25262 4 _0149_
rlabel metal2 s 5382 20162 5382 20162 4 _0150_
rlabel metal1 s 4814 22678 4814 22678 4 _0151_
rlabel metal1 s 9966 18326 9966 18326 4 _0152_
rlabel metal2 s 10718 16354 10718 16354 4 _0153_
rlabel metal1 s 10248 20910 10248 20910 4 _0154_
rlabel metal2 s 3910 18054 3910 18054 4 _0155_
rlabel metal2 s 6946 13464 6946 13464 4 _0156_
rlabel metal1 s 7390 7786 7390 7786 4 _0157_
rlabel metal2 s 10529 7854 10529 7854 4 _0158_
rlabel metal1 s 11806 13226 11806 13226 4 _0159_
rlabel metal1 s 20143 38250 20143 38250 4 _0160_
rlabel metal1 s 15762 29546 15762 29546 4 _0161_
rlabel metal1 s 13922 38250 13922 38250 4 _0162_
rlabel metal1 s 23184 33082 23184 33082 4 _0163_
rlabel metal2 s 22126 36006 22126 36006 4 _0164_
rlabel metal2 s 21569 27438 21569 27438 4 _0165_
rlabel metal2 s 13018 20706 13018 20706 4 _0166_
rlabel metal1 s 14393 23766 14393 23766 4 _0167_
rlabel metal2 s 12829 18734 12829 18734 4 _0168_
rlabel metal1 s 12082 16150 12082 16150 4 _0169_
rlabel metal1 s 13248 22202 13248 22202 4 _0170_
rlabel metal2 s 12558 15266 12558 15266 4 _0171_
rlabel metal2 s 14577 12818 14577 12818 4 _0172_
rlabel metal1 s 13473 7786 13473 7786 4 _0173_
rlabel metal1 s 13565 7446 13565 7446 4 _0174_
rlabel metal1 s 14296 10030 14296 10030 4 _0175_
rlabel metal2 s 19361 37910 19361 37910 4 _0176_
rlabel metal1 s 15302 29206 15302 29206 4 _0177_
rlabel metal2 s 13841 37842 13841 37842 4 _0178_
rlabel metal2 s 22126 31994 22126 31994 4 _0179_
rlabel metal1 s 21012 35054 21012 35054 4 _0180_
rlabel metal1 s 20235 27370 20235 27370 4 _0181_
rlabel metal2 s 14766 20706 14766 20706 4 _0182_
rlabel metal1 s 16038 24106 16038 24106 4 _0183_
rlabel metal1 s 13749 18326 13749 18326 4 _0184_
rlabel metal2 s 14761 16082 14761 16082 4 _0185_
rlabel metal1 s 15865 23086 15865 23086 4 _0186_
rlabel metal1 s 14888 15402 14888 15402 4 _0187_
rlabel metal2 s 15037 13294 15037 13294 4 _0188_
rlabel metal1 s 16008 7514 16008 7514 4 _0189_
rlabel metal1 s 15072 8534 15072 8534 4 _0190_
rlabel metal2 s 15221 10710 15221 10710 4 _0191_
rlabel metal1 s 24502 41174 24502 41174 4 _0192_
rlabel metal1 s 19448 32878 19448 32878 4 _0193_
rlabel metal2 s 18630 40732 18630 40732 4 _0194_
rlabel metal2 s 29210 32198 29210 32198 4 _0195_
rlabel metal1 s 28561 40086 28561 40086 4 _0196_
rlabel metal1 s 29026 28186 29026 28186 4 _0197_
rlabel metal1 s 32123 18632 32123 18632 4 _0198_
rlabel metal2 s 30217 23086 30217 23086 4 _0199_
rlabel metal1 s 28147 19414 28147 19414 4 _0200_
rlabel metal1 s 32052 13294 32052 13294 4 _0201_
rlabel metal2 s 28750 21726 28750 21726 4 _0202_
rlabel metal1 s 27692 12682 27692 12682 4 _0203_
rlabel metal2 s 29205 3026 29205 3026 4 _0204_
rlabel metal1 s 30631 5678 30631 5678 4 _0205_
rlabel metal1 s 14428 3094 14428 3094 4 _0206_
rlabel metal2 s 26542 6562 26542 6562 4 _0207_
rlabel metal2 s 22126 38318 22126 38318 4 _0208_
rlabel metal1 s 18768 28730 18768 28730 4 _0209_
rlabel metal1 s 16872 35666 16872 35666 4 _0210_
rlabel metal1 s 24191 30634 24191 30634 4 _0211_
rlabel metal2 s 23961 34578 23961 34578 4 _0212_
rlabel metal1 s 24600 27438 24600 27438 4 _0213_
rlabel metal1 s 17142 20502 17142 20502 4 _0214_
rlabel metal1 s 18625 24786 18625 24786 4 _0215_
rlabel metal2 s 16330 17986 16330 17986 4 _0216_
rlabel metal2 s 17250 16354 17250 16354 4 _0217_
rlabel metal1 s 17694 23018 17694 23018 4 _0218_
rlabel metal2 s 17245 15062 17245 15062 4 _0219_
rlabel metal1 s 16928 12954 16928 12954 4 _0220_
rlabel metal1 s 19304 6698 19304 6698 4 _0221_
rlabel metal1 s 17112 5882 17112 5882 4 _0222_
rlabel metal1 s 17429 10030 17429 10030 4 _0223_
rlabel metal1 s 34541 46614 34541 46614 4 _0224_
rlabel metal2 s 36381 45934 36381 45934 4 _0225_
rlabel metal2 s 30861 42194 30861 42194 4 _0226_
rlabel metal1 s 32200 46682 32200 46682 4 _0227_
rlabel metal2 s 36570 42942 36570 42942 4 _0228_
rlabel metal1 s 13524 41786 13524 41786 4 _0229_
rlabel metal2 s 13294 42466 13294 42466 4 _0230_
rlabel metal2 s 2806 25058 2806 25058 4 _0231_
rlabel metal1 s 7958 28730 7958 28730 4 _0232_
rlabel metal1 s 11254 24106 11254 24106 4 _0233_
rlabel metal2 s 2065 30702 2065 30702 4 _0234_
rlabel metal1 s 4538 28458 4538 28458 4 _0235_
rlabel metal1 s 2146 40426 2146 40426 4 _0236_
rlabel metal2 s 38778 43554 38778 43554 4 _0237_
rlabel metal1 s 2525 17578 2525 17578 4 _0238_
rlabel metal1 s 20649 41174 20649 41174 4 _0239_
rlabel metal2 s 25530 43554 25530 43554 4 _0240_
rlabel metal1 s 30222 46138 30222 46138 4 _0241_
rlabel metal1 s 27457 42670 27457 42670 4 _0242_
rlabel metal1 s 27324 46138 27324 46138 4 _0243_
rlabel metal2 s 22402 46818 22402 46818 4 _0244_
rlabel metal2 s 22586 43078 22586 43078 4 _0245_
rlabel metal2 s 20557 43758 20557 43758 4 _0246_
rlabel metal1 s 20695 46614 20695 46614 4 _0247_
rlabel metal2 s 25346 46342 25346 46342 4 _0248_
rlabel metal1 s 32517 42262 32517 42262 4 _0256_
rlabel metal1 s 34684 36346 34684 36346 4 _0257_
rlabel metal1 s 14388 31790 14388 31790 4 _0258_
rlabel metal1 s 12650 38216 12650 38216 4 _0259_
rlabel metal2 s 33994 31518 33994 31518 4 _0260_
rlabel metal1 s 31885 33898 31885 33898 4 _0261_
rlabel metal1 s 35266 27370 35266 27370 4 _0262_
rlabel metal2 s 35737 18734 35737 18734 4 _0263_
rlabel metal1 s 36294 23290 36294 23290 4 _0264_
rlabel metal2 s 36662 18530 36662 18530 4 _0265_
rlabel metal2 s 36110 13634 36110 13634 4 _0266_
rlabel metal1 s 37198 21590 37198 21590 4 _0267_
rlabel metal1 s 35726 13974 35726 13974 4 _0268_
rlabel metal2 s 35093 5270 35093 5270 4 _0269_
rlabel metal1 s 35266 7786 35266 7786 4 _0270_
rlabel metal1 s 21482 5304 21482 5304 4 _0271_
rlabel metal1 s 27508 3978 27508 3978 4 _0272_
rlabel metal1 s 24671 38216 24671 38216 4 _0273_
rlabel metal1 s 16544 32470 16544 32470 4 _0274_
rlabel metal2 s 17526 39066 17526 39066 4 _0275_
rlabel metal2 s 26082 33286 26082 33286 4 _0276_
rlabel metal1 s 27170 36822 27170 36822 4 _0277_
rlabel metal1 s 27963 27370 27963 27370 4 _0278_
rlabel metal1 s 29256 18938 29256 18938 4 _0279_
rlabel metal1 s 27232 24378 27232 24378 4 _0280_
rlabel metal1 s 26848 17238 26848 17238 4 _0281_
rlabel metal1 s 29516 15402 29516 15402 4 _0282_
rlabel metal2 s 24697 24174 24697 24174 4 _0283_
rlabel metal2 s 26358 15266 26358 15266 4 _0284_
rlabel metal1 s 27860 9962 27860 9962 4 _0285_
rlabel metal1 s 27262 7446 27262 7446 4 _0286_
rlabel metal2 s 13938 5304 13938 5304 4 _0287_
rlabel metal1 s 24502 8534 24502 8534 4 _0288_
rlabel metal2 s 23046 40290 23046 40290 4 _0289_
rlabel metal1 s 16366 31790 16366 31790 4 _0290_
rlabel metal1 s 16008 38522 16008 38522 4 _0291_
rlabel metal2 s 24794 32674 24794 32674 4 _0292_
rlabel metal1 s 26588 37978 26588 37978 4 _0293_
rlabel metal1 s 26894 27030 26894 27030 4 _0294_
rlabel metal1 s 29205 17238 29205 17238 4 _0295_
rlabel metal2 s 26082 24582 26082 24582 4 _0296_
rlabel metal2 s 24886 17000 24886 17000 4 _0297_
rlabel metal2 s 29113 12818 29113 12818 4 _0298_
rlabel metal1 s 24564 21658 24564 21658 4 _0299_
rlabel metal2 s 25433 13974 25433 13974 4 _0300_
rlabel metal1 s 27084 9554 27084 9554 4 _0301_
rlabel metal1 s 27360 6766 27360 6766 4 _0302_
rlabel metal1 s 12875 5270 12875 5270 4 _0303_
rlabel metal2 s 22857 7854 22857 7854 4 _0304_
rlabel metal1 s 37888 34646 37888 34646 4 _0305_
rlabel metal1 s 37520 33558 37520 33558 4 _0306_
rlabel metal1 s 34530 33898 34530 33898 4 _0307_
rlabel metal2 s 34086 40290 34086 40290 4 _0308_
rlabel metal2 s 14122 28934 14122 28934 4 _0309_
rlabel metal1 s 16958 43690 16958 43690 4 _0310_
rlabel metal1 s 16636 43350 16636 43350 4 _0311_
rlabel metal2 s 15410 44642 15410 44642 4 _0312_
rlabel metal2 s 16974 46342 16974 46342 4 _0313_
rlabel metal1 s 6946 26554 6946 26554 4 _0314_
rlabel metal2 s 6573 24174 6573 24174 4 _0315_
rlabel metal2 s 5474 30498 5474 30498 4 _0316_
rlabel metal1 s 5285 29206 5285 29206 4 _0317_
rlabel metal1 s 10897 29206 10897 29206 4 _0318_
rlabel metal2 s 11633 29614 11633 29614 4 _0319_
rlabel metal1 s 9793 26350 9793 26350 4 _0320_
rlabel metal1 s 10892 26350 10892 26350 4 _0321_
rlabel metal1 s 36427 35054 36427 35054 4 _0322_
rlabel metal1 s 36197 35734 36197 35734 4 _0323_
rlabel metal1 s 33713 38930 33713 38930 4 _0324_
rlabel metal2 s 34546 37026 34546 37026 4 _0325_
rlabel metal2 s 8878 40290 8878 40290 4 _0326_
rlabel metal2 s 26174 46546 26174 46546 4 _0327_
rlabel metal2 s 16969 3026 16969 3026 4 _0328_
rlabel metal1 s 33662 3026 33662 3026 4 _0329_
rlabel metal1 s 39187 36822 39187 36822 4 _0330_
rlabel metal1 s 13738 43350 13738 43350 4 _0331_
rlabel metal2 s 8602 30022 8602 30022 4 _0332_
rlabel metal2 s 10718 4998 10718 4998 4 _0333_
rlabel metal1 s 35236 43962 35236 43962 4 _0334_
rlabel metal1 s 35880 43418 35880 43418 4 _0335_
rlabel metal1 s 34449 43350 34449 43350 4 _0336_
rlabel metal2 s 33626 43010 33626 43010 4 _0337_
rlabel metal1 s 34730 18054 34730 18054 4 _0338_
rlabel metal2 s 30498 19754 30498 19754 4 _0339_
rlabel metal1 s 21482 24378 21482 24378 4 _0340_
rlabel metal1 s 30038 24174 30038 24174 4 _0341_
rlabel metal2 s 21298 23647 21298 23647 4 _0342_
rlabel metal1 s 21505 23562 21505 23562 4 _0343_
rlabel metal1 s 29716 23834 29716 23834 4 _0344_
rlabel metal2 s 29762 24378 29762 24378 4 _0345_
rlabel metal3 s 35282 23851 35282 23851 4 _0346_
rlabel metal2 s 29854 24378 29854 24378 4 _0347_
rlabel metal1 s 20792 18734 20792 18734 4 _0348_
rlabel metal1 s 20884 18802 20884 18802 4 _0349_
rlabel metal1 s 15042 18632 15042 18632 4 _0350_
rlabel metal2 s 21666 18530 21666 18530 4 _0351_
rlabel metal1 s 37858 19720 37858 19720 4 _0352_
rlabel metal2 s 21482 15878 21482 15878 4 _0353_
rlabel metal2 s 21206 16320 21206 16320 4 _0354_
rlabel metal1 s 22310 15946 22310 15946 4 _0355_
rlabel metal1 s 24886 15946 24886 15946 4 _0356_
rlabel metal1 s 31326 14042 31326 14042 4 _0357_
rlabel metal2 s 35282 14178 35282 14178 4 _0358_
rlabel metal1 s 29808 14586 29808 14586 4 _0359_
rlabel metal2 s 11362 21760 11362 21760 4 _0360_
rlabel metal1 s 22862 21522 22862 21522 4 _0361_
rlabel metal1 s 21804 22066 21804 22066 4 _0362_
rlabel metal1 s 22724 21386 22724 21386 4 _0363_
rlabel metal2 s 27370 21760 27370 21760 4 _0364_
rlabel metal1 s 35052 20570 35052 20570 4 _0365_
rlabel metal2 s 22570 21522 22570 21522 4 _0366_
rlabel metal2 s 24242 14824 24242 14824 4 _0367_
rlabel metal1 s 22770 16116 22770 16116 4 _0368_
rlabel metal2 s 27830 14722 27830 14722 4 _0369_
rlabel metal1 s 22908 15130 22908 15130 4 _0370_
rlabel metal2 s 20470 18190 20470 18190 4 _0371_
rlabel metal2 s 21114 17510 21114 17510 4 _0372_
rlabel metal1 s 21758 15606 21758 15606 4 _0373_
rlabel metal1 s 22310 15674 22310 15674 4 _0374_
rlabel metal1 s 19688 12070 19688 12070 4 _0375_
rlabel metal1 s 29762 11798 29762 11798 4 _0376_
rlabel metal3 s 8234 12597 8234 12597 4 _0377_
rlabel metal1 s 21413 13430 21413 13430 4 _0378_
rlabel metal2 s 30498 11016 30498 11016 4 _0379_
rlabel metal1 s 29670 11322 29670 11322 4 _0380_
rlabel metal1 s 32936 4794 32936 4794 4 _0381_
rlabel metal1 s 29486 11696 29486 11696 4 _0382_
rlabel metal2 s 9798 9248 9798 9248 4 _0383_
rlabel metal1 s 22954 8976 22954 8976 4 _0384_
rlabel metal2 s 20930 8840 20930 8840 4 _0385_
rlabel metal1 s 22264 9078 22264 9078 4 _0386_
rlabel metal1 s 31096 8058 31096 8058 4 _0387_
rlabel metal1 s 33810 8058 33810 8058 4 _0388_
rlabel metal1 s 22678 8908 22678 8908 4 _0389_
rlabel metal2 s 20102 9911 20102 9911 4 _0390_
rlabel metal2 s 21482 9724 21482 9724 4 _0391_
rlabel metal1 s 20838 8024 20838 8024 4 _0392_
rlabel metal1 s 22264 8602 22264 8602 4 _0393_
rlabel metal1 s 16882 6086 16882 6086 4 _0394_
rlabel metal2 s 23690 6936 23690 6936 4 _0395_
rlabel metal2 s 22034 8228 22034 8228 4 _0396_
rlabel metal2 s 25162 10982 25162 10982 4 _0397_
rlabel metal1 s 25944 11118 25944 11118 4 _0398_
rlabel metal1 s 14490 12614 14490 12614 4 _0399_
rlabel metal1 s 21988 12614 21988 12614 4 _0400_
rlabel metal1 s 26128 9622 26128 9622 4 _0401_
rlabel metal1 s 25622 11152 25622 11152 4 _0402_
rlabel metal2 s 27462 7888 27462 7888 4 _0403_
rlabel metal1 s 25714 11084 25714 11084 4 _0404_
rlabel metal2 s 11914 21488 11914 21488 4 _0405_
rlabel metal2 s 9246 37978 9246 37978 4 _0406_
rlabel metal1 s 11546 22032 11546 22032 4 _0407_
rlabel metal2 s 12466 37060 12466 37060 4 _0408_
rlabel metal1 s 11684 34578 11684 34578 4 _0409_
rlabel metal1 s 13340 13974 13340 13974 4 _0410_
rlabel metal2 s 12466 34782 12466 34782 4 _0411_
rlabel metal1 s 11638 34510 11638 34510 4 _0412_
rlabel metal2 s 16054 34782 16054 34782 4 _0413_
rlabel metal1 s 15778 19278 15778 19278 4 _0414_
rlabel metal1 s 19228 23562 19228 23562 4 _0415_
rlabel metal1 s 18400 21862 18400 21862 4 _0416_
rlabel metal1 s 19366 21556 19366 21556 4 _0417_
rlabel metal2 s 23046 37230 23046 37230 4 _0418_
rlabel metal2 s 23506 35632 23506 35632 4 _0419_
rlabel metal1 s 20838 19244 20838 19244 4 _0420_
rlabel metal2 s 20562 16286 20562 16286 4 _0421_
rlabel metal1 s 16652 21522 16652 21522 4 _0422_
rlabel metal1 s 20332 22542 20332 22542 4 _0423_
rlabel metal1 s 16836 14382 16836 14382 4 _0424_
rlabel metal1 s 21068 21114 21068 21114 4 _0425_
rlabel metal1 s 25944 34714 25944 34714 4 _0426_
rlabel metal1 s 15502 20774 15502 20774 4 _0427_
rlabel metal2 s 16146 16167 16146 16167 4 _0428_
rlabel metal1 s 32683 36006 32683 36006 4 _0429_
rlabel metal2 s 21666 23902 21666 23902 4 _0430_
rlabel metal1 s 24288 34714 24288 34714 4 _0431_
rlabel metal1 s 6946 32776 6946 32776 4 _0432_
rlabel metal1 s 12558 16626 12558 16626 4 _0433_
rlabel metal1 s 21390 32402 21390 32402 4 _0434_
rlabel metal2 s 19274 29682 19274 29682 4 _0435_
rlabel metal1 s 20102 30362 20102 30362 4 _0436_
rlabel metal2 s 20838 32640 20838 32640 4 _0437_
rlabel metal1 s 21206 33014 21206 33014 4 _0438_
rlabel metal1 s 21206 32368 21206 32368 4 _0439_
rlabel metal1 s 13294 35802 13294 35802 4 _0440_
rlabel metal1 s 14582 35054 14582 35054 4 _0441_
rlabel metal2 s 18722 36958 18722 36958 4 _0442_
rlabel metal1 s 16698 35258 16698 35258 4 _0443_
rlabel metal2 s 32798 30566 32798 30566 4 _0444_
rlabel metal2 s 11822 21913 11822 21913 4 _0445_
rlabel metal1 s 13570 35020 13570 35020 4 _0446_
rlabel metal1 s 13248 31994 13248 31994 4 _0447_
rlabel metal1 s 14076 35054 14076 35054 4 _0448_
rlabel metal1 s 11822 20978 11822 20978 4 _0449_
rlabel metal1 s 16284 35598 16284 35598 4 _0450_
rlabel metal1 s 14674 35530 14674 35530 4 _0451_
rlabel metal2 s 14398 35258 14398 35258 4 _0452_
rlabel metal1 s 25714 31178 25714 31178 4 _0453_
rlabel metal1 s 28106 31348 28106 31348 4 _0454_
rlabel metal1 s 11822 31858 11822 31858 4 _0455_
rlabel metal2 s 12558 31535 12558 31535 4 _0456_
rlabel metal2 s 14582 15980 14582 15980 4 _0457_
rlabel metal1 s 28658 31926 28658 31926 4 _0458_
rlabel metal2 s 29026 31416 29026 31416 4 _0459_
rlabel metal1 s 33902 30906 33902 30906 4 _0460_
rlabel metal1 s 19872 10030 19872 10030 4 _0461_
rlabel metal1 s 27830 31280 27830 31280 4 _0462_
rlabel metal1 s 26450 35190 26450 35190 4 _0463_
rlabel metal1 s 27922 34578 27922 34578 4 _0464_
rlabel metal1 s 12006 35122 12006 35122 4 _0465_
rlabel metal2 s 17342 34952 17342 34952 4 _0466_
rlabel metal1 s 28842 34442 28842 34442 4 _0467_
rlabel metal1 s 27646 34612 27646 34612 4 _0468_
rlabel metal1 s 29578 34646 29578 34646 4 _0469_
rlabel metal1 s 27738 34544 27738 34544 4 _0470_
rlabel metal1 s 5014 20332 5014 20332 4 _0471_
rlabel metal1 s 5474 17102 5474 17102 4 _0472_
rlabel metal2 s 9890 25636 9890 25636 4 _0473_
rlabel metal1 s 12144 20570 12144 20570 4 _0474_
rlabel metal1 s 23598 25874 23598 25874 4 _0475_
rlabel metal1 s 24288 26486 24288 26486 4 _0476_
rlabel metal1 s 23690 25806 23690 25806 4 _0477_
rlabel metal1 s 30314 17782 30314 17782 4 _0478_
rlabel metal2 s 31050 17374 31050 17374 4 _0479_
rlabel metal2 s 30590 26554 30590 26554 4 _0480_
rlabel metal2 s 33350 26520 33350 26520 4 _0481_
rlabel metal1 s 31970 14450 31970 14450 4 _0482_
rlabel metal2 s 23414 25891 23414 25891 4 _0483_
rlabel metal2 s 6210 20128 6210 20128 4 _0484_
rlabel metal1 s 16790 20230 16790 20230 4 _0485_
rlabel metal1 s 19274 21386 19274 21386 4 _0486_
rlabel metal2 s 20838 21216 20838 21216 4 _0487_
rlabel metal2 s 31694 18564 31694 18564 4 _0488_
rlabel metal1 s 33626 19278 33626 19278 4 _0489_
rlabel metal1 s 20654 20876 20654 20876 4 _0490_
rlabel metal2 s 21942 24446 21942 24446 4 _0491_
rlabel metal1 s 22678 24174 22678 24174 4 _0492_
rlabel metal1 s 7728 23154 7728 23154 4 _0493_
rlabel metal1 s 21298 24208 21298 24208 4 _0494_
rlabel metal1 s 28106 24038 28106 24038 4 _0495_
rlabel metal2 s 22448 24174 22448 24174 4 _0496_
rlabel metal2 s 33258 24480 33258 24480 4 _0497_
rlabel metal1 s 22494 24140 22494 24140 4 _0498_
rlabel metal1 s 26128 18598 26128 18598 4 _0499_
rlabel metal2 s 24886 18972 24886 18972 4 _0500_
rlabel metal1 s 23966 18598 23966 18598 4 _0501_
rlabel metal1 s 16100 18394 16100 18394 4 _0502_
rlabel metal1 s 13386 17714 13386 17714 4 _0503_
rlabel metal1 s 15410 19448 15410 19448 4 _0504_
rlabel metal1 s 20148 19482 20148 19482 4 _0505_
rlabel metal1 s 10856 16150 10856 16150 4 _0506_
rlabel metal1 s 20976 16558 20976 16558 4 _0507_
rlabel metal1 s 20056 16558 20056 16558 4 _0508_
rlabel metal1 s 18354 17034 18354 17034 4 _0509_
rlabel metal2 s 19274 17187 19274 17187 4 _0510_
rlabel metal2 s 20102 16830 20102 16830 4 _0511_
rlabel metal1 s 20424 16694 20424 16694 4 _0512_
rlabel metal1 s 31832 13498 31832 13498 4 _0513_
rlabel metal2 s 33350 12682 33350 12682 4 _0514_
rlabel metal1 s 34224 12750 34224 12750 4 _0515_
rlabel metal1 s 34822 12954 34822 12954 4 _0516_
rlabel metal1 s 20654 16626 20654 16626 4 _0517_
rlabel metal2 s 21574 22984 21574 22984 4 _0518_
rlabel metal1 s 23138 23154 23138 23154 4 _0519_
rlabel metal2 s 12926 23188 12926 23188 4 _0520_
rlabel metal1 s 21206 22984 21206 22984 4 _0521_
rlabel metal1 s 25714 21658 25714 21658 4 _0522_
rlabel metal1 s 23092 22746 23092 22746 4 _0523_
rlabel metal2 s 33534 21216 33534 21216 4 _0524_
rlabel metal1 s 22862 23052 22862 23052 4 _0525_
rlabel metal2 s 12374 16830 12374 16830 4 _0526_
rlabel metal2 s 21298 16354 21298 16354 4 _0527_
rlabel metal1 s 21206 14858 21206 14858 4 _0528_
rlabel metal1 s 21827 15130 21827 15130 4 _0529_
rlabel metal1 s 26818 14042 26818 14042 4 _0530_
rlabel metal2 s 24886 13600 24886 13600 4 _0531_
rlabel metal1 s 24242 14586 24242 14586 4 _0532_
rlabel metal1 s 9384 12342 9384 12342 4 _0533_
rlabel metal1 s 16054 13838 16054 13838 4 _0534_
rlabel metal1 s 19596 12682 19596 12682 4 _0535_
rlabel metal1 s 20056 12410 20056 12410 4 _0536_
rlabel metal1 s 31648 9962 31648 9962 4 _0537_
rlabel metal1 s 33672 5338 33672 5338 4 _0538_
rlabel metal2 s 19550 12036 19550 12036 4 _0539_
rlabel metal2 s 12834 10778 12834 10778 4 _0540_
rlabel metal2 s 23230 10676 23230 10676 4 _0541_
rlabel metal2 s 21114 8738 21114 8738 4 _0542_
rlabel metal2 s 23138 9792 23138 9792 4 _0543_
rlabel metal2 s 31326 9078 31326 9078 4 _0544_
rlabel metal2 s 34822 9010 34822 9010 4 _0545_
rlabel metal1 s 29946 9690 29946 9690 4 _0546_
rlabel metal2 s 13662 10268 13662 10268 4 _0547_
rlabel metal1 s 21298 10098 21298 10098 4 _0548_
rlabel metal1 s 19550 8602 19550 8602 4 _0549_
rlabel metal1 s 20286 9520 20286 9520 4 _0550_
rlabel metal1 s 17710 6698 17710 6698 4 _0551_
rlabel metal1 s 23460 5882 23460 5882 4 _0552_
rlabel metal1 s 20976 7514 20976 7514 4 _0553_
rlabel metal2 s 14490 11628 14490 11628 4 _0554_
rlabel metal2 s 16330 10472 16330 10472 4 _0555_
rlabel metal2 s 19734 10438 19734 10438 4 _0556_
rlabel metal1 s 20424 10234 20424 10234 4 _0557_
rlabel metal1 s 25806 7854 25806 7854 4 _0558_
rlabel metal2 s 26818 6528 26818 6528 4 _0559_
rlabel metal1 s 25070 7990 25070 7990 4 _0560_
rlabel metal1 s 38686 37094 38686 37094 4 _0561_
rlabel metal1 s 13432 29070 13432 29070 4 _0562_
rlabel metal1 s 33442 40052 33442 40052 4 _0563_
rlabel metal1 s 19458 42194 19458 42194 4 _0564_
rlabel metal1 s 15962 31722 15962 31722 4 _0565_
rlabel metal2 s 19090 41786 19090 41786 4 _0566_
rlabel metal2 s 16146 36516 16146 36516 4 _0567_
rlabel metal1 s 17940 46002 17940 46002 4 _0568_
rlabel metal1 s 16790 44370 16790 44370 4 _0569_
rlabel metal1 s 4462 43690 4462 43690 4 _0570_
rlabel metal2 s 18078 45764 18078 45764 4 _0571_
rlabel metal1 s 45034 31450 45034 31450 4 _0572_
rlabel metal1 s 44758 32402 44758 32402 4 _0573_
rlabel metal1 s 44988 31790 44988 31790 4 _0574_
rlabel metal1 s 46230 32368 46230 32368 4 _0575_
rlabel metal2 s 45496 33490 45496 33490 4 _0576_
rlabel metal1 s 45770 32266 45770 32266 4 _0577_
rlabel metal1 s 44482 33082 44482 33082 4 _0578_
rlabel metal2 s 41814 31552 41814 31552 4 _0579_
rlabel metal1 s 44482 33456 44482 33456 4 _0580_
rlabel metal1 s 44206 33524 44206 33524 4 _0581_
rlabel metal1 s 44482 32334 44482 32334 4 _0582_
rlabel metal1 s 44390 32538 44390 32538 4 _0583_
rlabel metal1 s 42826 33354 42826 33354 4 _0584_
rlabel metal2 s 45402 33694 45402 33694 4 _0585_
rlabel metal2 s 45034 33694 45034 33694 4 _0586_
rlabel metal1 s 46506 33422 46506 33422 4 _0587_
rlabel metal1 s 46414 33286 46414 33286 4 _0588_
rlabel metal1 s 40526 30736 40526 30736 4 _0589_
rlabel metal1 s 41452 32402 41452 32402 4 _0590_
rlabel metal2 s 41262 32844 41262 32844 4 _0591_
rlabel metal1 s 40986 33932 40986 33932 4 _0592_
rlabel metal1 s 42366 33490 42366 33490 4 _0593_
rlabel metal2 s 42090 33762 42090 33762 4 _0594_
rlabel metal2 s 41906 33252 41906 33252 4 _0595_
rlabel metal1 s 42458 33626 42458 33626 4 _0596_
rlabel metal2 s 41078 33796 41078 33796 4 _0597_
rlabel metal2 s 40342 33660 40342 33660 4 _0598_
rlabel metal1 s 41814 29580 41814 29580 4 _0599_
rlabel metal1 s 42090 29648 42090 29648 4 _0600_
rlabel metal1 s 41032 29682 41032 29682 4 _0601_
rlabel metal1 s 41722 26894 41722 26894 4 _0602_
rlabel metal1 s 41101 29818 41101 29818 4 _0603_
rlabel metal1 s 40940 29138 40940 29138 4 _0604_
rlabel metal1 s 42090 26962 42090 26962 4 _0605_
rlabel metal1 s 39238 26894 39238 26894 4 _0606_
rlabel metal2 s 42458 24191 42458 24191 4 _0607_
rlabel metal1 s 42826 26384 42826 26384 4 _0608_
rlabel metal1 s 42504 22950 42504 22950 4 _0609_
rlabel metal1 s 41262 27098 41262 27098 4 _0610_
rlabel metal1 s 41170 27438 41170 27438 4 _0611_
rlabel metal1 s 38962 26996 38962 26996 4 _0612_
rlabel metal1 s 44298 24786 44298 24786 4 _0613_
rlabel metal1 s 43930 24820 43930 24820 4 _0614_
rlabel metal1 s 43976 25670 43976 25670 4 _0615_
rlabel metal1 s 44390 25908 44390 25908 4 _0616_
rlabel metal1 s 45862 24140 45862 24140 4 _0617_
rlabel metal1 s 44114 24922 44114 24922 4 _0618_
rlabel metal2 s 45310 25534 45310 25534 4 _0619_
rlabel metal2 s 44758 24956 44758 24956 4 _0620_
rlabel metal2 s 39514 24140 39514 24140 4 _0621_
rlabel metal2 s 45770 23324 45770 23324 4 _0622_
rlabel metal1 s 45908 23698 45908 23698 4 _0623_
rlabel metal1 s 45678 23562 45678 23562 4 _0624_
rlabel metal2 s 46414 24174 46414 24174 4 _0625_
rlabel metal2 s 46598 24378 46598 24378 4 _0626_
rlabel metal1 s 46414 24106 46414 24106 4 _0627_
rlabel metal2 s 43562 20230 43562 20230 4 _0628_
rlabel metal2 s 43010 20230 43010 20230 4 _0629_
rlabel metal2 s 44574 19278 44574 19278 4 _0630_
rlabel metal1 s 44896 23086 44896 23086 4 _0631_
rlabel metal1 s 44022 15028 44022 15028 4 _0632_
rlabel metal1 s 38870 18870 38870 18870 4 _0633_
rlabel metal2 s 44298 19074 44298 19074 4 _0634_
rlabel metal1 s 43884 19482 43884 19482 4 _0635_
rlabel metal2 s 44390 19482 44390 19482 4 _0636_
rlabel metal1 s 45034 17170 45034 17170 4 _0637_
rlabel metal2 s 44574 17476 44574 17476 4 _0638_
rlabel metal2 s 42090 18462 42090 18462 4 _0639_
rlabel metal1 s 42734 17306 42734 17306 4 _0640_
rlabel metal1 s 43516 18190 43516 18190 4 _0641_
rlabel metal1 s 44436 18394 44436 18394 4 _0642_
rlabel metal1 s 44896 18190 44896 18190 4 _0643_
rlabel metal1 s 43010 16626 43010 16626 4 _0644_
rlabel metal1 s 43378 16218 43378 16218 4 _0645_
rlabel metal1 s 40848 16694 40848 16694 4 _0646_
rlabel metal2 s 45126 16490 45126 16490 4 _0647_
rlabel metal2 s 43194 17102 43194 17102 4 _0648_
rlabel metal1 s 43240 14994 43240 14994 4 _0649_
rlabel metal2 s 38962 16286 38962 16286 4 _0650_
rlabel metal2 s 45034 17034 45034 17034 4 _0651_
rlabel metal1 s 44068 16014 44068 16014 4 _0652_
rlabel metal2 s 43746 15436 43746 15436 4 _0653_
rlabel metal1 s 43700 12206 43700 12206 4 _0654_
rlabel metal1 s 40158 9996 40158 9996 4 _0655_
rlabel metal2 s 43194 9554 43194 9554 4 _0656_
rlabel metal1 s 43976 11118 43976 11118 4 _0657_
rlabel metal1 s 43654 11254 43654 11254 4 _0658_
rlabel metal1 s 40526 10778 40526 10778 4 _0659_
rlabel metal2 s 43424 9622 43424 9622 4 _0660_
rlabel metal1 s 42274 11832 42274 11832 4 _0661_
rlabel metal1 s 43286 12410 43286 12410 4 _0662_
rlabel metal2 s 43010 14416 43010 14416 4 _0663_
rlabel metal2 s 43102 14076 43102 14076 4 _0664_
rlabel metal2 s 42274 13056 42274 13056 4 _0665_
rlabel metal1 s 42044 12750 42044 12750 4 _0666_
rlabel metal1 s 42918 11866 42918 11866 4 _0667_
rlabel metal2 s 38870 10948 38870 10948 4 _0668_
rlabel metal1 s 38226 11628 38226 11628 4 _0669_
rlabel metal1 s 40204 12818 40204 12818 4 _0670_
rlabel metal1 s 41676 11866 41676 11866 4 _0671_
rlabel metal1 s 40526 12716 40526 12716 4 _0672_
rlabel metal1 s 38410 12138 38410 12138 4 _0673_
rlabel metal1 s 38732 12206 38732 12206 4 _0674_
rlabel metal1 s 38502 12274 38502 12274 4 _0675_
rlabel metal1 s 39422 12410 39422 12410 4 _0676_
rlabel metal1 s 39790 12852 39790 12852 4 _0677_
rlabel metal1 s 38594 11798 38594 11798 4 _0678_
rlabel metal1 s 38813 11798 38813 11798 4 _0679_
rlabel metal2 s 39606 12619 39606 12619 4 _0680_
rlabel metal2 s 34684 30804 34684 30804 4 _0681_
rlabel metal1 s 36846 32198 36846 32198 4 _0682_
rlabel metal2 s 38916 17170 38916 17170 4 _0683_
rlabel metal1 s 37030 31314 37030 31314 4 _0684_
rlabel metal1 s 36458 12206 36458 12206 4 _0685_
rlabel metal1 s 38042 19210 38042 19210 4 _0686_
rlabel metal2 s 39974 23596 39974 23596 4 _0687_
rlabel metal1 s 40388 27438 40388 27438 4 _0688_
rlabel metal1 s 43286 29580 43286 29580 4 _0689_
rlabel metal1 s 40871 28050 40871 28050 4 _0690_
rlabel metal1 s 39468 28186 39468 28186 4 _0691_
rlabel metal1 s 36110 29172 36110 29172 4 _0692_
rlabel metal2 s 21482 38216 21482 38216 4 _0693_
rlabel metal1 s 32752 37978 32752 37978 4 _0694_
rlabel metal1 s 16698 26418 16698 26418 4 _0695_
rlabel metal2 s 13846 28288 13846 28288 4 _0696_
rlabel metal1 s 12006 28492 12006 28492 4 _0697_
rlabel metal1 s 15318 27030 15318 27030 4 _0698_
rlabel metal1 s 10856 27030 10856 27030 4 _0699_
rlabel metal1 s 16836 9350 16836 9350 4 _0700_
rlabel metal1 s 13156 33422 13156 33422 4 _0701_
rlabel metal2 s 30866 39508 30866 39508 4 _0702_
rlabel metal1 s 45678 29580 45678 29580 4 _0703_
rlabel metal2 s 45494 29818 45494 29818 4 _0704_
rlabel metal1 s 45034 28594 45034 28594 4 _0705_
rlabel metal2 s 40986 16490 40986 16490 4 _0706_
rlabel metal1 s 44344 32470 44344 32470 4 _0707_
rlabel metal2 s 40066 12512 40066 12512 4 _0708_
rlabel metal2 s 41262 17952 41262 17952 4 _0709_
rlabel metal2 s 44942 28356 44942 28356 4 _0710_
rlabel metal1 s 37996 28390 37996 28390 4 _0711_
rlabel metal2 s 38410 19958 38410 19958 4 _0712_
rlabel metal1 s 37674 17646 37674 17646 4 _0713_
rlabel metal1 s 14352 29274 14352 29274 4 _0714_
rlabel metal1 s 38272 18734 38272 18734 4 _0715_
rlabel metal1 s 37536 28526 37536 28526 4 _0716_
rlabel metal1 s 36432 28730 36432 28730 4 _0717_
rlabel metal1 s 13156 33558 13156 33558 4 _0718_
rlabel metal1 s 12558 33490 12558 33490 4 _0719_
rlabel metal1 s 40204 16082 40204 16082 4 _0720_
rlabel metal2 s 42734 33966 42734 33966 4 _0721_
rlabel metal1 s 42826 33524 42826 33524 4 _0722_
rlabel metal1 s 43378 32368 43378 32368 4 _0723_
rlabel metal1 s 40710 21522 40710 21522 4 _0724_
rlabel metal2 s 42366 31790 42366 31790 4 _0725_
rlabel metal2 s 42182 32691 42182 32691 4 _0726_
rlabel metal1 s 41676 32198 41676 32198 4 _0727_
rlabel metal1 s 40894 30192 40894 30192 4 _0728_
rlabel metal2 s 18630 3553 18630 3553 4 _0729_
rlabel metal1 s 36432 30226 36432 30226 4 _0730_
rlabel metal2 s 16882 37536 16882 37536 4 _0731_
rlabel metal2 s 13662 39610 13662 39610 4 _0732_
rlabel metal1 s 11592 39542 11592 39542 4 _0733_
rlabel metal1 s 42090 31858 42090 31858 4 _0734_
rlabel metal2 s 42458 32640 42458 32640 4 _0735_
rlabel metal1 s 42458 31314 42458 31314 4 _0736_
rlabel metal1 s 41354 31246 41354 31246 4 _0737_
rlabel metal2 s 40434 30906 40434 30906 4 _0738_
rlabel metal2 s 39422 30396 39422 30396 4 _0739_
rlabel metal1 s 36754 30362 36754 30362 4 _0740_
rlabel metal1 s 26818 32980 26818 32980 4 _0741_
rlabel metal1 s 31004 31926 31004 31926 4 _0742_
rlabel metal2 s 31234 30906 31234 30906 4 _0743_
rlabel metal1 s 38778 30226 38778 30226 4 _0744_
rlabel metal2 s 43470 32844 43470 32844 4 _0745_
rlabel metal2 s 43194 32521 43194 32521 4 _0746_
rlabel metal1 s 42780 32198 42780 32198 4 _0747_
rlabel metal1 s 44482 30158 44482 30158 4 _0748_
rlabel metal1 s 43286 31790 43286 31790 4 _0749_
rlabel metal1 s 43194 29648 43194 29648 4 _0750_
rlabel metal1 s 42734 29614 42734 29614 4 _0751_
rlabel metal2 s 40894 30005 40894 30005 4 _0752_
rlabel metal1 s 35696 31790 35696 31790 4 _0753_
rlabel metal1 s 32338 33422 32338 33422 4 _0754_
rlabel metal1 s 27922 39474 27922 39474 4 _0755_
rlabel metal2 s 29946 38284 29946 38284 4 _0756_
rlabel metal1 s 41814 27982 41814 27982 4 _0757_
rlabel metal1 s 42458 28152 42458 28152 4 _0758_
rlabel metal2 s 42650 28186 42650 28186 4 _0759_
rlabel metal1 s 38778 27472 38778 27472 4 _0760_
rlabel metal1 s 37306 27302 37306 27302 4 _0761_
rlabel metal1 s 39514 27098 39514 27098 4 _0762_
rlabel metal1 s 37214 27438 37214 27438 4 _0763_
rlabel metal1 s 33626 28016 33626 28016 4 _0764_
rlabel metal1 s 29716 28186 29716 28186 4 _0765_
rlabel metal2 s 31970 28220 31970 28220 4 _0766_
rlabel metal1 s 43654 30260 43654 30260 4 _0767_
rlabel metal1 s 42872 30294 42872 30294 4 _0768_
rlabel metal2 s 42826 26146 42826 26146 4 _0769_
rlabel metal1 s 42090 24310 42090 24310 4 _0770_
rlabel metal2 s 41538 24548 41538 24548 4 _0771_
rlabel metal1 s 41998 24786 41998 24786 4 _0772_
rlabel metal1 s 41630 24684 41630 24684 4 _0773_
rlabel metal2 s 41170 25432 41170 25432 4 _0774_
rlabel metal2 s 36570 27676 36570 27676 4 _0775_
rlabel metal1 s 18078 19958 18078 19958 4 _0776_
rlabel metal1 s 32200 19686 32200 19686 4 _0777_
rlabel metal1 s 34500 15538 34500 15538 4 _0778_
rlabel metal1 s 34500 15674 34500 15674 4 _0779_
rlabel metal1 s 41998 23834 41998 23834 4 _0780_
rlabel metal1 s 42550 23086 42550 23086 4 _0781_
rlabel metal1 s 40526 23528 40526 23528 4 _0782_
rlabel metal2 s 40618 23868 40618 23868 4 _0783_
rlabel metal2 s 39790 23868 39790 23868 4 _0784_
rlabel metal1 s 40710 23732 40710 23732 4 _0785_
rlabel metal1 s 39284 23834 39284 23834 4 _0786_
rlabel metal1 s 19412 24038 19412 24038 4 _0787_
rlabel metal1 s 34776 24038 34776 24038 4 _0788_
rlabel metal1 s 33488 24378 33488 24378 4 _0789_
rlabel metal1 s 38090 17646 38090 17646 4 _0790_
rlabel metal2 s 42918 22780 42918 22780 4 _0791_
rlabel metal1 s 43470 23120 43470 23120 4 _0792_
rlabel metal2 s 43562 23596 43562 23596 4 _0793_
rlabel metal1 s 42872 22542 42872 22542 4 _0794_
rlabel metal1 s 43010 22406 43010 22406 4 _0795_
rlabel metal1 s 41354 18224 41354 18224 4 _0796_
rlabel metal1 s 42918 22066 42918 22066 4 _0797_
rlabel metal1 s 42412 21522 42412 21522 4 _0798_
rlabel metal2 s 43930 21284 43930 21284 4 _0799_
rlabel metal1 s 38042 17544 38042 17544 4 _0800_
rlabel metal2 s 37766 17986 37766 17986 4 _0801_
rlabel metal1 s 20148 17850 20148 17850 4 _0802_
rlabel metal2 s 23230 17204 23230 17204 4 _0803_
rlabel metal1 s 42090 19822 42090 19822 4 _0804_
rlabel metal2 s 41538 20026 41538 20026 4 _0805_
rlabel metal1 s 41492 20026 41492 20026 4 _0806_
rlabel metal1 s 37766 19856 37766 19856 4 _0807_
rlabel metal1 s 37766 19482 37766 19482 4 _0808_
rlabel metal1 s 19504 16218 19504 16218 4 _0809_
rlabel metal2 s 32522 14688 32522 14688 4 _0810_
rlabel metal2 s 34454 11322 34454 11322 4 _0811_
rlabel metal1 s 40772 18734 40772 18734 4 _0812_
rlabel metal2 s 41722 17680 41722 17680 4 _0813_
rlabel metal1 s 40710 18394 40710 18394 4 _0814_
rlabel metal1 s 40802 18632 40802 18632 4 _0815_
rlabel metal1 s 40940 18870 40940 18870 4 _0816_
rlabel metal2 s 40526 18462 40526 18462 4 _0817_
rlabel metal1 s 38594 20400 38594 20400 4 _0818_
rlabel metal1 s 18124 21998 18124 21998 4 _0819_
rlabel metal1 s 34086 20978 34086 20978 4 _0820_
rlabel metal1 s 33672 20910 33672 20910 4 _0821_
rlabel metal2 s 38502 16762 38502 16762 4 _0822_
rlabel metal1 s 40710 16524 40710 16524 4 _0823_
rlabel metal2 s 40802 16252 40802 16252 4 _0824_
rlabel metal1 s 40526 16014 40526 16014 4 _0825_
rlabel metal2 s 38318 16388 38318 16388 4 _0826_
rlabel metal1 s 18768 15470 18768 15470 4 _0827_
rlabel metal2 s 29302 12988 29302 12988 4 _0828_
rlabel metal2 s 23046 11084 23046 11084 4 _0829_
rlabel metal1 s 40388 17034 40388 17034 4 _0830_
rlabel metal1 s 42780 16558 42780 16558 4 _0831_
rlabel metal2 s 42366 16762 42366 16762 4 _0832_
rlabel metal1 s 42734 20978 42734 20978 4 _0833_
rlabel metal1 s 42688 11118 42688 11118 4 _0834_
rlabel metal1 s 43424 11322 43424 11322 4 _0835_
rlabel metal1 s 42918 10982 42918 10982 4 _0836_
rlabel metal2 s 43562 11900 43562 11900 4 _0837_
rlabel metal2 s 38778 12087 38778 12087 4 _0838_
rlabel metal1 s 19642 12818 19642 12818 4 _0839_
rlabel metal2 s 19274 4590 19274 4590 4 _0840_
rlabel metal1 s 32752 3502 32752 3502 4 _0841_
rlabel metal1 s 43194 9418 43194 9418 4 _0842_
rlabel metal1 s 42642 9996 42642 9996 4 _0843_
rlabel metal2 s 43102 9826 43102 9826 4 _0844_
rlabel metal1 s 43332 10098 43332 10098 4 _0845_
rlabel metal2 s 39790 9248 39790 9248 4 _0846_
rlabel metal1 s 38272 8398 38272 8398 4 _0847_
rlabel metal2 s 19642 7582 19642 7582 4 _0848_
rlabel metal1 s 20930 6154 20930 6154 4 _0849_
rlabel metal1 s 32200 8058 32200 8058 4 _0850_
rlabel metal1 s 42734 10574 42734 10574 4 _0851_
rlabel metal1 s 40480 9554 40480 9554 4 _0852_
rlabel metal1 s 40618 10234 40618 10234 4 _0853_
rlabel metal1 s 40388 10506 40388 10506 4 _0854_
rlabel metal1 s 39100 11254 39100 11254 4 _0855_
rlabel metal1 s 39836 9486 39836 9486 4 _0856_
rlabel metal1 s 40158 10098 40158 10098 4 _0857_
rlabel metal1 s 36386 8976 36386 8976 4 _0858_
rlabel metal1 s 17848 6630 17848 6630 4 _0859_
rlabel metal1 s 20470 3638 20470 3638 4 _0860_
rlabel metal1 s 21574 4114 21574 4114 4 _0861_
rlabel metal1 s 38640 9554 38640 9554 4 _0862_
rlabel metal2 s 38410 10812 38410 10812 4 _0863_
rlabel metal1 s 39238 10778 39238 10778 4 _0864_
rlabel metal1 s 38502 10676 38502 10676 4 _0865_
rlabel metal1 s 39146 14960 39146 14960 4 _0866_
rlabel metal2 s 38686 12682 38686 12682 4 _0867_
rlabel metal2 s 38410 10030 38410 10030 4 _0868_
rlabel metal2 s 17342 8976 17342 8976 4 _0869_
rlabel metal2 s 21390 3978 21390 3978 4 _0870_
rlabel metal2 s 25162 3468 25162 3468 4 _0871_
rlabel metal2 s 16330 25602 16330 25602 4 _0872_
rlabel metal1 s 13754 26214 13754 26214 4 _0873_
rlabel metal2 s 16974 27234 16974 27234 4 _0874_
rlabel metal1 s 15410 25330 15410 25330 4 _0875_
rlabel metal3 s 33971 13804 33971 13804 4 _0876_
rlabel metal2 s 15134 34969 15134 34969 4 _0877_
rlabel metal2 s 31602 38148 31602 38148 4 _0878_
rlabel metal1 s 14076 33966 14076 33966 4 _0879_
rlabel metal2 s 13202 40324 13202 40324 4 _0880_
rlabel metal2 s 32154 32708 32154 32708 4 _0881_
rlabel metal2 s 29946 37434 29946 37434 4 _0882_
rlabel metal1 s 34086 28458 34086 28458 4 _0883_
rlabel metal2 s 34362 13260 34362 13260 4 _0884_
rlabel metal1 s 35098 17170 35098 17170 4 _0885_
rlabel metal2 s 35374 24548 35374 24548 4 _0886_
rlabel metal2 s 24426 20230 24426 20230 4 _0887_
rlabel metal1 s 33764 13294 33764 13294 4 _0888_
rlabel metal2 s 35742 22100 35742 22100 4 _0889_
rlabel metal1 s 25162 12852 25162 12852 4 _0890_
rlabel metal1 s 32338 3706 32338 3706 4 _0891_
rlabel metal2 s 34362 6970 34362 6970 4 _0892_
rlabel metal1 s 22862 3502 22862 3502 4 _0893_
rlabel metal2 s 25806 3638 25806 3638 4 _0894_
rlabel metal2 s 16054 27132 16054 27132 4 _0895_
rlabel metal1 s 18538 3502 18538 3502 4 _0896_
rlabel metal1 s 13202 41038 13202 41038 4 _0897_
rlabel metal1 s 30774 40052 30774 40052 4 _0898_
rlabel metal1 s 12144 31654 12144 31654 4 _0899_
rlabel metal2 s 10718 40732 10718 40732 4 _0900_
rlabel metal1 s 31096 31314 31096 31314 4 _0901_
rlabel metal2 s 29762 35258 29762 35258 4 _0902_
rlabel metal1 s 32108 26962 32108 26962 4 _0903_
rlabel metal1 s 33166 21454 33166 21454 4 _0904_
rlabel metal2 s 32890 16762 32890 16762 4 _0905_
rlabel metal2 s 32430 24310 32430 24310 4 _0906_
rlabel metal2 s 22126 18700 22126 18700 4 _0907_
rlabel metal2 s 32706 11322 32706 11322 4 _0908_
rlabel metal1 s 32476 21522 32476 21522 4 _0909_
rlabel metal1 s 22678 11730 22678 11730 4 _0910_
rlabel metal2 s 31050 3638 31050 3638 4 _0911_
rlabel metal1 s 32016 6970 32016 6970 4 _0912_
rlabel metal1 s 19964 3502 19964 3502 4 _0913_
rlabel metal2 s 23506 3910 23506 3910 4 _0914_
rlabel metal2 s 15870 27642 15870 27642 4 _0915_
rlabel metal2 s 19596 17204 19596 17204 4 _0916_
rlabel metal1 s 16100 40562 16100 40562 4 _0917_
rlabel metal2 s 21850 41140 21850 41140 4 _0918_
rlabel metal2 s 16330 34374 16330 34374 4 _0919_
rlabel metal1 s 14858 40052 14858 40052 4 _0920_
rlabel metal1 s 27002 29818 27002 29818 4 _0921_
rlabel metal1 s 26450 40052 26450 40052 4 _0922_
rlabel metal1 s 27232 28050 27232 28050 4 _0923_
rlabel metal2 s 19826 18462 19826 18462 4 _0924_
rlabel metal2 s 31418 20230 31418 20230 4 _0925_
rlabel metal1 s 30958 24378 30958 24378 4 _0926_
rlabel metal1 s 19090 18258 19090 18258 4 _0927_
rlabel metal1 s 32177 15470 32177 15470 4 _0928_
rlabel metal2 s 23506 22406 23506 22406 4 _0929_
rlabel metal1 s 20470 13328 20470 13328 4 _0930_
rlabel metal1 s 17572 4590 17572 4590 4 _0931_
rlabel metal1 s 19688 6290 19688 6290 4 _0932_
rlabel metal2 s 16698 3740 16698 3740 4 _0933_
rlabel metal2 s 18630 4284 18630 4284 4 _0934_
rlabel metal1 s 14582 28050 14582 28050 4 _0935_
rlabel metal2 s 14398 25670 14398 25670 4 _0936_
rlabel metal1 s 15410 4692 15410 4692 4 _0937_
rlabel metal1 s 19734 34476 19734 34476 4 _0938_
rlabel metal2 s 24058 40630 24058 40630 4 _0939_
rlabel metal2 s 18538 34170 18538 34170 4 _0940_
rlabel metal1 s 17158 40154 17158 40154 4 _0941_
rlabel metal2 s 30406 32708 30406 32708 4 _0942_
rlabel metal2 s 27922 40018 27922 40018 4 _0943_
rlabel metal1 s 30222 29172 30222 29172 4 _0944_
rlabel metal1 s 31786 22100 31786 22100 4 _0945_
rlabel metal2 s 31326 16524 31326 16524 4 _0946_
rlabel metal2 s 31234 22304 31234 22304 4 _0947_
rlabel metal1 s 27324 18938 27324 18938 4 _0948_
rlabel metal2 s 31418 11084 31418 11084 4 _0949_
rlabel metal1 s 27646 22406 27646 22406 4 _0950_
rlabel metal2 s 26818 11900 26818 11900 4 _0951_
rlabel metal1 s 29394 4590 29394 4590 4 _0952_
rlabel metal2 s 30866 6970 30866 6970 4 _0953_
rlabel metal2 s 14766 3978 14766 3978 4 _0954_
rlabel metal1 s 24702 5610 24702 5610 4 _0955_
rlabel metal2 s 20194 38692 20194 38692 4 _0956_
rlabel metal1 s 13064 26010 13064 26010 4 _0957_
rlabel metal2 s 6578 16865 6578 16865 4 _0958_
rlabel metal1 s 3634 34476 3634 34476 4 _0959_
rlabel metal2 s 6670 37060 6670 37060 4 _0960_
rlabel metal2 s 16054 30498 16054 30498 4 _0961_
rlabel metal2 s 1702 32708 1702 32708 4 _0962_
rlabel metal1 s 14536 37094 14536 37094 4 _0963_
rlabel metal1 s 6486 35020 6486 35020 4 _0964_
rlabel metal1 s 16790 30804 16790 30804 4 _0965_
rlabel metal1 s 7038 32402 7038 32402 4 _0966_
rlabel metal1 s 20470 36754 20470 36754 4 _0967_
rlabel metal1 s 3450 34714 3450 34714 4 _0968_
rlabel metal1 s 4186 27302 4186 27302 4 _0969_
rlabel metal1 s 2346 25874 2346 25874 4 _0970_
rlabel metal1 s 4232 20502 4232 20502 4 _0971_
rlabel metal1 s 3542 20978 3542 20978 4 _0972_
rlabel metal1 s 2484 20910 2484 20910 4 _0973_
rlabel metal2 s 5842 21760 5842 21760 4 _0974_
rlabel metal2 s 3266 23222 3266 23222 4 _0975_
rlabel metal2 s 12006 17850 12006 17850 4 _0976_
rlabel metal1 s 6578 18190 6578 18190 4 _0977_
rlabel metal1 s 7130 15980 7130 15980 4 _0978_
rlabel metal2 s 5750 15708 5750 15708 4 _0979_
rlabel metal2 s 14858 22338 14858 22338 4 _0980_
rlabel metal1 s 8096 20910 8096 20910 4 _0981_
rlabel metal1 s 4968 15334 4968 15334 4 _0982_
rlabel metal1 s 3266 16422 3266 16422 4 _0983_
rlabel metal1 s 5474 11730 5474 11730 4 _0984_
rlabel metal1 s 4830 12954 4830 12954 4 _0985_
rlabel metal1 s 7682 10098 7682 10098 4 _0986_
rlabel metal1 s 6118 10132 6118 10132 4 _0987_
rlabel metal1 s 11040 8806 11040 8806 4 _0988_
rlabel metal1 s 10166 9078 10166 9078 4 _0989_
rlabel metal1 s 10948 12886 10948 12886 4 _0990_
rlabel metal2 s 9706 13158 9706 13158 4 _0991_
rlabel metal1 s 5796 11662 5796 11662 4 _0992_
rlabel metal2 s 7682 35904 7682 35904 4 _0993_
rlabel metal1 s 6578 37366 6578 37366 4 _0994_
rlabel metal1 s 2530 33490 2530 33490 4 _0995_
rlabel metal1 s 7084 35666 7084 35666 4 _0996_
rlabel metal1 s 6992 32878 6992 32878 4 _0997_
rlabel metal2 s 3358 35836 3358 35836 4 _0998_
rlabel metal2 s 2346 28220 2346 28220 4 _0999_
rlabel metal1 s 3864 21998 3864 21998 4 _1000_
rlabel metal1 s 2576 19482 2576 19482 4 _1001_
rlabel metal1 s 2484 21998 2484 21998 4 _1002_
rlabel metal2 s 7590 18054 7590 18054 4 _1003_
rlabel metal2 s 6578 15334 6578 15334 4 _1004_
rlabel metal1 s 7406 22406 7406 22406 4 _1005_
rlabel metal1 s 3404 15470 3404 15470 4 _1006_
rlabel metal1 s 4600 11730 4600 11730 4 _1007_
rlabel metal1 s 6670 10642 6670 10642 4 _1008_
rlabel metal1 s 9430 10064 9430 10064 4 _1009_
rlabel metal1 s 10074 11118 10074 11118 4 _1010_
rlabel metal1 s 7912 20434 7912 20434 4 _1011_
rlabel metal1 s 5290 34034 5290 34034 4 _1012_
rlabel metal2 s 7682 38012 7682 38012 4 _1013_
rlabel metal2 s 3910 33660 3910 33660 4 _1014_
rlabel metal2 s 8970 35462 8970 35462 4 _1015_
rlabel metal1 s 8602 31790 8602 31790 4 _1016_
rlabel metal1 s 3910 36890 3910 36890 4 _1017_
rlabel metal1 s 3588 27438 3588 27438 4 _1018_
rlabel metal2 s 4094 19890 4094 19890 4 _1019_
rlabel metal1 s 3864 19822 3864 19822 4 _1020_
rlabel metal1 s 4462 23120 4462 23120 4 _1021_
rlabel metal2 s 8786 17748 8786 17748 4 _1022_
rlabel metal1 s 8004 15470 8004 15470 4 _1023_
rlabel metal2 s 8786 23290 8786 23290 4 _1024_
rlabel metal2 s 4094 14637 4094 14637 4 _1025_
rlabel metal1 s 6210 11730 6210 11730 4 _1026_
rlabel metal1 s 8648 8058 8648 8058 4 _1027_
rlabel metal1 s 11086 6766 11086 6766 4 _1028_
rlabel metal2 s 10442 13124 10442 13124 4 _1029_
rlabel metal1 s 16238 25330 16238 25330 4 _1030_
rlabel metal1 s 8510 19856 8510 19856 4 _1031_
rlabel metal3 s 8188 31756 8188 31756 4 _1032_
rlabel metal2 s 10534 38454 10534 38454 4 _1033_
rlabel metal1 s 4048 30702 4048 30702 4 _1034_
rlabel metal2 s 9614 35836 9614 35836 4 _1035_
rlabel metal1 s 9706 32844 9706 32844 4 _1036_
rlabel metal2 s 5290 37876 5290 37876 4 _1037_
rlabel metal2 s 4002 26554 4002 26554 4 _1038_
rlabel metal2 s 6302 18292 6302 18292 4 _1039_
rlabel metal1 s 6026 19346 6026 19346 4 _1040_
rlabel metal2 s 5382 22406 5382 22406 4 _1041_
rlabel metal1 s 10718 18258 10718 18258 4 _1042_
rlabel metal1 s 10258 15130 10258 15130 4 _1043_
rlabel metal1 s 10304 21522 10304 21522 4 _1044_
rlabel metal1 s 4968 16762 4968 16762 4 _1045_
rlabel metal1 s 7452 12410 7452 12410 4 _1046_
rlabel metal2 s 7314 8092 7314 8092 4 _1047_
rlabel metal2 s 11730 8262 11730 8262 4 _1048_
rlabel metal2 s 11730 13124 11730 13124 4 _1049_
rlabel metal1 s 14306 26350 14306 26350 4 _1050_
rlabel metal1 s 14904 17714 14904 17714 4 _1051_
rlabel metal1 s 16468 37774 16468 37774 4 _1052_
rlabel metal2 s 20930 38522 20930 38522 4 _1053_
rlabel metal2 s 15686 29818 15686 29818 4 _1054_
rlabel metal1 s 14352 37978 14352 37978 4 _1055_
rlabel metal1 s 22908 32878 22908 32878 4 _1056_
rlabel metal1 s 21896 36142 21896 36142 4 _1057_
rlabel metal2 s 21850 28356 21850 28356 4 _1058_
rlabel metal1 s 14628 21862 14628 21862 4 _1059_
rlabel metal1 s 13248 20434 13248 20434 4 _1060_
rlabel metal1 s 14766 23290 14766 23290 4 _1061_
rlabel metal2 s 13110 18598 13110 18598 4 _1062_
rlabel metal1 s 12213 16082 12213 16082 4 _1063_
rlabel metal1 s 13708 21998 13708 21998 4 _1064_
rlabel metal1 s 12788 14994 12788 14994 4 _1065_
rlabel metal1 s 14628 12410 14628 12410 4 _1066_
rlabel metal2 s 14306 8092 14306 8092 4 _1067_
rlabel metal2 s 14582 8466 14582 8466 4 _1068_
rlabel metal1 s 14076 10642 14076 10642 4 _1069_
rlabel metal1 s 16468 12750 16468 12750 4 _1070_
rlabel metal1 s 15410 37298 15410 37298 4 _1071_
rlabel metal2 s 19550 38012 19550 38012 4 _1072_
rlabel metal2 s 15410 29818 15410 29818 4 _1073_
rlabel metal1 s 14122 37434 14122 37434 4 _1074_
rlabel metal1 s 22126 31178 22126 31178 4 _1075_
rlabel metal1 s 20884 35666 20884 35666 4 _1076_
rlabel metal1 s 21574 27098 21574 27098 4 _1077_
rlabel metal1 s 15916 16626 15916 16626 4 _1078_
rlabel metal1 s 14996 20434 14996 20434 4 _1079_
rlabel metal1 s 16330 23834 16330 23834 4 _1080_
rlabel metal1 s 14260 17306 14260 17306 4 _1081_
rlabel metal1 s 14904 16558 14904 16558 4 _1082_
rlabel metal1 s 16146 22746 16146 22746 4 _1083_
rlabel metal2 s 15318 15266 15318 15266 4 _1084_
rlabel metal1 s 15548 12954 15548 12954 4 _1085_
rlabel metal2 s 16146 8092 16146 8092 4 _1086_
rlabel metal2 s 14858 8636 14858 8636 4 _1087_
rlabel metal1 s 15456 11118 15456 11118 4 _1088_
rlabel metal1 s 16054 3570 16054 3570 4 _1089_
rlabel metal2 s 18906 35343 18906 35343 4 _1090_
rlabel metal1 s 24656 40154 24656 40154 4 _1091_
rlabel metal1 s 18262 32876 18262 32876 4 _1092_
rlabel metal1 s 18814 40562 18814 40562 4 _1093_
rlabel metal2 s 29394 32266 29394 32266 4 _1094_
rlabel metal2 s 29394 40324 29394 40324 4 _1095_
rlabel metal1 s 29210 28050 29210 28050 4 _1096_
rlabel metal2 s 32706 13362 32706 13362 4 _1097_
rlabel metal1 s 31970 18394 31970 18394 4 _1098_
rlabel metal2 s 30498 23222 30498 23222 4 _1099_
rlabel metal2 s 28934 19652 28934 19652 4 _1100_
rlabel metal1 s 32062 13906 32062 13906 4 _1101_
rlabel metal1 s 28980 22406 28980 22406 4 _1102_
rlabel metal1 s 28428 12818 28428 12818 4 _1103_
rlabel metal1 s 29486 3366 29486 3366 4 _1104_
rlabel metal1 s 30590 5338 30590 5338 4 _1105_
rlabel metal1 s 14490 3468 14490 3468 4 _1106_
rlabel metal2 s 26726 6222 26726 6222 4 _1107_
rlabel metal1 s 18170 18224 18170 18224 4 _1108_
rlabel metal2 s 19182 36261 19182 36261 4 _1109_
rlabel metal1 s 21666 37910 21666 37910 4 _1110_
rlabel metal2 s 18446 29274 18446 29274 4 _1111_
rlabel metal2 s 16518 36758 16518 36758 4 _1112_
rlabel metal1 s 25438 30770 25438 30770 4 _1113_
rlabel metal2 s 24058 35258 24058 35258 4 _1114_
rlabel metal1 s 23230 27438 23230 27438 4 _1115_
rlabel metal1 s 18538 19890 18538 19890 4 _1116_
rlabel metal1 s 17342 20026 17342 20026 4 _1117_
rlabel metal1 s 18814 24378 18814 24378 4 _1118_
rlabel metal1 s 16514 17748 16514 17748 4 _1119_
rlabel metal1 s 17480 16082 17480 16082 4 _1120_
rlabel metal1 s 17986 22746 17986 22746 4 _1121_
rlabel metal1 s 17480 15470 17480 15470 4 _1122_
rlabel metal1 s 17066 12886 17066 12886 4 _1123_
rlabel metal2 s 19090 6970 19090 6970 4 _1124_
rlabel metal2 s 17342 6154 17342 6154 4 _1125_
rlabel metal2 s 17802 10812 17802 10812 4 _1126_
rlabel metal1 s 35742 46478 35742 46478 4 _1127_
rlabel metal1 s 35236 46682 35236 46682 4 _1128_
rlabel metal2 s 37306 45934 37306 45934 4 _1129_
rlabel metal2 s 32154 42228 32154 42228 4 _1130_
rlabel metal2 s 31970 46852 31970 46852 4 _1131_
rlabel metal1 s 37030 43282 37030 43282 4 _1132_
rlabel metal1 s 3036 18190 3036 18190 4 _1133_
rlabel metal2 s 2530 25469 2530 25469 4 _1134_
rlabel metal1 s 13018 30906 13018 30906 4 _1135_
rlabel metal1 s 13018 30090 13018 30090 4 _1136_
rlabel metal1 s 2369 24650 2369 24650 4 _1137_
rlabel metal1 s 8602 28526 8602 28526 4 _1138_
rlabel metal1 s 11178 24276 11178 24276 4 _1139_
rlabel metal1 s 2116 30362 2116 30362 4 _1140_
rlabel metal1 s 5060 27642 5060 27642 4 _1141_
rlabel metal1 s 2162 40154 2162 40154 4 _1142_
rlabel metal1 s 38962 43316 38962 43316 4 _1143_
rlabel metal2 s 3358 17884 3358 17884 4 _1144_
rlabel metal1 s 20562 40698 20562 40698 4 _1145_
rlabel metal1 s 34178 44302 34178 44302 4 _1146_
rlabel metal2 s 29486 46274 29486 46274 4 _1147_
rlabel metal1 s 29624 44710 29624 44710 4 _1148_
rlabel metal1 s 30452 44846 30452 44846 4 _1149_
rlabel metal2 s 25990 43724 25990 43724 4 _1150_
rlabel metal1 s 26358 43418 26358 43418 4 _1151_
rlabel metal2 s 26450 43996 26450 43996 4 _1152_
rlabel metal1 s 33304 44506 33304 44506 4 _1153_
rlabel metal2 s 27738 44625 27738 44625 4 _1154_
rlabel metal1 s 25898 43316 25898 43316 4 _1155_
rlabel metal1 s 25898 43214 25898 43214 4 _1156_
rlabel metal1 s 26956 43350 26956 43350 4 _1157_
rlabel metal1 s 27048 43418 27048 43418 4 _1158_
rlabel metal1 s 29900 42738 29900 42738 4 _1159_
rlabel metal3 s 28658 44965 28658 44965 4 _1160_
rlabel metal1 s 26772 44370 26772 44370 4 _1161_
rlabel metal1 s 30774 45900 30774 45900 4 _1162_
rlabel metal1 s 29946 44438 29946 44438 4 _1163_
rlabel metal2 s 31142 45254 31142 45254 4 _1164_
rlabel metal2 s 31050 45152 31050 45152 4 _1165_
rlabel metal1 s 31004 44982 31004 44982 4 _1166_
rlabel metal2 s 33442 45662 33442 45662 4 _1167_
rlabel metal1 s 33764 45594 33764 45594 4 _1168_
rlabel metal1 s 33350 44914 33350 44914 4 _1169_
rlabel metal2 s 32338 45050 32338 45050 4 _1170_
rlabel metal1 s 32798 45050 32798 45050 4 _1171_
rlabel metal1 s 31142 45594 31142 45594 4 _1172_
rlabel metal1 s 30130 42670 30130 42670 4 _1173_
rlabel metal1 s 29992 42874 29992 42874 4 _1174_
rlabel metal1 s 29532 42670 29532 42670 4 _1175_
rlabel metal1 s 29670 42806 29670 42806 4 _1176_
rlabel metal1 s 30268 42534 30268 42534 4 _1177_
rlabel metal2 s 30406 43520 30406 43520 4 _1178_
rlabel metal2 s 29854 43996 29854 43996 4 _1179_
rlabel metal1 s 29992 43758 29992 43758 4 _1180_
rlabel metal1 s 29440 43826 29440 43826 4 _1181_
rlabel metal1 s 28566 43792 28566 43792 4 _1182_
rlabel metal1 s 28658 45424 28658 45424 4 _1183_
rlabel metal2 s 29210 46206 29210 46206 4 _1184_
rlabel metal2 s 29302 46240 29302 46240 4 _1185_
rlabel metal1 s 29210 45798 29210 45798 4 _1186_
rlabel metal2 s 29854 46852 29854 46852 4 _1187_
rlabel metal1 s 29348 46546 29348 46546 4 _1188_
rlabel metal1 s 29026 45492 29026 45492 4 _1189_
rlabel metal1 s 28244 45594 28244 45594 4 _1190_
rlabel metal2 s 22770 46240 22770 46240 4 _1191_
rlabel metal1 s 22954 46478 22954 46478 4 _1192_
rlabel metal2 s 23322 46002 23322 46002 4 _1193_
rlabel metal1 s 22862 46580 22862 46580 4 _1194_
rlabel metal1 s 21666 45832 21666 45832 4 _1195_
rlabel metal1 s 21712 43418 21712 43418 4 _1196_
rlabel metal1 s 21298 43350 21298 43350 4 _1197_
rlabel metal1 s 23506 45968 23506 45968 4 _1198_
rlabel metal1 s 21942 43792 21942 43792 4 _1199_
rlabel metal1 s 22816 43962 22816 43962 4 _1200_
rlabel metal2 s 21390 43588 21390 43588 4 _1201_
rlabel metal1 s 23092 42670 23092 42670 4 _1202_
rlabel metal1 s 20608 43690 20608 43690 4 _1203_
rlabel metal1 s 19412 43690 19412 43690 4 _1204_
rlabel metal1 s 21206 43282 21206 43282 4 _1205_
rlabel metal1 s 20976 44370 20976 44370 4 _1206_
rlabel metal1 s 25024 44506 25024 44506 4 _1207_
rlabel metal1 s 20654 44404 20654 44404 4 _1208_
rlabel metal2 s 21390 45050 21390 45050 4 _1209_
rlabel metal1 s 20838 44506 20838 44506 4 _1210_
rlabel metal2 s 20930 45458 20930 45458 4 _1211_
rlabel metal1 s 21022 45050 21022 45050 4 _1212_
rlabel metal2 s 21390 46580 21390 46580 4 _1213_
rlabel metal1 s 22494 45900 22494 45900 4 _1214_
rlabel metal1 s 36294 40494 36294 40494 4 _1215_
rlabel metal1 s 35052 41242 35052 41242 4 _1216_
rlabel metal1 s 35282 41480 35282 41480 4 _1217_
rlabel metal1 s 33856 41106 33856 41106 4 _1218_
rlabel metal1 s 16974 28594 16974 28594 4 _1219_
rlabel metal1 s 36386 15470 36386 15470 4 _1220_
rlabel metal1 s 13754 37264 13754 37264 4 _1221_
rlabel metal1 s 34316 36142 34316 36142 4 _1222_
rlabel metal1 s 14398 31450 14398 31450 4 _1223_
rlabel metal1 s 13294 37434 13294 37434 4 _1224_
rlabel metal1 s 34408 31790 34408 31790 4 _1225_
rlabel metal2 s 31694 33796 31694 33796 4 _1226_
rlabel metal1 s 35236 27098 35236 27098 4 _1227_
rlabel metal1 s 37858 18156 37858 18156 4 _1228_
rlabel metal1 s 35880 18394 35880 18394 4 _1229_
rlabel metal1 s 36248 23086 36248 23086 4 _1230_
rlabel metal1 s 37076 18258 37076 18258 4 _1231_
rlabel metal1 s 36800 12818 36800 12818 4 _1232_
rlabel metal2 s 36386 21692 36386 21692 4 _1233_
rlabel metal1 s 36248 13498 36248 13498 4 _1234_
rlabel metal1 s 35236 4794 35236 4794 4 _1235_
rlabel metal1 s 35558 7514 35558 7514 4 _1236_
rlabel metal2 s 21666 4998 21666 4998 4 _1237_
rlabel metal2 s 27554 4556 27554 4556 4 _1238_
rlabel metal2 s 14996 17204 14996 17204 4 _1239_
rlabel metal1 s 17434 32946 17434 32946 4 _1240_
rlabel metal2 s 24150 38522 24150 38522 4 _1241_
rlabel metal1 s 16882 32402 16882 32402 4 _1242_
rlabel metal2 s 16422 38760 16422 38760 4 _1243_
rlabel metal1 s 26312 32878 26312 32878 4 _1244_
rlabel metal1 s 27278 37876 27278 37876 4 _1245_
rlabel metal2 s 28750 27642 28750 27642 4 _1246_
rlabel metal1 s 29302 18802 29302 18802 4 _1247_
rlabel metal1 s 29486 18734 29486 18734 4 _1248_
rlabel metal2 s 27094 24004 27094 24004 4 _1249_
rlabel metal1 s 26542 16762 26542 16762 4 _1250_
rlabel metal1 s 29348 15130 29348 15130 4 _1251_
rlabel metal2 s 25254 24310 25254 24310 4 _1252_
rlabel metal1 s 26772 14994 26772 14994 4 _1253_
rlabel metal1 s 28106 9690 28106 9690 4 _1254_
rlabel metal1 s 26818 7446 26818 7446 4 _1255_
rlabel metal2 s 14122 5644 14122 5644 4 _1256_
rlabel metal1 s 24242 9044 24242 9044 4 _1257_
rlabel metal1 s 14536 17170 14536 17170 4 _1258_
rlabel metal2 s 17342 39168 17342 39168 4 _1259_
rlabel metal2 s 23230 39814 23230 39814 4 _1260_
rlabel metal1 s 16330 32402 16330 32402 4 _1261_
rlabel metal1 s 16468 38318 16468 38318 4 _1262_
rlabel metal1 s 25024 32402 25024 32402 4 _1263_
rlabel metal1 s 26634 37434 26634 37434 4 _1264_
rlabel metal1 s 26220 27438 26220 27438 4 _1265_
rlabel metal1 s 26680 17102 26680 17102 4 _1266_
rlabel metal1 s 29762 17714 29762 17714 4 _1267_
rlabel metal1 s 26312 24174 26312 24174 4 _1268_
rlabel metal1 s 25530 16558 25530 16558 4 _1269_
rlabel metal2 s 28658 14790 28658 14790 4 _1270_
rlabel metal2 s 24518 21692 24518 21692 4 _1271_
rlabel metal1 s 25576 13498 25576 13498 4 _1272_
rlabel metal1 s 27048 9146 27048 9146 4 _1273_
rlabel metal2 s 27186 7548 27186 7548 4 _1274_
rlabel metal1 s 13662 5882 13662 5882 4 _1275_
rlabel metal2 s 23138 7990 23138 7990 4 _1276_
rlabel metal1 s 37674 34714 37674 34714 4 _1277_
rlabel metal1 s 36478 36346 36478 36346 4 _1278_
rlabel metal1 s 37490 36346 37490 36346 4 _1279_
rlabel metal2 s 36432 34204 36432 34204 4 _1280_
rlabel metal1 s 17480 43418 17480 43418 4 _1281_
rlabel metal2 s 16606 43078 16606 43078 4 _1282_
rlabel metal2 s 15594 44812 15594 44812 4 _1283_
rlabel metal2 s 17158 46410 17158 46410 4 _1284_
rlabel metal2 s 7222 26826 7222 26826 4 _1285_
rlabel metal2 s 6854 25466 6854 25466 4 _1286_
rlabel metal1 s 6026 30226 6026 30226 4 _1287_
rlabel metal2 s 6394 29444 6394 29444 4 _1288_
rlabel metal1 s 10074 28594 10074 28594 4 _1289_
rlabel metal1 s 10442 28730 10442 28730 4 _1290_
rlabel metal2 s 12742 28560 12742 28560 4 _1291_
rlabel metal1 s 11960 28186 11960 28186 4 _1292_
rlabel metal2 s 10166 29036 10166 29036 4 _1293_
rlabel metal1 s 10120 26962 10120 26962 4 _1294_
rlabel metal1 s 10810 27506 10810 27506 4 _1295_
rlabel metal2 s 10810 27132 10810 27132 4 _1296_
rlabel metal1 s 37122 36176 37122 36176 4 _1297_
rlabel metal1 s 36570 36108 36570 36108 4 _1298_
rlabel metal1 s 36340 38318 36340 38318 4 _1299_
rlabel metal2 s 17802 39406 17802 39406 4 _1300_
rlabel metal1 s 9062 40052 9062 40052 4 _1301_
rlabel metal2 s 26358 46138 26358 46138 4 _1302_
rlabel metal1 s 12190 5168 12190 5168 4 _1303_
rlabel metal1 s 17664 3706 17664 3706 4 _1304_
rlabel metal1 s 34178 2414 34178 2414 4 _1305_
rlabel metal1 s 38916 37230 38916 37230 4 _1306_
rlabel metal1 s 15594 42568 15594 42568 4 _1307_
rlabel metal1 s 9108 29614 9108 29614 4 _1308_
rlabel metal1 s 11224 4590 11224 4590 4 _1309_
rlabel metal1 s 36340 43282 36340 43282 4 _1310_
rlabel metal1 s 35374 42874 35374 42874 4 _1311_
rlabel metal1 s 33810 42092 33810 42092 4 _1312_
rlabel metal1 s 39606 15402 39606 15402 4 _1313_
rlabel metal1 s 38318 19176 38318 19176 4 _1314_
rlabel metal1 s 38272 33966 38272 33966 4 _1315_
rlabel metal1 s 40112 26962 40112 26962 4 _1316_
rlabel metal1 s 39514 16082 39514 16082 4 _1317_
rlabel metal1 s 39422 15946 39422 15946 4 _1318_
rlabel metal1 s 38180 32878 38180 32878 4 _1319_
rlabel metal1 s 39606 25262 39606 25262 4 _1320_
rlabel metal2 s 39698 26044 39698 26044 4 _1321_
rlabel metal2 s 38318 27132 38318 27132 4 _1322_
rlabel metal1 s 39238 29648 39238 29648 4 _1323_
rlabel metal1 s 39146 33082 39146 33082 4 _1324_
rlabel metal2 s 41262 15028 41262 15028 4 _1325_
rlabel metal2 s 45862 16966 45862 16966 4 _1326_
rlabel metal2 s 45218 15232 45218 15232 4 _1327_
rlabel metal1 s 45678 17646 45678 17646 4 _1328_
rlabel metal2 s 46230 26996 46230 26996 4 _1329_
rlabel metal1 s 45908 26010 45908 26010 4 _1330_
rlabel metal2 s 46782 26758 46782 26758 4 _1331_
rlabel metal2 s 46782 21318 46782 21318 4 _1332_
rlabel metal2 s 46230 20230 46230 20230 4 _1333_
rlabel metal1 s 46184 17850 46184 17850 4 _1334_
rlabel metal1 s 46046 15130 46046 15130 4 _1335_
rlabel metal2 s 45494 13498 45494 13498 4 _1336_
rlabel metal2 s 44206 14076 44206 14076 4 _1337_
rlabel metal2 s 42182 14790 42182 14790 4 _1338_
rlabel metal2 s 40710 14076 40710 14076 4 _1339_
rlabel metal1 s 38686 29172 38686 29172 4 _1340_
rlabel metal1 s 43930 28050 43930 28050 4 _1341_
rlabel metal1 s 45218 27982 45218 27982 4 _1342_
rlabel metal1 s 45540 28050 45540 28050 4 _1343_
rlabel metal1 s 38594 40154 38594 40154 4 _1344_
rlabel metal2 s 38962 41242 38962 41242 4 _1345_
rlabel metal1 s 36432 41106 36432 41106 4 _1346_
rlabel metal1 s 37950 25194 37950 25194 4 _1347_
rlabel metal3 s 39261 40052 39261 40052 4 _1348_
rlabel metal1 s 38134 14586 38134 14586 4 _1349_
rlabel metal1 s 38594 22202 38594 22202 4 _1350_
rlabel metal1 s 38410 25228 38410 25228 4 _1351_
rlabel metal1 s 38180 32198 38180 32198 4 _1352_
rlabel metal1 s 38870 25296 38870 25296 4 _1353_
rlabel metal1 s 38180 38930 38180 38930 4 _1354_
rlabel metal1 s 34960 40494 34960 40494 4 _1355_
rlabel metal1 s 35604 41106 35604 41106 4 _1356_
rlabel metal1 s 35328 38318 35328 38318 4 _1357_
rlabel metal1 s 39100 40970 39100 40970 4 _1358_
rlabel metal1 s 37444 40494 37444 40494 4 _1359_
rlabel metal1 s 37444 40086 37444 40086 4 _1360_
rlabel metal1 s 34868 38318 34868 38318 4 _1361_
rlabel metal1 s 39698 40052 39698 40052 4 _1362_
rlabel metal1 s 37628 38930 37628 38930 4 _1363_
rlabel metal1 s 37674 39338 37674 39338 4 _1364_
rlabel metal1 s 36432 39950 36432 39950 4 _1365_
rlabel metal1 s 36386 39372 36386 39372 4 _1366_
rlabel metal2 s 33810 39202 33810 39202 4 _1367_
rlabel metal2 s 34454 38743 34454 38743 4 _1368_
rlabel metal1 s 37076 38386 37076 38386 4 _1369_
rlabel metal1 s 37398 38454 37398 38454 4 _1370_
rlabel metal1 s 36110 36788 36110 36788 4 _1371_
rlabel metal1 s 33534 38488 33534 38488 4 _1372_
rlabel metal1 s 7590 29682 7590 29682 4 _1373_
rlabel metal2 s 8602 26180 8602 26180 4 _1374_
rlabel metal1 s 7636 24174 7636 24174 4 _1375_
rlabel metal1 s 7176 28050 7176 28050 4 _1376_
rlabel metal1 s 7682 28084 7682 28084 4 _1377_
rlabel metal2 s 21758 16881 21758 16881 4 _1378_
rlabel metal1 s 18722 26962 18722 26962 4 _1379_
rlabel metal3 s 19320 15164 19320 15164 4 _1380_
rlabel metal1 s 18400 28050 18400 28050 4 _1381_
rlabel metal2 s 18446 38148 18446 38148 4 _1382_
rlabel metal2 s 23690 36958 23690 36958 4 _1383_
rlabel metal1 s 27554 35700 27554 35700 4 _1384_
rlabel metal2 s 11178 19652 11178 19652 4 _1385_
rlabel metal2 s 4922 17714 4922 17714 4 _1386_
rlabel metal2 s 11730 19006 11730 19006 4 _1387_
rlabel metal1 s 5934 19890 5934 19890 4 _1388_
rlabel metal1 s 19688 36074 19688 36074 4 _1389_
rlabel metal2 s 20930 29920 20930 29920 4 _1390_
rlabel metal1 s 20516 18734 20516 18734 4 _1391_
rlabel metal1 s 21160 20434 21160 20434 4 _1392_
rlabel metal1 s 21160 20502 21160 20502 4 _1393_
rlabel metal1 s 27002 35530 27002 35530 4 _1394_
rlabel metal1 s 30544 19890 30544 19890 4 _1395_
rlabel metal4 s 20355 16524 20355 16524 4 _1396_
rlabel metal3 s 20999 16524 20999 16524 4 _1397_
rlabel metal2 s 26450 36584 26450 36584 4 _1398_
rlabel metal1 s 26910 35666 26910 35666 4 _1399_
rlabel metal1 s 33672 18122 33672 18122 4 _1400_
rlabel metal2 s 33350 35360 33350 35360 4 _1401_
rlabel metal1 s 32867 35802 32867 35802 4 _1402_
rlabel metal1 s 31142 19346 31142 19346 4 _1403_
rlabel metal1 s 29670 34578 29670 34578 4 _1404_
rlabel metal1 s 27416 35258 27416 35258 4 _1405_
rlabel metal1 s 7038 12648 7038 12648 4 _1406_
rlabel metal1 s 7682 12750 7682 12750 4 _1407_
rlabel metal1 s 16882 32538 16882 32538 4 _1408_
rlabel metal1 s 21758 16082 21758 16082 4 _1409_
rlabel metal1 s 21068 31314 21068 31314 4 _1410_
rlabel metal1 s 21298 30702 21298 30702 4 _1411_
rlabel metal1 s 19044 15946 19044 15946 4 _1412_
rlabel metal1 s 19826 16014 19826 16014 4 _1413_
rlabel metal2 s 21022 31246 21022 31246 4 _1414_
rlabel metal2 s 21114 31008 21114 31008 4 _1415_
rlabel metal2 s 21574 31909 21574 31909 4 _1416_
rlabel metal1 s 20424 31314 20424 31314 4 _1417_
rlabel metal1 s 21482 23698 21482 23698 4 _1418_
rlabel metal2 s 10166 22015 10166 22015 4 _1419_
rlabel metal3 s 10718 21981 10718 21981 4 _1420_
rlabel metal1 s 19826 29750 19826 29750 4 _1421_
rlabel metal2 s 20746 30566 20746 30566 4 _1422_
rlabel metal1 s 19504 36618 19504 36618 4 _1423_
rlabel metal2 s 19734 36108 19734 36108 4 _1424_
rlabel metal1 s 19780 36006 19780 36006 4 _1425_
rlabel metal1 s 20056 35530 20056 35530 4 _1426_
rlabel metal1 s 17664 20978 17664 20978 4 _1427_
rlabel metal1 s 18630 12274 18630 12274 4 _1428_
rlabel metal1 s 17664 36074 17664 36074 4 _1429_
rlabel metal3 s 21574 33915 21574 33915 4 _1430_
rlabel metal1 s 19366 6800 19366 6800 4 _1431_
rlabel metal2 s 13754 35700 13754 35700 4 _1432_
rlabel metal1 s 21206 19856 21206 19856 4 _1433_
rlabel metal2 s 19458 36006 19458 36006 4 _1434_
rlabel metal1 s 19182 30056 19182 30056 4 _1435_
rlabel metal1 s 21436 13498 21436 13498 4 _1436_
rlabel metal2 s 21206 29920 21206 29920 4 _1437_
rlabel metal2 s 25530 29886 25530 29886 4 _1438_
rlabel metal2 s 25714 29920 25714 29920 4 _1439_
rlabel metal1 s 21942 8908 21942 8908 4 _1440_
rlabel metal1 s 28750 32198 28750 32198 4 _1441_
rlabel metal1 s 33672 20366 33672 20366 4 _1442_
rlabel metal2 s 34638 14943 34638 14943 4 _1443_
rlabel metal1 s 32062 30056 32062 30056 4 _1444_
rlabel metal1 s 27876 21454 27876 21454 4 _1445_
rlabel metal2 s 25898 30396 25898 30396 4 _1446_
rlabel metal1 s 27048 35190 27048 35190 4 _1447_
rlabel metal1 s 29394 35122 29394 35122 4 _1448_
rlabel metal2 s 20194 35411 20194 35411 4 _1449_
rlabel metal1 s 25162 35156 25162 35156 4 _1450_
rlabel metal1 s 28842 35564 28842 35564 4 _1451_
rlabel metal2 s 29026 35258 29026 35258 4 _1452_
rlabel metal2 s 29762 34816 29762 34816 4 _1453_
rlabel metal1 s 29256 34714 29256 34714 4 _1454_
rlabel metal2 s 21482 26639 21482 26639 4 _1455_
rlabel metal1 s 21597 27030 21597 27030 4 _1456_
rlabel metal1 s 25254 27914 25254 27914 4 _1457_
rlabel metal1 s 25668 26894 25668 26894 4 _1458_
rlabel metal1 s 31004 27642 31004 27642 4 _1459_
rlabel metal2 s 34546 27744 34546 27744 4 _1460_
rlabel metal1 s 25530 26894 25530 26894 4 _1461_
rlabel metal2 s 19274 20536 19274 20536 4 _1462_
rlabel metal1 s 30130 20502 30130 20502 4 _1463_
rlabel metal2 s 6394 19550 6394 19550 4 _1464_
rlabel metal3 s 23322 20315 23322 20315 4 _1465_
rlabel metal2 s 31142 19176 31142 19176 4 _1466_
rlabel metal1 s 30360 20026 30360 20026 4 _1467_
rlabel metal1 s 46046 27098 46046 27098 4 _1468_
rlabel metal1 s 45862 26860 45862 26860 4 _1469_
rlabel metal2 s 46230 28866 46230 28866 4 _1470_
rlabel metal1 s 39606 33388 39606 33388 4 _1471_
rlabel metal1 s 39376 29818 39376 29818 4 _1472_
rlabel metal1 s 38272 27098 38272 27098 4 _1473_
rlabel metal2 s 40342 25466 40342 25466 4 _1474_
rlabel metal2 s 40066 24650 40066 24650 4 _1475_
rlabel metal2 s 45770 21148 45770 21148 4 _1476_
rlabel metal1 s 45494 20332 45494 20332 4 _1477_
rlabel metal2 s 45862 18428 45862 18428 4 _1478_
rlabel metal1 s 46000 15674 46000 15674 4 _1479_
rlabel metal2 s 45126 12988 45126 12988 4 _1480_
rlabel metal1 s 43746 13906 43746 13906 4 _1481_
rlabel metal2 s 41170 14348 41170 14348 4 _1482_
rlabel metal2 s 40158 14212 40158 14212 4 _1483_
rlabel metal1 s 38824 47634 38824 47634 4 clock
rlabel metal1 s 3404 47770 3404 47770 4 led_clock
rlabel metal2 s 10626 48739 10626 48739 4 leds[0]
rlabel metal2 s 32246 1520 32246 1520 4 leds[1]
rlabel metal3 s 820 14348 820 14348 4 leds[2]
rlabel metal3 s 820 44268 820 44268 4 leds[3]
rlabel metal1 s 36202 19482 36202 19482 4 net1
rlabel metal2 s 6118 47906 6118 47906 4 net10
rlabel metal1 s 18998 6154 18998 6154 4 net100
rlabel metal2 s 16790 7072 16790 7072 4 net101
rlabel metal1 s 14766 8398 14766 8398 4 net102
rlabel metal1 s 19780 13906 19780 13906 4 net103
rlabel metal1 s 16790 13294 16790 13294 4 net104
rlabel metal2 s 10258 14280 10258 14280 4 net105
rlabel metal1 s 2254 16966 2254 16966 4 net106
rlabel metal1 s 6210 17578 6210 17578 4 net107
rlabel metal1 s 4922 20910 4922 20910 4 net108
rlabel metal2 s 7222 21794 7222 21794 4 net109
rlabel metal3 s 1702 31875 1702 31875 4 net11
rlabel metal2 s 5704 21828 5704 21828 4 net110
rlabel metal1 s 9890 18190 9890 18190 4 net111
rlabel metal1 s 12834 18258 12834 18258 4 net112
rlabel metal2 s 16974 15776 16974 15776 4 net113
rlabel metal1 s 13524 20910 13524 20910 4 net114
rlabel metal1 s 17434 20434 17434 20434 4 net115
rlabel metal1 s 18308 19346 18308 19346 4 net116
rlabel metal1 s 18446 14382 18446 14382 4 net117
rlabel metal2 s 21850 4080 21850 4080 4 net118
rlabel metal1 s 29440 5746 29440 5746 4 net119
rlabel metal1 s 32890 30804 32890 30804 4 net12
rlabel metal1 s 24104 7378 24104 7378 4 net120
rlabel metal1 s 27508 13294 27508 13294 4 net121
rlabel metal1 s 28750 12750 28750 12750 4 net122
rlabel metal1 s 29348 13430 29348 13430 4 net123
rlabel metal1 s 32200 8942 32200 8942 4 net124
rlabel metal2 s 34822 4624 34822 4624 4 net125
rlabel metal1 s 38640 8806 38640 8806 4 net126
rlabel metal2 s 35742 13821 35742 13821 4 net127
rlabel metal1 s 27554 15470 27554 15470 4 net128
rlabel metal1 s 29532 19822 29532 19822 4 net129
rlabel metal3 s 1702 29699 1702 29699 4 net13
rlabel metal1 s 27692 21998 27692 21998 4 net130
rlabel metal1 s 29348 19890 29348 19890 4 net131
rlabel metal1 s 31878 16082 31878 16082 4 net132
rlabel metal2 s 31970 20366 31970 20366 4 net133
rlabel metal1 s 30314 24718 30314 24718 4 net134
rlabel metal1 s 37076 21454 37076 21454 4 net135
rlabel metal1 s 36340 14994 36340 14994 4 net136
rlabel metal1 s 1794 25262 1794 25262 4 net137
rlabel metal2 s 9982 29648 9982 29648 4 net138
rlabel metal1 s 4738 29070 4738 29070 4 net139
rlabel metal3 s 46230 2499 46230 2499 4 net14
rlabel metal1 s 2346 36210 2346 36210 4 net140
rlabel metal2 s 6578 34816 6578 34816 4 net141
rlabel metal2 s 4002 34816 4002 34816 4 net142
rlabel metal1 s 12880 34510 12880 34510 4 net143
rlabel metal1 s 16652 32334 16652 32334 4 net144
rlabel metal1 s 19044 33286 19044 33286 4 net145
rlabel metal2 s 18538 35326 18538 35326 4 net146
rlabel metal2 s 11546 40460 11546 40460 4 net147
rlabel metal1 s 9062 38284 9062 38284 4 net148
rlabel metal1 s 3956 47022 3956 47022 4 net149
rlabel metal2 s 45678 2329 45678 2329 4 net15
rlabel metal1 s 13570 37876 13570 37876 4 net150
rlabel metal1 s 19182 38318 19182 38318 4 net151
rlabel metal1 s 20286 43860 20286 43860 4 net152
rlabel metal1 s 18860 46002 18860 46002 4 net153
rlabel metal1 s 17066 35734 17066 35734 4 net154
rlabel metal1 s 11086 41514 11086 41514 4 net155
rlabel metal1 s 20562 27438 20562 27438 4 net156
rlabel metal1 s 29072 28662 29072 28662 4 net157
rlabel metal1 s 21850 35564 21850 35564 4 net158
rlabel metal1 s 29072 35666 29072 35666 4 net159
rlabel metal3 s 35075 23188 35075 23188 4 net16
rlabel metal1 s 29578 36074 29578 36074 4 net160
rlabel metal1 s 38134 34442 38134 34442 4 net161
rlabel metal2 s 36018 34272 36018 34272 4 net162
rlabel metal2 s 36294 35972 36294 35972 4 net163
rlabel metal1 s 21804 41038 21804 41038 4 net164
rlabel metal1 s 29026 38386 29026 38386 4 net165
rlabel metal1 s 21022 47090 21022 47090 4 net166
rlabel metal1 s 27048 46546 27048 46546 4 net167
rlabel metal1 s 26680 38318 26680 38318 4 net168
rlabel metal1 s 34730 37264 34730 37264 4 net169
rlabel metal2 s 45678 46954 45678 46954 4 net17
rlabel metal2 s 33074 39678 33074 39678 4 net170
rlabel metal1 s 32246 43758 32246 43758 4 net171
rlabel metal1 s 35926 46002 35926 46002 4 net172
rlabel metal1 s 38364 38998 38364 38998 4 net173
rlabel metal1 s 39146 35054 39146 35054 4 net174
rlabel metal1 s 18170 25908 18170 25908 4 net175
rlabel metal2 s 39606 43078 39606 43078 4 net176
rlabel metal1 s 39233 8534 39233 8534 4 net177
rlabel metal1 s 18844 46954 18844 46954 4 net178
rlabel metal1 s 38221 4182 38221 4182 4 net179
rlabel metal1 s 1932 37094 1932 37094 4 net18
rlabel metal1 s 4968 46546 4968 46546 4 net180
rlabel metal1 s 27503 3094 27503 3094 4 net181
rlabel metal1 s 24456 46954 24456 46954 4 net182
rlabel metal1 s 6256 2618 6256 2618 4 net19
rlabel metal2 s 43102 35880 43102 35880 4 net2
rlabel metal1 s 2576 2550 2576 2550 4 net20
rlabel metal2 s 46598 45322 46598 45322 4 net21
rlabel metal1 s 1840 17306 1840 17306 4 net22
rlabel metal3 s 20769 2652 20769 2652 4 net23
rlabel metal1 s 37766 45356 37766 45356 4 net24
rlabel metal4 s 32637 41412 32637 41412 4 net25
rlabel metal1 s 15295 47498 15295 47498 4 net26
rlabel metal4 s 37789 42908 37789 42908 4 net27
rlabel metal3 s 11569 2652 11569 2652 4 net28
rlabel metal1 s 16974 2380 16974 2380 4 net29
rlabel metal2 s 1610 20893 1610 20893 4 net3
rlabel metal1 s 1932 21862 1932 21862 4 net30
rlabel metal3 s 9430 28475 9430 28475 4 net31
rlabel metal1 s 21022 2516 21022 2516 4 net32
rlabel metal2 s 38870 46138 38870 46138 4 net33
rlabel metal2 s 46874 36215 46874 36215 4 net34
rlabel metal1 s 36294 34714 36294 34714 4 net35
rlabel metal1 s 38456 21930 38456 21930 4 net36
rlabel metal1 s 44068 33082 44068 33082 4 net37
rlabel metal1 s 38456 14382 38456 14382 4 net38
rlabel metal1 s 38272 14314 38272 14314 4 net39
rlabel metal3 s 1702 12733 1702 12733 4 net4
rlabel metal1 s 46690 35666 46690 35666 4 net40
rlabel metal1 s 1426 2380 1426 2380 4 net41
rlabel metal1 s 43746 32810 43746 32810 4 net42
rlabel metal2 s 42182 34391 42182 34391 4 net43
rlabel metal1 s 39882 31926 39882 31926 4 net44
rlabel metal1 s 36248 33286 36248 33286 4 net45
rlabel metal3 s 2254 9979 2254 9979 4 net46
rlabel metal1 s 46046 40494 46046 40494 4 net47
rlabel metal1 s 1702 41582 1702 41582 4 net48
rlabel metal2 s 21206 19737 21206 19737 4 net49
rlabel metal2 s 37674 5508 37674 5508 4 net5
rlabel metal2 s 2208 20332 2208 20332 4 net50
rlabel metal1 s 4646 2482 4646 2482 4 net51
rlabel metal1 s 27324 47226 27324 47226 4 net52
rlabel metal1 s 18768 2414 18768 2414 4 net53
rlabel metal1 s 35098 3162 35098 3162 4 net54
rlabel metal2 s 44206 37366 44206 37366 4 net55
rlabel metal1 s 15180 43418 15180 43418 4 net56
rlabel metal2 s 4140 21420 4140 21420 4 net57
rlabel metal2 s 11362 3706 11362 3706 4 net58
rlabel metal3 s 36823 2652 36823 2652 4 net59
rlabel metal2 s 36478 5780 36478 5780 4 net6
rlabel metal1 s 34408 39066 34408 39066 4 net60
rlabel metal1 s 28428 43962 28428 43962 4 net61
rlabel metal1 s 25852 46342 25852 46342 4 net62
rlabel metal2 s 6026 46750 6026 46750 4 net63
rlabel metal3 s 39238 3995 39238 3995 4 net64
rlabel metal1 s 18998 47226 18998 47226 4 net65
rlabel metal2 s 39882 9571 39882 9571 4 net66
rlabel metal2 s 40434 43367 40434 43367 4 net67
rlabel metal2 s 30866 44812 30866 44812 4 net68
rlabel metal2 s 1518 37128 1518 37128 4 net69
rlabel metal1 s 39100 2618 39100 2618 4 net7
rlabel metal1 s 18630 47600 18630 47600 4 net70
rlabel metal1 s 22034 43248 22034 43248 4 net71
rlabel metal1 s 1426 5270 1426 5270 4 net72
rlabel metal3 s 2254 2907 2254 2907 4 net73
rlabel metal2 s 2668 40052 2668 40052 4 net74
rlabel metal2 s 20378 46784 20378 46784 4 net75
rlabel metal2 s 32246 47430 32246 47430 4 net76
rlabel metal1 s 41446 47600 41446 47600 4 net77
rlabel metal2 s 3082 47430 3082 47430 4 net78
rlabel metal2 s 2622 40256 2622 40256 4 net79
rlabel metal3 s 40181 2652 40181 2652 4 net8
rlabel metal1 s 32338 2448 32338 2448 4 net80
rlabel metal1 s 3082 18326 3082 18326 4 net81
rlabel metal1 s 35742 41718 35742 41718 4 net82
rlabel metal2 s 2070 31212 2070 31212 4 net83
rlabel metal2 s 38410 25976 38410 25976 4 net84
rlabel metal1 s 20102 17102 20102 17102 4 net85
rlabel metal2 s 37306 15997 37306 15997 4 net86
rlabel metal1 s 35926 31790 35926 31790 4 net87
rlabel metal1 s 37858 20026 37858 20026 4 net88
rlabel metal2 s 38042 18938 38042 18938 4 net89
rlabel metal1 s 36202 30804 36202 30804 4 net9
rlabel metal1 s 38778 34578 38778 34578 4 net90
rlabel metal2 s 35834 34170 35834 34170 4 net91
rlabel metal3 s 34339 2516 34339 2516 4 net92
rlabel metal1 s 2254 39542 2254 39542 4 net93
rlabel metal2 s 1426 43316 1426 43316 4 net94
rlabel metal2 s 3082 18207 3082 18207 4 net95
rlabel metal1 s 3772 12274 3772 12274 4 net96
rlabel metal1 s 6486 13430 6486 13430 4 net97
rlabel metal1 s 9936 5202 9936 5202 4 net98
rlabel metal1 s 13892 4046 13892 4046 4 net99
rlabel metal2 s 44206 34374 44206 34374 4 po_0._1_\[0\]
rlabel metal2 s 41078 19278 41078 19278 4 po_0._1_\[10\]
rlabel metal1 s 40250 17136 40250 17136 4 po_0._1_\[11\]
rlabel metal2 s 38594 11390 38594 11390 4 po_0._1_\[12\]
rlabel metal2 s 40802 9316 40802 9316 4 po_0._1_\[13\]
rlabel metal2 s 38134 9996 38134 9996 4 po_0._1_\[14\]
rlabel metal2 s 37950 10948 37950 10948 4 po_0._1_\[15\]
rlabel metal2 s 45034 32164 45034 32164 4 po_0._1_\[1\]
rlabel metal2 s 41262 35020 41262 35020 4 po_0._1_\[2\]
rlabel metal1 s 40480 32402 40480 32402 4 po_0._1_\[3\]
rlabel metal2 s 41538 27438 41538 27438 4 po_0._1_\[4\]
rlabel metal2 s 37122 26520 37122 26520 4 po_0._1_\[5\]
rlabel metal1 s 41262 21862 41262 21862 4 po_0._1_\[6\]
rlabel metal2 s 43746 23324 43746 23324 4 po_0._1_\[7\]
rlabel metal1 s 40894 19380 40894 19380 4 po_0._1_\[8\]
rlabel metal2 s 40526 19333 40526 19333 4 po_0._1_\[9\]
rlabel metal2 s 45494 27676 45494 27676 4 po_0.alu_0._10_\[0\]
rlabel metal1 s 45540 18190 45540 18190 4 po_0.alu_0._10_\[10\]
rlabel metal2 s 45402 16422 45402 16422 4 po_0.alu_0._10_\[11\]
rlabel metal1 s 44712 11662 44712 11662 4 po_0.alu_0._10_\[12\]
rlabel metal1 s 43010 12954 43010 12954 4 po_0.alu_0._10_\[13\]
rlabel metal1 s 40894 12750 40894 12750 4 po_0.alu_0._10_\[14\]
rlabel metal1 s 39790 12954 39790 12954 4 po_0.alu_0._10_\[15\]
rlabel metal1 s 45724 26962 45724 26962 4 po_0.alu_0._10_\[1\]
rlabel metal1 s 45816 30226 45816 30226 4 po_0.alu_0._10_\[2\]
rlabel metal1 s 39790 33490 39790 33490 4 po_0.alu_0._10_\[3\]
rlabel metal1 s 40250 29274 40250 29274 4 po_0.alu_0._10_\[4\]
rlabel metal2 s 38778 27574 38778 27574 4 po_0.alu_0._10_\[5\]
rlabel metal1 s 44160 24650 44160 24650 4 po_0.alu_0._10_\[6\]
rlabel metal1 s 42366 24276 42366 24276 4 po_0.alu_0._10_\[7\]
rlabel metal1 s 45218 20978 45218 20978 4 po_0.alu_0._10_\[8\]
rlabel metal1 s 44988 19278 44988 19278 4 po_0.alu_0._10_\[9\]
rlabel metal1 s 45770 27642 45770 27642 4 po_0.alu_0._11_\[0\]
rlabel metal1 s 41170 18292 41170 18292 4 po_0.alu_0._11_\[10\]
rlabel metal1 s 42642 15980 42642 15980 4 po_0.alu_0._11_\[11\]
rlabel metal1 s 44942 12614 44942 12614 4 po_0.alu_0._11_\[12\]
rlabel metal2 s 43286 13498 43286 13498 4 po_0.alu_0._11_\[13\]
rlabel metal2 s 40986 14212 40986 14212 4 po_0.alu_0._11_\[14\]
rlabel metal2 s 39698 14688 39698 14688 4 po_0.alu_0._11_\[15\]
rlabel metal1 s 44758 28084 44758 28084 4 po_0.alu_0._11_\[1\]
rlabel metal1 s 42573 30226 42573 30226 4 po_0.alu_0._11_\[2\]
rlabel metal2 s 40066 31994 40066 31994 4 po_0.alu_0._11_\[3\]
rlabel metal1 s 40618 30192 40618 30192 4 po_0.alu_0._11_\[4\]
rlabel metal1 s 38134 27506 38134 27506 4 po_0.alu_0._11_\[5\]
rlabel metal2 s 40894 24956 40894 24956 4 po_0.alu_0._11_\[6\]
rlabel metal1 s 39882 24378 39882 24378 4 po_0.alu_0._11_\[7\]
rlabel metal1 s 43746 20978 43746 20978 4 po_0.alu_0._11_\[8\]
rlabel metal1 s 41170 20468 41170 20468 4 po_0.alu_0._11_\[9\]
rlabel metal1 s 39100 33286 39100 33286 4 po_0.alu_0.s0
rlabel metal1 s 39790 21318 39790 21318 4 po_0.alu_0.s1
rlabel metal1 s 35098 45934 35098 45934 4 po_0.muxf_0.rf_w_data\[0\]
rlabel metal2 s 36754 45662 36754 45662 4 po_0.muxf_0.rf_w_data\[1\]
rlabel metal1 s 30590 41514 30590 41514 4 po_0.muxf_0.rf_w_data\[2\]
rlabel metal2 s 34684 17068 34684 17068 4 po_0.muxf_0.rf_w_data\[3\]
rlabel metal2 s 23138 45390 23138 45390 4 po_0.muxf_0.rf_w_data\[4\]
rlabel metal1 s 16376 42194 16376 42194 4 po_0.muxf_0.rf_w_data\[5\]
rlabel metal1 s 15318 43758 15318 43758 4 po_0.muxf_0.rf_w_data\[6\]
rlabel metal1 s 3588 43690 3588 43690 4 po_0.muxf_0.rf_w_data\[7\]
rlabel metal2 s 37398 35700 37398 35700 4 po_0.muxf_0.s0
rlabel metal1 s 36984 35802 36984 35802 4 po_0.muxf_0.s1
rlabel metal2 s 33074 34731 33074 34731 4 po_0.regf_0._3_\[0\]
rlabel metal1 s 25576 22678 25576 22678 4 po_0.regf_0._3_\[10\]
rlabel metal2 s 37582 16031 37582 16031 4 po_0.regf_0._3_\[11\]
rlabel metal1 s 20194 12172 20194 12172 4 po_0.regf_0._3_\[12\]
rlabel metal1 s 34086 11016 34086 11016 4 po_0.regf_0._3_\[13\]
rlabel metal1 s 34178 10098 34178 10098 4 po_0.regf_0._3_\[14\]
rlabel metal2 s 20102 10438 20102 10438 4 po_0.regf_0._3_\[15\]
rlabel metal2 s 36018 32589 36018 32589 4 po_0.regf_0._3_\[1\]
rlabel metal3 s 14122 35003 14122 35003 4 po_0.regf_0._3_\[2\]
rlabel metal2 s 31878 31008 31878 31008 4 po_0.regf_0._3_\[3\]
rlabel metal1 s 32430 33524 32430 33524 4 po_0.regf_0._3_\[4\]
rlabel metal2 s 23414 25466 23414 25466 4 po_0.regf_0._3_\[5\]
rlabel metal1 s 33534 20910 33534 20910 4 po_0.regf_0._3_\[6\]
rlabel metal1 s 22310 24378 22310 24378 4 po_0.regf_0._3_\[7\]
rlabel metal1 s 20470 19788 20470 19788 4 po_0.regf_0._3_\[8\]
rlabel metal2 s 20378 17000 20378 17000 4 po_0.regf_0._3_\[9\]
rlabel metal2 s 39882 35139 39882 35139 4 po_0.regf_0._5_\[0\]
rlabel metal2 s 40158 21165 40158 21165 4 po_0.regf_0._5_\[10\]
rlabel metal1 s 37214 15436 37214 15436 4 po_0.regf_0._5_\[11\]
rlabel metal2 s 35926 11356 35926 11356 4 po_0.regf_0._5_\[12\]
rlabel metal1 s 36570 9384 36570 9384 4 po_0.regf_0._5_\[13\]
rlabel metal2 s 21758 8670 21758 8670 4 po_0.regf_0._5_\[14\]
rlabel metal2 s 36018 10863 36018 10863 4 po_0.regf_0._5_\[15\]
rlabel metal1 s 37858 31790 37858 31790 4 po_0.regf_0._5_\[1\]
rlabel metal3 s 19182 35581 19182 35581 4 po_0.regf_0._5_\[2\]
rlabel metal2 s 28290 29920 28290 29920 4 po_0.regf_0._5_\[3\]
rlabel metal2 s 40158 35105 40158 35105 4 po_0.regf_0._5_\[4\]
rlabel metal1 s 33074 26520 33074 26520 4 po_0.regf_0._5_\[5\]
rlabel metal1 s 32062 20264 32062 20264 4 po_0.regf_0._5_\[6\]
rlabel metal1 s 38364 23698 38364 23698 4 po_0.regf_0._5_\[7\]
rlabel metal1 s 38870 19380 38870 19380 4 po_0.regf_0._5_\[8\]
rlabel metal1 s 32154 15946 32154 15946 4 po_0.regf_0._5_\[9\]
rlabel metal1 s 25622 40154 25622 40154 4 po_0.regf_0.rf\[0\]\[0\]
rlabel metal2 s 29486 21216 29486 21216 4 po_0.regf_0.rf\[0\]\[10\]
rlabel metal1 s 27140 13838 27140 13838 4 po_0.regf_0.rf\[0\]\[11\]
rlabel metal1 s 29486 10030 29486 10030 4 po_0.regf_0.rf\[0\]\[12\]
rlabel metal1 s 29716 7854 29716 7854 4 po_0.regf_0.rf\[0\]\[13\]
rlabel metal2 s 15502 3264 15502 3264 4 po_0.regf_0.rf\[0\]\[14\]
rlabel metal2 s 24610 9248 24610 9248 4 po_0.regf_0.rf\[0\]\[15\]
rlabel metal1 s 19734 32742 19734 32742 4 po_0.regf_0.rf\[0\]\[1\]
rlabel metal2 s 18262 40732 18262 40732 4 po_0.regf_0.rf\[0\]\[2\]
rlabel metal2 s 27186 32096 27186 32096 4 po_0.regf_0.rf\[0\]\[3\]
rlabel metal1 s 29302 39916 29302 39916 4 po_0.regf_0.rf\[0\]\[4\]
rlabel metal1 s 29900 28186 29900 28186 4 po_0.regf_0.rf\[0\]\[5\]
rlabel metal2 s 32614 18496 32614 18496 4 po_0.regf_0.rf\[0\]\[6\]
rlabel metal1 s 28106 23596 28106 23596 4 po_0.regf_0.rf\[0\]\[7\]
rlabel metal1 s 25760 19822 25760 19822 4 po_0.regf_0.rf\[0\]\[8\]
rlabel metal1 s 32936 13906 32936 13906 4 po_0.regf_0.rf\[0\]\[9\]
rlabel metal2 s 20470 37434 20470 37434 4 po_0.regf_0.rf\[10\]\[0\]
rlabel metal2 s 20758 22066 20758 22066 4 po_0.regf_0.rf\[10\]\[10\]
rlabel metal1 s 20493 14926 20493 14926 4 po_0.regf_0.rf\[10\]\[11\]
rlabel metal2 s 16146 13056 16146 13056 4 po_0.regf_0.rf\[10\]\[12\]
rlabel metal2 s 17158 8466 17158 8466 4 po_0.regf_0.rf\[10\]\[13\]
rlabel metal1 s 15962 8602 15962 8602 4 po_0.regf_0.rf\[10\]\[14\]
rlabel metal1 s 16100 10778 16100 10778 4 po_0.regf_0.rf\[10\]\[15\]
rlabel metal1 s 16238 29274 16238 29274 4 po_0.regf_0.rf\[10\]\[1\]
rlabel metal1 s 14812 37230 14812 37230 4 po_0.regf_0.rf\[10\]\[2\]
rlabel metal2 s 24622 31246 24622 31246 4 po_0.regf_0.rf\[10\]\[3\]
rlabel metal1 s 22080 35190 22080 35190 4 po_0.regf_0.rf\[10\]\[4\]
rlabel metal1 s 22402 26962 22402 26962 4 po_0.regf_0.rf\[10\]\[5\]
rlabel metal2 s 15870 20672 15870 20672 4 po_0.regf_0.rf\[10\]\[6\]
rlabel metal2 s 17434 23936 17434 23936 4 po_0.regf_0.rf\[10\]\[7\]
rlabel metal1 s 15801 18190 15801 18190 4 po_0.regf_0.rf\[10\]\[8\]
rlabel metal2 s 19378 16082 19378 16082 4 po_0.regf_0.rf\[10\]\[9\]
rlabel metal2 s 20654 38726 20654 38726 4 po_0.regf_0.rf\[11\]\[0\]
rlabel metal1 s 20470 22508 20470 22508 4 po_0.regf_0.rf\[11\]\[10\]
rlabel metal2 s 20102 15266 20102 15266 4 po_0.regf_0.rf\[11\]\[11\]
rlabel metal1 s 17986 12750 17986 12750 4 po_0.regf_0.rf\[11\]\[12\]
rlabel metal2 s 13938 8262 13938 8262 4 po_0.regf_0.rf\[11\]\[13\]
rlabel metal2 s 13846 8160 13846 8160 4 po_0.regf_0.rf\[11\]\[14\]
rlabel metal1 s 15410 10166 15410 10166 4 po_0.regf_0.rf\[11\]\[15\]
rlabel metal1 s 17112 29818 17112 29818 4 po_0.regf_0.rf\[11\]\[1\]
rlabel metal1 s 15456 37978 15456 37978 4 po_0.regf_0.rf\[11\]\[2\]
rlabel metal2 s 24472 31246 24472 31246 4 po_0.regf_0.rf\[11\]\[3\]
rlabel metal1 s 22770 35802 22770 35802 4 po_0.regf_0.rf\[11\]\[4\]
rlabel metal1 s 22632 27642 22632 27642 4 po_0.regf_0.rf\[11\]\[5\]
rlabel metal2 s 18032 20910 18032 20910 4 po_0.regf_0.rf\[11\]\[6\]
rlabel metal2 s 15134 23256 15134 23256 4 po_0.regf_0.rf\[11\]\[7\]
rlabel metal2 s 13938 18122 13938 18122 4 po_0.regf_0.rf\[11\]\[8\]
rlabel metal1 s 19044 16014 19044 16014 4 po_0.regf_0.rf\[11\]\[9\]
rlabel metal2 s 10902 38080 10902 38080 4 po_0.regf_0.rf\[12\]\[0\]
rlabel metal2 s 10718 21318 10718 21318 4 po_0.regf_0.rf\[12\]\[10\]
rlabel metal1 s 4462 17714 4462 17714 4 po_0.regf_0.rf\[12\]\[11\]
rlabel metal1 s 6302 12750 6302 12750 4 po_0.regf_0.rf\[12\]\[12\]
rlabel metal1 s 8004 9554 8004 9554 4 po_0.regf_0.rf\[12\]\[13\]
rlabel metal1 s 11546 10098 11546 10098 4 po_0.regf_0.rf\[12\]\[14\]
rlabel metal1 s 11822 12818 11822 12818 4 po_0.regf_0.rf\[12\]\[15\]
rlabel metal1 s 4462 32334 4462 32334 4 po_0.regf_0.rf\[12\]\[1\]
rlabel metal1 s 10258 35020 10258 35020 4 po_0.regf_0.rf\[12\]\[2\]
rlabel metal1 s 9798 32402 9798 32402 4 po_0.regf_0.rf\[12\]\[3\]
rlabel metal1 s 5428 37230 5428 37230 4 po_0.regf_0.rf\[12\]\[4\]
rlabel metal1 s 4370 25806 4370 25806 4 po_0.regf_0.rf\[12\]\[5\]
rlabel metal1 s 6624 19822 6624 19822 4 po_0.regf_0.rf\[12\]\[6\]
rlabel metal1 s 4922 23154 4922 23154 4 po_0.regf_0.rf\[12\]\[7\]
rlabel metal2 s 10718 18224 10718 18224 4 po_0.regf_0.rf\[12\]\[8\]
rlabel metal2 s 10166 15742 10166 15742 4 po_0.regf_0.rf\[12\]\[9\]
rlabel metal1 s 8556 37842 8556 37842 4 po_0.regf_0.rf\[13\]\[0\]
rlabel metal1 s 9338 22610 9338 22610 4 po_0.regf_0.rf\[13\]\[10\]
rlabel metal1 s 4186 17068 4186 17068 4 po_0.regf_0.rf\[13\]\[11\]
rlabel metal2 s 6762 11526 6762 11526 4 po_0.regf_0.rf\[13\]\[12\]
rlabel metal1 s 7820 9486 7820 9486 4 po_0.regf_0.rf\[13\]\[13\]
rlabel metal2 s 11270 10336 11270 10336 4 po_0.regf_0.rf\[13\]\[14\]
rlabel metal1 s 10764 12954 10764 12954 4 po_0.regf_0.rf\[13\]\[15\]
rlabel metal1 s 5106 33898 5106 33898 4 po_0.regf_0.rf\[13\]\[1\]
rlabel metal1 s 9706 35054 9706 35054 4 po_0.regf_0.rf\[13\]\[2\]
rlabel metal1 s 9338 32300 9338 32300 4 po_0.regf_0.rf\[13\]\[3\]
rlabel metal2 s 4462 36992 4462 36992 4 po_0.regf_0.rf\[13\]\[4\]
rlabel metal1 s 4094 27438 4094 27438 4 po_0.regf_0.rf\[13\]\[5\]
rlabel metal2 s 4554 19652 4554 19652 4 po_0.regf_0.rf\[13\]\[6\]
rlabel metal2 s 4554 22865 4554 22865 4 po_0.regf_0.rf\[13\]\[7\]
rlabel metal1 s 9844 17646 9844 17646 4 po_0.regf_0.rf\[13\]\[8\]
rlabel metal2 s 8970 15300 8970 15300 4 po_0.regf_0.rf\[13\]\[9\]
rlabel metal2 s 7038 37706 7038 37706 4 po_0.regf_0.rf\[14\]\[0\]
rlabel metal2 s 10546 22066 10546 22066 4 po_0.regf_0.rf\[14\]\[10\]
rlabel metal2 s 5267 17102 5267 17102 4 po_0.regf_0.rf\[14\]\[11\]
rlabel metal1 s 5244 11866 5244 11866 4 po_0.regf_0.rf\[14\]\[12\]
rlabel metal2 s 8706 10642 8706 10642 4 po_0.regf_0.rf\[14\]\[13\]
rlabel metal1 s 10902 10778 10902 10778 4 po_0.regf_0.rf\[14\]\[14\]
rlabel metal1 s 10672 11866 10672 11866 4 po_0.regf_0.rf\[14\]\[15\]
rlabel metal1 s 3082 33082 3082 33082 4 po_0.regf_0.rf\[14\]\[1\]
rlabel metal2 s 7958 35428 7958 35428 4 po_0.regf_0.rf\[14\]\[2\]
rlabel metal2 s 7774 32640 7774 32640 4 po_0.regf_0.rf\[14\]\[3\]
rlabel metal2 s 4186 35904 4186 35904 4 po_0.regf_0.rf\[14\]\[4\]
rlabel metal1 s 3036 27642 3036 27642 4 po_0.regf_0.rf\[14\]\[5\]
rlabel metal2 s 5578 19890 5578 19890 4 po_0.regf_0.rf\[14\]\[6\]
rlabel metal1 s 3082 22406 3082 22406 4 po_0.regf_0.rf\[14\]\[7\]
rlabel metal1 s 8372 18598 8372 18598 4 po_0.regf_0.rf\[14\]\[8\]
rlabel metal2 s 7774 14552 7774 14552 4 po_0.regf_0.rf\[14\]\[9\]
rlabel metal2 s 7774 37298 7774 37298 4 po_0.regf_0.rf\[15\]\[0\]
rlabel metal1 s 8740 21658 8740 21658 4 po_0.regf_0.rf\[15\]\[10\]
rlabel metal1 s 4922 17102 4922 17102 4 po_0.regf_0.rf\[15\]\[11\]
rlabel metal1 s 5566 12750 5566 12750 4 po_0.regf_0.rf\[15\]\[12\]
rlabel metal1 s 8464 9962 8464 9962 4 po_0.regf_0.rf\[15\]\[13\]
rlabel metal1 s 11132 9894 11132 9894 4 po_0.regf_0.rf\[15\]\[14\]
rlabel metal2 s 10350 12410 10350 12410 4 po_0.regf_0.rf\[15\]\[15\]
rlabel metal2 s 5014 32470 5014 32470 4 po_0.regf_0.rf\[15\]\[1\]
rlabel metal2 s 10442 34646 10442 34646 4 po_0.regf_0.rf\[15\]\[2\]
rlabel metal2 s 8234 32368 8234 32368 4 po_0.regf_0.rf\[15\]\[3\]
rlabel metal2 s 5198 35360 5198 35360 4 po_0.regf_0.rf\[15\]\[4\]
rlabel metal3 s 4922 25891 4922 25891 4 po_0.regf_0.rf\[15\]\[5\]
rlabel metal1 s 3036 20570 3036 20570 4 po_0.regf_0.rf\[15\]\[6\]
rlabel metal1 s 3726 22746 3726 22746 4 po_0.regf_0.rf\[15\]\[7\]
rlabel metal2 s 11270 18224 11270 18224 4 po_0.regf_0.rf\[15\]\[8\]
rlabel metal1 s 7176 15606 7176 15606 4 po_0.regf_0.rf\[15\]\[9\]
rlabel metal1 s 24426 40052 24426 40052 4 po_0.regf_0.rf\[1\]\[0\]
rlabel metal1 s 25346 21964 25346 21964 4 po_0.regf_0.rf\[1\]\[10\]
rlabel metal2 s 27002 14042 27002 14042 4 po_0.regf_0.rf\[1\]\[11\]
rlabel metal1 s 29302 10098 29302 10098 4 po_0.regf_0.rf\[1\]\[12\]
rlabel metal1 s 30176 7446 30176 7446 4 po_0.regf_0.rf\[1\]\[13\]
rlabel metal2 s 15134 4216 15134 4216 4 po_0.regf_0.rf\[1\]\[14\]
rlabel metal2 s 24426 9282 24426 9282 4 po_0.regf_0.rf\[1\]\[15\]
rlabel metal1 s 19274 34646 19274 34646 4 po_0.regf_0.rf\[1\]\[1\]
rlabel metal2 s 17710 40256 17710 40256 4 po_0.regf_0.rf\[1\]\[2\]
rlabel metal1 s 26818 32334 26818 32334 4 po_0.regf_0.rf\[1\]\[3\]
rlabel metal2 s 28290 39882 28290 39882 4 po_0.regf_0.rf\[1\]\[4\]
rlabel metal2 s 29578 29308 29578 29308 4 po_0.regf_0.rf\[1\]\[5\]
rlabel metal2 s 32154 17000 32154 17000 4 po_0.regf_0.rf\[1\]\[6\]
rlabel metal1 s 30774 21862 30774 21862 4 po_0.regf_0.rf\[1\]\[7\]
rlabel metal1 s 27232 19142 27232 19142 4 po_0.regf_0.rf\[1\]\[8\]
rlabel metal1 s 29992 13294 29992 13294 4 po_0.regf_0.rf\[1\]\[9\]
rlabel metal2 s 23598 39882 23598 39882 4 po_0.regf_0.rf\[2\]\[0\]
rlabel metal2 s 25818 21522 25818 21522 4 po_0.regf_0.rf\[2\]\[10\]
rlabel metal2 s 26542 13498 26542 13498 4 po_0.regf_0.rf\[2\]\[11\]
rlabel metal2 s 28382 9146 28382 9146 4 po_0.regf_0.rf\[2\]\[12\]
rlabel metal2 s 30602 7922 30602 7922 4 po_0.regf_0.rf\[2\]\[13\]
rlabel metal2 s 14490 5304 14490 5304 4 po_0.regf_0.rf\[2\]\[14\]
rlabel metal2 s 23966 7616 23966 7616 4 po_0.regf_0.rf\[2\]\[15\]
rlabel metal2 s 18538 32198 18538 32198 4 po_0.regf_0.rf\[2\]\[1\]
rlabel metal1 s 16790 38930 16790 38930 4 po_0.regf_0.rf\[2\]\[2\]
rlabel metal2 s 25438 32640 25438 32640 4 po_0.regf_0.rf\[2\]\[3\]
rlabel metal2 s 28394 37298 28394 37298 4 po_0.regf_0.rf\[2\]\[4\]
rlabel metal2 s 26634 27200 26634 27200 4 po_0.regf_0.rf\[2\]\[5\]
rlabel metal1 s 29486 17306 29486 17306 4 po_0.regf_0.rf\[2\]\[6\]
rlabel metal2 s 26726 24378 26726 24378 4 po_0.regf_0.rf\[2\]\[7\]
rlabel metal1 s 26508 19890 26508 19890 4 po_0.regf_0.rf\[2\]\[8\]
rlabel metal2 s 30786 13906 30786 13906 4 po_0.regf_0.rf\[2\]\[9\]
rlabel metal2 s 25806 38726 25806 38726 4 po_0.regf_0.rf\[3\]\[0\]
rlabel metal1 s 26174 22066 26174 22066 4 po_0.regf_0.rf\[3\]\[10\]
rlabel metal2 s 26910 14144 26910 14144 4 po_0.regf_0.rf\[3\]\[11\]
rlabel metal2 s 29210 9758 29210 9758 4 po_0.regf_0.rf\[3\]\[12\]
rlabel metal1 s 29118 7310 29118 7310 4 po_0.regf_0.rf\[3\]\[13\]
rlabel metal2 s 14030 6052 14030 6052 4 po_0.regf_0.rf\[3\]\[14\]
rlabel metal1 s 25254 9010 25254 9010 4 po_0.regf_0.rf\[3\]\[15\]
rlabel metal2 s 18078 32674 18078 32674 4 po_0.regf_0.rf\[3\]\[1\]
rlabel metal2 s 16790 38794 16790 38794 4 po_0.regf_0.rf\[3\]\[2\]
rlabel metal1 s 26634 32878 26634 32878 4 po_0.regf_0.rf\[3\]\[3\]
rlabel metal1 s 28382 37774 28382 37774 4 po_0.regf_0.rf\[3\]\[4\]
rlabel metal2 s 28474 27846 28474 27846 4 po_0.regf_0.rf\[3\]\[5\]
rlabel metal1 s 30130 18190 30130 18190 4 po_0.regf_0.rf\[3\]\[6\]
rlabel metal1 s 28566 23630 28566 23630 4 po_0.regf_0.rf\[3\]\[7\]
rlabel metal2 s 26496 18802 26496 18802 4 po_0.regf_0.rf\[3\]\[8\]
rlabel metal1 s 30314 15130 30314 15130 4 po_0.regf_0.rf\[3\]\[9\]
rlabel metal2 s 34086 36312 34086 36312 4 po_0.regf_0.rf\[4\]\[0\]
rlabel metal1 s 36846 21998 36846 21998 4 po_0.regf_0.rf\[4\]\[10\]
rlabel metal1 s 36156 13294 36156 13294 4 po_0.regf_0.rf\[4\]\[11\]
rlabel metal2 s 35466 4794 35466 4794 4 po_0.regf_0.rf\[4\]\[12\]
rlabel metal1 s 32936 7922 32936 7922 4 po_0.regf_0.rf\[4\]\[13\]
rlabel metal1 s 21965 5746 21965 5746 4 po_0.regf_0.rf\[4\]\[14\]
rlabel metal1 s 28336 5202 28336 5202 4 po_0.regf_0.rf\[4\]\[15\]
rlabel metal1 s 15456 31926 15456 31926 4 po_0.regf_0.rf\[4\]\[1\]
rlabel metal2 s 12558 37536 12558 37536 4 po_0.regf_0.rf\[4\]\[2\]
rlabel metal1 s 35328 31178 35328 31178 4 po_0.regf_0.rf\[4\]\[3\]
rlabel metal2 s 32522 33728 32522 33728 4 po_0.regf_0.rf\[4\]\[4\]
rlabel metal1 s 36156 27098 36156 27098 4 po_0.regf_0.rf\[4\]\[5\]
rlabel metal2 s 33718 18768 33718 18768 4 po_0.regf_0.rf\[4\]\[6\]
rlabel metal1 s 36800 23086 36800 23086 4 po_0.regf_0.rf\[4\]\[7\]
rlabel metal1 s 35052 18938 35052 18938 4 po_0.regf_0.rf\[4\]\[8\]
rlabel metal1 s 33580 13838 33580 13838 4 po_0.regf_0.rf\[4\]\[9\]
rlabel metal2 s 32522 38080 32522 38080 4 po_0.regf_0.rf\[5\]\[0\]
rlabel metal1 s 35144 21998 35144 21998 4 po_0.regf_0.rf\[5\]\[10\]
rlabel metal1 s 25300 13158 25300 13158 4 po_0.regf_0.rf\[5\]\[11\]
rlabel metal2 s 32154 4896 32154 4896 4 po_0.regf_0.rf\[5\]\[12\]
rlabel metal1 s 33994 7310 33994 7310 4 po_0.regf_0.rf\[5\]\[13\]
rlabel metal1 s 21666 5610 21666 5610 4 po_0.regf_0.rf\[5\]\[14\]
rlabel metal1 s 25300 4658 25300 4658 4 po_0.regf_0.rf\[5\]\[15\]
rlabel metal1 s 14720 34714 14720 34714 4 po_0.regf_0.rf\[5\]\[1\]
rlabel metal2 s 13570 40256 13570 40256 4 po_0.regf_0.rf\[5\]\[2\]
rlabel metal1 s 32614 32538 32614 32538 4 po_0.regf_0.rf\[5\]\[3\]
rlabel metal1 s 30682 37842 30682 37842 4 po_0.regf_0.rf\[5\]\[4\]
rlabel metal1 s 34776 29002 34776 29002 4 po_0.regf_0.rf\[5\]\[5\]
rlabel metal1 s 35236 17578 35236 17578 4 po_0.regf_0.rf\[5\]\[6\]
rlabel metal1 s 35926 23698 35926 23698 4 po_0.regf_0.rf\[5\]\[7\]
rlabel metal1 s 23092 19278 23092 19278 4 po_0.regf_0.rf\[5\]\[8\]
rlabel metal1 s 35144 13226 35144 13226 4 po_0.regf_0.rf\[5\]\[9\]
rlabel metal1 s 33005 36210 33005 36210 4 po_0.regf_0.rf\[6\]\[0\]
rlabel metal2 s 33350 21284 33350 21284 4 po_0.regf_0.rf\[6\]\[10\]
rlabel metal2 s 23460 12070 23460 12070 4 po_0.regf_0.rf\[6\]\[11\]
rlabel metal1 s 32522 3638 32522 3638 4 po_0.regf_0.rf\[6\]\[12\]
rlabel metal2 s 33534 6970 33534 6970 4 po_0.regf_0.rf\[6\]\[13\]
rlabel metal2 s 22690 5746 22690 5746 4 po_0.regf_0.rf\[6\]\[14\]
rlabel metal2 s 24886 3264 24886 3264 4 po_0.regf_0.rf\[6\]\[15\]
rlabel metal1 s 14214 32538 14214 32538 4 po_0.regf_0.rf\[6\]\[1\]
rlabel metal2 s 12190 40902 12190 40902 4 po_0.regf_0.rf\[6\]\[2\]
rlabel metal2 s 31970 31110 31970 31110 4 po_0.regf_0.rf\[6\]\[3\]
rlabel metal1 s 30636 35802 30636 35802 4 po_0.regf_0.rf\[6\]\[4\]
rlabel metal1 s 33592 27506 33592 27506 4 po_0.regf_0.rf\[6\]\[5\]
rlabel metal2 s 34558 18258 34558 18258 4 po_0.regf_0.rf\[6\]\[6\]
rlabel metal1 s 34328 23630 34328 23630 4 po_0.regf_0.rf\[6\]\[7\]
rlabel metal2 s 24162 19278 24162 19278 4 po_0.regf_0.rf\[6\]\[8\]
rlabel metal2 s 34466 13838 34466 13838 4 po_0.regf_0.rf\[6\]\[9\]
rlabel metal1 s 32568 39270 32568 39270 4 po_0.regf_0.rf\[7\]\[0\]
rlabel metal2 s 34454 20196 34454 20196 4 po_0.regf_0.rf\[7\]\[10\]
rlabel metal1 s 23644 12750 23644 12750 4 po_0.regf_0.rf\[7\]\[11\]
rlabel metal1 s 33442 3162 33442 3162 4 po_0.regf_0.rf\[7\]\[12\]
rlabel metal1 s 33534 7922 33534 7922 4 po_0.regf_0.rf\[7\]\[13\]
rlabel metal2 s 22586 5950 22586 5950 4 po_0.regf_0.rf\[7\]\[14\]
rlabel metal2 s 25898 4896 25898 4896 4 po_0.regf_0.rf\[7\]\[15\]
rlabel metal1 s 13156 33082 13156 33082 4 po_0.regf_0.rf\[7\]\[1\]
rlabel metal2 s 12466 39967 12466 39967 4 po_0.regf_0.rf\[7\]\[2\]
rlabel metal1 s 32798 30158 32798 30158 4 po_0.regf_0.rf\[7\]\[3\]
rlabel metal2 s 30958 38726 30958 38726 4 po_0.regf_0.rf\[7\]\[4\]
rlabel metal1 s 33534 28152 33534 28152 4 po_0.regf_0.rf\[7\]\[5\]
rlabel metal1 s 34362 18190 34362 18190 4 po_0.regf_0.rf\[7\]\[6\]
rlabel metal2 s 34362 24956 34362 24956 4 po_0.regf_0.rf\[7\]\[7\]
rlabel metal2 s 24012 18258 24012 18258 4 po_0.regf_0.rf\[7\]\[8\]
rlabel metal2 s 34178 13328 34178 13328 4 po_0.regf_0.rf\[7\]\[9\]
rlabel metal1 s 23368 38318 23368 38318 4 po_0.regf_0.rf\[8\]\[0\]
rlabel metal1 s 19504 22950 19504 22950 4 po_0.regf_0.rf\[8\]\[10\]
rlabel metal2 s 19366 15266 19366 15266 4 po_0.regf_0.rf\[8\]\[11\]
rlabel metal1 s 18722 13158 18722 13158 4 po_0.regf_0.rf\[8\]\[12\]
rlabel metal2 s 19550 7174 19550 7174 4 po_0.regf_0.rf\[8\]\[13\]
rlabel metal2 s 17710 6528 17710 6528 4 po_0.regf_0.rf\[8\]\[14\]
rlabel metal2 s 18078 10846 18078 10846 4 po_0.regf_0.rf\[8\]\[15\]
rlabel metal1 s 17618 29206 17618 29206 4 po_0.regf_0.rf\[8\]\[1\]
rlabel metal1 s 17526 36754 17526 36754 4 po_0.regf_0.rf\[8\]\[2\]
rlabel metal1 s 24012 30906 24012 30906 4 po_0.regf_0.rf\[8\]\[3\]
rlabel metal1 s 24702 35054 24702 35054 4 po_0.regf_0.rf\[8\]\[4\]
rlabel metal1 s 23966 27370 23966 27370 4 po_0.regf_0.rf\[8\]\[5\]
rlabel metal2 s 17250 21216 17250 21216 4 po_0.regf_0.rf\[8\]\[6\]
rlabel metal1 s 19596 24242 19596 24242 4 po_0.regf_0.rf\[8\]\[7\]
rlabel metal1 s 17158 17646 17158 17646 4 po_0.regf_0.rf\[8\]\[8\]
rlabel metal1 s 18308 16762 18308 16762 4 po_0.regf_0.rf\[8\]\[9\]
rlabel metal2 s 22034 40698 22034 40698 4 po_0.regf_0.rf\[9\]\[0\]
rlabel metal1 s 19734 21930 19734 21930 4 po_0.regf_0.rf\[9\]\[10\]
rlabel metal2 s 19734 14756 19734 14756 4 po_0.regf_0.rf\[9\]\[11\]
rlabel metal1 s 17066 12750 17066 12750 4 po_0.regf_0.rf\[9\]\[12\]
rlabel metal1 s 19182 7922 19182 7922 4 po_0.regf_0.rf\[9\]\[13\]
rlabel metal1 s 17664 4182 17664 4182 4 po_0.regf_0.rf\[9\]\[14\]
rlabel metal2 s 17894 10064 17894 10064 4 po_0.regf_0.rf\[9\]\[15\]
rlabel metal2 s 16698 34170 16698 34170 4 po_0.regf_0.rf\[9\]\[1\]
rlabel metal1 s 15548 36142 15548 36142 4 po_0.regf_0.rf\[9\]\[2\]
rlabel metal1 s 23552 30226 23552 30226 4 po_0.regf_0.rf\[9\]\[3\]
rlabel metal1 s 27232 40154 27232 40154 4 po_0.regf_0.rf\[9\]\[4\]
rlabel metal1 s 23092 27982 23092 27982 4 po_0.regf_0.rf\[9\]\[5\]
rlabel metal1 s 17112 20910 17112 20910 4 po_0.regf_0.rf\[9\]\[6\]
rlabel metal2 s 19550 24004 19550 24004 4 po_0.regf_0.rf\[9\]\[7\]
rlabel metal1 s 19366 18870 19366 18870 4 po_0.regf_0.rf\[9\]\[8\]
rlabel metal2 s 18354 15997 18354 15997 4 po_0.regf_0.rf\[9\]\[9\]
rlabel metal2 s 7958 27064 7958 27064 4 po_0.regf_0.rp_addr\[0\]
rlabel metal1 s 7636 25330 7636 25330 4 po_0.regf_0.rp_addr\[1\]
rlabel metal2 s 6854 30464 6854 30464 4 po_0.regf_0.rp_addr\[2\]
rlabel metal1 s 6854 29036 6854 29036 4 po_0.regf_0.rp_addr\[3\]
rlabel metal2 s 33608 40018 33608 40018 4 po_0.regf_0.rp_rd
rlabel metal1 s 19090 43282 19090 43282 4 po_0.regf_0.rq_addr\[0\]
rlabel metal2 s 18078 42704 18078 42704 4 po_0.regf_0.rq_addr\[1\]
rlabel metal2 s 16882 45152 16882 45152 4 po_0.regf_0.rq_addr\[2\]
rlabel metal1 s 17802 46682 17802 46682 4 po_0.regf_0.rq_addr\[3\]
rlabel metal2 s 36110 34374 36110 34374 4 po_0.regf_0.rq_rd
rlabel metal1 s 11546 28594 11546 28594 4 po_0.regf_0.w_addr\[0\]
rlabel metal2 s 12650 29036 12650 29036 4 po_0.regf_0.w_addr\[1\]
rlabel metal1 s 11086 25874 11086 25874 4 po_0.regf_0.w_addr\[2\]
rlabel metal2 s 14122 25534 14122 25534 4 po_0.regf_0.w_addr\[3\]
rlabel metal1 s 15188 28458 15188 28458 4 po_0.regf_0.w_wr
rlabel metal2 s 46598 23137 46598 23137 4 reset
rlabel metal2 s 32982 42500 32982 42500 4 uc_0._00_
rlabel metal1 s 33304 44370 33304 44370 4 uc_0._01_
rlabel metal1 s 34178 44370 34178 44370 4 uc_0._02_
rlabel metal1 s 37398 43962 37398 43962 4 uc_0._03_
rlabel metal1 s 2553 30226 2553 30226 4 uc_0._20_\[10\]
rlabel metal1 s 7406 28526 7406 28526 4 uc_0._20_\[11\]
rlabel metal1 s 8050 27370 8050 27370 4 uc_0._20_\[8\]
rlabel metal2 s 13110 27302 13110 27302 4 uc_0._20_\[9\]
rlabel metal2 s 36846 38046 36846 38046 4 uc_0.bc_0._54_\[0\]
rlabel metal1 s 36800 39542 36800 39542 4 uc_0.bc_0._54_\[1\]
rlabel metal2 s 37498 37978 37498 37978 4 uc_0.bc_0._54_\[2\]
rlabel metal2 s 37858 39610 37858 39610 4 uc_0.bc_0._54_\[3\]
rlabel metal2 s 39422 39440 39422 39440 4 uc_0.bc_0._55_\[0\]
rlabel metal2 s 38870 40358 38870 40358 4 uc_0.bc_0._55_\[1\]
rlabel metal1 s 39698 39950 39698 39950 4 uc_0.bc_0._55_\[2\]
rlabel metal1 s 39790 39610 39790 39610 4 uc_0.bc_0._55_\[3\]
flabel metal3 s 47480 8168 48280 8288 0 FreeSans 600 0 0 0 D_R_data[0]
port 1 nsew
flabel metal2 s 43166 49624 43222 50424 0 FreeSans 280 90 0 0 D_R_data[10]
port 2 nsew
flabel metal3 s 0 24488 800 24608 0 FreeSans 600 0 0 0 D_R_data[11]
port 3 nsew
flabel metal3 s 0 12248 800 12368 0 FreeSans 600 0 0 0 D_R_data[12]
port 4 nsew
flabel metal2 s 13542 0 13598 800 0 FreeSans 280 90 0 0 D_R_data[13]
port 5 nsew
flabel metal2 s 23202 0 23258 800 0 FreeSans 280 90 0 0 D_R_data[14]
port 6 nsew
flabel metal2 s 39302 0 39358 800 0 FreeSans 280 90 0 0 D_R_data[15]
port 7 nsew
flabel metal2 s 41878 0 41934 800 0 FreeSans 280 90 0 0 D_R_data[1]
port 8 nsew
flabel metal3 s 47480 47608 48280 47728 0 FreeSans 600 0 0 0 D_R_data[2]
port 9 nsew
flabel metal2 s 5814 49624 5870 50424 0 FreeSans 280 90 0 0 D_R_data[3]
port 10 nsew
flabel metal3 s 0 31968 800 32088 0 FreeSans 600 0 0 0 D_R_data[4]
port 11 nsew
flabel metal2 s 24490 49624 24546 50424 0 FreeSans 280 90 0 0 D_R_data[5]
port 12 nsew
flabel metal3 s 0 29248 800 29368 0 FreeSans 600 0 0 0 D_R_data[6]
port 13 nsew
flabel metal3 s 47480 688 48280 808 0 FreeSans 600 0 0 0 D_R_data[7]
port 14 nsew
flabel metal2 s 46386 0 46442 800 0 FreeSans 280 90 0 0 D_R_data[8]
port 15 nsew
flabel metal2 s 27066 49624 27122 50424 0 FreeSans 280 90 0 0 D_R_data[9]
port 16 nsew
flabel metal2 s 36082 49624 36138 50424 0 FreeSans 280 90 0 0 D_W_data[0]
port 17 nsew
flabel metal3 s 47480 5448 48280 5568 0 FreeSans 600 0 0 0 D_W_data[10]
port 18 nsew
flabel metal3 s 47480 32648 48280 32768 0 FreeSans 600 0 0 0 D_W_data[11]
port 19 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 D_W_data[12]
port 20 nsew
flabel metal3 s 47480 15648 48280 15768 0 FreeSans 600 0 0 0 D_W_data[13]
port 21 nsew
flabel metal3 s 47480 35368 48280 35488 0 FreeSans 600 0 0 0 D_W_data[14]
port 22 nsew
flabel metal3 s 0 2048 800 2168 0 FreeSans 600 0 0 0 D_W_data[15]
port 23 nsew
flabel metal3 s 47480 42848 48280 42968 0 FreeSans 600 0 0 0 D_W_data[1]
port 24 nsew
flabel metal3 s 47480 17688 48280 17808 0 FreeSans 600 0 0 0 D_W_data[2]
port 25 nsew
flabel metal3 s 47480 29928 48280 30048 0 FreeSans 600 0 0 0 D_W_data[3]
port 26 nsew
flabel metal3 s 47480 12928 48280 13048 0 FreeSans 600 0 0 0 D_W_data[4]
port 27 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 D_W_data[5]
port 28 nsew
flabel metal3 s 47480 40128 48280 40248 0 FreeSans 600 0 0 0 D_W_data[6]
port 29 nsew
flabel metal3 s 0 41488 800 41608 0 FreeSans 600 0 0 0 D_W_data[7]
port 30 nsew
flabel metal3 s 0 46928 800 47048 0 FreeSans 600 0 0 0 D_W_data[8]
port 31 nsew
flabel metal3 s 0 48968 800 49088 0 FreeSans 600 0 0 0 D_W_data[9]
port 32 nsew
flabel metal2 s 4526 0 4582 800 0 FreeSans 280 90 0 0 D_addr[0]
port 33 nsew
flabel metal2 s 28998 49624 29054 50424 0 FreeSans 280 90 0 0 D_addr[1]
port 34 nsew
flabel metal2 s 18694 0 18750 800 0 FreeSans 280 90 0 0 D_addr[2]
port 35 nsew
flabel metal2 s 30286 0 30342 800 0 FreeSans 280 90 0 0 D_addr[3]
port 36 nsew
flabel metal3 s 47480 37408 48280 37528 0 FreeSans 600 0 0 0 D_addr[4]
port 37 nsew
flabel metal2 s 15474 49624 15530 50424 0 FreeSans 280 90 0 0 D_addr[5]
port 38 nsew
flabel metal3 s 0 19728 800 19848 0 FreeSans 600 0 0 0 D_addr[6]
port 39 nsew
flabel metal2 s 11610 0 11666 800 0 FreeSans 280 90 0 0 D_addr[7]
port 40 nsew
flabel metal2 s 37370 0 37426 800 0 FreeSans 280 90 0 0 D_rd
port 41 nsew
flabel metal2 s 34150 49624 34206 50424 0 FreeSans 280 90 0 0 D_wr
port 42 nsew
flabel metal3 s 0 39448 800 39568 0 FreeSans 600 0 0 0 I_addr[0]
port 43 nsew
flabel metal2 s 27710 0 27766 800 0 FreeSans 280 90 0 0 I_addr[10]
port 44 nsew
flabel metal2 s 1306 49624 1362 50424 0 FreeSans 280 90 0 0 I_addr[11]
port 45 nsew
flabel metal2 s 44454 0 44510 800 0 FreeSans 280 90 0 0 I_addr[12]
port 46 nsew
flabel metal2 s 17406 49624 17462 50424 0 FreeSans 280 90 0 0 I_addr[13]
port 47 nsew
flabel metal3 s 47480 10208 48280 10328 0 FreeSans 600 0 0 0 I_addr[14]
port 48 nsew
flabel metal3 s 47480 20408 48280 20528 0 FreeSans 600 0 0 0 I_addr[15]
port 49 nsew
flabel metal2 s 34794 0 34850 800 0 FreeSans 280 90 0 0 I_addr[1]
port 50 nsew
flabel metal3 s 0 34008 800 34128 0 FreeSans 600 0 0 0 I_addr[2]
port 51 nsew
flabel metal2 s 12898 49624 12954 50424 0 FreeSans 280 90 0 0 I_addr[3]
port 52 nsew
flabel metal2 s 22558 49624 22614 50424 0 FreeSans 280 90 0 0 I_addr[4]
port 53 nsew
flabel metal3 s 0 4768 800 4888 0 FreeSans 600 0 0 0 I_addr[5]
port 54 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 I_addr[6]
port 55 nsew
flabel metal3 s 0 26528 800 26648 0 FreeSans 600 0 0 0 I_addr[7]
port 56 nsew
flabel metal2 s 19982 49624 20038 50424 0 FreeSans 280 90 0 0 I_addr[8]
port 57 nsew
flabel metal2 s 31574 49624 31630 50424 0 FreeSans 280 90 0 0 I_addr[9]
port 58 nsew
flabel metal2 s 45742 49624 45798 50424 0 FreeSans 280 90 0 0 I_data[0]
port 59 nsew
flabel metal3 s 0 36728 800 36848 0 FreeSans 600 0 0 0 I_data[10]
port 60 nsew
flabel metal2 s 6458 0 6514 800 0 FreeSans 280 90 0 0 I_data[11]
port 61 nsew
flabel metal2 s 1950 0 2006 800 0 FreeSans 280 90 0 0 I_data[12]
port 62 nsew
flabel metal2 s 47674 49624 47730 50424 0 FreeSans 280 90 0 0 I_data[13]
port 63 nsew
flabel metal3 s 0 17008 800 17128 0 FreeSans 600 0 0 0 I_data[14]
port 64 nsew
flabel metal2 s 20626 0 20682 800 0 FreeSans 280 90 0 0 I_data[15]
port 65 nsew
flabel metal3 s 47480 44888 48280 45008 0 FreeSans 600 0 0 0 I_data[1]
port 66 nsew
flabel metal3 s 47480 2728 48280 2848 0 FreeSans 600 0 0 0 I_data[2]
port 67 nsew
flabel metal2 s 8390 49624 8446 50424 0 FreeSans 280 90 0 0 I_data[3]
port 68 nsew
flabel metal3 s 47480 25168 48280 25288 0 FreeSans 600 0 0 0 I_data[4]
port 69 nsew
flabel metal2 s 9034 0 9090 800 0 FreeSans 280 90 0 0 I_data[5]
port 70 nsew
flabel metal2 s 16118 0 16174 800 0 FreeSans 280 90 0 0 I_data[6]
port 71 nsew
flabel metal3 s 0 21768 800 21888 0 FreeSans 600 0 0 0 I_data[7]
port 72 nsew
flabel metal3 s 47480 27888 48280 28008 0 FreeSans 600 0 0 0 I_data[8]
port 73 nsew
flabel metal2 s 25134 0 25190 800 0 FreeSans 280 90 0 0 I_data[9]
port 74 nsew
flabel metal2 s 41234 49624 41290 50424 0 FreeSans 280 90 0 0 I_rd
port 75 nsew
flabel metal5 s 1056 36642 47152 36962 0 FreeSans 3200 0 0 0 VGND
port 76 nsew
flabel metal5 s 1056 6006 47152 6326 0 FreeSans 3200 0 0 0 VGND
port 76 nsew
flabel metal4 s 35588 2128 35908 47920 0 FreeSans 2400 90 0 0 VGND
port 76 nsew
flabel metal4 s 4868 2128 5188 47920 0 FreeSans 2400 90 0 0 VGND
port 76 nsew
flabel metal5 s 1056 35982 47152 36302 0 FreeSans 3200 0 0 0 VPWR
port 77 nsew
flabel metal5 s 1056 5346 47152 5666 0 FreeSans 3200 0 0 0 VPWR
port 77 nsew
flabel metal4 s 34928 2128 35248 47920 0 FreeSans 2400 90 0 0 VPWR
port 77 nsew
flabel metal4 s 4208 2128 4528 47920 0 FreeSans 2400 90 0 0 VPWR
port 77 nsew
flabel metal2 s 38658 49624 38714 50424 0 FreeSans 280 90 0 0 clock
port 78 nsew
flabel metal2 s 3238 49624 3294 50424 0 FreeSans 280 90 0 0 led_clock
port 79 nsew
flabel metal2 s 10322 49624 10378 50424 0 FreeSans 280 90 0 0 leds[0]
port 80 nsew
flabel metal2 s 32218 0 32274 800 0 FreeSans 280 90 0 0 leds[1]
port 81 nsew
flabel metal3 s 0 14288 800 14408 0 FreeSans 600 0 0 0 leds[2]
port 82 nsew
flabel metal3 s 0 44208 800 44328 0 FreeSans 600 0 0 0 leds[3]
port 83 nsew
flabel metal3 s 47480 23128 48280 23248 0 FreeSans 600 0 0 0 reset
port 84 nsew
<< properties >>
string FIXED_BBOX 0 0 48280 50424
<< end >>
