* NGSPICE file created from vahid6i.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt vahid6i D_R_data[0] D_R_data[10] D_R_data[11] D_R_data[12] D_R_data[13] D_R_data[14]
+ D_R_data[15] D_R_data[1] D_R_data[2] D_R_data[3] D_R_data[4] D_R_data[5] D_R_data[6]
+ D_R_data[7] D_R_data[8] D_R_data[9] D_W_data[0] D_W_data[10] D_W_data[11] D_W_data[12]
+ D_W_data[13] D_W_data[14] D_W_data[15] D_W_data[1] D_W_data[2] D_W_data[3] D_W_data[4]
+ D_W_data[5] D_W_data[6] D_W_data[7] D_W_data[8] D_W_data[9] D_addr[0] D_addr[1]
+ D_addr[2] D_addr[3] D_addr[4] D_addr[5] D_addr[6] D_addr[7] D_rd D_wr I_addr[0]
+ I_addr[10] I_addr[11] I_addr[12] I_addr[13] I_addr[14] I_addr[15] I_addr[1] I_addr[2]
+ I_addr[3] I_addr[4] I_addr[5] I_addr[6] I_addr[7] I_addr[8] I_addr[9] I_data[0]
+ I_data[10] I_data[11] I_data[12] I_data[13] I_data[14] I_data[15] I_data[1] I_data[2]
+ I_data[3] I_data[4] I_data[5] I_data[6] I_data[7] I_data[8] I_data[9] I_rd VGND
+ VPWR clock led_clock leds[0] leds[1] leds[2] leds[3] reset
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3155_ net142 _0130_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3086_ net109 _0009_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__dfxtp_1
X_2106_ _0721_ _0722_ _0723_ _0726_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__o31a_1
X_2037_ _0632_ _0649_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__nand2_1
XFILLER_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2939_ net91 _1219_ _0563_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__a21o_1
XFILLER_45_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2724_ _1133_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__buf_2
X_2655_ _1096_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__clkbuf_1
X_1606_ _1390_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__clkbuf_2
X_2586_ _1051_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__buf_2
Xfanout105 net117 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlymetal6s2s_1
X_1537_ net39 net38 net41 net40 VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__nor4_1
Xfanout127 net136 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout116 net117 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout138 net139 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout149 net155 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlymetal6s2s_1
X_3207_ net114 _0182_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3138_ net140 _0113_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3069_ net169 _0048_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2440_ _0975_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
X_2371_ _0932_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2707_ _1124_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__clkbuf_1
X_2638_ po_0.regf_0.rf\[10\]\[14\] _0988_ _1070_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__mux2_1
X_2569_ po_0.regf_0.rf\[12\]\[15\] _0990_ _1031_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__mux2_1
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1940_ _0572_ _0577_ VGND VGND VPWR VPWR po_0.alu_0._10_\[1\] sky130_fd_sc_hd__xor2_1
X_1871_ _0430_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__and2b_1
X_2423_ po_0.regf_0.rf\[15\]\[2\] _0963_ _0959_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__mux2_1
X_2354_ _0923_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
X_2285_ _0885_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2070_ _0681_ _0683_ _0685_ net1 _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__a221o_2
XFILLER_78_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2972_ _1296_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__clkbuf_1
X_1923_ _0564_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
X_1854_ _0502_ _0503_ _0414_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__mux2_1
X_1785_ _0440_ _0411_ _0420_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__a21o_1
X_2406_ _0952_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_3386_ po_0.alu_0._10_\[7\] _1475_ VGND VGND VPWR VPWR po_0.alu_0._11_\[7\] sky130_fd_sc_hd__ebufn_1
X_2337_ _0913_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
X_2268_ po_0.regf_0.w_addr\[2\] VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2199_ net49 po_0._1_\[8\] po_0._1_\[9\] _0633_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__a22oi_2
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1570_ uc_0._20_\[10\] po_0.regf_0.rp_addr\[2\] _1373_ VGND VGND VPWR VPWR _1376_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_5 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ net115 _0215_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ net142 _0146_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2122_ _0741_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2053_ _0670_ _0672_ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2955_ uc_0._20_\[9\] po_0.regf_0.rp_addr\[1\] _1373_ VGND VGND VPWR VPWR _1286_
+ sky130_fd_sc_hd__mux2_1
X_1906_ _0508_ _0549_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__and2b_1
X_2886_ _1250_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__clkbuf_1
X_1837_ po_0.regf_0.rf\[4\]\[6\] po_0.regf_0.rf\[5\]\[6\] po_0.regf_0.rf\[6\]\[6\]
+ po_0.regf_0.rf\[7\]\[6\] _0427_ _0428_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__mux4_1
X_1768_ po_0.regf_0.rf\[0\]\[0\] po_0.regf_0.rf\[1\]\[0\] po_0.regf_0.rf\[2\]\[0\]
+ po_0.regf_0.rf\[3\]\[0\] _0423_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux4_1
X_1699_ _1378_ _0362_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__and2b_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ net170 uc_0.bc_0._54_\[2\] VGND VGND VPWR VPWR uc_0.bc_0._55_\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput42 net42 VGND VGND VPWR VPWR D_W_data[1] sky130_fd_sc_hd__buf_2
Xoutput75 net75 VGND VGND VPWR VPWR I_addr[8] sky130_fd_sc_hd__buf_2
Xoutput53 net53 VGND VGND VPWR VPWR D_addr[2] sky130_fd_sc_hd__buf_2
Xoutput64 net64 VGND VGND VPWR VPWR I_addr[12] sky130_fd_sc_hd__buf_2
XFILLER_48_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2740_ _1142_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__clkbuf_1
X_2671_ _0849_ po_0.regf_0.rf\[0\]\[13\] _1089_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__mux2_1
X_1622_ _1378_ _1423_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__and2b_1
X_1553_ _1362_ uc_0.bc_0._55_\[1\] uc_0.bc_0._55_\[0\] uc_0.bc_0._55_\[2\] uc_0.bc_0._55_\[3\]
+ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__a311oi_4
X_1484_ po_0.alu_0.s0 VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3223_ net132 _0198_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3154_ net142 _0129_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3085_ net109 _0008_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__dfxtp_1
X_2105_ _0593_ _0723_ _0725_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__a21oi_1
X_2036_ _0654_ _0658_ _0660_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__o211a_1
XFILLER_35_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2938_ _1315_ _0563_ _1370_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__o21ba_1
X_2869_ _1241_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__clkbuf_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2723_ uc_0._03_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__buf_4
X_2654_ _0765_ po_0.regf_0.rf\[0\]\[5\] _1090_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__mux2_1
X_2585_ _1058_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
X_1605_ po_0.regf_0.rf\[4\]\[1\] po_0.regf_0.rf\[5\]\[1\] po_0.regf_0.rf\[6\]\[1\]
+ po_0.regf_0.rf\[7\]\[1\] _1406_ _1407_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__mux4_1
X_1536_ uc_0.bc_0._55_\[1\] uc_0.bc_0._55_\[2\] uc_0.bc_0._55_\[3\] uc_0.bc_0._55_\[0\]
+ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__and4bb_1
Xfanout106 net107 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
Xfanout128 net129 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
Xfanout117 net175 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout139 net146 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlymetal6s2s_1
X_3206_ net156 _0181_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3137_ net147 _0112_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3068_ po_0.regf_0._3_\[15\] net85 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlxtp_1
X_2019_ _0637_ _0643_ _0638_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__o21ai_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2370_ po_0.regf_0.rf\[9\]\[13\] _0849_ _0916_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__mux2_1
XFILLER_68_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2706_ po_0.regf_0.rf\[8\]\[13\] _0848_ _1108_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__mux2_1
X_2637_ _1086_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__clkbuf_1
X_2568_ _1048_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2499_ _1010_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
X_1519_ _1325_ _1327_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__or2b_1
XFILLER_67_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1870_ po_0.regf_0.rf\[8\]\[10\] po_0.regf_0.rf\[9\]\[10\] po_0.regf_0.rf\[10\]\[10\]
+ po_0.regf_0.rf\[11\]\[10\] _0423_ _0425_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__mux4_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2422_ _0731_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__clkbuf_2
X_2353_ po_0.regf_0.rf\[9\]\[5\] _0765_ _0917_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__mux2_1
X_2284_ po_0.regf_0.rf\[5\]\[6\] _0777_ _0884_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__mux2_1
X_1999_ _0628_ _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__nand2_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2971_ _0915_ _1295_ _1280_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__mux2_1
X_1922_ po_0.regf_0.rq_addr\[0\] _0561_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__mux2_1
X_1853_ po_0.regf_0.rf\[12\]\[8\] po_0.regf_0.rf\[13\]\[8\] po_0.regf_0.rf\[14\]\[8\]
+ po_0.regf_0.rf\[15\]\[8\] _0000_ _0001_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__mux4_1
X_1784_ po_0.regf_0.rf\[4\]\[2\] po_0.regf_0.rf\[5\]\[2\] po_0.regf_0.rf\[6\]\[2\]
+ po_0.regf_0.rf\[7\]\[2\] _0406_ _0408_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__mux4_1
X_2405_ po_0.regf_0.rf\[1\]\[12\] _0840_ _0937_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__mux2_1
X_3385_ po_0.alu_0._10_\[6\] _1474_ VGND VGND VPWR VPWR po_0.alu_0._11_\[6\] sky130_fd_sc_hd__ebufn_1
XFILLER_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2336_ po_0.regf_0.rf\[6\]\[14\] _0860_ _0896_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__mux2_1
XFILLER_57_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2267_ po_0.regf_0.w_addr\[1\] po_0.regf_0.w_addr\[0\] VGND VGND VPWR VPWR _0874_
+ sky130_fd_sc_hd__and2b_1
XFILLER_57_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2198_ _0811_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_6 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ net140 _0145_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2121_ po_0.muxf_0.rf_w_data\[3\] _0683_ _0685_ net10 _0740_ VGND VGND VPWR VPWR
+ _0741_ sky130_fd_sc_hd__a221o_2
X_2052_ _0673_ _0674_ _0675_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__or3b_1
XFILLER_47_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2954_ _1285_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__clkbuf_1
X_1905_ po_0.regf_0.rf\[8\]\[14\] po_0.regf_0.rf\[9\]\[14\] po_0.regf_0.rf\[10\]\[14\]
+ po_0.regf_0.rf\[11\]\[14\] _0509_ _0510_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__mux4_1
X_2885_ po_0.regf_0.rf\[3\]\[8\] _0801_ _1247_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__mux2_1
X_1836_ po_0.regf_0.rf\[0\]\[6\] po_0.regf_0.rf\[1\]\[6\] po_0.regf_0.rf\[2\]\[6\]
+ po_0.regf_0.rf\[3\]\[6\] _0478_ _0479_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux4_1
X_1767_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__buf_2
X_1698_ po_0.regf_0.rf\[8\]\[10\] po_0.regf_0.rf\[9\]\[10\] po_0.regf_0.rf\[10\]\[10\]
+ po_0.regf_0.rf\[11\]\[10\] _1412_ _1413_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__mux4_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ net173 uc_0.bc_0._54_\[1\] VGND VGND VPWR VPWR uc_0.bc_0._55_\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _0896_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__clkbuf_4
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3299_ net125 _0270_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput43 net43 VGND VGND VPWR VPWR D_W_data[2] sky130_fd_sc_hd__clkbuf_4
Xoutput76 net76 VGND VGND VPWR VPWR I_addr[9] sky130_fd_sc_hd__clkbuf_4
Xoutput65 net65 VGND VGND VPWR VPWR I_addr[13] sky130_fd_sc_hd__buf_2
Xoutput54 net54 VGND VGND VPWR VPWR D_addr[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2670_ _1104_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__clkbuf_1
X_1621_ po_0.regf_0.rf\[0\]\[2\] po_0.regf_0.rf\[1\]\[2\] po_0.regf_0.rf\[2\]\[2\]
+ po_0.regf_0.rf\[3\]\[2\] _1380_ _1382_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__mux4_1
X_1552_ net95 net94 net80 VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__or3b_1
X_3222_ net157 _0197_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3153_ net148 _0128_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2104_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__buf_2
X_3084_ net118 _0063_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2035_ po_0._1_\[12\] _0655_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__or2b_1
XFILLER_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2937_ _1277_ _1319_ _1370_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__a21o_1
X_2868_ po_0.regf_0.rf\[3\]\[0\] _0693_ _1240_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__mux2_1
X_2799_ _1191_ _1192_ _1193_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__o21ai_1
X_1819_ _0407_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__buf_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2722_ _1132_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2653_ _1095_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__clkbuf_1
X_1604_ _1381_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__clkbuf_4
X_2584_ po_0.regf_0.rf\[11\]\[5\] _0969_ _1052_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__mux2_1
X_1535_ net47 VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__buf_2
Xfanout118 net120 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout107 net111 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout129 net131 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlymetal6s2s_1
X_3205_ net158 _0180_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3136_ net97 _0111_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3067_ po_0.regf_0._3_\[14\] net86 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlxtp_1
X_2018_ _0644_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__nor2_2
XFILLER_23_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2705_ _1123_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__clkbuf_1
X_2636_ po_0.regf_0.rf\[10\]\[13\] _0986_ _1070_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__mux2_1
X_2567_ po_0.regf_0.rf\[12\]\[14\] _0988_ _1031_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__mux2_1
X_2498_ po_0.regf_0.rf\[14\]\[15\] _0990_ _0992_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__mux2_1
X_1518_ _1335_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3119_ net99 _0094_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2421_ _0962_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
X_2352_ _0922_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_2283_ _0876_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__buf_2
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1998_ net83 po_0._1_\[8\] VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__or2_1
X_2619_ po_0.regf_0.rf\[10\]\[5\] _0969_ _1071_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__mux2_1
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2970_ uc_0._20_\[11\] po_0.muxf_0.rf_w_data\[3\] _0562_ VGND VGND VPWR VPWR _1295_
+ sky130_fd_sc_hd__mux2_1
X_1921_ _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__buf_2
X_1852_ po_0.regf_0.rf\[8\]\[8\] po_0.regf_0.rf\[9\]\[8\] po_0.regf_0.rf\[10\]\[8\]
+ po_0.regf_0.rf\[11\]\[8\] _0000_ _0001_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__mux4_1
X_1783_ _0434_ _0436_ _0421_ _0439_ VGND VGND VPWR VPWR po_0.regf_0._3_\[1\] sky130_fd_sc_hd__o22a_1
X_2404_ _0951_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
X_3384_ po_0.alu_0._10_\[5\] _1473_ VGND VGND VPWR VPWR po_0.alu_0._11_\[5\] sky130_fd_sc_hd__ebufn_1
X_2335_ _0912_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
X_2266_ _0872_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__clkbuf_2
X_2197_ po_0.regf_0.rf\[7\]\[9\] _0810_ _0778_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__mux2_1
XFILLER_25_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_7 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2120_ _0589_ _0686_ _1314_ _0687_ _0739_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__o311a_1
X_2051_ po_0._1_\[14\] net40 VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__or2b_1
XFILLER_54_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2953_ uc_0._20_\[8\] po_0.regf_0.rp_addr\[0\] _1373_ VGND VGND VPWR VPWR _1285_
+ sky130_fd_sc_hd__mux2_1
X_1904_ _0547_ _0457_ _0003_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__a21bo_1
XFILLER_30_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2884_ _1249_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__clkbuf_1
X_1835_ _0415_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__and2b_1
X_1766_ _0001_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__buf_2
X_1697_ _0360_ _1409_ _1392_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__a21o_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ net170 uc_0.bc_0._54_\[0\] VGND VGND VPWR VPWR uc_0.bc_0._55_\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _0903_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3298_ net125 _0269_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_2249_ _0855_ _0856_ _0857_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__o21ai_1
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput66 net66 VGND VGND VPWR VPWR I_addr[14] sky130_fd_sc_hd__buf_2
Xoutput44 net44 VGND VGND VPWR VPWR D_W_data[3] sky130_fd_sc_hd__buf_2
Xoutput55 net55 VGND VGND VPWR VPWR D_addr[4] sky130_fd_sc_hd__buf_2
Xoutput77 net77 VGND VGND VPWR VPWR I_rd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1620_ _1410_ _1415_ _1417_ _1422_ VGND VGND VPWR VPWR po_0.regf_0._5_\[1\] sky130_fd_sc_hd__o22a_1
X_1551_ _1357_ _1361_ VGND VGND VPWR VPWR uc_0.bc_0._54_\[0\] sky130_fd_sc_hd__nor2_1
X_3221_ net165 _0196_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3152_ net97 _0127_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2103_ po_0.alu_0.s1 _1313_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__or2b_1
X_3083_ net100 _0062_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_2034_ _0659_ po_0._1_\[13\] VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__xor2_2
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2936_ _1215_ _1359_ _1365_ _1366_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__or4_1
X_2867_ _1239_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__clkbuf_4
X_1818_ _0405_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__clkbuf_4
X_2798_ _1186_ _1184_ _1185_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__a21boi_1
X_1749_ _0001_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__clkbuf_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2721_ _0561_ net27 _1127_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__mux2_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2652_ _0755_ po_0.regf_0.rf\[0\]\[4\] _1090_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__mux2_1
X_1603_ _1379_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__clkbuf_4
X_2583_ _1057_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
X_1534_ net80 net94 _1345_ net95 VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__and4bb_1
Xfanout119 net120 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout108 net110 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlymetal6s2s_1
X_3204_ net158 _0179_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3135_ net96 _0110_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_3066_ po_0.regf_0._3_\[13\] net86 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlxtp_1
X_2017_ net37 po_0._1_\[11\] VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__and2_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2919_ _1268_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2704_ po_0.regf_0.rf\[8\]\[12\] _0839_ _1108_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__mux2_1
X_2635_ _1085_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__clkbuf_1
X_2566_ _1047_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
X_2497_ _1009_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
X_1517_ _1325_ _1327_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__or2b_1
XFILLER_74_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3118_ net125 _0093_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3049_ po_0.regf_0._5_\[12\] net88 VGND VGND VPWR VPWR po_0._1_\[12\] sky130_fd_sc_hd__dlxtp_1
XFILLER_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout90 net91 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
X_2420_ po_0.regf_0.rf\[15\]\[1\] _0961_ _0959_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__mux2_1
X_2351_ po_0.regf_0.rf\[9\]\[4\] _0755_ _0917_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__mux2_1
X_2282_ _0883_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1997_ net83 po_0._1_\[8\] VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__nand2_1
X_2618_ _1076_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
X_2549_ _1038_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1920_ _1371_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__clkbuf_4
X_1851_ _0499_ _0500_ _0414_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__mux2_1
X_1782_ _0437_ _0438_ _0430_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__mux2_1
X_2403_ po_0.regf_0.rf\[1\]\[11\] _0828_ _0945_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__mux2_1
X_3383_ po_0.alu_0._10_\[4\] _1472_ VGND VGND VPWR VPWR po_0.alu_0._11_\[4\] sky130_fd_sc_hd__ebufn_1
X_2334_ po_0.regf_0.rf\[6\]\[13\] _0849_ _0896_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__mux2_1
XFILLER_69_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2265_ po_0.regf_0.w_wr VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2196_ _0809_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_8 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2050_ net41 po_0._1_\[15\] VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__nor2_1
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2952_ _1284_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__clkbuf_1
X_1903_ po_0.regf_0.rf\[12\]\[14\] po_0.regf_0.rf\[13\]\[14\] po_0.regf_0.rf\[14\]\[14\]
+ po_0.regf_0.rf\[15\]\[14\] _0449_ _0450_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__mux4_1
X_2883_ po_0.regf_0.rf\[3\]\[7\] _0787_ _1247_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__mux2_1
X_1834_ po_0.regf_0.rf\[8\]\[6\] po_0.regf_0.rf\[9\]\[6\] po_0.regf_0.rf\[10\]\[6\]
+ po_0.regf_0.rf\[11\]\[6\] _0416_ _0417_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux4_1
X_1765_ _0422_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__clkbuf_4
X_1696_ po_0.regf_0.rf\[12\]\[10\] po_0.regf_0.rf\[13\]\[10\] po_0.regf_0.rf\[14\]\[10\]
+ po_0.regf_0.rf\[15\]\[10\] _1419_ _1420_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__mux4_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ net171 _0337_ VGND VGND VPWR VPWR uc_0._01_ sky130_fd_sc_hd__dfxtp_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ net127 _0268_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_2317_ po_0.regf_0.rf\[6\]\[5\] _0765_ _0897_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__mux2_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _0686_ po_0.alu_0._11_\[14\] _0720_ net40 VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__a22oi_1
X_2179_ _0621_ po_0._1_\[7\] _0792_ _0793_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__o22a_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput56 net56 VGND VGND VPWR VPWR D_addr[5] sky130_fd_sc_hd__buf_2
Xoutput45 net84 VGND VGND VPWR VPWR D_W_data[4] sky130_fd_sc_hd__buf_2
Xoutput67 net67 VGND VGND VPWR VPWR I_addr[15] sky130_fd_sc_hd__buf_2
Xoutput78 net78 VGND VGND VPWR VPWR led_clock sky130_fd_sc_hd__buf_2
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1550_ _1360_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__clkbuf_2
X_3220_ net159 _0195_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3151_ net97 _0126_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2102_ _0582_ _0578_ _0707_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__o21ai_2
X_3082_ net124 _0061_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_2033_ net39 VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__buf_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2935_ _1276_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2866_ _0696_ _0697_ _0873_ _0936_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__and4_4
X_1817_ _0464_ _0466_ _0468_ _0470_ VGND VGND VPWR VPWR po_0.regf_0._3_\[4\] sky130_fd_sc_hd__o22a_1
X_2797_ net71 po_0.muxf_0.rf_w_data\[4\] VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__nor2_1
X_1748_ _0405_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__clkbuf_4
X_1679_ po_0.regf_0.rf\[4\]\[7\] po_0.regf_0.rf\[5\]\[7\] po_0.regf_0.rf\[6\]\[7\]
+ po_0.regf_0.rf\[7\]\[7\] _1400_ _1401_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__mux4_1
XFILLER_77_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3349_ net138 _0320_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2720_ _1131_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2651_ _1094_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1602_ _1384_ _1394_ _1399_ _1405_ VGND VGND VPWR VPWR po_0.regf_0._5_\[0\] sky130_fd_sc_hd__o22a_1
X_2582_ po_0.regf_0.rf\[11\]\[4\] _0967_ _1052_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__mux2_1
X_1533_ uc_0.bc_0._55_\[0\] uc_0.bc_0._55_\[1\] _1344_ VGND VGND VPWR VPWR _1345_
+ sky130_fd_sc_hd__and3_1
Xfanout109 net110 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlymetal6s2s_1
X_3203_ net150 _0178_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3134_ net96 _0109_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3065_ po_0.regf_0._3_\[12\] net85 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlxtp_1
X_2016_ net37 po_0._1_\[11\] VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__nor2_1
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2918_ po_0.regf_0.rf\[2\]\[7\] _0787_ _1266_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__mux2_1
X_2849_ _1230_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2703_ _1122_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__clkbuf_1
X_2634_ po_0.regf_0.rf\[10\]\[12\] _0984_ _1070_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__mux2_1
X_2565_ po_0.regf_0.rf\[12\]\[13\] _0986_ _1031_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__mux2_1
X_1516_ _1334_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__clkbuf_1
X_2496_ po_0.regf_0.rf\[14\]\[14\] _0988_ _0992_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__mux2_1
XFILLER_59_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3117_ net119 _0092_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3048_ po_0.regf_0._5_\[11\] net88 VGND VGND VPWR VPWR po_0._1_\[11\] sky130_fd_sc_hd__dlxtp_1
XFILLER_70_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout91 po_0.regf_0.rq_rd VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2350_ _0921_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
X_2281_ po_0.regf_0.rf\[5\]\[5\] _0765_ _0877_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__mux2_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1996_ _0626_ _0627_ VGND VGND VPWR VPWR po_0.alu_0._10_\[7\] sky130_fd_sc_hd__nor2_1
X_2617_ po_0.regf_0.rf\[10\]\[4\] _0967_ _1071_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__mux2_1
X_2548_ po_0.regf_0.rf\[12\]\[5\] _0969_ _1032_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__mux2_1
X_2479_ _0992_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__buf_2
XFILLER_75_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1850_ po_0.regf_0.rf\[4\]\[8\] po_0.regf_0.rf\[5\]\[8\] po_0.regf_0.rf\[6\]\[8\]
+ po_0.regf_0.rf\[7\]\[8\] _0422_ _0424_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__mux4_1
X_1781_ po_0.regf_0.rf\[4\]\[1\] po_0.regf_0.rf\[5\]\[1\] po_0.regf_0.rf\[6\]\[1\]
+ po_0.regf_0.rf\[7\]\[1\] _0427_ _0428_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__mux4_1
XFILLER_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2402_ _0950_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
X_3382_ po_0.alu_0._10_\[3\] _1471_ VGND VGND VPWR VPWR po_0.alu_0._11_\[3\] sky130_fd_sc_hd__ebufn_1
X_2333_ _0911_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
X_2264_ _0871_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__clkbuf_1
X_2195_ net16 _0790_ _0807_ _0808_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__a22o_2
XFILLER_77_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1979_ _0612_ VGND VGND VPWR VPWR po_0.alu_0._10_\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2951_ po_0.regf_0.rq_addr\[3\] _0570_ _0568_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__mux2_1
XFILLER_22_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1902_ _0541_ _0543_ _0461_ _0546_ VGND VGND VPWR VPWR po_0.regf_0._3_\[13\] sky130_fd_sc_hd__o22a_1
XFILLER_30_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2882_ _1248_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_1
X_1833_ _0484_ _0433_ _0474_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a21bo_1
X_1764_ _0000_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__buf_2
X_1695_ _0354_ _0356_ _1440_ _0359_ VGND VGND VPWR VPWR po_0.regf_0._5_\[9\] sky130_fd_sc_hd__o22a_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ net171 _0336_ VGND VGND VPWR VPWR uc_0._02_ sky130_fd_sc_hd__dfxtp_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ net135 _0267_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_2316_ _0902_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _0670_ _0852_ _0854_ _0725_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__a31o_1
XFILLER_38_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2178_ _0607_ _0613_ _0614_ _0769_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__nor4b_1
XFILLER_53_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput35 net35 VGND VGND VPWR VPWR D_W_data[0] sky130_fd_sc_hd__buf_2
Xoutput46 net46 VGND VGND VPWR VPWR D_W_data[5] sky130_fd_sc_hd__clkbuf_4
Xoutput57 net57 VGND VGND VPWR VPWR D_addr[6] sky130_fd_sc_hd__buf_2
Xoutput79 net79 VGND VGND VPWR VPWR leds[0] sky130_fd_sc_hd__buf_2
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput68 net92 VGND VGND VPWR VPWR I_addr[1] sky130_fd_sc_hd__buf_2
XFILLER_48_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3150_ net96 _0125_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3081_ net124 _0060_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2101_ _0579_ po_0._1_\[2\] VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__and2b_1
X_2032_ _0654_ _0658_ VGND VGND VPWR VPWR po_0.alu_0._10_\[12\] sky130_fd_sc_hd__xor2_1
XFILLER_35_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2934_ po_0.regf_0.rf\[2\]\[15\] _0869_ _1258_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__mux2_1
X_2865_ _1238_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__clkbuf_1
X_1816_ _0469_ _0447_ _0461_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a21o_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2796_ net71 po_0.muxf_0.rf_w_data\[4\] VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__and2_1
X_1747_ _0000_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__clkbuf_2
X_1678_ _1395_ _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__and2b_1
X_3348_ net145 _0319_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ net119 net181 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfxtp_1
XFILLER_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2650_ _0742_ po_0.regf_0.rf\[0\]\[3\] _1090_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__mux2_1
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1601_ _1402_ _1403_ _1404_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__a21o_1
X_2581_ _1056_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
X_1532_ uc_0.bc_0._55_\[2\] uc_0.bc_0._55_\[3\] VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__nor2_1
X_3202_ net145 _0177_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3133_ net96 _0108_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3064_ po_0.regf_0._3_\[11\] net86 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlxtp_1
XFILLER_67_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2015_ _0639_ _0643_ VGND VGND VPWR VPWR po_0.alu_0._10_\[10\] sky130_fd_sc_hd__xor2_1
XFILLER_35_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2917_ _1267_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2848_ po_0.regf_0.rf\[4\]\[7\] _0787_ _1228_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__mux2_1
X_2779_ _1173_ _1174_ _1175_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__or3b_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2702_ po_0.regf_0.rf\[8\]\[11\] _0827_ _1116_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__mux2_1
XFILLER_9_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2633_ _1084_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__clkbuf_1
X_2564_ _1046_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
X_1515_ _1326_ _1328_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__or2b_1
X_2495_ _1008_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
X_3116_ net121 _0091_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3047_ po_0.regf_0._5_\[10\] net89 VGND VGND VPWR VPWR po_0._1_\[10\] sky130_fd_sc_hd__dlxtp_1
XFILLER_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout92 net68 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_2
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3279__181 VGND VGND VPWR VPWR _3279__181/HI net181 sky130_fd_sc_hd__conb_1
XFILLER_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2280_ _0882_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1995_ _0617_ _0622_ _0623_ _0624_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__nor4_1
X_2616_ _1075_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
X_2547_ _1037_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
X_2478_ _0999_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1780_ po_0.regf_0.rf\[0\]\[1\] po_0.regf_0.rf\[1\]\[1\] po_0.regf_0.rf\[2\]\[1\]
+ po_0.regf_0.rf\[3\]\[1\] _0423_ _0425_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__mux4_1
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2401_ po_0.regf_0.rf\[1\]\[10\] _0820_ _0945_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__mux2_1
X_3381_ po_0.alu_0._10_\[2\] _1470_ VGND VGND VPWR VPWR po_0.alu_0._11_\[2\] sky130_fd_sc_hd__ebufn_1
X_2332_ po_0.regf_0.rf\[6\]\[12\] _0840_ _0896_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__mux2_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2263_ po_0.regf_0.rf\[7\]\[15\] _0870_ _0700_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__mux2_1
X_2194_ _0633_ _0686_ _1314_ _0712_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__o31a_1
XFILLER_65_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1978_ _0610_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__or2_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283__177 VGND VGND VPWR VPWR _3283__177/HI net177 sky130_fd_sc_hd__conb_1
XFILLER_62_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2950_ _1283_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__clkbuf_1
X_1901_ _0544_ _0545_ _0482_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__mux2_1
X_2881_ po_0.regf_0.rf\[3\]\[6\] _0776_ _1247_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__mux2_1
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1832_ po_0.regf_0.rf\[12\]\[6\] po_0.regf_0.rf\[13\]\[6\] po_0.regf_0.rf\[14\]\[6\]
+ po_0.regf_0.rf\[15\]\[6\] _0471_ _0472_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__mux4_1
X_1763_ _0420_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__buf_2
X_1694_ _0357_ _0358_ _1445_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ net173 _0335_ VGND VGND VPWR VPWR uc_0._03_ sky130_fd_sc_hd__dfxtp_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ net127 _0266_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_2315_ po_0.regf_0.rf\[6\]\[4\] _0755_ _0897_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__mux2_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _0852_ _0854_ _0670_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__a21oi_1
X_2177_ _1347_ po_0._1_\[6\] po_0._1_\[7\] _0621_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__a22o_1
XFILLER_53_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput36 net36 VGND VGND VPWR VPWR D_W_data[10] sky130_fd_sc_hd__clkbuf_4
Xoutput58 net58 VGND VGND VPWR VPWR D_addr[7] sky130_fd_sc_hd__buf_2
Xoutput47 net47 VGND VGND VPWR VPWR D_W_data[6] sky130_fd_sc_hd__buf_2
Xoutput69 net69 VGND VGND VPWR VPWR I_addr[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_56_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3080_ net121 _0059_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_2100_ po_0._1_\[2\] net43 VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__and2b_1
X_2031_ _0656_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__and2_1
XFILLER_47_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2933_ _1275_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2864_ po_0.regf_0.rf\[4\]\[15\] _0869_ _1220_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__mux2_1
X_2795_ net70 _1153_ _1147_ _1162_ _1190_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__o311a_1
X_1815_ po_0.regf_0.rf\[4\]\[4\] po_0.regf_0.rf\[5\]\[4\] po_0.regf_0.rf\[6\]\[4\]
+ po_0.regf_0.rf\[7\]\[4\] _0444_ _0445_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__mux4_1
X_1746_ _0398_ _0400_ _0402_ _0404_ VGND VGND VPWR VPWR po_0.regf_0._5_\[15\] sky130_fd_sc_hd__o22a_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1677_ po_0.regf_0.rf\[0\]\[7\] po_0.regf_0.rf\[1\]\[7\] po_0.regf_0.rf\[2\]\[7\]
+ po_0.regf_0.rf\[3\]\[7\] _1396_ _1397_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__mux4_1
X_3347_ net138 _0318_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ net167 net182 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfxtp_1
X_2229_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__clkbuf_2
XFILLER_26_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1600_ _0007_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__buf_2
X_2580_ po_0.regf_0.rf\[11\]\[3\] _0965_ _1052_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__mux2_1
X_1531_ _1343_ VGND VGND VPWR VPWR po_0.alu_0._10_\[0\] sky130_fd_sc_hd__clkbuf_1
X_3201_ net151 _0176_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3132_ net106 _0107_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3063_ po_0.regf_0._3_\[10\] net86 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlxtp_1
X_2014_ _0630_ _0632_ _0634_ _0642_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__a31oi_2
X_2916_ po_0.regf_0.rf\[2\]\[6\] _0776_ _1266_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2847_ _1229_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__clkbuf_1
X_2778_ net69 _0729_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__nand2_1
X_1729_ _0384_ _0386_ _1440_ _0389_ VGND VGND VPWR VPWR po_0.regf_0._5_\[13\] sky130_fd_sc_hd__o22a_1
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2701_ _1121_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2632_ po_0.regf_0.rf\[10\]\[11\] _0982_ _1078_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__mux2_1
X_2563_ po_0.regf_0.rf\[12\]\[12\] _0984_ _1031_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__mux2_1
X_1514_ _1333_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__clkbuf_1
X_2494_ po_0.regf_0.rf\[14\]\[13\] _0986_ _0992_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__mux2_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3115_ net130 _0090_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_3046_ po_0.regf_0._5_\[9\] net89 VGND VGND VPWR VPWR po_0._1_\[9\] sky130_fd_sc_hd__dlxtp_1
XFILLER_67_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout93 net61 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_2
XFILLER_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1994_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__inv_2
XFILLER_60_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2615_ po_0.regf_0.rf\[10\]\[3\] _0965_ _1071_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__mux2_1
X_2546_ po_0.regf_0.rf\[12\]\[4\] _0967_ _1032_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__mux2_1
X_2477_ po_0.regf_0.rf\[14\]\[5\] _0969_ _0993_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__mux2_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3029_ net130 _0040_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2400_ _0949_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
X_3380_ po_0.alu_0._10_\[1\] _1469_ VGND VGND VPWR VPWR po_0.alu_0._11_\[1\] sky130_fd_sc_hd__ebufn_1
X_2331_ _0910_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
X_2262_ _0869_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__clkbuf_2
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2193_ po_0.alu_0._11_\[9\] _0725_ _0720_ _0806_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__a211o_1
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1977_ _0602_ _0609_ _0605_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__nor3_1
XFILLER_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2529_ po_0.regf_0.rf\[13\]\[13\] _0986_ _1011_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__mux2_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1900_ po_0.regf_0.rf\[4\]\[13\] po_0.regf_0.rf\[5\]\[13\] po_0.regf_0.rf\[6\]\[13\]
+ po_0.regf_0.rf\[7\]\[13\] _0514_ _0515_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__mux4_1
X_2880_ _1239_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__buf_2
X_1831_ _0475_ _0477_ _0421_ _0483_ VGND VGND VPWR VPWR po_0.regf_0._3_\[5\] sky130_fd_sc_hd__o22a_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1762_ _0003_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__buf_2
X_1693_ po_0.regf_0.rf\[4\]\[9\] po_0.regf_0.rf\[5\]\[9\] po_0.regf_0.rf\[6\]\[9\]
+ po_0.regf_0.rf\[7\]\[9\] _1442_ _1443_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__mux4_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ net172 _0334_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfxtp_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ net135 _0265_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_2314_ _0901_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _0659_ po_0._1_\[13\] _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2176_ _0603_ _0609_ _0618_ _0781_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__nand4_1
XFILLER_80_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput37 net37 VGND VGND VPWR VPWR D_W_data[11] sky130_fd_sc_hd__buf_2
Xoutput48 net48 VGND VGND VPWR VPWR D_W_data[7] sky130_fd_sc_hd__buf_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput59 net59 VGND VGND VPWR VPWR D_rd sky130_fd_sc_hd__buf_2
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2030_ _0655_ po_0._1_\[12\] VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__or2_1
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2932_ po_0.regf_0.rf\[2\]\[14\] _0859_ _1258_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__mux2_1
X_2863_ _1237_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__clkbuf_1
X_2794_ _1146_ _1160_ _1183_ _1189_ _1148_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__a311o_1
X_1814_ _0457_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__and2b_1
X_1745_ _0403_ _1403_ _1404_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__a21o_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1676_ _0342_ _1418_ _1436_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__a21o_1
X_3346_ net139 _0317_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ net166 _0248_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfxtp_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ net4 _0685_ _0838_ _0713_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__a22o_2
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2159_ _0774_ _0713_ _0775_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__a21o_2
XFILLER_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1530_ _1341_ _1342_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__and2_1
X_3200_ net103 _0175_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_3131_ net109 _0106_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_3062_ po_0.regf_0._3_\[9\] net85 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlxtp_1
X_2013_ _0635_ _0640_ _0641_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__o21ai_1
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2915_ _1258_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__buf_2
XFILLER_50_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2846_ po_0.regf_0.rf\[4\]\[6\] _0776_ _1228_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__mux2_1
X_2777_ net69 po_0.muxf_0.rf_w_data\[2\] VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nor2_1
X_1728_ _0387_ _0388_ _1445_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__mux2_1
X_1659_ _1411_ _1457_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__and2b_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ net122 _0300_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2700_ po_0.regf_0.rf\[8\]\[10\] _0819_ _1116_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__mux2_1
X_2631_ _1083_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__clkbuf_1
X_2562_ _1045_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1513_ _1326_ _1328_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__or2b_1
X_2493_ _1007_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
X_3114_ net126 _0089_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_3045_ po_0.regf_0._5_\[8\] net88 VGND VGND VPWR VPWR po_0._1_\[8\] sky130_fd_sc_hd__dlxtp_1
XFILLER_55_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2829_ _1218_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__buf_2
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout83 net49 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout94 net82 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_2
XFILLER_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1993_ _0622_ _0623_ _0624_ _0617_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__o22ai_4
X_2614_ _1074_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
X_2545_ _1036_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
X_2476_ _0998_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3028_ net134 _0039_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2330_ po_0.regf_0.rf\[6\]\[11\] _0828_ _0904_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__mux2_1
X_2261_ _0862_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__nand2_2
X_2192_ _0804_ _0805_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__nor2_1
XFILLER_77_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1976_ _0602_ _0605_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__o21a_1
X_2528_ _1026_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
X_2459_ _0859_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__clkbuf_2
XFILLER_56_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1830_ _0480_ _0481_ _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__mux2_1
XFILLER_51_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1761_ _0415_ _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__and2b_1
X_1692_ po_0.regf_0.rf\[0\]\[9\] po_0.regf_0.rf\[1\]\[9\] po_0.regf_0.rf\[2\]\[9\]
+ po_0.regf_0.rf\[3\]\[9\] _1430_ _1431_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__mux4_1
X_3362_ net98 _0333_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfxtp_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ po_0.regf_0.rf\[6\]\[3\] _0742_ _0897_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__mux2_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ net134 _0264_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _0659_ po_0._1_\[13\] po_0._1_\[12\] _0655_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__o211a_1
X_2175_ _0715_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__buf_2
XFILLER_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1959_ _0589_ po_0._1_\[3\] VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__nand2_1
Xoutput49 net83 VGND VGND VPWR VPWR D_W_data[8] sky130_fd_sc_hd__buf_2
Xoutput38 net38 VGND VGND VPWR VPWR D_W_data[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2931_ _1274_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2862_ po_0.regf_0.rf\[4\]\[14\] _0859_ _1220_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__mux2_1
X_2793_ _1187_ _1188_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__nor2_1
XFILLER_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1813_ po_0.regf_0.rf\[0\]\[4\] po_0.regf_0.rf\[1\]\[4\] po_0.regf_0.rf\[2\]\[4\]
+ po_0.regf_0.rf\[3\]\[4\] _0449_ _0450_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux4_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1744_ po_0.regf_0.rf\[4\]\[15\] po_0.regf_0.rf\[5\]\[15\] po_0.regf_0.rf\[6\]\[15\]
+ po_0.regf_0.rf\[7\]\[15\] _1400_ _1401_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__mux4_1
X_1675_ po_0.regf_0.rf\[12\]\[7\] po_0.regf_0.rf\[13\]\[7\] po_0.regf_0.rf\[14\]\[7\]
+ po_0.regf_0.rf\[15\]\[7\] _1406_ _1407_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__mux4_1
X_3345_ net139 _0316_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ net166 _0247_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfxtp_2
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _0835_ _0836_ _0706_ _0837_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__a31o_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2158_ _0567_ _0682_ _0715_ net13 VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__a22o_1
X_2089_ _0705_ _0706_ _0707_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__a31o_1
XFILLER_83_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3130_ net106 _0105_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3061_ po_0.regf_0._3_\[8\] net85 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlxtp_1
X_2012_ po_0._1_\[9\] _0633_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__or2b_1
XFILLER_35_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2914_ _1265_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__clkbuf_1
X_2845_ _1220_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__buf_2
XFILLER_31_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2776_ net92 _0714_ _1169_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__a21oi_1
X_1727_ po_0.regf_0.rf\[4\]\[13\] po_0.regf_0.rf\[5\]\[13\] po_0.regf_0.rf\[6\]\[13\]
+ po_0.regf_0.rf\[7\]\[13\] _1442_ _1443_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__mux4_1
X_1658_ po_0.regf_0.rf\[8\]\[5\] po_0.regf_0.rf\[9\]\[5\] po_0.regf_0.rf\[10\]\[5\]
+ po_0.regf_0.rf\[11\]\[5\] _1412_ _1413_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__mux4_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ _1392_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__clkbuf_2
X_3328_ net130 _0299_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ net140 _0234_ VGND VGND VPWR VPWR uc_0._20_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2630_ po_0.regf_0.rf\[10\]\[10\] _0980_ _1078_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__mux2_1
X_2561_ po_0.regf_0.rf\[12\]\[11\] _0982_ _1039_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__mux2_1
X_2492_ po_0.regf_0.rf\[14\]\[12\] _0984_ _0992_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__mux2_1
X_1512_ _1332_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3113_ net128 _0088_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_3044_ po_0.regf_0._5_\[7\] net90 VGND VGND VPWR VPWR po_0._1_\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2828_ _1216_ _1217_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__nor2_1
X_2759_ net67 net64 _1156_ _1157_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__or4_1
XFILLER_78_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout95 net81 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_4
Xfanout84 net45 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1992_ po_0._1_\[6\] _1347_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__and2b_1
XFILLER_9_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2613_ po_0.regf_0.rf\[10\]\[2\] _0963_ _1071_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__mux2_1
X_2544_ po_0.regf_0.rf\[12\]\[3\] _0965_ _1032_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__mux2_1
X_2475_ po_0.regf_0.rf\[14\]\[4\] _0967_ _0993_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__mux2_1
XFILLER_83_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3027_ net132 _0038_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2260_ _0863_ _0865_ _0867_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__o21ai_1
X_2191_ _0628_ _0634_ _0796_ _0724_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__a31o_1
XFILLER_45_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1975_ _0607_ _0608_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__nor2_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2527_ po_0.regf_0.rf\[13\]\[12\] _0984_ _1011_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2458_ _0987_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2389_ _0943_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1760_ po_0.regf_0.rf\[8\]\[0\] po_0.regf_0.rf\[9\]\[0\] po_0.regf_0.rf\[10\]\[0\]
+ po_0.regf_0.rf\[11\]\[0\] _0416_ _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux4_1
X_1691_ _1411_ _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__and2b_1
X_3361_ net139 _0332_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2312_ _0900_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ net135 _0263_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _0834_ _0851_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__nand2_1
XFILLER_57_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2174_ _0789_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
X_1958_ _0585_ _0576_ _0586_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__a21oi_1
X_1889_ po_0.regf_0.rf\[8\]\[12\] po_0.regf_0.rf\[9\]\[12\] po_0.regf_0.rf\[10\]\[12\]
+ po_0.regf_0.rf\[11\]\[12\] _0509_ _0510_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__mux4_1
Xoutput39 net39 VGND VGND VPWR VPWR D_W_data[13] sky130_fd_sc_hd__buf_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2930_ po_0.regf_0.rf\[2\]\[13\] _0848_ _1258_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__mux2_1
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2861_ _1236_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__clkbuf_1
X_2792_ _1186_ _1185_ _1184_ _1147_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__a31o_1
X_1812_ _0465_ _0411_ _0412_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__a21bo_1
X_1743_ _1411_ _0401_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__and2b_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1674_ _1433_ _0340_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__and2b_1
X_3344_ net110 _0315_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ net152 _0246_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfxtp_2
X_2226_ _0708_ po_0.alu_0._11_\[12\] _0709_ _0655_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__a22o_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2157_ _0771_ _0772_ _0706_ _0773_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__a31o_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2088_ _0708_ po_0.alu_0._11_\[1\] _0709_ _0574_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__a22o_1
XFILLER_5_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3060_ po_0.regf_0._3_\[7\] net85 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlxtp_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2011_ net50 po_0._1_\[9\] VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__xor2_2
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2913_ po_0.regf_0.rf\[2\]\[5\] _0764_ _1259_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__mux2_1
X_2844_ _1227_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__clkbuf_1
X_2775_ _1163_ _1153_ _1147_ _1172_ _1162_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__o311a_1
X_1726_ po_0.regf_0.rf\[0\]\[13\] po_0.regf_0.rf\[1\]\[13\] po_0.regf_0.rf\[2\]\[13\]
+ po_0.regf_0.rf\[3\]\[13\] _1430_ _1431_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__mux4_1
XFILLER_7_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1657_ _1455_ _1409_ _1436_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__a21o_1
X_1588_ _0007_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__clkinv_2
X_3327_ net122 _0298_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ net114 _0233_ VGND VGND VPWR VPWR uc_0._20_\[9\] sky130_fd_sc_hd__dfxtp_1
X_2209_ _0821_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
X_3189_ net158 _0164_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2560_ _1044_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
X_2491_ _1006_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
X_1511_ _1326_ _1328_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__or2b_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3112_ net133 _0087_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3043_ po_0.regf_0._5_\[6\] net89 VGND VGND VPWR VPWR po_0._1_\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_63_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2827_ _1215_ _1366_ uc_0.bc_0._54_\[1\] _1361_ _1356_ VGND VGND VPWR VPWR _1217_
+ sky130_fd_sc_hd__o2111a_1
X_2758_ net63 net62 net76 net75 VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__or4_1
X_1709_ _0371_ _1391_ _1393_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a21o_1
X_2689_ po_0.regf_0.rf\[8\]\[5\] _0764_ _1109_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__mux2_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout96 net105 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout85 net87 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1991_ _0621_ po_0._1_\[7\] VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__and2_1
XFILLER_9_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2612_ _1073_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2543_ _1035_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
X_2474_ _0997_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3026_ net163 _0037_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2190_ _0628_ _0796_ _0634_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1974_ _0606_ po_0._1_\[5\] VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__and2_1
X_2526_ _1025_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
X_2457_ po_0.regf_0.rf\[15\]\[13\] _0986_ _0958_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__mux2_1
X_2388_ po_0.regf_0.rf\[1\]\[4\] _0755_ _0938_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__mux2_1
XFILLER_83_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3009_ net165 _0020_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1690_ po_0.regf_0.rf\[8\]\[9\] po_0.regf_0.rf\[9\]\[9\] po_0.regf_0.rf\[10\]\[9\]
+ po_0.regf_0.rf\[11\]\[9\] _1412_ _1413_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux4_1
X_3360_ net153 _0331_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfxtp_1
X_2311_ po_0.regf_0.rf\[6\]\[2\] _0732_ _0897_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__mux2_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ net163 _0262_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ _0660_ _0657_ _0656_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__and3_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2173_ po_0.regf_0.rf\[7\]\[7\] _0788_ _0778_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__mux2_1
XFILLER_80_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1957_ _0580_ _0581_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__nand2_1
X_1888_ _0533_ _0433_ _0474_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2509_ _1016_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2860_ po_0.regf_0.rf\[4\]\[13\] _0848_ _1220_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__mux2_1
X_1811_ po_0.regf_0.rf\[12\]\[4\] po_0.regf_0.rf\[13\]\[4\] po_0.regf_0.rf\[14\]\[4\]
+ po_0.regf_0.rf\[15\]\[4\] _0406_ _0408_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__mux4_1
X_2791_ _1184_ _1185_ _1186_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__a21oi_1
X_1742_ po_0.regf_0.rf\[0\]\[15\] po_0.regf_0.rf\[1\]\[15\] po_0.regf_0.rf\[2\]\[15\]
+ po_0.regf_0.rf\[3\]\[15\] _1412_ _1413_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__mux4_1
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1673_ po_0.regf_0.rf\[8\]\[7\] po_0.regf_0.rf\[9\]\[7\] po_0.regf_0.rf\[10\]\[7\]
+ po_0.regf_0.rf\[11\]\[7\] _1427_ _1428_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__mux4_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ net138 _0314_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ net166 _0245_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfxtp_2
X_2225_ _0834_ _0658_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__nand2_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2156_ _0708_ po_0.alu_0._11_\[6\] _0709_ _1347_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__a22o_1
X_2087_ _0688_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__buf_2
XFILLER_41_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2989_ _1305_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2010_ _0637_ _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__nand2b_2
XFILLER_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2912_ _1264_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2843_ po_0.regf_0.rf\[4\]\[5\] _0764_ _1221_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__mux2_1
X_2774_ _1164_ _1165_ _1166_ _1171_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__o31ai_1
X_1725_ _1378_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__and2b_1
X_1656_ po_0.regf_0.rf\[12\]\[5\] po_0.regf_0.rf\[13\]\[5\] po_0.regf_0.rf\[14\]\[5\]
+ po_0.regf_0.rf\[15\]\[5\] _1406_ _1407_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__mux4_1
X_1587_ _1390_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__clkbuf_2
X_3326_ net129 _0297_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ net138 _0232_ VGND VGND VPWR VPWR uc_0._20_\[8\] sky130_fd_sc_hd__dfxtp_1
X_2208_ po_0.regf_0.rf\[7\]\[10\] _0820_ _0778_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__mux2_1
X_3188_ net158 _0163_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2139_ _0746_ _0750_ _0603_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__o21a_1
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2490_ po_0.regf_0.rf\[14\]\[11\] _0982_ _1000_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__mux2_1
X_1510_ _1331_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3111_ net132 _0086_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3042_ po_0.regf_0._5_\[5\] net90 VGND VGND VPWR VPWR po_0._1_\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2826_ _1215_ _1366_ _1368_ _1356_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__o211a_1
X_2757_ net74 net73 net72 net71 VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__or4_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1708_ po_0.regf_0.rf\[12\]\[11\] po_0.regf_0.rf\[13\]\[11\] po_0.regf_0.rf\[14\]\[11\]
+ po_0.regf_0.rf\[15\]\[11\] _1386_ _1388_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__mux4_1
X_2688_ _1114_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__clkbuf_1
X_1639_ _0007_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__buf_2
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ net131 _0280_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout97 net98 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout86 net87 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1990_ _0621_ po_0._1_\[7\] VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__nor2_2
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2611_ po_0.regf_0.rf\[10\]\[1\] _0961_ _1071_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__mux2_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2542_ po_0.regf_0.rf\[12\]\[2\] _0963_ _1032_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__mux2_1
X_2473_ po_0.regf_0.rf\[14\]\[3\] _0965_ _0993_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__mux2_1
XFILLER_68_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3025_ net169 _0036_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2809_ _1202_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1973_ _0606_ po_0._1_\[5\] VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__nor2_2
X_2525_ po_0.regf_0.rf\[13\]\[11\] _0982_ _1019_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__mux2_1
X_2456_ _0848_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__clkbuf_2
X_2387_ _0942_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3008_ net161 _0019_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2310_ _0899_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
X_3290_ net161 _0261_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _0850_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2172_ _0787_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1956_ _0580_ _0584_ _0590_ _0591_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__o2bb2ai_1
X_1887_ po_0.regf_0.rf\[12\]\[12\] po_0.regf_0.rf\[13\]\[12\] po_0.regf_0.rf\[14\]\[12\]
+ po_0.regf_0.rf\[15\]\[12\] _0471_ _0472_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__mux4_1
X_2508_ po_0.regf_0.rf\[13\]\[3\] _0965_ _1012_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__mux2_1
X_2439_ po_0.regf_0.rf\[15\]\[7\] _0974_ _0972_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__mux2_1
XFILLER_29_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1810_ _0430_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__and2b_1
X_2790_ _1173_ _1174_ _1175_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__o21ai_1
X_1741_ _0399_ _1418_ _1436_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__a21o_1
XFILLER_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1672_ _1463_ _1465_ _1467_ _0339_ VGND VGND VPWR VPWR po_0.regf_0._5_\[6\] sky130_fd_sc_hd__o22a_1
X_3342_ net153 _0313_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ net166 _0244_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfxtp_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _0656_ _0657_ _0834_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__a21o_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _0606_ po_0._1_\[5\] _0769_ _0757_ _0618_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__o221ai_2
XFILLER_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2086_ _1316_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__buf_2
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2988_ po_0.muxf_0.rf_w_data\[3\] net54 _1303_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__mux2_1
XFILLER_21_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1939_ _0575_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__nand2_1
XFILLER_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2911_ po_0.regf_0.rf\[2\]\[4\] _0754_ _1259_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__mux2_1
XFILLER_31_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2842_ _1226_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__clkbuf_1
X_2773_ uc_0._00_ uc_0._02_ _1169_ _1170_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__or4b_1
X_1724_ po_0.regf_0.rf\[8\]\[13\] po_0.regf_0.rf\[9\]\[13\] po_0.regf_0.rf\[10\]\[13\]
+ po_0.regf_0.rf\[11\]\[13\] _1380_ _1382_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__mux4_1
X_1655_ _1448_ _1450_ _1452_ _1454_ VGND VGND VPWR VPWR po_0.regf_0._5_\[4\] sky130_fd_sc_hd__o22a_1
X_1586_ _0006_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ net131 _0296_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ net137 _0231_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[7\] sky130_fd_sc_hd__dfxtp_2
X_2207_ _0819_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__clkbuf_2
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ net150 _0162_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2138_ _0756_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
X_2069_ _1340_ _0686_ _1314_ _0687_ _0691_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__o311a_1
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3110_ net156 _0085_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3041_ po_0.regf_0._5_\[4\] net90 VGND VGND VPWR VPWR po_0._1_\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2825_ _1357_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2756_ _1151_ _1152_ _1153_ _1154_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__and4_1
X_1707_ _1378_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__and2b_1
X_2687_ po_0.regf_0.rf\[8\]\[4\] _0754_ _1109_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__mux2_1
X_1638_ _1411_ _1438_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__and2b_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ _1375_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__clkbuf_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ net128 _0279_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ net115 _0214_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout98 net105 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
Xfanout87 po_0.regf_0.rp_rd VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
XFILLER_10_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2610_ _1072_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__clkbuf_1
X_2541_ _1034_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
X_2472_ _0996_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3024_ net161 _0035_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2808_ _1200_ _1195_ _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__and3_1
X_2739_ net79 net20 _1133_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__mux2_1
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1972_ net46 VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__clkbuf_2
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2524_ _1024_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
X_2455_ _0985_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
X_2386_ po_0.regf_0.rf\[1\]\[3\] _0742_ _0938_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__mux2_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3007_ net147 _0018_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ po_0.regf_0.rf\[7\]\[13\] _0849_ _0700_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__mux2_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2171_ po_0.muxf_0.rf_w_data\[7\] _0683_ _0685_ net14 _0786_ VGND VGND VPWR VPWR
+ _0787_ sky130_fd_sc_hd__a221o_2
XFILLER_46_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1955_ _0589_ po_0._1_\[3\] VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__nor2_1
X_1886_ _0527_ _0529_ _0421_ _0532_ VGND VGND VPWR VPWR po_0.regf_0._3_\[11\] sky130_fd_sc_hd__o22a_1
X_2507_ _1015_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
X_2438_ _0787_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__clkbuf_2
X_2369_ _0931_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1740_ po_0.regf_0.rf\[12\]\[15\] po_0.regf_0.rf\[13\]\[15\] po_0.regf_0.rf\[14\]\[15\]
+ po_0.regf_0.rf\[15\]\[15\] _1406_ _1407_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__mux4_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1671_ _0338_ _1403_ _1404_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a21o_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3341_ net153 _0312_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ net167 _0243_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfxtp_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _0644_ _0831_ _0832_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__o22ai_2
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _0613_ _0614_ _0770_ _0607_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__o22ai_1
XFILLER_38_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2085_ _0586_ _0704_ _0703_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__o21ai_2
X_2987_ _1304_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1938_ net42 po_0._1_\[1\] VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__or2b_1
X_1869_ _0507_ _0512_ _0421_ _0517_ VGND VGND VPWR VPWR po_0.regf_0._3_\[9\] sky130_fd_sc_hd__o22a_1
XFILLER_67_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2910_ _1263_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2841_ po_0.regf_0.rf\[4\]\[4\] _0754_ _1221_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__mux2_1
X_2772_ net93 po_0.muxf_0.rf_w_data\[0\] _1168_ _1167_ VGND VGND VPWR VPWR _1170_
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1723_ _0383_ _1395_ _1392_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__a21o_1
X_1654_ _1453_ _1403_ _1404_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__a21o_1
X_1585_ po_0.regf_0.rf\[12\]\[0\] po_0.regf_0.rf\[13\]\[0\] po_0.regf_0.rf\[14\]\[0\]
+ po_0.regf_0.rf\[15\]\[0\] _1386_ _1388_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__mux4_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ net129 _0295_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3255_ net153 _0230_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[6\] sky130_fd_sc_hd__dfxtp_1
X_2206_ net2 _0790_ _0818_ _0713_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__a22o_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ net145 _0161_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2137_ po_0.regf_0.rf\[7\]\[4\] _0755_ _0701_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__mux2_1
X_2068_ _1317_ po_0.alu_0._11_\[0\] _0688_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__a211o_1
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3040_ po_0.regf_0._5_\[3\] net90 VGND VGND VPWR VPWR po_0._1_\[3\] sky130_fd_sc_hd__dlxtp_1
X_2824_ _1214_ _1211_ _1154_ _1153_ _1162_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__o2111a_1
X_2755_ uc_0._00_ uc_0._02_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__nor2_1
X_1706_ po_0.regf_0.rf\[0\]\[11\] po_0.regf_0.rf\[1\]\[11\] po_0.regf_0.rf\[2\]\[11\]
+ po_0.regf_0.rf\[3\]\[11\] _1380_ _1382_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux4_1
X_2686_ _1113_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__clkbuf_1
X_1637_ po_0.regf_0.rf\[8\]\[3\] po_0.regf_0.rf\[9\]\[3\] po_0.regf_0.rf\[10\]\[3\]
+ po_0.regf_0.rf\[11\]\[3\] _1412_ _1413_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__mux4_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ uc_0._20_\[9\] po_0.regf_0.rp_addr\[1\] _1373_ VGND VGND VPWR VPWR _1375_
+ sky130_fd_sc_hd__mux2_1
X_3307_ net157 _0278_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1315_ _1319_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__or2b_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ net156 _0213_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3169_ net148 _0144_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout99 net102 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout88 net91 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2540_ po_0.regf_0.rf\[12\]\[1\] _0961_ _1032_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__mux2_1
XFILLER_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2471_ po_0.regf_0.rf\[14\]\[2\] _0963_ _0993_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__mux2_1
XFILLER_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3023_ net150 _0034_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2807_ _1191_ _1199_ _1196_ _1197_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__o211ai_2
X_2738_ _1141_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__clkbuf_1
X_2669_ _0840_ po_0.regf_0.rf\[0\]\[12\] _1089_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__mux2_1
XFILLER_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1971_ po_0._1_\[4\] net84 VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__and2b_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2523_ po_0.regf_0.rf\[13\]\[10\] _0980_ _1019_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__mux2_1
X_2454_ po_0.regf_0.rf\[15\]\[12\] _0984_ _0958_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__mux2_1
XFILLER_68_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2385_ _0941_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 D_R_data[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3006_ net143 _0017_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _0725_ _0782_ _0783_ _0785_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__o31a_1
XFILLER_65_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1954_ _0589_ po_0._1_\[3\] VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__and2_1
X_1885_ _0530_ _0531_ _0482_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2506_ po_0.regf_0.rf\[13\]\[2\] _0963_ _1012_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__mux2_1
X_2437_ _0973_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
X_2368_ po_0.regf_0.rf\[9\]\[12\] _0840_ _0916_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__mux2_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2299_ _0892_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1670_ po_0.regf_0.rf\[4\]\[6\] po_0.regf_0.rf\[5\]\[6\] po_0.regf_0.rf\[6\]\[6\]
+ po_0.regf_0.rf\[7\]\[6\] _1400_ _1401_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__mux4_1
X_3340_ net152 _0311_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ net167 _0242_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfxtp_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2222_ _0768_ _0797_ _0794_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__a21oi_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2153_ _0768_ _0603_ _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2084_ _0689_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__buf_2
XFILLER_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2986_ _0729_ net53 _1303_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__mux2_1
X_1937_ _0573_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__or2b_1
X_1868_ _0513_ _0516_ _0482_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__mux2_1
X_1799_ _0430_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__and2b_1
XFILLER_67_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2840_ _1225_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2771_ _1167_ po_0.muxf_0.rf_w_data\[0\] net93 _1168_ VGND VGND VPWR VPWR _1169_
+ sky130_fd_sc_hd__and4_1
X_1722_ po_0.regf_0.rf\[12\]\[13\] po_0.regf_0.rf\[13\]\[13\] po_0.regf_0.rf\[14\]\[13\]
+ po_0.regf_0.rf\[15\]\[13\] _1419_ _1420_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__mux4_1
X_1653_ po_0.regf_0.rf\[4\]\[4\] po_0.regf_0.rf\[5\]\[4\] po_0.regf_0.rf\[6\]\[4\]
+ po_0.regf_0.rf\[7\]\[4\] _1400_ _1401_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__mux4_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1584_ _1387_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__buf_2
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ net157 _0294_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ net153 _0229_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[5\] sky130_fd_sc_hd__dfxtp_1
X_2205_ _0814_ _0725_ _0816_ _0817_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__o31ai_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ net151 _0160_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2136_ _0754_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__clkbuf_2
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2067_ _1341_ _1342_ _0689_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__and3_1
XFILLER_81_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2969_ _1294_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2823_ net74 _0570_ net75 VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__a21o_1
X_2754_ uc_0._01_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__clkbuf_2
X_1705_ _0367_ _1409_ _0007_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__a21o_1
X_2685_ po_0.regf_0.rf\[8\]\[3\] _0741_ _1109_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__mux2_1
X_1636_ _1435_ _1409_ _1436_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__a21o_1
X_1567_ _1374_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ net168 _0277_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1323_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__clkbuf_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ net159 _0212_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3168_ net97 _0143_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2119_ _1317_ po_0.alu_0._11_\[3\] _0688_ _0738_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__a211o_1
XFILLER_54_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3099_ net130 _0074_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout89 net91 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2470_ _0995_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3022_ net143 _0033_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2806_ net71 _0561_ _1196_ _1197_ _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__a221o_1
X_2737_ uc_0._20_\[11\] net19 _1133_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__mux2_1
X_2668_ _1103_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__clkbuf_1
X_1619_ _1418_ _1421_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__and2b_1
X_2599_ po_0.regf_0.rf\[11\]\[12\] _0984_ _1051_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__mux2_1
XFILLER_75_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1970_ _0602_ _0604_ VGND VGND VPWR VPWR po_0.alu_0._10_\[4\] sky130_fd_sc_hd__nor2_1
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2522_ _1023_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2453_ _0839_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__clkbuf_2
X_2384_ po_0.regf_0.rf\[1\]\[2\] _0732_ _0938_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__mux2_1
XFILLER_68_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput2 D_R_data[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3005_ net169 _0016_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1953_ net44 VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1884_ po_0.regf_0.rf\[4\]\[11\] po_0.regf_0.rf\[5\]\[11\] po_0.regf_0.rf\[6\]\[11\]
+ po_0.regf_0.rf\[7\]\[11\] _0514_ _0515_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__mux4_1
X_2505_ _1014_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
X_2436_ po_0.regf_0.rf\[15\]\[6\] _0971_ _0972_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__mux2_1
X_2367_ _0930_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
X_2298_ po_0.regf_0.rf\[5\]\[13\] _0849_ _0876_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__mux2_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3270_ net172 _0241_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfxtp_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _0648_ _0640_ _0639_ _0646_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__nand4_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2152_ net45 po_0._1_\[4\] po_0._1_\[5\] _0606_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__a22o_1
X_2083_ _0703_ _0586_ _0704_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__or3_1
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2985_ _1299_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__clkbuf_8
X_1936_ net42 VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__clkbuf_2
X_1867_ po_0.regf_0.rf\[4\]\[9\] po_0.regf_0.rf\[5\]\[9\] po_0.regf_0.rf\[6\]\[9\]
+ po_0.regf_0.rf\[7\]\[9\] _0514_ _0515_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__mux4_1
X_1798_ po_0.regf_0.rf\[8\]\[3\] po_0.regf_0.rf\[9\]\[3\] po_0.regf_0.rf\[10\]\[3\]
+ po_0.regf_0.rf\[11\]\[3\] _0423_ _0425_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__mux4_1
X_2419_ _0717_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__clkbuf_2
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2770_ net92 po_0.muxf_0.rf_w_data\[1\] VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__nand2_1
X_1721_ _0376_ _0378_ _0380_ _0382_ VGND VGND VPWR VPWR po_0.regf_0._5_\[12\] sky130_fd_sc_hd__o22a_1
X_1652_ _1395_ _1451_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__and2b_1
X_1583_ _0005_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__buf_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ net168 _0293_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3253_ net166 _0228_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[4\] sky130_fd_sc_hd__dfxtp_1
X_3184_ net103 _0159_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_2204_ _0686_ po_0.alu_0._11_\[10\] _0709_ net36 VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__a22oi_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _0561_ _0683_ _0685_ net11 _0753_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__a221o_2
XFILLER_26_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2066_ _1316_ po_0.alu_0.s0 VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__and2b_1
XFILLER_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2968_ _0699_ _1293_ _1280_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__mux2_1
X_1919_ po_0.muxf_0.rf_w_data\[4\] VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__buf_2
X_2899_ po_0.regf_0.rf\[3\]\[15\] _0869_ _1239_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__mux2_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2822_ _1213_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__clkbuf_1
X_2753_ _1149_ _0681_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__nand2_1
X_1704_ po_0.regf_0.rf\[4\]\[11\] po_0.regf_0.rf\[5\]\[11\] po_0.regf_0.rf\[6\]\[11\]
+ po_0.regf_0.rf\[7\]\[11\] _1419_ _1420_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__mux4_1
X_2684_ _1112_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__clkbuf_1
X_1635_ _1392_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__clkbuf_2
X_1566_ uc_0._20_\[8\] po_0.regf_0.rp_addr\[0\] _1373_ VGND VGND VPWR VPWR _1374_
+ sky130_fd_sc_hd__mux2_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ net159 _0276_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ _1315_ _1319_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__or2b_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3236_ net158 _0211_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3167_ net98 _0142_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3098_ net132 _0073_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_2118_ _0734_ _0736_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__a21oi_1
X_2049_ net41 po_0._1_\[15\] VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__and2_1
XFILLER_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3021_ net169 _0032_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2805_ _1198_ _1193_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__nor2_1
X_2736_ _1140_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__clkbuf_1
X_2667_ _0828_ po_0.regf_0.rf\[0\]\[11\] _1097_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__mux2_1
X_1618_ po_0.regf_0.rf\[8\]\[1\] po_0.regf_0.rf\[9\]\[1\] po_0.regf_0.rf\[10\]\[1\]
+ po_0.regf_0.rf\[11\]\[1\] _1419_ _1420_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__mux4_1
X_2598_ _1065_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__clkbuf_1
X_1549_ _1344_ _1354_ _1359_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__o21ba_1
X_3219_ net151 _0194_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2521_ po_0.regf_0.rf\[13\]\[9\] _0978_ _1019_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__mux2_1
X_2452_ _0983_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2383_ _0940_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 D_R_data[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
X_3004_ _1312_ _1355_ _1153_ _1219_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2719_ po_0.muxf_0.rf_w_data\[3\] net26 _1127_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__mux2_1
XFILLER_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1952_ _0588_ VGND VGND VPWR VPWR po_0.alu_0._10_\[2\] sky130_fd_sc_hd__clkbuf_1
X_1883_ po_0.regf_0.rf\[0\]\[11\] po_0.regf_0.rf\[1\]\[11\] po_0.regf_0.rf\[2\]\[11\]
+ po_0.regf_0.rf\[3\]\[11\] _0478_ _0479_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__mux4_1
X_2504_ po_0.regf_0.rf\[13\]\[1\] _0961_ _1012_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__mux2_1
X_2435_ _0958_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__buf_2
X_2366_ po_0.regf_0.rf\[9\]\[11\] _0828_ _0924_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__mux2_1
X_2297_ _0891_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_30 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _0812_ _0813_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__o21a_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2151_ _0749_ _0767_ _0746_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__o21bai_2
X_2082_ _0574_ _0573_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__and2b_1
XFILLER_19_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2984_ _1302_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__clkbuf_1
X_1935_ po_0._1_\[1\] VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__clkbuf_2
X_1866_ _0424_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__buf_2
X_1797_ _0441_ _0443_ _0448_ _0452_ VGND VGND VPWR VPWR po_0.regf_0._3_\[2\] sky130_fd_sc_hd__o22a_1
X_2418_ _0960_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2349_ po_0.regf_0.rf\[9\]\[3\] _0742_ _0917_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__mux2_1
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1720_ _0381_ _1403_ _1404_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__a21o_1
X_1651_ po_0.regf_0.rf\[0\]\[4\] po_0.regf_0.rf\[1\]\[4\] po_0.regf_0.rf\[2\]\[4\]
+ po_0.regf_0.rf\[3\]\[4\] _1396_ _1397_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__mux4_1
X_1582_ _1385_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__clkbuf_4
X_3321_ net158 _0292_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ net171 _0227_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[3\] sky130_fd_sc_hd__dfxtp_4
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ net98 _0158_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_2203_ _0639_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__nor2_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2134_ _0744_ _0752_ _0712_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__o21a_1
XFILLER_81_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2065_ _1316_ _1313_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__nor2_2
X_2967_ uc_0._20_\[10\] _0729_ _0562_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__mux2_1
X_1918_ _0555_ _0557_ _0461_ _0560_ VGND VGND VPWR VPWR po_0.regf_0._3_\[15\] sky130_fd_sc_hd__o22a_1
X_2898_ _1256_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1849_ po_0.regf_0.rf\[0\]\[8\] po_0.regf_0.rf\[1\]\[8\] po_0.regf_0.rf\[2\]\[8\]
+ po_0.regf_0.rf\[3\]\[8\] _0422_ _0424_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__mux4_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2821_ _1211_ _1212_ _1195_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__and3b_1
X_2752_ _1149_ _0681_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__or2_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1703_ _0361_ _0363_ _1440_ _0366_ VGND VGND VPWR VPWR po_0.regf_0._5_\[10\] sky130_fd_sc_hd__o22a_1
X_2683_ po_0.regf_0.rf\[8\]\[2\] _0731_ _1109_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__mux2_1
X_1634_ po_0.regf_0.rf\[12\]\[3\] po_0.regf_0.rf\[13\]\[3\] po_0.regf_0.rf\[14\]\[3\]
+ po_0.regf_0.rf\[15\]\[3\] _1406_ _1407_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__mux4_1
X_1565_ _1372_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__clkbuf_2
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ net150 _0275_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _1322_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__clkbuf_1
X_3235_ net154 _0210_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3166_ net98 _0141_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3097_ net113 _0072_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_2117_ _0734_ _0736_ _0689_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__o21ai_1
XFILLER_54_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2048_ _0670_ _0672_ VGND VGND VPWR VPWR po_0.alu_0._10_\[14\] sky130_fd_sc_hd__xor2_1
XFILLER_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3020_ net118 _0031_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2804_ _1191_ _1192_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__or2_1
XFILLER_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2735_ uc_0._20_\[10\] net18 _1134_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__mux2_1
X_2666_ _1102_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__clkbuf_1
X_1617_ _1381_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__clkbuf_4
X_2597_ po_0.regf_0.rf\[11\]\[11\] _0982_ _1059_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__mux2_1
X_1548_ net79 net94 _1358_ _1344_ uc_0.bc_0._55_\[1\] VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__o311a_1
X_3218_ net144 _0193_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3149_ net96 _0124_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2520_ _1022_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
X_2451_ po_0.regf_0.rf\[15\]\[11\] _0982_ _0972_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__mux2_1
XFILLER_5_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2382_ po_0.regf_0.rf\[1\]\[1\] _0718_ _0938_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__mux2_1
XFILLER_83_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput4 D_R_data[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
X_3003_ _1215_ _1359_ _1365_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__or3_1
XFILLER_76_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2718_ _1130_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__clkbuf_1
X_2649_ _1093_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1951_ _0584_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__and2_1
X_1882_ _0508_ _0528_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__and2b_1
X_2503_ _1013_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
X_2434_ _0776_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__clkbuf_2
X_2365_ _0929_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
X_2296_ po_0.regf_0.rf\[5\]\[12\] _0840_ _0876_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__mux2_1
XFILLER_37_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_20 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2150_ _0577_ _0703_ _0748_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__a21boi_1
X_2081_ po_0._1_\[0\] _1340_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__and2_1
XFILLER_19_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2983_ _0714_ net52 _1300_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__mux2_1
XFILLER_61_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1934_ _1340_ po_0._1_\[0\] VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__and2b_1
X_1865_ _0422_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__clkbuf_4
X_1796_ _0411_ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__and2b_1
X_2417_ po_0.regf_0.rf\[15\]\[0\] _0956_ _0959_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__mux2_1
X_2348_ _0920_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
X_2279_ po_0.regf_0.rf\[5\]\[4\] _0755_ _0877_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__mux2_1
XFILLER_32_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1650_ _1449_ _1391_ _1393_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__a21o_1
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1581_ _0004_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__buf_2
X_3320_ net151 _0291_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ net171 _0226_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[2\] sky130_fd_sc_hd__dfxtp_1
X_3182_ net98 _0157_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2202_ _0812_ _0796_ po_0._1_\[9\] _0633_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__o2bb2a_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2133_ _0599_ _0600_ _0747_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__o31a_1
X_2064_ _0682_ _0684_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__nor2_2
XFILLER_22_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2966_ _1292_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__clkbuf_1
X_1917_ _0558_ _0559_ _0410_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__mux2_1
X_2897_ po_0.regf_0.rf\[3\]\[14\] _0859_ _1239_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__mux2_1
X_1848_ _0492_ _0494_ _0496_ _0498_ VGND VGND VPWR VPWR po_0.regf_0._3_\[7\] sky130_fd_sc_hd__o22a_1
X_1779_ _0415_ _0435_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__and2b_1
XFILLER_1_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2820_ net73 _0567_ _1209_ _1210_ _1206_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__a221o_1
X_2751_ _1146_ _1148_ _1149_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__mux2_1
X_1702_ _0364_ _0365_ _1445_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__mux2_1
X_2682_ _1111_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__clkbuf_1
X_1633_ _1424_ _1426_ _1393_ _1434_ VGND VGND VPWR VPWR po_0.regf_0._5_\[2\] sky130_fd_sc_hd__o22a_1
X_1564_ _1367_ _1368_ _1371_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__a21oi_4
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _1315_ _1319_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__or2b_1
X_3303_ net144 _0274_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ net145 _0209_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ net96 _0140_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3096_ net134 _0071_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2116_ _0593_ _0723_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__a21bo_1
X_2047_ _0671_ po_0._1_\[13\] _0665_ _0654_ _0667_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__o221ai_4
XFILLER_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2949_ po_0.regf_0.rq_addr\[2\] _0567_ _0568_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__mux2_1
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2803_ net72 po_0.muxf_0.rf_w_data\[5\] VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__or2_1
X_2734_ _1139_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__clkbuf_1
X_2665_ _0820_ po_0.regf_0.rf\[0\]\[10\] _1097_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__mux2_1
X_2596_ _1064_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__clkbuf_1
X_1616_ _1379_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__clkbuf_4
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1547_ net80 net95 uc_0.bc_0._55_\[0\] VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__a21bo_1
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3217_ net164 _0192_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3148_ net106 _0123_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3079_ net133 _0058_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2450_ _0827_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__clkbuf_2
X_2381_ _0939_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
Xinput5 D_R_data[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_3002_ _1311_ _1367_ _1216_ _1146_ _1300_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__o221a_1
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2717_ _0729_ net25 _1127_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__mux2_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2648_ _0732_ po_0.regf_0.rf\[0\]\[2\] _1090_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__mux2_1
X_2579_ _1055_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1950_ _0585_ _0576_ _0580_ _0581_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__a221o_1
XFILLER_14_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1881_ po_0.regf_0.rf\[8\]\[11\] po_0.regf_0.rf\[9\]\[11\] po_0.regf_0.rf\[10\]\[11\]
+ po_0.regf_0.rf\[11\]\[11\] _0509_ _0510_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__mux4_1
X_2502_ po_0.regf_0.rf\[13\]\[0\] _0956_ _1012_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__mux2_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2433_ _0970_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
X_2364_ po_0.regf_0.rf\[9\]\[10\] _0820_ _0924_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__mux2_1
X_2295_ _0890_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_10 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2080_ _0702_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2982_ _1301_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__clkbuf_1
X_1933_ _0571_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1864_ po_0.regf_0.rf\[0\]\[9\] po_0.regf_0.rf\[1\]\[9\] po_0.regf_0.rf\[2\]\[9\]
+ po_0.regf_0.rf\[3\]\[9\] _0478_ _0479_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__mux4_1
Xinput30 I_data[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
X_1795_ po_0.regf_0.rf\[8\]\[2\] po_0.regf_0.rf\[9\]\[2\] po_0.regf_0.rf\[10\]\[2\]
+ po_0.regf_0.rf\[11\]\[2\] _0449_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__mux4_1
X_2416_ _0958_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__buf_2
X_2347_ po_0.regf_0.rf\[9\]\[2\] _0732_ _0917_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__mux2_1
X_2278_ _0881_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1580_ _1378_ _1383_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__and2b_1
XFILLER_3_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ net172 _0225_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ net97 _0156_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_2201_ _0796_ _0812_ _0813_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__a21oi_2
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2132_ _0603_ _0746_ _0750_ _0689_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__o31a_1
X_2063_ _1316_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__clkbuf_2
XFILLER_34_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2965_ _0696_ _1291_ _1280_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__mux2_1
X_2896_ _1255_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__clkbuf_1
X_1916_ po_0.regf_0.rf\[4\]\[15\] po_0.regf_0.rf\[5\]\[15\] po_0.regf_0.rf\[6\]\[15\]
+ po_0.regf_0.rf\[7\]\[15\] _0514_ _0515_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__mux4_1
X_1847_ _0497_ _0447_ _0420_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__a21o_1
X_1778_ po_0.regf_0.rf\[8\]\[1\] po_0.regf_0.rf\[9\]\[1\] po_0.regf_0.rf\[10\]\[1\]
+ po_0.regf_0.rf\[11\]\[1\] _0416_ _0417_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__mux4_1
X_3379_ po_0.alu_0._10_\[0\] _1468_ VGND VGND VPWR VPWR po_0.alu_0._11_\[0\] sky130_fd_sc_hd__ebufn_1
XFILLER_69_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2750_ net93 VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__clkbuf_2
X_1701_ po_0.regf_0.rf\[4\]\[10\] po_0.regf_0.rf\[5\]\[10\] po_0.regf_0.rf\[6\]\[10\]
+ po_0.regf_0.rf\[7\]\[10\] _1442_ _1443_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux4_1
X_2681_ po_0.regf_0.rf\[8\]\[1\] _0717_ _1109_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__mux2_1
X_1632_ _1429_ _1432_ _1433_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__mux2_1
X_1563_ _1361_ uc_0.bc_0._54_\[1\] _1369_ _1370_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__a31o_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _1321_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__clkbuf_1
X_3302_ net164 _0273_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3233_ net164 _0208_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3164_ net106 _0139_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_3095_ net133 _0070_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2115_ _0579_ po_0._1_\[2\] VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__nand2_1
X_2046_ _0659_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__inv_2
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2948_ _1282_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__clkbuf_1
X_2879_ _1246_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2802_ net72 _0565_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__nand2_1
X_3278__182 VGND VGND VPWR VPWR _3278__182/HI net182 sky130_fd_sc_hd__conb_1
X_2733_ uc_0._20_\[9\] net32 _1134_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__mux2_1
X_2664_ _1101_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__clkbuf_1
X_2595_ po_0.regf_0.rf\[11\]\[10\] _0980_ _1059_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__mux2_1
X_1615_ _1390_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__clkbuf_2
X_1546_ net34 VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__clkbuf_2
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3216_ net103 _0191_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3147_ net109 _0122_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3078_ net126 _0057_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_2029_ _0655_ po_0._1_\[12\] VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__nand2_1
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2380_ po_0.regf_0.rf\[1\]\[0\] _0694_ _0938_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__mux2_1
Xinput6 D_R_data[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_3001_ uc_0.bc_0._54_\[1\] VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__inv_2
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2716_ _1129_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2647_ _1092_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2578_ po_0.regf_0.rf\[11\]\[2\] _0963_ _1052_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__mux2_1
X_1529_ po_0._1_\[0\] _1340_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__nand2_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _0526_ _0433_ _0474_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__a21bo_1
X_2501_ _1011_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__buf_2
X_2432_ po_0.regf_0.rf\[15\]\[5\] _0969_ _0959_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__mux2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2363_ _0928_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
X_2294_ po_0.regf_0.rf\[5\]\[11\] _0828_ _0884_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__mux2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3282__178 VGND VGND VPWR VPWR _3282__178/HI net178 sky130_fd_sc_hd__conb_1
XFILLER_52_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_11 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2981_ _0681_ net51 _1300_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__mux2_1
X_1932_ po_0.regf_0.rq_addr\[3\] _0570_ _0568_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__mux2_1
X_1863_ _0508_ _0511_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__and2b_1
Xinput20 I_data[12] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
Xinput31 I_data[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
X_1794_ _0407_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__clkbuf_4
X_2415_ _0696_ _0697_ _0957_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__and3_2
XFILLER_69_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2346_ _0919_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2277_ po_0.regf_0.rf\[5\]\[3\] _0742_ _0877_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__mux2_1
XFILLER_37_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _0633_ po_0._1_\[9\] _0639_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__o21ai_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ net106 _0155_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_2131_ _0707_ _0748_ _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__a21oi_1
X_2062_ _0684_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__buf_2
XFILLER_19_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2964_ uc_0._20_\[9\] _0714_ _0562_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__mux2_1
X_1915_ po_0.regf_0.rf\[0\]\[15\] po_0.regf_0.rf\[1\]\[15\] po_0.regf_0.rf\[2\]\[15\]
+ po_0.regf_0.rf\[3\]\[15\] _0427_ _0428_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__mux4_1
X_2895_ po_0.regf_0.rf\[3\]\[13\] _0848_ _1239_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__mux2_1
X_1846_ po_0.regf_0.rf\[4\]\[7\] po_0.regf_0.rf\[5\]\[7\] po_0.regf_0.rf\[6\]\[7\]
+ po_0.regf_0.rf\[7\]\[7\] _0444_ _0445_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__mux4_1
X_1777_ _0432_ _0433_ _0412_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a21bo_1
X_3378_ net149 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2329_ _0909_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1700_ po_0.regf_0.rf\[0\]\[10\] po_0.regf_0.rf\[1\]\[10\] po_0.regf_0.rf\[2\]\[10\]
+ po_0.regf_0.rf\[3\]\[10\] _1430_ _1431_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__mux4_1
X_2680_ _1110_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1631_ _0006_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__buf_2
X_3301_ net119 _0272_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_1562_ uc_0.bc_0._54_\[3\] _1360_ _1364_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__and3_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _1315_ _1319_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__or2b_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ net120 _0207_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ net110 _0138_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_2114_ _0590_ _0591_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__nor2_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3094_ net156 _0069_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2045_ _0668_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__or2_1
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2947_ po_0.regf_0.rq_addr\[1\] _0565_ _0568_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__mux2_1
X_2878_ po_0.regf_0.rf\[3\]\[5\] _0764_ _1240_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__mux2_1
X_1829_ _0414_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__clkbuf_4
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2801_ _1191_ _1192_ _1193_ _1194_ _1195_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__o311a_1
X_2732_ _1138_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2663_ _0810_ po_0.regf_0.rf\[0\]\[9\] _1097_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__mux2_1
X_2594_ _1063_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_1
X_1614_ _1416_ _1391_ _1393_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__a21o_1
X_1545_ _1356_ VGND VGND VPWR VPWR uc_0.bc_0._54_\[3\] sky130_fd_sc_hd__inv_2
X_3215_ net102 _0190_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3146_ net106 _0121_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3077_ net129 _0056_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2028_ net38 VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 D_R_data[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3000_ _1127_ _1217_ _1300_ _1310_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o211a_1
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2715_ _0714_ net24 _1127_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__mux2_1
X_2646_ _0718_ po_0.regf_0.rf\[0\]\[1\] _1090_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__mux2_1
X_2577_ _1054_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
X_1528_ po_0._1_\[0\] _1340_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__or2_1
XFILLER_59_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3129_ net107 _0104_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2500_ _0699_ _0915_ _0935_ _0874_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__and4_2
X_2431_ _0764_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__clkbuf_2
X_2362_ po_0.regf_0.rf\[9\]\[9\] _0810_ _0924_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__mux2_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2293_ _0889_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_12 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2629_ _1082_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2980_ _1300_ uc_0.bc_0._54_\[0\] net59 _1219_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1931_ po_0.muxf_0.rf_w_data\[7\] VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__clkbuf_4
X_1862_ po_0.regf_0.rf\[8\]\[9\] po_0.regf_0.rf\[9\]\[9\] po_0.regf_0.rf\[10\]\[9\]
+ po_0.regf_0.rf\[11\]\[9\] _0509_ _0510_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__mux4_1
Xinput10 D_R_data[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 I_data[13] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 I_data[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
X_1793_ _0405_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__buf_4
X_2414_ po_0.regf_0.w_addr\[2\] po_0.regf_0.w_addr\[3\] _0872_ VGND VGND VPWR VPWR
+ _0957_ sky130_fd_sc_hd__and3_1
X_3394_ po_0.alu_0._10_\[15\] _1483_ VGND VGND VPWR VPWR po_0.alu_0._11_\[15\] sky130_fd_sc_hd__ebufn_1
X_2345_ po_0.regf_0.rf\[9\]\[1\] _0718_ _0917_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__mux2_1
X_2276_ _0880_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2130_ _0721_ _0722_ _0734_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__o21ai_1
XFILLER_66_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2061_ po_0.muxf_0.s1 po_0.muxf_0.s0 VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__and2b_1
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2963_ _1290_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__clkbuf_1
X_1914_ _0508_ _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__and2b_1
X_2894_ _1254_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1845_ _0457_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__and2b_1
X_1776_ _0410_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__clkbuf_2
X_2328_ po_0.regf_0.rf\[6\]\[10\] _0820_ _0904_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__mux2_1
XFILLER_69_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2259_ net41 _0686_ _1314_ _0866_ _0687_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__o311a_1
XFILLER_25_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1630_ po_0.regf_0.rf\[12\]\[2\] po_0.regf_0.rf\[13\]\[2\] po_0.regf_0.rf\[14\]\[2\]
+ po_0.regf_0.rf\[15\]\[2\] _1430_ _1431_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__mux4_1
X_3300_ net118 _0271_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_1561_ net81 net94 _1345_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__nor3b_2
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _1320_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ net99 _0206_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ net107 _0137_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_2113_ _0733_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
X_3093_ net165 _0068_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2044_ net40 po_0._1_\[14\] VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__nor2_1
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2946_ _1281_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__clkbuf_1
X_2877_ _1245_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_1
X_1828_ po_0.regf_0.rf\[4\]\[5\] po_0.regf_0.rf\[5\]\[5\] po_0.regf_0.rf\[6\]\[5\]
+ po_0.regf_0.rf\[7\]\[5\] _0427_ _0428_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__mux4_1
X_1759_ _0407_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__buf_2
XFILLER_57_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2800_ uc_0._01_ _1154_ _1162_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__and3_1
X_2731_ uc_0._20_\[8\] net31 _1134_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__mux2_1
X_2662_ _1100_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2593_ po_0.regf_0.rf\[11\]\[9\] _0978_ _1059_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__mux2_1
X_1613_ po_0.regf_0.rf\[12\]\[1\] po_0.regf_0.rf\[13\]\[1\] po_0.regf_0.rf\[14\]\[1\]
+ po_0.regf_0.rf\[15\]\[1\] _1386_ _1388_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__mux4_1
X_1544_ net34 _1355_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__or2_1
X_3214_ net101 _0189_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3145_ net107 _0120_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3076_ net133 _0055_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2027_ _0632_ _0649_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__a21oi_2
XFILLER_35_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2929_ _1273_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 D_R_data[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2714_ _1128_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__clkbuf_1
X_2645_ _1091_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2576_ po_0.regf_0.rf\[11\]\[1\] _0961_ _1052_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__mux2_1
X_1527_ net35 VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__clkbuf_2
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3128_ net108 _0103_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3059_ po_0.regf_0._3_\[6\] net86 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlxtp_1
XFILLER_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2430_ _0968_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
X_2361_ _0927_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
X_2292_ po_0.regf_0.rf\[5\]\[10\] _0820_ _0884_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__mux2_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_13 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2628_ po_0.regf_0.rf\[10\]\[9\] _0978_ _1078_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__mux2_1
X_2559_ po_0.regf_0.rf\[12\]\[10\] _0980_ _1039_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__mux2_1
XFILLER_46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1930_ _0569_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
X_1861_ _0407_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__clkbuf_2
Xinput22 I_data[14] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 D_R_data[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput33 clock VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
X_1792_ _0446_ _0447_ _0420_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__a21bo_1
X_3393_ po_0.alu_0._10_\[14\] _1482_ VGND VGND VPWR VPWR po_0.alu_0._11_\[14\] sky130_fd_sc_hd__ebufn_1
X_2413_ _0693_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__clkbuf_2
X_2344_ _0918_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
X_2275_ po_0.regf_0.rf\[5\]\[2\] _0732_ _0877_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__mux2_1
XFILLER_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__clkbuf_2
XFILLER_66_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2962_ _0697_ _1289_ _1280_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__mux2_1
X_1913_ po_0.regf_0.rf\[8\]\[15\] po_0.regf_0.rf\[9\]\[15\] po_0.regf_0.rf\[10\]\[15\]
+ po_0.regf_0.rf\[11\]\[15\] _0509_ _0510_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__mux4_1
X_2893_ po_0.regf_0.rf\[3\]\[12\] _0839_ _1239_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__mux2_1
X_1844_ po_0.regf_0.rf\[0\]\[7\] po_0.regf_0.rf\[1\]\[7\] po_0.regf_0.rf\[2\]\[7\]
+ po_0.regf_0.rf\[3\]\[7\] _0449_ _0450_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__mux4_1
X_1775_ po_0.regf_0.rf\[12\]\[1\] po_0.regf_0.rf\[13\]\[1\] po_0.regf_0.rf\[14\]\[1\]
+ po_0.regf_0.rf\[15\]\[1\] _0406_ _0408_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__mux4_1
X_2327_ _0908_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2258_ po_0.alu_0._11_\[15\] _1317_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__or2b_1
XFILLER_69_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2189_ _0803_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1560_ _1357_ _1354_ _1361_ _1363_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__nor4_4
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ _1315_ _1319_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__or2b_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ net119 _0205_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ net107 _0136_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2112_ po_0.regf_0.rf\[7\]\[2\] _0732_ _0701_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__mux2_1
X_3092_ net156 _0067_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2043_ net40 po_0._1_\[14\] VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__and2_1
XFILLER_62_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2945_ po_0.regf_0.rq_addr\[0\] _0561_ _0568_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__mux2_1
X_2876_ po_0.regf_0.rf\[3\]\[4\] _0754_ _1240_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__mux2_1
X_1827_ po_0.regf_0.rf\[0\]\[5\] po_0.regf_0.rf\[1\]\[5\] po_0.regf_0.rf\[2\]\[5\]
+ po_0.regf_0.rf\[3\]\[5\] _0478_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__mux4_1
X_1758_ _0405_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__clkbuf_4
X_1689_ _0353_ _1409_ _1436_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__a21o_1
X_3359_ net170 _0330_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dfxtp_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2730_ _1137_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__clkbuf_1
X_2661_ _0802_ po_0.regf_0.rf\[0\]\[8\] _1097_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__mux2_1
X_1612_ _1411_ _1414_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__and2b_1
X_2592_ _1062_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
X_1543_ _1346_ _1354_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__nor2_1
X_3213_ net103 _0188_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3144_ net108 _0119_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3075_ net132 _0054_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2026_ _0650_ po_0._1_\[11\] _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2928_ po_0.regf_0.rf\[2\]\[12\] _0839_ _1258_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__mux2_1
XFILLER_10_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2859_ _1235_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput9 D_R_data[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2713_ _0681_ net17 _1127_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__mux2_1
X_2644_ _0694_ po_0.regf_0.rf\[0\]\[0\] _1090_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__mux2_1
X_2575_ _1053_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
X_1526_ _1339_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__clkbuf_1
X_3127_ net108 _0102_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3058_ po_0.regf_0._3_\[5\] net85 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlxtp_1
X_2009_ po_0._1_\[10\] net36 VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__or2b_1
XFILLER_2_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2360_ po_0.regf_0.rf\[9\]\[8\] _0802_ _0924_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__mux2_1
X_2291_ _0888_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_14 _0714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2627_ _1081_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__clkbuf_1
X_2558_ _1043_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
X_2489_ _1005_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
X_1509_ _1326_ _1328_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__or2b_1
XFILLER_28_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1860_ _0405_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__buf_2
Xinput12 D_R_data[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
X_1791_ _0410_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__buf_2
Xinput23 I_data[15] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xinput34 reset VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2412_ _0955_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
X_3392_ po_0.alu_0._10_\[13\] _1481_ VGND VGND VPWR VPWR po_0.alu_0._11_\[13\] sky130_fd_sc_hd__ebufn_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2343_ po_0.regf_0.rf\[9\]\[0\] _0694_ _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__mux2_1
X_2274_ _0879_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1989_ net48 VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__clkbuf_2
XFILLER_57_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2961_ uc_0._20_\[8\] _0681_ _0562_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__mux2_1
X_1912_ _0554_ _0457_ _0003_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2892_ _1253_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1843_ _0493_ _0411_ _0412_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__a21bo_1
X_1774_ _0413_ _0419_ _0421_ _0431_ VGND VGND VPWR VPWR po_0.regf_0._3_\[0\] sky130_fd_sc_hd__o22a_1
X_2326_ po_0.regf_0.rf\[6\]\[9\] _0810_ _0904_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__mux2_1
XFILLER_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2257_ _0668_ _0864_ _0855_ _0706_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__o31ai_1
X_2188_ po_0.regf_0.rf\[7\]\[8\] _0802_ _0778_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__mux2_1
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1318_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ net110 _0135_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2111_ _0731_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__clkbuf_2
X_3091_ net150 _0066_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2042_ _0662_ _0666_ _0667_ VGND VGND VPWR VPWR po_0.alu_0._10_\[13\] sky130_fd_sc_hd__nor3b_1
XFILLER_66_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2944_ _0935_ _1219_ _1280_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__a21o_1
X_2875_ _1244_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__clkbuf_1
X_1826_ _0424_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__buf_2
X_1757_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__clkbuf_2
X_1688_ po_0.regf_0.rf\[12\]\[9\] po_0.regf_0.rf\[13\]\[9\] po_0.regf_0.rf\[14\]\[9\]
+ po_0.regf_0.rf\[15\]\[9\] _1419_ _1420_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__mux4_1
X_3358_ net124 _0329_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ po_0.regf_0.rf\[6\]\[1\] _0718_ _0897_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__mux2_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ net161 _0260_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2660_ _1099_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__clkbuf_1
X_1611_ po_0.regf_0.rf\[0\]\[1\] po_0.regf_0.rf\[1\]\[1\] po_0.regf_0.rf\[2\]\[1\]
+ po_0.regf_0.rf\[3\]\[1\] _1412_ _1413_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__mux4_1
XFILLER_5_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2591_ po_0.regf_0.rf\[11\]\[8\] _0976_ _1059_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__mux2_1
X_1542_ _1347_ _1351_ _1352_ _1353_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__nor4_4
X_3212_ net112 _0187_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3143_ net108 _0118_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3074_ net163 _0053_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2025_ _0637_ _0646_ _0651_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or3_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2927_ _1272_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__clkbuf_1
X_2858_ po_0.regf_0.rf\[4\]\[12\] _0839_ _1220_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__mux2_1
X_2789_ net70 po_0.muxf_0.rf_w_data\[3\] VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__nand2_1
X_1809_ po_0.regf_0.rf\[8\]\[4\] po_0.regf_0.rf\[9\]\[4\] po_0.regf_0.rf\[10\]\[4\]
+ po_0.regf_0.rf\[11\]\[4\] _0423_ _0425_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__mux4_1
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2712_ uc_0._03_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__buf_2
X_2643_ _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__clkbuf_4
X_2574_ po_0.regf_0.rf\[11\]\[0\] _0956_ _1052_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__mux2_1
X_1525_ _1325_ _1327_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__or2b_1
XFILLER_67_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3126_ net137 _0101_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3057_ po_0.regf_0._3_\[4\] net87 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlxtp_1
X_2008_ net36 po_0._1_\[10\] VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__and2b_1
XFILLER_70_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2290_ po_0.regf_0.rf\[5\]\[9\] _0810_ _0884_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__mux2_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_15 _0714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2626_ po_0.regf_0.rf\[10\]\[8\] _0976_ _1078_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__mux2_1
X_2557_ po_0.regf_0.rf\[12\]\[9\] _0978_ _1039_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__mux2_1
X_2488_ po_0.regf_0.rf\[14\]\[10\] _0980_ _1000_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__mux2_1
X_1508_ _1330_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3109_ net165 _0084_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 D_R_data[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1790_ po_0.regf_0.rf\[12\]\[2\] po_0.regf_0.rf\[13\]\[2\] po_0.regf_0.rf\[14\]\[2\]
+ po_0.regf_0.rf\[15\]\[2\] _0444_ _0445_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__mux4_1
Xinput24 I_data[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2411_ po_0.regf_0.rf\[1\]\[15\] _0870_ _0937_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__mux2_1
X_3391_ po_0.alu_0._10_\[12\] _1480_ VGND VGND VPWR VPWR po_0.alu_0._11_\[12\] sky130_fd_sc_hd__ebufn_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2342_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__clkbuf_4
X_2273_ po_0.regf_0.rf\[5\]\[1\] _0718_ _0877_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__mux2_1
XFILLER_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1988_ _0620_ VGND VGND VPWR VPWR po_0.alu_0._10_\[6\] sky130_fd_sc_hd__clkbuf_1
X_2609_ po_0.regf_0.rf\[10\]\[0\] _0956_ _1071_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__mux2_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2960_ _1288_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__clkbuf_1
X_1911_ po_0.regf_0.rf\[12\]\[15\] po_0.regf_0.rf\[13\]\[15\] po_0.regf_0.rf\[14\]\[15\]
+ po_0.regf_0.rf\[15\]\[15\] _0449_ _0450_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__mux4_1
X_2891_ po_0.regf_0.rf\[3\]\[11\] _0827_ _1247_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__mux2_1
XFILLER_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1842_ po_0.regf_0.rf\[12\]\[7\] po_0.regf_0.rf\[13\]\[7\] po_0.regf_0.rf\[14\]\[7\]
+ po_0.regf_0.rf\[15\]\[7\] _0406_ _0408_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__mux4_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1773_ _0426_ _0429_ _0430_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__mux2_1
X_2325_ _0907_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2256_ _0673_ _0674_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__or2_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2187_ _0801_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__clkbuf_2
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2110_ _0728_ _0713_ _0730_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__a21o_2
X_3090_ net143 _0065_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2041_ po_0._1_\[12\] _0660_ _0655_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__or3b_2
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2943_ _1278_ _1279_ _1371_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__or3_4
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2874_ po_0.regf_0.rf\[3\]\[3\] _0741_ _1240_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__mux2_1
X_1825_ _0422_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__clkbuf_4
X_1756_ _0002_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__buf_2
X_1687_ _0352_ VGND VGND VPWR VPWR po_0.regf_0._5_\[8\] sky130_fd_sc_hd__clkbuf_1
X_3357_ net100 _0328_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dfxtp_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _0898_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3288_ net150 _0259_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2239_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__clkbuf_2
XFILLER_53_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1610_ _1381_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__buf_2
X_2590_ _1061_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1541_ net46 net84 net48 VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__or3_1
X_3211_ net115 _0186_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3142_ net137 _0117_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3073_ net159 _0052_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2024_ _0635_ _0640_ _0641_ _0638_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__o211a_1
X_2926_ po_0.regf_0.rf\[2\]\[11\] _0827_ _1266_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__mux2_1
X_2857_ _1234_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1808_ _0454_ _0456_ _0459_ _0462_ VGND VGND VPWR VPWR po_0.regf_0._3_\[3\] sky130_fd_sc_hd__o22a_1
X_2788_ net70 po_0.muxf_0.rf_w_data\[3\] VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__or2_1
X_1739_ _1433_ _0397_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__and2b_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2711_ _1126_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__clkbuf_1
X_2642_ _0699_ _0695_ _0935_ _1030_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__or4bb_4
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2573_ _1051_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__clkbuf_4
X_1524_ _1338_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3125_ net140 _0100_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3056_ po_0.regf_0._3_\[3\] net87 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlxtp_1
X_2007_ _0634_ _0636_ VGND VGND VPWR VPWR po_0.alu_0._10_\[9\] sky130_fd_sc_hd__xor2_1
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2909_ po_0.regf_0.rf\[2\]\[3\] _0741_ _1259_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__mux2_1
XFILLER_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_16 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_27 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2625_ _1080_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
X_2556_ _1042_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
X_2487_ _1004_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
X_1507_ _1326_ _1328_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__or2b_1
X_3108_ net159 _0083_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3039_ po_0.regf_0._5_\[2\] net90 VGND VGND VPWR VPWR po_0._1_\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_62_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 D_R_data[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput25 I_data[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2410_ _0954_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
X_3390_ po_0.alu_0._10_\[11\] _1479_ VGND VGND VPWR VPWR po_0.alu_0._11_\[11\] sky130_fd_sc_hd__ebufn_2
X_2341_ _0875_ _0915_ _0873_ _0874_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__and4b_4
X_2272_ _0878_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1987_ _0617_ _0619_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__and2b_1
X_2608_ _1070_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__clkbuf_4
X_2539_ _1033_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1910_ _0548_ _0550_ _0461_ _0553_ VGND VGND VPWR VPWR po_0.regf_0._3_\[14\] sky130_fd_sc_hd__o22a_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2890_ _1252_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1841_ _0430_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__and2b_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1772_ _0414_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__clkbuf_2
X_2324_ po_0.regf_0.rf\[6\]\[8\] _0802_ _0904_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__mux2_1
X_2255_ _0673_ _0674_ _0855_ _0668_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__o22a_1
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2186_ net15 _0790_ _0800_ _0713_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__a22o_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2040_ _0663_ _0664_ _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__a21oi_1
XFILLER_74_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2942_ _1361_ _1365_ uc_0.bc_0._54_\[2\] VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__and3_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2873_ _1243_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1824_ _0415_ _0476_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__and2b_1
X_1755_ _0409_ _0411_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__a21bo_1
X_1686_ _0348_ _0349_ _0350_ _0351_ _1392_ _1418_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__mux4_1
X_3356_ net167 _0327_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dfxtp_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3287_ net143 _0258_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ po_0.regf_0.rf\[6\]\[0\] _0694_ _0897_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__mux2_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2238_ _0846_ _0847_ _0712_ _0790_ net5 VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__a32o_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2169_ _0621_ _1317_ _1313_ _0784_ _0687_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__o311a_1
XFILLER_70_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1540_ net35 net42 net44 net43 VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__or4_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3210_ net112 _0185_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3141_ net140 _0116_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3072_ net161 _0051_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2023_ net37 VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__inv_2
XFILLER_35_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2925_ _1271_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__clkbuf_1
X_2856_ po_0.regf_0.rf\[4\]\[11\] _0827_ _1228_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__mux2_1
X_1807_ _0460_ _0447_ _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__a21o_1
X_2787_ _1159_ _1163_ _1149_ net70 VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__a31o_1
X_1738_ po_0.regf_0.rf\[8\]\[15\] po_0.regf_0.rf\[9\]\[15\] po_0.regf_0.rf\[10\]\[15\]
+ po_0.regf_0.rf\[11\]\[15\] _1427_ _1428_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__mux4_1
X_1669_ _1395_ _1466_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__and2b_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ net152 _0310_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2710_ po_0.regf_0.rf\[8\]\[15\] _0869_ _1108_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__mux2_1
XFILLER_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2641_ _1088_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__clkbuf_1
X_2572_ _0696_ _0697_ _1050_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__and3_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1523_ _1325_ _1327_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__or2b_1
X_3124_ net141 _0099_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3055_ po_0.regf_0._3_\[2\] net87 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlxtp_1
X_2006_ _0630_ _0632_ _0635_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__a21bo_1
XFILLER_23_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2908_ _1262_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__clkbuf_1
X_2839_ po_0.regf_0.rf\[4\]\[3\] _0741_ _1221_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__mux2_1
XFILLER_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_17 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2624_ po_0.regf_0.rf\[10\]\[7\] _0974_ _1078_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__mux2_1
X_2555_ po_0.regf_0.rf\[12\]\[8\] _0976_ _1039_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__mux2_1
X_2486_ po_0.regf_0.rf\[14\]\[9\] _0978_ _1000_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__mux2_1
X_1506_ _1329_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__clkbuf_1
X_3107_ net151 _0082_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3038_ po_0.regf_0._5_\[1\] net91 VGND VGND VPWR VPWR po_0._1_\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 I_data[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput15 D_R_data[8] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
X_2340_ po_0.regf_0.w_addr\[3\] VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2271_ po_0.regf_0.rf\[5\]\[0\] _0694_ _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__mux2_1
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1986_ _0616_ _0618_ _0615_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__nand3_1
XFILLER_60_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2607_ _0875_ _0915_ _0872_ _0895_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__and4b_2
X_2538_ po_0.regf_0.rf\[12\]\[0\] _0956_ _1032_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__mux2_1
X_2469_ po_0.regf_0.rf\[14\]\[1\] _0961_ _0993_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__mux2_1
XFILLER_28_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout170 net173 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1840_ po_0.regf_0.rf\[8\]\[7\] po_0.regf_0.rf\[9\]\[7\] po_0.regf_0.rf\[10\]\[7\]
+ po_0.regf_0.rf\[11\]\[7\] _0423_ _0425_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__mux4_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1771_ po_0.regf_0.rf\[4\]\[0\] po_0.regf_0.rf\[5\]\[0\] po_0.regf_0.rf\[6\]\[0\]
+ po_0.regf_0.rf\[7\]\[0\] _0427_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__mux4_1
XFILLER_6_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2323_ _0906_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2254_ net7 _0790_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__nand2_1
X_2185_ _0796_ _0706_ _0798_ _0799_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__a31o_1
XFILLER_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1969_ _0592_ _0603_ _0601_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__and3_1
XFILLER_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2941_ _1354_ _1363_ _1369_ uc_0.bc_0._54_\[0\] VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__o211a_1
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2872_ po_0.regf_0.rf\[3\]\[2\] _0731_ _1240_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__mux2_1
X_1823_ po_0.regf_0.rf\[8\]\[5\] po_0.regf_0.rf\[9\]\[5\] po_0.regf_0.rf\[10\]\[5\]
+ po_0.regf_0.rf\[11\]\[5\] _0416_ _0417_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__mux4_1
X_1754_ _0003_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__clkbuf_2
X_1685_ po_0.regf_0.rf\[4\]\[8\] po_0.regf_0.rf\[5\]\[8\] po_0.regf_0.rf\[6\]\[8\]
+ po_0.regf_0.rf\[7\]\[8\] _1385_ _1387_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__mux4_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ net148 _0326_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfxtp_1
X_2306_ _0896_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__clkbuf_4
X_3286_ net169 _0257_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ _0659_ _0708_ _1313_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__or3_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2168_ po_0.alu_0._11_\[7\] _1316_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__or2b_1
XFILLER_53_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2099_ _0688_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__buf_2
XFILLER_65_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3140_ net141 _0115_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3071_ net148 _0050_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2022_ _0648_ _0640_ _0639_ _0646_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__nor4_1
XFILLER_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2924_ po_0.regf_0.rf\[2\]\[10\] _0819_ _1266_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__mux2_1
X_2855_ _1233_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__clkbuf_1
X_1806_ _0003_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__buf_2
X_2786_ _1159_ _1153_ _1147_ _1162_ _1182_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__o311a_1
X_1737_ _0391_ _0393_ _1440_ _0396_ VGND VGND VPWR VPWR po_0.regf_0._5_\[14\] sky130_fd_sc_hd__o22a_1
X_1668_ po_0.regf_0.rf\[0\]\[6\] po_0.regf_0.rf\[1\]\[6\] po_0.regf_0.rf\[2\]\[6\]
+ po_0.regf_0.rf\[3\]\[6\] _1396_ _1397_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__mux4_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ net145 _0309_ VGND VGND VPWR VPWR po_0.regf_0.w_wr sky130_fd_sc_hd__dfxtp_1
X_1599_ _1390_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__buf_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3269_ net166 _0240_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfxtp_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2640_ po_0.regf_0.rf\[10\]\[15\] _0990_ _1070_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__mux2_1
XFILLER_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2571_ po_0.regf_0.w_addr\[2\] po_0.regf_0.w_addr\[3\] _0872_ VGND VGND VPWR VPWR
+ _1050_ sky130_fd_sc_hd__and3b_1
X_1522_ _1337_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3123_ net141 _0098_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3054_ po_0.regf_0._3_\[1\] net87 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlxtp_1
X_2005_ po_0._1_\[8\] net83 VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__or2b_1
XFILLER_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2907_ po_0.regf_0.rf\[2\]\[2\] _0731_ _1259_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__mux2_1
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2838_ _1224_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__clkbuf_1
X_2769_ net92 po_0.muxf_0.rf_w_data\[1\] VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__or2_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_18 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_29 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2623_ _1079_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
X_2554_ _1041_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
X_1505_ _1326_ _1328_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__or2b_1
X_2485_ _1003_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3106_ net143 _0081_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3037_ po_0.regf_0._5_\[0\] net90 VGND VGND VPWR VPWR po_0._1_\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput16 D_R_data[9] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
Xinput27 I_data[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2270_ _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1985_ _0613_ _0614_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__nor2_1
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2606_ _1069_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_1
X_2537_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__buf_2
X_2468_ _0994_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
X_2399_ po_0.regf_0.rf\[1\]\[9\] _0810_ _0945_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__mux2_1
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout171 net172 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout160 net174 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1770_ _0424_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__buf_4
XFILLER_6_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2322_ po_0.regf_0.rf\[6\]\[7\] _0788_ _0904_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__mux2_1
X_2253_ _0861_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2184_ _0708_ po_0.alu_0._11_\[8\] _0709_ net83 VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__a22o_1
XFILLER_18_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1968_ _0599_ _0600_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__nor2_2
X_1899_ po_0.regf_0.rf\[0\]\[13\] po_0.regf_0.rf\[1\]\[13\] po_0.regf_0.rf\[2\]\[13\]
+ po_0.regf_0.rf\[3\]\[13\] _0478_ _0479_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__mux4_1
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2940_ _1367_ _1368_ _1218_ po_0.regf_0.rp_rd _0563_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__a221o_1
X_2871_ _1242_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__clkbuf_1
X_1822_ _0473_ _0433_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__a21bo_1
X_1753_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__clkbuf_2
X_1684_ po_0.regf_0.rf\[12\]\[8\] po_0.regf_0.rf\[13\]\[8\] po_0.regf_0.rf\[14\]\[8\]
+ po_0.regf_0.rf\[15\]\[8\] _1385_ _1387_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__mux4_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ net169 _0325_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfxtp_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _0695_ _0873_ _0895_ _0875_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__and4b_4
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ net171 _0256_ VGND VGND VPWR VPWR uc_0._00_ sky130_fd_sc_hd__dfxtp_1
X_2236_ _0843_ _0844_ _0845_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__o21ai_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ _0607_ _0614_ _0770_ _0781_ _0780_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__o311a_1
XFILLER_53_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2098_ _0719_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3070_ net143 _0049_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2021_ _0628_ _0629_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__and2_1
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2923_ _1270_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__clkbuf_1
X_2854_ po_0.regf_0.rf\[4\]\[10\] _0819_ _1228_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__mux2_1
X_1805_ po_0.regf_0.rf\[4\]\[3\] po_0.regf_0.rf\[5\]\[3\] po_0.regf_0.rf\[6\]\[3\]
+ po_0.regf_0.rf\[7\]\[3\] _0444_ _0445_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__mux4_1
X_2785_ _1176_ _1178_ _1154_ _1181_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__a31o_1
X_1736_ _0394_ _0395_ _1445_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux2_1
X_1667_ _1464_ _1391_ _1393_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__a21o_1
X_1598_ po_0.regf_0.rf\[4\]\[0\] po_0.regf_0.rf\[5\]\[0\] po_0.regf_0.rf\[6\]\[0\]
+ po_0.regf_0.rf\[7\]\[0\] _1400_ _1401_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__mux4_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3337_ net170 _0308_ VGND VGND VPWR VPWR po_0.regf_0.rp_rd sky130_fd_sc_hd__dfxtp_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3268_ net152 _0015_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__dfxtp_2
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3199_ net99 _0174_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_2219_ net37 po_0._1_\[11\] _0823_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2570_ _1049_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
X_1521_ _1325_ _1327_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__or2b_1
X_3122_ net140 _0097_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3053_ po_0.regf_0._3_\[0\] po_0.regf_0.rp_rd VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlxtp_1
XFILLER_82_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2004_ _0633_ po_0._1_\[9\] VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__xnor2_2
XFILLER_48_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2906_ _1261_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__clkbuf_1
X_2837_ po_0.regf_0.rf\[4\]\[2\] _0731_ _1221_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__mux2_1
X_2768_ _1163_ _1149_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__nor2_1
X_1719_ po_0.regf_0.rf\[4\]\[12\] po_0.regf_0.rf\[5\]\[12\] po_0.regf_0.rf\[6\]\[12\]
+ po_0.regf_0.rf\[7\]\[12\] _1400_ _1401_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__mux4_1
X_2699_ _1120_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__clkbuf_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2622_ po_0.regf_0.rf\[10\]\[6\] _0971_ _1078_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__mux2_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2553_ po_0.regf_0.rf\[12\]\[7\] _0974_ _1039_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__mux2_1
X_1504_ _1327_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2484_ po_0.regf_0.rf\[14\]\[8\] _0976_ _1000_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__mux2_1
X_3105_ net164 _0080_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3036_ net119 _0047_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput17 I_data[0] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput28 I_data[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1984_ _0613_ _0614_ _0615_ _0616_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__a2bb2oi_2
X_2605_ po_0.regf_0.rf\[11\]\[15\] _0990_ _1051_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__mux2_1
X_2536_ _0699_ _0915_ _0873_ _1030_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__and4_2
X_2467_ po_0.regf_0.rf\[14\]\[0\] _0956_ _0993_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__mux2_1
X_2398_ _0948_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3019_ net118 _0030_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout161 net163 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
Xfanout150 net151 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout172 net173 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3370_ net173 uc_0.bc_0._54_\[3\] VGND VGND VPWR VPWR uc_0.bc_0._55_\[3\] sky130_fd_sc_hd__dfxtp_1
X_2321_ _0905_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
X_2252_ po_0.regf_0.rf\[7\]\[14\] _0860_ _0700_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2183_ _0768_ _0797_ _0794_ _0648_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__a211o_1
XFILLER_65_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1967_ _0599_ _0600_ _0601_ _0592_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__a2bb2oi_2
X_1898_ _0508_ _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__and2b_1
X_2519_ po_0.regf_0.rf\[13\]\[8\] _0976_ _1019_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__mux2_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2870_ po_0.regf_0.rf\[3\]\[1\] _0717_ _1240_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__mux2_1
X_1821_ _0003_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__clkbuf_2
X_1752_ _0002_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__buf_2
XFILLER_7_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1683_ po_0.regf_0.rf\[0\]\[8\] po_0.regf_0.rf\[1\]\[8\] po_0.regf_0.rf\[2\]\[8\]
+ po_0.regf_0.rf\[3\]\[8\] _1385_ _1387_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__mux4_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ net170 _0324_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfxtp_1
X_2304_ po_0.regf_0.w_addr\[0\] po_0.regf_0.w_addr\[1\] VGND VGND VPWR VPWR _0895_
+ sky130_fd_sc_hd__and2b_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ net172 net176 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfxtp_1
X_2235_ _1318_ po_0.alu_0._11_\[13\] _0709_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__a21oi_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2166_ _0780_ _0772_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2097_ po_0.regf_0.rf\[7\]\[1\] _0718_ _0701_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__mux2_1
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2999_ net77 _1216_ _1217_ _1300_ _1310_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__o311a_1
XFILLER_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2020_ _0646_ _0647_ VGND VGND VPWR VPWR po_0.alu_0._10_\[11\] sky130_fd_sc_hd__xnor2_1
X_2922_ po_0.regf_0.rf\[2\]\[9\] _0809_ _1266_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__mux2_1
XFILLER_50_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2853_ _1232_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__clkbuf_1
X_1804_ _0457_ _0458_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__and2b_1
X_2784_ _1146_ _1179_ _1180_ _1148_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__a31o_1
X_1735_ po_0.regf_0.rf\[4\]\[14\] po_0.regf_0.rf\[5\]\[14\] po_0.regf_0.rf\[6\]\[14\]
+ po_0.regf_0.rf\[7\]\[14\] _1442_ _1443_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__mux4_1
X_1666_ po_0.regf_0.rf\[12\]\[6\] po_0.regf_0.rf\[13\]\[6\] po_0.regf_0.rf\[14\]\[6\]
+ po_0.regf_0.rf\[15\]\[6\] _1386_ _1388_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__mux4_1
X_1597_ _1387_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__clkbuf_4
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ net162 _0307_ VGND VGND VPWR VPWR po_0.regf_0.rq_rd sky130_fd_sc_hd__dfxtp_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ net152 _0014_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__dfxtp_1
X_2218_ _0829_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
X_3198_ net99 _0173_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2149_ _0766_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1520_ _1336_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__clkbuf_1
X_3121_ net147 _0096_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3052_ po_0.regf_0._5_\[15\] net88 VGND VGND VPWR VPWR po_0._1_\[15\] sky130_fd_sc_hd__dlxtp_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2003_ net50 VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__buf_2
XFILLER_23_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2905_ po_0.regf_0.rf\[2\]\[1\] _0717_ _1259_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__mux2_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2836_ _1223_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__clkbuf_1
X_2767_ _1163_ _1149_ _1146_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__and3_1
X_1718_ _1411_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__and2b_1
X_2698_ po_0.regf_0.rf\[8\]\[9\] _0809_ _1116_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__mux2_1
X_1649_ po_0.regf_0.rf\[12\]\[4\] po_0.regf_0.rf\[13\]\[4\] po_0.regf_0.rf\[14\]\[4\]
+ po_0.regf_0.rf\[15\]\[4\] _1386_ _1388_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__mux4_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ net144 _0290_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2621_ _1070_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__buf_2
X_2552_ _1040_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1503_ _1318_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__clkbuf_1
X_2483_ _1002_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
X_3104_ net100 _0079_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_3035_ net118 _0046_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2819_ _1203_ _1206_ _1209_ _1210_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__o211a_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 I_data[10] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 I_data[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1983_ _0607_ _0608_ _0605_ _0602_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__o22ai_2
X_2604_ _1068_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__clkbuf_1
X_2535_ _0696_ _0697_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__nor2_1
X_2466_ _0992_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__buf_2
X_2397_ po_0.regf_0.rf\[1\]\[8\] _0802_ _0945_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__mux2_1
XFILLER_83_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3018_ net124 _0029_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout140 net142 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout162 net163 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
Xfanout151 net154 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout173 net174 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2320_ po_0.regf_0.rf\[6\]\[6\] _0777_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__mux2_1
X_2251_ _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2182_ _0603_ _0609_ _0618_ _0781_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__and4_1
XFILLER_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1966_ po_0._1_\[3\] _0589_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__or2b_1
X_1897_ po_0.regf_0.rf\[8\]\[13\] po_0.regf_0.rf\[9\]\[13\] po_0.regf_0.rf\[10\]\[13\]
+ po_0.regf_0.rf\[11\]\[13\] _0509_ _0510_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__mux4_1
X_2518_ _1021_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2449_ _0981_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1820_ po_0.regf_0.rf\[12\]\[5\] po_0.regf_0.rf\[13\]\[5\] po_0.regf_0.rf\[14\]\[5\]
+ po_0.regf_0.rf\[15\]\[5\] _0471_ _0472_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux4_1
X_1751_ po_0.regf_0.rf\[12\]\[0\] po_0.regf_0.rf\[13\]\[0\] po_0.regf_0.rf\[14\]\[0\]
+ po_0.regf_0.rf\[15\]\[0\] _0406_ _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__mux4_1
XFILLER_7_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1682_ po_0.regf_0.rf\[8\]\[8\] po_0.regf_0.rf\[9\]\[8\] po_0.regf_0.rf\[10\]\[8\]
+ po_0.regf_0.rf\[11\]\[8\] _1385_ _1387_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__mux4_1
X_3352_ net162 _0323_ VGND VGND VPWR VPWR po_0.muxf_0.s1 sky130_fd_sc_hd__dfxtp_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _0894_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ net126 net177 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfxtp_2
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _0656_ _0842_ _0836_ _0725_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__a31o_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ _0622_ _0623_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__nor2_1
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2096_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__clkbuf_2
XFILLER_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2998_ _1215_ _1361_ _1365_ _1367_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__or4_1
X_1949_ _0573_ net42 VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__and2b_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2921_ _1269_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__clkbuf_1
X_2852_ po_0.regf_0.rf\[4\]\[9\] _0809_ _1228_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__mux2_1
X_1803_ po_0.regf_0.rf\[0\]\[3\] po_0.regf_0.rf\[1\]\[3\] po_0.regf_0.rf\[2\]\[3\]
+ po_0.regf_0.rf\[3\]\[3\] _0449_ _0450_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__mux4_1
X_2783_ net68 net61 _1159_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__a21o_1
X_1734_ po_0.regf_0.rf\[0\]\[14\] po_0.regf_0.rf\[1\]\[14\] po_0.regf_0.rf\[2\]\[14\]
+ po_0.regf_0.rf\[3\]\[14\] _1430_ _1431_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__mux4_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1665_ _1433_ _1462_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__and2b_1
X_1596_ _1385_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__clkbuf_4
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ net162 _0306_ VGND VGND VPWR VPWR po_0.alu_0.s0 sky130_fd_sc_hd__dfxtp_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ net154 _0013_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__dfxtp_1
X_2217_ po_0.regf_0.rf\[7\]\[11\] _0828_ _0778_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__mux2_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ net103 _0172_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2148_ po_0.regf_0.rf\[7\]\[5\] _0765_ _0701_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__mux2_1
X_2079_ po_0.regf_0.rf\[7\]\[0\] _0694_ _0701_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__mux2_1
XFILLER_14_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3120_ net118 _0095_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_3051_ po_0.regf_0._5_\[14\] net88 VGND VGND VPWR VPWR po_0._1_\[14\] sky130_fd_sc_hd__dlxtp_1
X_2002_ _0630_ _0632_ VGND VGND VPWR VPWR po_0.alu_0._10_\[8\] sky130_fd_sc_hd__xor2_1
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2904_ _1260_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__clkbuf_1
X_2835_ po_0.regf_0.rf\[4\]\[1\] _0717_ _1221_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__mux2_1
X_2766_ uc_0._01_ uc_0._00_ _1146_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__o21ba_1
X_1717_ po_0.regf_0.rf\[0\]\[12\] po_0.regf_0.rf\[1\]\[12\] po_0.regf_0.rf\[2\]\[12\]
+ po_0.regf_0.rf\[3\]\[12\] _1396_ _1397_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__mux4_1
X_2697_ _1119_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__clkbuf_1
X_1648_ _1433_ _1447_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__and2b_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ po_0.regf_0.rf\[8\]\[0\] po_0.regf_0.rf\[9\]\[0\] po_0.regf_0.rf\[10\]\[0\]
+ po_0.regf_0.rf\[11\]\[0\] _1380_ _1382_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__mux4_1
X_3318_ net165 _0289_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3249_ net171 _0224_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2620_ _1077_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2551_ po_0.regf_0.rf\[12\]\[6\] _0971_ _1039_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__mux2_1
X_1502_ _1325_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2482_ po_0.regf_0.rf\[14\]\[7\] _0974_ _1000_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__mux2_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3103_ net100 _0078_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_3034_ net125 _0045_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2818_ net74 po_0.muxf_0.rf_w_data\[7\] VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__or2_1
X_2749_ uc_0._01_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__nor2_1
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 I_data[11] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1982_ po_0._1_\[5\] _0606_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__or2b_1
XFILLER_60_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2603_ po_0.regf_0.rf\[11\]\[14\] _0988_ _1051_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__mux2_1
X_2534_ _1029_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2465_ _0699_ _0915_ _0935_ _0895_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__and4_2
X_2396_ _0947_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3017_ net124 _0028_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout130 net131 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout152 net153 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout141 net142 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout163 net174 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
Xfanout174 net175 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2250_ net6 _0685_ _0858_ _0712_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__a22o_2
XFILLER_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2181_ _0795_ _0648_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__nand2_2
XFILLER_65_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1965_ net84 po_0._1_\[4\] VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__nor2_1
X_1896_ _0540_ _0457_ _0474_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__a21bo_1
X_2517_ po_0.regf_0.rf\[13\]\[7\] _0974_ _1019_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__mux2_1
X_2448_ po_0.regf_0.rf\[15\]\[10\] _0980_ _0972_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__mux2_1
X_2379_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__clkbuf_4
XFILLER_56_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1750_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__buf_2
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1681_ _0341_ _0343_ _0345_ _0347_ VGND VGND VPWR VPWR po_0.regf_0._5_\[7\] sky130_fd_sc_hd__o22a_1
X_3351_ net162 _0322_ VGND VGND VPWR VPWR po_0.muxf_0.s0 sky130_fd_sc_hd__dfxtp_1
X_2302_ po_0.regf_0.rf\[5\]\[15\] _0870_ _0876_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__mux2_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ net154 net178 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfxtp_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _0656_ _0836_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2164_ _1347_ po_0._1_\[6\] VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__nand2_1
X_2095_ _0711_ _0713_ _0716_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__a21o_2
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2997_ _1309_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__clkbuf_1
X_1948_ _1340_ po_0._1_\[0\] VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__or2b_1
X_1879_ po_0.regf_0.rf\[12\]\[11\] po_0.regf_0.rf\[13\]\[11\] po_0.regf_0.rf\[14\]\[11\]
+ po_0.regf_0.rf\[15\]\[11\] _0471_ _0472_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__mux4_1
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2920_ po_0.regf_0.rf\[2\]\[8\] _0801_ _1266_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__mux2_1
X_2851_ _1231_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1802_ _0410_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__buf_2
X_2782_ _1159_ _1163_ net93 VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__nand3_1
X_1733_ _1378_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__and2b_1
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1664_ po_0.regf_0.rf\[8\]\[6\] po_0.regf_0.rf\[9\]\[6\] po_0.regf_0.rf\[10\]\[6\]
+ po_0.regf_0.rf\[11\]\[6\] _1427_ _1428_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__mux4_1
X_1595_ _1395_ _1398_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__and2b_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ net161 _0305_ VGND VGND VPWR VPWR po_0.alu_0.s1 sky130_fd_sc_hd__dfxtp_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3265_ net152 _0012_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__dfxtp_1
X_2216_ _0827_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__clkbuf_2
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ net112 _0171_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2147_ _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2078_ _0700_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__clkbuf_4
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3050_ po_0.regf_0._5_\[13\] net88 VGND VGND VPWR VPWR po_0._1_\[13\] sky130_fd_sc_hd__dlxtp_1
X_2001_ _0631_ po_0._1_\[7\] _0625_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__o21ai_4
XFILLER_48_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2903_ po_0.regf_0.rf\[2\]\[0\] _0693_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__mux2_1
XFILLER_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2834_ _1222_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__clkbuf_1
X_2765_ net92 VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1716_ _0377_ _1418_ _1436_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__a21o_1
X_2696_ po_0.regf_0.rf\[8\]\[8\] _0801_ _1116_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__mux2_1
X_1647_ po_0.regf_0.rf\[8\]\[4\] po_0.regf_0.rf\[9\]\[4\] po_0.regf_0.rf\[10\]\[4\]
+ po_0.regf_0.rf\[11\]\[4\] _1380_ _1382_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__mux4_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ net121 _0288_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_1578_ _1381_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__clkbuf_4
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ net104 _0223_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3179_ net109 _0154_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2550_ _1031_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__buf_2
X_1501_ _1314_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2481_ _1001_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
X_3102_ net100 _0077_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3033_ net124 _0044_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2817_ net74 _0570_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__nand2_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2748_ uc_0._00_ uc_0._02_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__or2_2
X_2679_ po_0.regf_0.rf\[8\]\[0\] _0693_ _1109_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__mux2_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1981_ _1347_ po_0._1_\[6\] VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__nor2_2
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2602_ _1067_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2533_ po_0.regf_0.rf\[13\]\[15\] _0990_ _1011_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__mux2_1
X_2464_ _0991_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
X_2395_ po_0.regf_0.rf\[1\]\[7\] _0788_ _0945_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__mux2_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3016_ net121 _0027_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout120 net123 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout131 net136 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
Xfanout153 net154 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
Xfanout142 net146 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout164 net165 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout175 net33 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_2
XFILLER_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2180_ _0791_ _0747_ _0794_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__o21bai_1
XFILLER_65_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1964_ net84 po_0._1_\[4\] VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__and2_1
X_1895_ po_0.regf_0.rf\[12\]\[13\] po_0.regf_0.rf\[13\]\[13\] po_0.regf_0.rf\[14\]\[13\]
+ po_0.regf_0.rf\[15\]\[13\] _0471_ _0472_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__mux4_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2516_ _1020_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
X_2447_ _0819_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__clkbuf_2
X_2378_ _0935_ _0874_ _0936_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__and3_4
XFILLER_68_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1680_ _0346_ _1403_ _1404_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__a21o_1
X_3350_ net138 _0321_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[3\] sky130_fd_sc_hd__dfxtp_1
X_2301_ _0893_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ net125 net179 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfxtp_2
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ _0659_ po_0._1_\[13\] VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2163_ _0779_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2094_ _0714_ _0683_ _0715_ net8 VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__a22o_1
XFILLER_21_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2996_ _0570_ net58 _1303_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__mux2_1
X_1947_ _0574_ _0578_ _0580_ _0581_ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__o2111ai_2
X_1878_ _0519_ _0521_ _0523_ _0525_ VGND VGND VPWR VPWR po_0.regf_0._3_\[10\] sky130_fd_sc_hd__o22a_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2850_ po_0.regf_0.rf\[4\]\[8\] _0801_ _1228_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__mux2_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1801_ _0455_ _0447_ _0412_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a21bo_1
X_2781_ _1163_ _0714_ _1177_ _1175_ _1169_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__a221o_1
X_1732_ po_0.regf_0.rf\[8\]\[14\] po_0.regf_0.rf\[9\]\[14\] po_0.regf_0.rf\[10\]\[14\]
+ po_0.regf_0.rf\[11\]\[14\] _1380_ _1382_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__mux4_1
XFILLER_7_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1663_ _1456_ _1458_ _1440_ _1461_ VGND VGND VPWR VPWR po_0.regf_0._5_\[5\] sky130_fd_sc_hd__o22a_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ po_0.regf_0.rf\[0\]\[0\] po_0.regf_0.rf\[1\]\[0\] po_0.regf_0.rf\[2\]\[0\]
+ po_0.regf_0.rf\[3\]\[0\] _1396_ _1397_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__mux4_1
X_3333_ net120 _0304_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ net164 _0239_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_1
X_2215_ net3 _0790_ _0822_ _0826_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__o2bb2ai_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ net114 _0170_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2146_ _0761_ _0712_ _0762_ _0763_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__a31o_2
XFILLER_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2077_ _0695_ _0698_ _0699_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__and3b_4
XFILLER_53_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2979_ _1299_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__clkbuf_4
XFILLER_69_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3284__176 VGND VGND VPWR VPWR _3284__176/HI net176 sky130_fd_sc_hd__conb_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2000_ _0621_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__inv_2
XFILLER_48_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2902_ _1258_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__clkbuf_4
XFILLER_50_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2833_ po_0.regf_0.rf\[4\]\[0\] _0693_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__mux2_1
X_2764_ _1150_ _1155_ _1162_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__o21a_1
X_1715_ po_0.regf_0.rf\[12\]\[12\] po_0.regf_0.rf\[13\]\[12\] po_0.regf_0.rf\[14\]\[12\]
+ po_0.regf_0.rf\[15\]\[12\] _1406_ _1407_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__mux4_1
X_2695_ _1118_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__clkbuf_1
X_1646_ _1437_ _1439_ _1440_ _1446_ VGND VGND VPWR VPWR po_0.regf_0._5_\[3\] sky130_fd_sc_hd__o22a_1
X_1577_ _0005_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ net99 _0287_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ net101 _0222_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ net111 _0153_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2129_ _0574_ _0573_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__nand2_1
XFILLER_81_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2480_ po_0.regf_0.rf\[14\]\[6\] _0971_ _1000_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__mux2_1
X_1500_ _1324_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__clkbuf_1
X_3101_ net100 _0076_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3032_ net121 _0043_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2816_ _1206_ _1208_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__nor2_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2747_ uc_0._02_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2678_ _1108_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__buf_2
X_1629_ _0005_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__clkbuf_4
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3281__179 VGND VGND VPWR VPWR _3281__179/HI net179 sky130_fd_sc_hd__conb_1
XFILLER_27_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1980_ net47 po_0._1_\[6\] VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__and2_1
XFILLER_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2601_ po_0.regf_0.rf\[11\]\[13\] _0986_ _1051_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__mux2_1
XFILLER_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2532_ _1028_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
X_2463_ po_0.regf_0.rf\[15\]\[15\] _0990_ _0958_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__mux2_1
X_2394_ _0946_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3015_ net133 _0026_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout121 net123 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
Xfanout110 net111 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout154 net155 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout132 net135 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout143 net146 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
Xfanout165 net168 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1963_ _0598_ VGND VGND VPWR VPWR po_0.alu_0._10_\[3\] sky130_fd_sc_hd__clkbuf_1
X_1894_ _0534_ _0536_ _0461_ _0539_ VGND VGND VPWR VPWR po_0.regf_0._3_\[12\] sky130_fd_sc_hd__o22a_1
X_2515_ po_0.regf_0.rf\[13\]\[6\] _0971_ _1019_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__mux2_1
X_2446_ _0979_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
X_2377_ po_0.regf_0.w_addr\[2\] po_0.regf_0.w_addr\[3\] VGND VGND VPWR VPWR _0936_
+ sky130_fd_sc_hd__nor2_1
XFILLER_56_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3280_ net149 net180 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfxtp_1
X_2300_ po_0.regf_0.rf\[5\]\[14\] _0860_ _0876_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__mux2_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _0841_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2162_ po_0.regf_0.rf\[7\]\[6\] _0777_ _0778_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__mux2_1
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2093_ _0684_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2995_ _1308_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1946_ _0573_ _0582_ _0572_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__o21ai_1
X_1877_ _0524_ _0447_ _0420_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__a21o_1
X_2429_ po_0.regf_0.rf\[15\]\[4\] _0967_ _0959_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__mux2_1
XFILLER_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1800_ po_0.regf_0.rf\[12\]\[3\] po_0.regf_0.rf\[13\]\[3\] po_0.regf_0.rf\[14\]\[3\]
+ po_0.regf_0.rf\[15\]\[3\] _0444_ _0445_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__mux4_1
X_2780_ _1159_ _0729_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__or2_1
X_1731_ _0390_ _1395_ _1392_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__a21o_1
X_1662_ _1459_ _1460_ _1445_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__mux2_1
X_3332_ net99 _0303_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_1593_ _1381_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__clkbuf_4
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ net107 _0238_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfxtp_2
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ net112 _0169_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_2214_ _1318_ po_0.alu_0._11_\[11\] _0824_ _0825_ _0720_ VGND VGND VPWR VPWR _0826_
+ sky130_fd_sc_hd__a221oi_4
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ _0565_ _0682_ _0715_ net12 VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__a22o_1
XFILLER_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2076_ po_0.regf_0.w_addr\[2\] VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2978_ _1357_ _1363_ _1366_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__or3_1
X_1929_ po_0.regf_0.rq_addr\[2\] _0567_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__mux2_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2901_ _0935_ _0895_ _0936_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__and3_4
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2832_ _1220_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__clkbuf_4
X_2763_ _1161_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__clkbuf_2
X_1714_ _1433_ _0375_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__and2b_1
X_2694_ po_0.regf_0.rf\[8\]\[7\] _0787_ _1116_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__mux2_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1645_ _1441_ _1444_ _1445_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__mux2_1
X_1576_ _1379_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__clkbuf_4
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ net120 _0286_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ net101 _0221_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3177_ net111 _0152_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_2128_ _0723_ _0745_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__a21oi_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2059_ po_0.muxf_0.s0 po_0.muxf_0.s1 VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__and2b_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput80 net80 VGND VGND VPWR VPWR leds[1] sky130_fd_sc_hd__buf_2
X_3100_ net103 _0075_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_3031_ net134 _0042_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2815_ _1196_ _1201_ _1205_ _1207_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__a31o_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2746_ _1145_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__clkbuf_1
X_2677_ _0875_ _0695_ _0872_ _1030_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__and4b_4
X_1628_ _0004_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__buf_4
X_1559_ _1355_ _1366_ _1357_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__a21oi_2
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ net119 _0204_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2600_ _1066_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__clkbuf_1
X_2531_ po_0.regf_0.rf\[13\]\[14\] _0988_ _1011_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__mux2_1
XFILLER_5_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2462_ _0869_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__clkbuf_2
XFILLER_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2393_ po_0.regf_0.rf\[1\]\[6\] _0777_ _0945_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__mux2_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3014_ net126 _0025_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3280__180 VGND VGND VPWR VPWR _3280__180/HI net180 sky130_fd_sc_hd__conb_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2729_ _0570_ net30 _1134_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__mux2_1
Xfanout100 net102 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout122 net123 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout111 net117 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout155 net175 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout133 net134 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout144 net145 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout166 net167 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1962_ _0592_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__and2_1
X_1893_ _0537_ _0538_ _0482_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__mux2_1
X_2514_ _1011_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__buf_2
X_2445_ po_0.regf_0.rf\[15\]\[9\] _0978_ _0972_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__mux2_1
X_2376_ _0872_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2230_ po_0.regf_0.rf\[7\]\[12\] _0840_ _0700_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__mux2_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2161_ _0700_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__buf_2
X_2092_ po_0.muxf_0.rf_w_data\[1\] VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__clkbuf_4
XFILLER_65_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2994_ _0567_ net57 _1303_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__mux2_1
X_1945_ _0574_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__inv_2
X_1876_ po_0.regf_0.rf\[4\]\[10\] po_0.regf_0.rf\[5\]\[10\] po_0.regf_0.rf\[6\]\[10\]
+ po_0.regf_0.rf\[7\]\[10\] _0444_ _0445_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__mux4_1
XFILLER_0_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2428_ _0754_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__clkbuf_2
X_2359_ _0926_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1730_ po_0.regf_0.rf\[12\]\[14\] po_0.regf_0.rf\[13\]\[14\] po_0.regf_0.rf\[14\]\[14\]
+ po_0.regf_0.rf\[15\]\[14\] _1419_ _1420_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux4_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1661_ po_0.regf_0.rf\[4\]\[5\] po_0.regf_0.rf\[5\]\[5\] po_0.regf_0.rf\[6\]\[5\]
+ po_0.regf_0.rf\[7\]\[5\] _1442_ _1443_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__mux4_1
X_3331_ net120 _0302_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_1592_ _1379_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__clkbuf_4
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ net172 _0237_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfxtp_2
X_2213_ _0823_ _0814_ _0646_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__o21ai_2
X_3193_ net112 _0168_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2144_ _0606_ _0708_ _1313_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__or3_1
XFILLER_19_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2075_ _0696_ _0697_ po_0.regf_0.w_wr VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__and3_1
XFILLER_53_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2977_ uc_0.bc_0._54_\[0\] _1365_ _1369_ _1219_ net60 VGND VGND VPWR VPWR _0324_
+ sky130_fd_sc_hd__a32o_1
X_1928_ _0562_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__clkbuf_2
X_1859_ _0414_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2900_ _1257_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2831_ _0695_ _0873_ _1030_ _0875_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__and4b_4
X_2762_ net66 net65 _1158_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__nor4b_1
X_1713_ po_0.regf_0.rf\[8\]\[12\] po_0.regf_0.rf\[9\]\[12\] po_0.regf_0.rf\[10\]\[12\]
+ po_0.regf_0.rf\[11\]\[12\] _1427_ _1428_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__mux4_1
X_2693_ _1117_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__clkbuf_1
X_1644_ _0006_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__clkbuf_4
X_1575_ _0004_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ net122 _0285_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ net104 _0220_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3176_ net110 _0151_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2127_ _0596_ po_0._1_\[2\] _0579_ _0590_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__a31o_1
XFILLER_66_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2058_ po_0.muxf_0.rf_w_data\[0\] VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__clkbuf_4
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput70 net70 VGND VGND VPWR VPWR I_addr[3] sky130_fd_sc_hd__buf_2
Xoutput81 net95 VGND VGND VPWR VPWR leds[2] sky130_fd_sc_hd__buf_2
X_3030_ net126 _0041_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2814_ uc_0._00_ uc_0._02_ _1161_ uc_0._01_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__or4bb_1
X_2745_ net82 net23 _1133_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__mux2_1
X_2676_ _1107_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__clkbuf_1
X_1627_ po_0.regf_0.rf\[8\]\[2\] po_0.regf_0.rf\[9\]\[2\] po_0.regf_0.rf\[10\]\[2\]
+ po_0.regf_0.rf\[11\]\[2\] _1427_ _1428_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__mux4_1
X_1558_ _1357_ _1366_ VGND VGND VPWR VPWR uc_0.bc_0._54_\[2\] sky130_fd_sc_hd__nor2_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ _1317_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__buf_2
X_3228_ net121 _0203_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3159_ net108 _0134_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2530_ _1027_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
X_2461_ _0989_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
X_2392_ _0937_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__buf_2
X_3013_ net129 _0024_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2728_ _1136_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__clkbuf_1
X_2659_ _0788_ po_0.regf_0.rf\[0\]\[7\] _1097_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__mux2_1
Xfanout101 net102 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
Xfanout112 net116 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout123 net136 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xfanout134 net135 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout156 net160 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
Xfanout145 net146 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
Xfanout167 net168 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1961_ _0593_ _0594_ _0595_ _0596_ _0580_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__o2111ai_1
X_1892_ po_0.regf_0.rf\[4\]\[12\] po_0.regf_0.rf\[5\]\[12\] po_0.regf_0.rf\[6\]\[12\]
+ po_0.regf_0.rf\[7\]\[12\] _0514_ _0515_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__mux4_1
X_2513_ _1018_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
X_2444_ _0809_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__clkbuf_2
X_2375_ _0934_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2091_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2993_ _1307_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__clkbuf_1
X_1944_ _0579_ po_0._1_\[2\] VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__or2b_1
X_1875_ _0415_ _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__and2b_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2427_ _0966_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2358_ po_0.regf_0.rf\[9\]\[7\] _0788_ _0924_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__mux2_1
XFILLER_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2289_ _0887_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1660_ po_0.regf_0.rf\[0\]\[5\] po_0.regf_0.rf\[1\]\[5\] po_0.regf_0.rf\[2\]\[5\]
+ po_0.regf_0.rf\[3\]\[5\] _1430_ _1431_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__mux4_1
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1591_ _1390_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__buf_2
X_3330_ net122 _0301_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ net147 _0236_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dfxtp_2
X_2212_ _0823_ _0646_ _0814_ _0706_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__o31a_1
X_3192_ net114 _0167_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _1318_ po_0.alu_0._11_\[5\] _0720_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__a211o_1
XFILLER_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2074_ po_0.regf_0.w_addr\[0\] VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2976_ po_0.muxf_0.s1 _1278_ _1298_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__o21a_1
X_1927_ po_0.muxf_0.rf_w_data\[6\] VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__buf_2
X_1858_ _0506_ _0433_ _0474_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__a21bo_1
X_1789_ _0407_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2830_ _1215_ uc_0._00_ _1219_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__o21a_1
X_2761_ net70 _1159_ net92 net93 VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__nand4_1
X_1712_ _0368_ _0370_ _0372_ _0374_ VGND VGND VPWR VPWR po_0.regf_0._5_\[11\] sky130_fd_sc_hd__o22a_1
X_2692_ po_0.regf_0.rf\[8\]\[6\] _0776_ _1116_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__mux2_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1643_ po_0.regf_0.rf\[4\]\[3\] po_0.regf_0.rf\[5\]\[3\] po_0.regf_0.rf\[6\]\[3\]
+ po_0.regf_0.rf\[7\]\[3\] _1442_ _1443_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__mux4_1
XANTENNA_1 _0681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1574_ _0006_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__clkbuf_2
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ net128 _0284_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ net113 _0219_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ net108 _0150_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2126_ _0721_ _0722_ _0595_ _0596_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__o211a_1
X_2057_ _0677_ _0680_ VGND VGND VPWR VPWR po_0.alu_0._10_\[15\] sky130_fd_sc_hd__nor2_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2959_ uc_0._20_\[11\] po_0.regf_0.rp_addr\[3\] _1372_ VGND VGND VPWR VPWR _1288_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput60 net60 VGND VGND VPWR VPWR D_wr sky130_fd_sc_hd__buf_2
Xoutput71 net71 VGND VGND VPWR VPWR I_addr[4] sky130_fd_sc_hd__buf_2
Xoutput82 net94 VGND VGND VPWR VPWR leds[3] sky130_fd_sc_hd__buf_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2813_ _1196_ _1201_ _1205_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__a21oi_1
X_2744_ _1144_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__clkbuf_1
X_2675_ _0870_ po_0.regf_0.rf\[0\]\[15\] _1089_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__mux2_1
X_1626_ _1381_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__buf_2
X_1557_ net95 net94 _1345_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__or3b_2
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ _1316_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__clkbuf_2
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ net130 _0202_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_3158_ net137 _0133_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2109_ _0729_ _0682_ _0715_ net9 VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__a22o_1
X_3089_ net164 _0064_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2460_ po_0.regf_0.rf\[15\]\[14\] _0988_ _0958_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__mux2_1
X_2391_ _0944_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
X_3012_ net133 _0023_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2727_ _0567_ net29 _1134_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__mux2_1
X_2658_ _1098_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__clkbuf_1
Xfanout102 net104 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout113 net116 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
X_2589_ po_0.regf_0.rf\[11\]\[7\] _0974_ _1059_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__mux2_1
X_1609_ _1379_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__clkbuf_4
Xfanout124 net125 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout135 net136 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout146 net155 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout168 net174 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout157 net160 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1960_ _0589_ po_0._1_\[3\] VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__or2_1
X_1891_ po_0.regf_0.rf\[0\]\[12\] po_0.regf_0.rf\[1\]\[12\] po_0.regf_0.rf\[2\]\[12\]
+ po_0.regf_0.rf\[3\]\[12\] _0478_ _0479_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__mux4_1
X_2512_ po_0.regf_0.rf\[13\]\[5\] _0969_ _1012_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__mux2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2443_ _0977_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_2374_ po_0.regf_0.rf\[9\]\[15\] _0870_ _0916_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__mux2_1
XFILLER_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2090_ _0687_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__clkbuf_2
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2992_ _0565_ net56 _1303_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__mux2_1
X_1943_ po_0._1_\[2\] _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__nand2b_2
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1874_ po_0.regf_0.rf\[0\]\[10\] po_0.regf_0.rf\[1\]\[10\] po_0.regf_0.rf\[2\]\[10\]
+ po_0.regf_0.rf\[3\]\[10\] _0416_ _0417_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__mux4_1
X_2426_ po_0.regf_0.rf\[15\]\[3\] _0965_ _0959_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__mux2_1
X_2357_ _0925_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
X_2288_ po_0.regf_0.rf\[5\]\[8\] _0802_ _0884_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__mux2_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1590_ _1389_ _1391_ _1393_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__a21o_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ net137 _0235_ VGND VGND VPWR VPWR uc_0._20_\[11\] sky130_fd_sc_hd__dfxtp_1
X_2211_ net36 po_0._1_\[10\] VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__and2_1
X_3191_ net114 _0166_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2142_ _0758_ _0689_ _0759_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__and3_1
XFILLER_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2073_ po_0.regf_0.w_addr\[1\] VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2975_ _1279_ _0563_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__nor2_1
X_1926_ _0566_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
X_1857_ po_0.regf_0.rf\[12\]\[9\] po_0.regf_0.rf\[13\]\[9\] po_0.regf_0.rf\[14\]\[9\]
+ po_0.regf_0.rf\[15\]\[9\] _0471_ _0472_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__mux4_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1788_ _0405_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__buf_4
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2409_ po_0.regf_0.rf\[1\]\[14\] _0860_ _0937_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__mux2_1
X_3389_ po_0.alu_0._10_\[10\] _1478_ VGND VGND VPWR VPWR po_0.alu_0._11_\[10\] sky130_fd_sc_hd__ebufn_1
XFILLER_57_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2760_ net69 VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__clkbuf_2
X_1711_ _1418_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__and2b_1
X_2691_ _1108_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__buf_2
XFILLER_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1642_ _0005_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_2 _0717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1573_ _1377_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ net130 _0283_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ net115 _0218_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3174_ net137 _0149_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2125_ _1317_ po_0.alu_0._11_\[4\] _0688_ net84 VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__a22o_1
X_2056_ _0673_ _0674_ _0675_ _0679_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__a2bb2oi_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2958_ _1287_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__clkbuf_1
X_1909_ _0551_ _0552_ _0410_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__mux2_1
X_2889_ po_0.regf_0.rf\[3\]\[10\] _0819_ _1247_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__mux2_1
XFILLER_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput50 net50 VGND VGND VPWR VPWR D_W_data[9] sky130_fd_sc_hd__clkbuf_4
Xoutput61 net93 VGND VGND VPWR VPWR I_addr[0] sky130_fd_sc_hd__buf_2
Xoutput72 net72 VGND VGND VPWR VPWR I_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2812_ _1203_ _1204_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__or2_1
X_2743_ net95 net22 _1133_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__mux2_1
X_2674_ _1106_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__clkbuf_1
X_1625_ _1379_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__clkbuf_4
X_1556_ net34 _1365_ VGND VGND VPWR VPWR uc_0.bc_0._54_\[1\] sky130_fd_sc_hd__nor2_2
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ po_0.alu_0.s1 VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__dlymetal6s2s_1
X_3226_ net126 _0201_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3157_ net147 _0132_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2108_ po_0.muxf_0.rf_w_data\[2\] VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__clkbuf_4
XFILLER_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3088_ net138 _0011_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__dfxtp_2
X_2039_ _0656_ _0657_ _0660_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__a21o_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2390_ po_0.regf_0.rf\[1\]\[5\] _0765_ _0938_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__mux2_1
X_3011_ net132 _0022_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2726_ _1135_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__clkbuf_1
X_2657_ _0777_ po_0.regf_0.rf\[0\]\[6\] _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__mux2_1
X_1608_ _1390_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__clkbuf_2
Xfanout103 net104 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
X_2588_ _1060_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
Xfanout125 net127 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
X_1539_ _1348_ _1349_ _1350_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__nand3_1
Xfanout114 net116 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout136 net175 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout147 net149 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
Xfanout158 net159 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout169 net170 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
X_3209_ net112 _0184_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1890_ _0508_ _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__and2b_1
X_2511_ _1017_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2442_ po_0.regf_0.rf\[15\]\[8\] _0976_ _0972_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__mux2_1
X_2373_ _0933_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2709_ _1125_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2991_ _1306_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1942_ net43 VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__clkbuf_2
X_1873_ _0520_ _0411_ _0412_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__a21bo_1
X_2425_ _0741_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__clkbuf_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2356_ po_0.regf_0.rf\[9\]\[6\] _0777_ _0924_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__mux2_1
X_2287_ _0886_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _0650_ _0720_ _0683_ _0715_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__a211o_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ net156 _0165_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2141_ _0599_ _0757_ _0609_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__o21ai_1
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2072_ po_0.regf_0.w_addr\[3\] VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2974_ po_0.muxf_0.s0 _1279_ _1297_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__o21a_1
X_1925_ po_0.regf_0.rq_addr\[1\] _0565_ _0563_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__mux2_1
X_1856_ _0505_ VGND VGND VPWR VPWR po_0.regf_0._3_\[8\] sky130_fd_sc_hd__clkbuf_1
X_1787_ _0415_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__and2b_1
X_2408_ _0953_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
X_3388_ po_0.alu_0._10_\[9\] _1477_ VGND VGND VPWR VPWR po_0.alu_0._11_\[9\] sky130_fd_sc_hd__ebufn_1
X_2339_ _0914_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1710_ po_0.regf_0.rf\[8\]\[11\] po_0.regf_0.rf\[9\]\[11\] po_0.regf_0.rf\[10\]\[11\]
+ po_0.regf_0.rf\[11\]\[11\] _1396_ _1397_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__mux4_1
X_2690_ _1115_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_3 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1641_ _0004_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__buf_4
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3311_ net128 _0282_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_1572_ uc_0._20_\[11\] po_0.regf_0.rp_addr\[3\] _1373_ VGND VGND VPWR VPWR _1377_
+ sky130_fd_sc_hd__mux2_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ net113 _0217_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ net147 _0148_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2124_ _0743_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2055_ _0668_ _0669_ _0678_ _0666_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__o22ai_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2957_ uc_0._20_\[10\] po_0.regf_0.rp_addr\[2\] _1372_ VGND VGND VPWR VPWR _1287_
+ sky130_fd_sc_hd__mux2_1
X_1908_ po_0.regf_0.rf\[4\]\[14\] po_0.regf_0.rf\[5\]\[14\] po_0.regf_0.rf\[6\]\[14\]
+ po_0.regf_0.rf\[7\]\[14\] _0514_ _0515_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__mux4_1
X_2888_ _1251_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__clkbuf_1
X_1839_ _0485_ _0487_ _0421_ _0490_ VGND VGND VPWR VPWR po_0.regf_0._3_\[6\] sky130_fd_sc_hd__o22a_1
XFILLER_9_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput51 net51 VGND VGND VPWR VPWR D_addr[0] sky130_fd_sc_hd__buf_2
Xoutput40 net40 VGND VGND VPWR VPWR D_W_data[14] sky130_fd_sc_hd__buf_2
Xoutput73 net73 VGND VGND VPWR VPWR I_addr[6] sky130_fd_sc_hd__clkbuf_4
Xoutput62 net62 VGND VGND VPWR VPWR I_addr[10] sky130_fd_sc_hd__buf_2
XFILLER_0_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2811_ net73 po_0.muxf_0.rf_w_data\[6\] VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__nor2_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2742_ _1143_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__clkbuf_1
X_2673_ _0860_ po_0.regf_0.rf\[0\]\[14\] _1089_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__mux2_1
X_1624_ _1425_ _1391_ _0007_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__a21o_1
X_1555_ _1364_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__clkbuf_2
X_3225_ net128 _0200_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1486_ _1314_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__clkbuf_2
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3156_ net141 _0131_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3087_ net109 _0010_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__dfxtp_1
X_2107_ _1318_ po_0.alu_0._11_\[2\] _0720_ _0579_ _0727_ VGND VGND VPWR VPWR _0728_
+ sky130_fd_sc_hd__a221o_1
XFILLER_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2038_ _0653_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__inv_2
XFILLER_50_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3010_ net163 _0021_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2725_ _0565_ net28 _1134_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__mux2_1
X_2656_ _1089_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__buf_2
X_1607_ _1408_ _1409_ _0007_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__a21o_1
Xfanout104 net105 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlymetal6s2s_1
X_2587_ po_0.regf_0.rf\[11\]\[6\] _0971_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__mux2_1
Xfanout126 net127 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
X_1538_ net50 net83 net37 net36 VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__nor4_1
Xfanout115 net116 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
Xfanout137 net139 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout159 net160 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
Xfanout148 net149 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
X_3208_ net114 _0183_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3139_ net141 _0114_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2510_ po_0.regf_0.rf\[13\]\[4\] _0967_ _1012_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__mux2_1
X_2441_ _0801_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2372_ po_0.regf_0.rf\[9\]\[14\] _0860_ _0916_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__mux2_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2708_ po_0.regf_0.rf\[8\]\[14\] _0859_ _1108_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__mux2_1
X_2639_ _1087_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2990_ _0561_ net55 _1303_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__mux2_1
X_1941_ _0573_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__inv_2
X_1872_ po_0.regf_0.rf\[12\]\[10\] po_0.regf_0.rf\[13\]\[10\] po_0.regf_0.rf\[14\]\[10\]
+ po_0.regf_0.rf\[15\]\[10\] _0406_ _0408_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__mux4_1
X_2424_ _0964_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
X_2355_ _0916_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__clkbuf_4
X_2286_ po_0.regf_0.rf\[5\]\[7\] _0788_ _0884_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__mux2_1
XFILLER_56_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _0599_ _0609_ _0757_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__or3_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2071_ _0693_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__clkbuf_2
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2973_ uc_0.bc_0._54_\[1\] _1369_ _1370_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__a21oi_1
X_1924_ po_0.muxf_0.rf_w_data\[5\] VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__buf_2
X_1855_ _0501_ _0504_ _0420_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__mux2_1
X_1786_ po_0.regf_0.rf\[0\]\[2\] po_0.regf_0.rf\[1\]\[2\] po_0.regf_0.rf\[2\]\[2\]
+ po_0.regf_0.rf\[3\]\[2\] _0416_ _0417_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__mux4_1
X_2407_ po_0.regf_0.rf\[1\]\[13\] _0849_ _0937_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__mux2_1
X_3387_ po_0.alu_0._10_\[8\] _1476_ VGND VGND VPWR VPWR po_0.alu_0._11_\[8\] sky130_fd_sc_hd__ebufn_1
XFILLER_69_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2338_ po_0.regf_0.rf\[6\]\[15\] _0870_ _0896_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__mux2_1
X_2269_ _0695_ _0873_ _0874_ _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__and4b_4
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1640_ po_0.regf_0.rf\[0\]\[3\] po_0.regf_0.rf\[1\]\[3\] po_0.regf_0.rf\[2\]\[3\]
+ po_0.regf_0.rf\[3\]\[3\] _1427_ _1428_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__mux4_1
XANTENNA_4 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1571_ _1376_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3310_ net128 _0281_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ net113 _0216_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3172_ net141 _0147_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2123_ po_0.regf_0.rf\[7\]\[3\] _0742_ _0701_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__mux2_1
XFILLER_81_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2054_ _0671_ po_0._1_\[13\] _0667_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__o21ai_1
XFILLER_66_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2956_ _1286_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__clkbuf_1
X_1907_ po_0.regf_0.rf\[0\]\[14\] po_0.regf_0.rf\[1\]\[14\] po_0.regf_0.rf\[2\]\[14\]
+ po_0.regf_0.rf\[3\]\[14\] _0427_ _0428_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__mux4_1
X_2887_ po_0.regf_0.rf\[3\]\[9\] _0809_ _1247_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__mux2_1
X_1838_ _0488_ _0489_ _0482_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__mux2_1
X_1769_ _0422_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__buf_4
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput52 net52 VGND VGND VPWR VPWR D_addr[1] sky130_fd_sc_hd__buf_2
Xoutput41 net41 VGND VGND VPWR VPWR D_W_data[15] sky130_fd_sc_hd__buf_2
Xoutput63 net63 VGND VGND VPWR VPWR I_addr[11] sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 VGND VGND VPWR VPWR I_addr[7] sky130_fd_sc_hd__buf_2
XFILLER_63_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2810_ net73 po_0.muxf_0.rf_w_data\[6\] VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__and2_1
XFILLER_31_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2741_ net80 net21 _1133_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__mux2_1
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2672_ _1105_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1623_ po_0.regf_0.rf\[4\]\[2\] po_0.regf_0.rf\[5\]\[2\] po_0.regf_0.rf\[6\]\[2\]
+ po_0.regf_0.rf\[7\]\[2\] _1386_ _1388_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__mux4_1
X_1554_ _1354_ _1363_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__nor2_1
X_1485_ _1313_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__clkbuf_2
X_3224_ net134 _0199_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
.ends

