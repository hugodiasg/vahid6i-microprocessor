module vahid6i (D_rd,
    D_wr,
    I_rd,
    clock,
    led_clock,
    reset,
    D_R_data,
    D_W_data,
    D_addr,
    I_addr,
    I_data,
    leds);
 output D_rd;
 output D_wr;
 output I_rd;
 input clock;
 output led_clock;
 input reset;
 input [7:0] D_R_data;
 output [7:0] D_W_data;
 output [7:0] D_addr;
 output [7:0] I_addr;
 input [7:0] I_data;
 output [3:0] leds;

 wire net110;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \po_0._1_[0] ;
 wire \po_0._1_[1] ;
 wire \po_0._1_[2] ;
 wire \po_0._1_[3] ;
 wire \po_0._1_[4] ;
 wire \po_0._1_[5] ;
 wire \po_0._1_[6] ;
 wire \po_0._1_[7] ;
 wire \po_0.alu_0._10_[0] ;
 wire \po_0.alu_0._10_[1] ;
 wire \po_0.alu_0._10_[2] ;
 wire \po_0.alu_0._10_[3] ;
 wire \po_0.alu_0._10_[4] ;
 wire \po_0.alu_0._10_[5] ;
 wire \po_0.alu_0._10_[6] ;
 wire \po_0.alu_0._10_[7] ;
 wire \po_0.alu_0._11_[0] ;
 wire \po_0.alu_0._11_[1] ;
 wire \po_0.alu_0._11_[2] ;
 wire \po_0.alu_0._11_[3] ;
 wire \po_0.alu_0._11_[4] ;
 wire \po_0.alu_0._11_[5] ;
 wire \po_0.alu_0._11_[6] ;
 wire \po_0.alu_0._11_[7] ;
 wire \po_0.alu_0.s0 ;
 wire \po_0.alu_0.s1 ;
 wire \po_0.muxf_0.rf_w_data[0] ;
 wire \po_0.muxf_0.rf_w_data[1] ;
 wire \po_0.muxf_0.rf_w_data[2] ;
 wire \po_0.muxf_0.rf_w_data[3] ;
 wire \po_0.muxf_0.rf_w_data[4] ;
 wire \po_0.muxf_0.rf_w_data[5] ;
 wire \po_0.muxf_0.rf_w_data[6] ;
 wire \po_0.muxf_0.rf_w_data[7] ;
 wire \po_0.muxf_0.s0 ;
 wire \po_0.muxf_0.s1 ;
 wire \po_0.regf_0._3_[0] ;
 wire \po_0.regf_0._3_[1] ;
 wire \po_0.regf_0._3_[2] ;
 wire \po_0.regf_0._3_[3] ;
 wire \po_0.regf_0._3_[4] ;
 wire \po_0.regf_0._3_[5] ;
 wire \po_0.regf_0._3_[6] ;
 wire \po_0.regf_0._3_[7] ;
 wire \po_0.regf_0._5_[0] ;
 wire \po_0.regf_0._5_[1] ;
 wire \po_0.regf_0._5_[2] ;
 wire \po_0.regf_0._5_[3] ;
 wire \po_0.regf_0._5_[4] ;
 wire \po_0.regf_0._5_[5] ;
 wire \po_0.regf_0._5_[6] ;
 wire \po_0.regf_0._5_[7] ;
 wire \po_0.regf_0.rf[0][0] ;
 wire \po_0.regf_0.rf[0][1] ;
 wire \po_0.regf_0.rf[0][2] ;
 wire \po_0.regf_0.rf[0][3] ;
 wire \po_0.regf_0.rf[0][4] ;
 wire \po_0.regf_0.rf[0][5] ;
 wire \po_0.regf_0.rf[0][6] ;
 wire \po_0.regf_0.rf[0][7] ;
 wire \po_0.regf_0.rf[10][0] ;
 wire \po_0.regf_0.rf[10][1] ;
 wire \po_0.regf_0.rf[10][2] ;
 wire \po_0.regf_0.rf[10][3] ;
 wire \po_0.regf_0.rf[10][4] ;
 wire \po_0.regf_0.rf[10][5] ;
 wire \po_0.regf_0.rf[10][6] ;
 wire \po_0.regf_0.rf[10][7] ;
 wire \po_0.regf_0.rf[11][0] ;
 wire \po_0.regf_0.rf[11][1] ;
 wire \po_0.regf_0.rf[11][2] ;
 wire \po_0.regf_0.rf[11][3] ;
 wire \po_0.regf_0.rf[11][4] ;
 wire \po_0.regf_0.rf[11][5] ;
 wire \po_0.regf_0.rf[11][6] ;
 wire \po_0.regf_0.rf[11][7] ;
 wire \po_0.regf_0.rf[12][0] ;
 wire \po_0.regf_0.rf[12][1] ;
 wire \po_0.regf_0.rf[12][2] ;
 wire \po_0.regf_0.rf[12][3] ;
 wire \po_0.regf_0.rf[12][4] ;
 wire \po_0.regf_0.rf[12][5] ;
 wire \po_0.regf_0.rf[12][6] ;
 wire \po_0.regf_0.rf[12][7] ;
 wire \po_0.regf_0.rf[13][0] ;
 wire \po_0.regf_0.rf[13][1] ;
 wire \po_0.regf_0.rf[13][2] ;
 wire \po_0.regf_0.rf[13][3] ;
 wire \po_0.regf_0.rf[13][4] ;
 wire \po_0.regf_0.rf[13][5] ;
 wire \po_0.regf_0.rf[13][6] ;
 wire \po_0.regf_0.rf[13][7] ;
 wire \po_0.regf_0.rf[14][0] ;
 wire \po_0.regf_0.rf[14][1] ;
 wire \po_0.regf_0.rf[14][2] ;
 wire \po_0.regf_0.rf[14][3] ;
 wire \po_0.regf_0.rf[14][4] ;
 wire \po_0.regf_0.rf[14][5] ;
 wire \po_0.regf_0.rf[14][6] ;
 wire \po_0.regf_0.rf[14][7] ;
 wire \po_0.regf_0.rf[15][0] ;
 wire \po_0.regf_0.rf[15][1] ;
 wire \po_0.regf_0.rf[15][2] ;
 wire \po_0.regf_0.rf[15][3] ;
 wire \po_0.regf_0.rf[15][4] ;
 wire \po_0.regf_0.rf[15][5] ;
 wire \po_0.regf_0.rf[15][6] ;
 wire \po_0.regf_0.rf[15][7] ;
 wire \po_0.regf_0.rf[1][0] ;
 wire \po_0.regf_0.rf[1][1] ;
 wire \po_0.regf_0.rf[1][2] ;
 wire \po_0.regf_0.rf[1][3] ;
 wire \po_0.regf_0.rf[1][4] ;
 wire \po_0.regf_0.rf[1][5] ;
 wire \po_0.regf_0.rf[1][6] ;
 wire \po_0.regf_0.rf[1][7] ;
 wire \po_0.regf_0.rf[2][0] ;
 wire \po_0.regf_0.rf[2][1] ;
 wire \po_0.regf_0.rf[2][2] ;
 wire \po_0.regf_0.rf[2][3] ;
 wire \po_0.regf_0.rf[2][4] ;
 wire \po_0.regf_0.rf[2][5] ;
 wire \po_0.regf_0.rf[2][6] ;
 wire \po_0.regf_0.rf[2][7] ;
 wire \po_0.regf_0.rf[3][0] ;
 wire \po_0.regf_0.rf[3][1] ;
 wire \po_0.regf_0.rf[3][2] ;
 wire \po_0.regf_0.rf[3][3] ;
 wire \po_0.regf_0.rf[3][4] ;
 wire \po_0.regf_0.rf[3][5] ;
 wire \po_0.regf_0.rf[3][6] ;
 wire \po_0.regf_0.rf[3][7] ;
 wire \po_0.regf_0.rf[4][0] ;
 wire \po_0.regf_0.rf[4][1] ;
 wire \po_0.regf_0.rf[4][2] ;
 wire \po_0.regf_0.rf[4][3] ;
 wire \po_0.regf_0.rf[4][4] ;
 wire \po_0.regf_0.rf[4][5] ;
 wire \po_0.regf_0.rf[4][6] ;
 wire \po_0.regf_0.rf[4][7] ;
 wire \po_0.regf_0.rf[5][0] ;
 wire \po_0.regf_0.rf[5][1] ;
 wire \po_0.regf_0.rf[5][2] ;
 wire \po_0.regf_0.rf[5][3] ;
 wire \po_0.regf_0.rf[5][4] ;
 wire \po_0.regf_0.rf[5][5] ;
 wire \po_0.regf_0.rf[5][6] ;
 wire \po_0.regf_0.rf[5][7] ;
 wire \po_0.regf_0.rf[6][0] ;
 wire \po_0.regf_0.rf[6][1] ;
 wire \po_0.regf_0.rf[6][2] ;
 wire \po_0.regf_0.rf[6][3] ;
 wire \po_0.regf_0.rf[6][4] ;
 wire \po_0.regf_0.rf[6][5] ;
 wire \po_0.regf_0.rf[6][6] ;
 wire \po_0.regf_0.rf[6][7] ;
 wire \po_0.regf_0.rf[7][0] ;
 wire \po_0.regf_0.rf[7][1] ;
 wire \po_0.regf_0.rf[7][2] ;
 wire \po_0.regf_0.rf[7][3] ;
 wire \po_0.regf_0.rf[7][4] ;
 wire \po_0.regf_0.rf[7][5] ;
 wire \po_0.regf_0.rf[7][6] ;
 wire \po_0.regf_0.rf[7][7] ;
 wire \po_0.regf_0.rf[8][0] ;
 wire \po_0.regf_0.rf[8][1] ;
 wire \po_0.regf_0.rf[8][2] ;
 wire \po_0.regf_0.rf[8][3] ;
 wire \po_0.regf_0.rf[8][4] ;
 wire \po_0.regf_0.rf[8][5] ;
 wire \po_0.regf_0.rf[8][6] ;
 wire \po_0.regf_0.rf[8][7] ;
 wire \po_0.regf_0.rf[9][0] ;
 wire \po_0.regf_0.rf[9][1] ;
 wire \po_0.regf_0.rf[9][2] ;
 wire \po_0.regf_0.rf[9][3] ;
 wire \po_0.regf_0.rf[9][4] ;
 wire \po_0.regf_0.rf[9][5] ;
 wire \po_0.regf_0.rf[9][6] ;
 wire \po_0.regf_0.rf[9][7] ;
 wire \po_0.regf_0.rp_addr[0] ;
 wire \po_0.regf_0.rp_addr[1] ;
 wire \po_0.regf_0.rp_addr[2] ;
 wire \po_0.regf_0.rp_addr[3] ;
 wire \po_0.regf_0.rp_rd ;
 wire \po_0.regf_0.rq_addr[0] ;
 wire \po_0.regf_0.rq_addr[1] ;
 wire \po_0.regf_0.rq_addr[2] ;
 wire \po_0.regf_0.rq_addr[3] ;
 wire \po_0.regf_0.rq_rd ;
 wire \po_0.regf_0.w_addr[0] ;
 wire \po_0.regf_0.w_addr[1] ;
 wire \po_0.regf_0.w_addr[2] ;
 wire \po_0.regf_0.w_addr[3] ;
 wire \po_0.regf_0.w_wr ;
 wire \uc_0._00_ ;
 wire \uc_0._01_ ;
 wire \uc_0._02_ ;
 wire \uc_0._21_[0] ;
 wire \uc_0._21_[1] ;
 wire \uc_0._21_[2] ;
 wire \uc_0._21_[3] ;
 wire \uc_0._21_[4] ;
 wire \uc_0._21_[5] ;
 wire \uc_0._21_[6] ;
 wire \uc_0._21_[7] ;
 wire \uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[0] ;
 wire \uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[1] ;
 wire \uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[2] ;
 wire \uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[3] ;
 wire \uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[4] ;
 wire \uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[5] ;
 wire \uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[6] ;
 wire \uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[7] ;
 wire \uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[0] ;
 wire \uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[1] ;
 wire \uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[2] ;
 wire \uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[3] ;
 wire \uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[4] ;
 wire \uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[5] ;
 wire \uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[6] ;
 wire \uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[7] ;
 wire \uc_0.bc_0._12_[0] ;
 wire \uc_0.bc_0._12_[1] ;
 wire \uc_0.bc_0._12_[2] ;
 wire \uc_0.bc_0._12_[3] ;
 wire \uc_0.bc_0._14_[0] ;
 wire \uc_0.bc_0._14_[1] ;
 wire \uc_0.bc_0._14_[2] ;
 wire \uc_0.bc_0._14_[3] ;
 wire \uc_0.bc_0._14_[4] ;
 wire \uc_0.bc_0._14_[5] ;
 wire \uc_0.bc_0._14_[6] ;
 wire \uc_0.bc_0._14_[7] ;
 wire \uc_0.bc_0._85_[0] ;
 wire \uc_0.bc_0._85_[1] ;
 wire \uc_0.bc_0._85_[2] ;
 wire \uc_0.bc_0._85_[3] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\po_0.muxf_0.rf_w_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\po_0.regf_0._5_[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net57));
 sky130_fd_sc_hd__decap_8 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_95 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 _0889_ (.A(\po_0.alu_0.s0 ),
    .X(_0447_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0890_ (.A(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0891_ (.A(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_2 _0892_ (.A(\po_0.alu_0.s1 ),
    .X(_0450_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0893_ (.A(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0894_ (.A(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0895_ (.A(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__or2b_1 _0896_ (.A(_0449_),
    .B_N(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _0897_ (.A(_0454_),
    .X(_0888_));
 sky130_fd_sc_hd__or2b_1 _0898_ (.A(_0449_),
    .B_N(_0453_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_1 _0899_ (.A(_0455_),
    .X(_0887_));
 sky130_fd_sc_hd__or2b_1 _0900_ (.A(_0449_),
    .B_N(_0453_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _0901_ (.A(_0456_),
    .X(_0886_));
 sky130_fd_sc_hd__or2b_1 _0902_ (.A(_0449_),
    .B_N(_0453_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _0903_ (.A(_0457_),
    .X(_0885_));
 sky130_fd_sc_hd__or2b_1 _0904_ (.A(_0449_),
    .B_N(_0453_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _0905_ (.A(_0458_),
    .X(_0884_));
 sky130_fd_sc_hd__or2b_1 _0906_ (.A(_0449_),
    .B_N(_0453_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_1 _0907_ (.A(_0459_),
    .X(_0883_));
 sky130_fd_sc_hd__or2b_1 _0908_ (.A(_0448_),
    .B_N(_0452_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _0909_ (.A(_0460_),
    .X(_0882_));
 sky130_fd_sc_hd__or2b_1 _0910_ (.A(_0448_),
    .B_N(_0452_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _0911_ (.A(_0461_),
    .X(_0881_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0912_ (.A(\uc_0.bc_0._12_[3] ),
    .X(_0462_));
 sky130_fd_sc_hd__and4bb_1 _0913_ (.A_N(\uc_0.bc_0._12_[1] ),
    .B_N(_0462_),
    .C(\uc_0.bc_0._12_[2] ),
    .D(\uc_0.bc_0._12_[0] ),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_2 _0914_ (.A(\uc_0.bc_0._14_[5] ),
    .X(_0464_));
 sky130_fd_sc_hd__nor2_1 _0915_ (.A(_0464_),
    .B(\uc_0.bc_0._14_[7] ),
    .Y(_0465_));
 sky130_fd_sc_hd__clkbuf_2 _0916_ (.A(\uc_0.bc_0._12_[2] ),
    .X(_0466_));
 sky130_fd_sc_hd__nor2_1 _0917_ (.A(_0462_),
    .B(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__clkbuf_2 _0918_ (.A(\uc_0.bc_0._12_[1] ),
    .X(_0468_));
 sky130_fd_sc_hd__nor2b_2 _0919_ (.A(_0468_),
    .B_N(\uc_0.bc_0._12_[0] ),
    .Y(_0469_));
 sky130_fd_sc_hd__clkbuf_2 _0920_ (.A(\uc_0.bc_0._12_[0] ),
    .X(_0470_));
 sky130_fd_sc_hd__nor4b_1 _0921_ (.A(_0470_),
    .B(_0462_),
    .C(_0466_),
    .D_N(_0468_),
    .Y(_0471_));
 sky130_fd_sc_hd__clkbuf_2 _0922_ (.A(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__a221oi_1 _0923_ (.A1(_0463_),
    .A2(_0465_),
    .B1(_0467_),
    .B2(_0469_),
    .C1(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__nor2_1 _0924_ (.A(net58),
    .B(_0473_),
    .Y(\uc_0.bc_0._85_[1] ));
 sky130_fd_sc_hd__or2_1 _0925_ (.A(\uc_0.bc_0._14_[5] ),
    .B(\uc_0.bc_0._14_[7] ),
    .X(_0474_));
 sky130_fd_sc_hd__or4bb_1 _0926_ (.A(\uc_0.bc_0._12_[1] ),
    .B(\uc_0.bc_0._12_[3] ),
    .C_N(\uc_0.bc_0._12_[2] ),
    .D_N(\uc_0.bc_0._12_[0] ),
    .X(_0475_));
 sky130_fd_sc_hd__and4b_1 _0927_ (.A_N(\uc_0.bc_0._12_[2] ),
    .B(\uc_0.bc_0._12_[3] ),
    .C(\uc_0.bc_0._12_[1] ),
    .D(\uc_0.bc_0._12_[0] ),
    .X(_0476_));
 sky130_fd_sc_hd__nor4_1 _0928_ (.A(net24),
    .B(net50),
    .C(net26),
    .D(net25),
    .Y(_0477_));
 sky130_fd_sc_hd__clkbuf_2 _0929_ (.A(net20),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_2 _0930_ (.A(net19),
    .X(_0479_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0931_ (.A(net21),
    .X(_0480_));
 sky130_fd_sc_hd__nor4_1 _0932_ (.A(_0478_),
    .B(_0479_),
    .C(net51),
    .D(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__nand3_1 _0933_ (.A(_0476_),
    .B(_0477_),
    .C(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__nor3b_1 _0934_ (.A(\uc_0.bc_0._12_[3] ),
    .B(\uc_0.bc_0._12_[2] ),
    .C_N(\uc_0.bc_0._12_[1] ),
    .Y(_0483_));
 sky130_fd_sc_hd__nor4b_1 _0935_ (.A(\uc_0.bc_0._12_[0] ),
    .B(\uc_0.bc_0._12_[1] ),
    .C(\uc_0.bc_0._12_[3] ),
    .D_N(\uc_0.bc_0._12_[2] ),
    .Y(_0484_));
 sky130_fd_sc_hd__a21oi_1 _0936_ (.A1(_0470_),
    .A2(_0483_),
    .B1(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__o311a_1 _0937_ (.A1(_0474_),
    .A2(\uc_0.bc_0._14_[6] ),
    .A3(_0475_),
    .B1(_0482_),
    .C1(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__nor2_1 _0938_ (.A(net58),
    .B(_0486_),
    .Y(\uc_0.bc_0._85_[2] ));
 sky130_fd_sc_hd__clkbuf_2 _0939_ (.A(net59),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_2 _0940_ (.A(_0484_),
    .X(_0488_));
 sky130_fd_sc_hd__a211oi_2 _0941_ (.A1(_0469_),
    .A2(_0467_),
    .B1(_0483_),
    .C1(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__a211o_1 _0942_ (.A1(_0464_),
    .A2(\uc_0.bc_0._14_[6] ),
    .B1(\uc_0.bc_0._14_[7] ),
    .C1(\uc_0.bc_0._14_[4] ),
    .X(_0490_));
 sky130_fd_sc_hd__a211o_1 _0943_ (.A1(_0463_),
    .A2(_0490_),
    .B1(_0488_),
    .C1(_0471_),
    .X(_0491_));
 sky130_fd_sc_hd__a31oi_2 _0944_ (.A1(_0475_),
    .A2(_0482_),
    .A3(_0489_),
    .B1(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__clkbuf_2 _0945_ (.A(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__nor2_1 _0946_ (.A(_0487_),
    .B(_0493_),
    .Y(\uc_0.bc_0._85_[0] ));
 sky130_fd_sc_hd__a21o_1 _0947_ (.A1(_0464_),
    .A2(\uc_0.bc_0._14_[6] ),
    .B1(\uc_0.bc_0._14_[7] ),
    .X(_0494_));
 sky130_fd_sc_hd__nor2_1 _0948_ (.A(_0464_),
    .B(\uc_0.bc_0._14_[6] ),
    .Y(_0495_));
 sky130_fd_sc_hd__o31a_2 _0949_ (.A1(_0494_),
    .A2(_0495_),
    .A3(_0475_),
    .B1(_0482_),
    .X(_0496_));
 sky130_fd_sc_hd__nor2_2 _0950_ (.A(net60),
    .B(_0496_),
    .Y(\uc_0.bc_0._85_[3] ));
 sky130_fd_sc_hd__or2_1 _0951_ (.A(net19),
    .B(\po_0._1_[0] ),
    .X(_0497_));
 sky130_fd_sc_hd__nand2_1 _0952_ (.A(_0479_),
    .B(\po_0._1_[0] ),
    .Y(_0498_));
 sky130_fd_sc_hd__and2_1 _0953_ (.A(_0497_),
    .B(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_1 _0954_ (.A(_0499_),
    .X(\po_0.alu_0._10_[0] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0955_ (.A(_0006_),
    .X(_0500_));
 sky130_fd_sc_hd__buf_2 _0956_ (.A(_0004_),
    .X(_0501_));
 sky130_fd_sc_hd__buf_2 _0957_ (.A(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__buf_2 _0958_ (.A(_0005_),
    .X(_0503_));
 sky130_fd_sc_hd__clkbuf_2 _0959_ (.A(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__mux4_1 _0960_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(\po_0.regf_0.rf[9][0] ),
    .A2(\po_0.regf_0.rf[10][0] ),
    .A3(\po_0.regf_0.rf[11][0] ),
    .S0(_0502_),
    .S1(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__and2b_1 _0961_ (.A_N(_0500_),
    .B(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__clkbuf_4 _0962_ (.A(_0501_),
    .X(_0507_));
 sky130_fd_sc_hd__buf_2 _0963_ (.A(_0503_),
    .X(_0508_));
 sky130_fd_sc_hd__mux4_1 _0964_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(\po_0.regf_0.rf[13][0] ),
    .A2(\po_0.regf_0.rf[14][0] ),
    .A3(\po_0.regf_0.rf[15][0] ),
    .S0(_0507_),
    .S1(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__buf_2 _0965_ (.A(_0006_),
    .X(_0510_));
 sky130_fd_sc_hd__clkbuf_2 _0966_ (.A(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__clkbuf_2 _0967_ (.A(_0007_),
    .X(_0512_));
 sky130_fd_sc_hd__a21bo_1 _0968_ (.A1(_0509_),
    .A2(_0511_),
    .B1_N(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_2 _0969_ (.A(_0006_),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_4 _0970_ (.A(_0501_),
    .X(_0515_));
 sky130_fd_sc_hd__buf_2 _0971_ (.A(_0503_),
    .X(_0516_));
 sky130_fd_sc_hd__mux4_1 _0972_ (.A0(\po_0.regf_0.rf[0][0] ),
    .A1(\po_0.regf_0.rf[1][0] ),
    .A2(\po_0.regf_0.rf[2][0] ),
    .A3(\po_0.regf_0.rf[3][0] ),
    .S0(_0515_),
    .S1(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__and2b_1 _0973_ (.A_N(_0514_),
    .B(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__mux4_1 _0974_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(\po_0.regf_0.rf[5][0] ),
    .A2(\po_0.regf_0.rf[6][0] ),
    .A3(\po_0.regf_0.rf[7][0] ),
    .S0(_0507_),
    .S1(_0508_),
    .X(_0519_));
 sky130_fd_sc_hd__clkbuf_2 _0975_ (.A(_0007_),
    .X(_0520_));
 sky130_fd_sc_hd__a21o_1 _0976_ (.A1(_0519_),
    .A2(_0511_),
    .B1(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__o22a_1 _0977_ (.A1(_0506_),
    .A2(_0513_),
    .B1(_0518_),
    .B2(_0521_),
    .X(\po_0.regf_0._5_[0] ));
 sky130_fd_sc_hd__clkbuf_4 _0978_ (.A(_0501_),
    .X(_0522_));
 sky130_fd_sc_hd__buf_2 _0979_ (.A(_0503_),
    .X(_0523_));
 sky130_fd_sc_hd__mux4_1 _0980_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(\po_0.regf_0.rf[13][1] ),
    .A2(\po_0.regf_0.rf[14][1] ),
    .A3(\po_0.regf_0.rf[15][1] ),
    .S0(_0522_),
    .S1(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__clkbuf_2 _0981_ (.A(_0510_),
    .X(_0525_));
 sky130_fd_sc_hd__a21bo_1 _0982_ (.A1(_0524_),
    .A2(_0525_),
    .B1_N(_0007_),
    .X(_0526_));
 sky130_fd_sc_hd__mux4_1 _0983_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(\po_0.regf_0.rf[9][1] ),
    .A2(\po_0.regf_0.rf[10][1] ),
    .A3(\po_0.regf_0.rf[11][1] ),
    .S0(_0515_),
    .S1(_0516_),
    .X(_0527_));
 sky130_fd_sc_hd__and2b_1 _0984_ (.A_N(_0514_),
    .B(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__clkbuf_4 _0985_ (.A(_0004_),
    .X(_0529_));
 sky130_fd_sc_hd__buf_2 _0986_ (.A(_0005_),
    .X(_0530_));
 sky130_fd_sc_hd__mux4_1 _0987_ (.A0(\po_0.regf_0.rf[0][1] ),
    .A1(\po_0.regf_0.rf[1][1] ),
    .A2(\po_0.regf_0.rf[2][1] ),
    .A3(\po_0.regf_0.rf[3][1] ),
    .S0(_0529_),
    .S1(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__mux4_1 _0988_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(\po_0.regf_0.rf[5][1] ),
    .A2(\po_0.regf_0.rf[6][1] ),
    .A3(\po_0.regf_0.rf[7][1] ),
    .S0(_0529_),
    .S1(_0530_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _0989_ (.A0(_0531_),
    .A1(_0532_),
    .S(_0510_),
    .X(_0533_));
 sky130_fd_sc_hd__o22a_1 _0990_ (.A1(_0526_),
    .A2(_0528_),
    .B1(_0520_),
    .B2(_0533_),
    .X(\po_0.regf_0._5_[1] ));
 sky130_fd_sc_hd__mux4_1 _0991_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(\po_0.regf_0.rf[9][2] ),
    .A2(\po_0.regf_0.rf[10][2] ),
    .A3(\po_0.regf_0.rf[11][2] ),
    .S0(_0502_),
    .S1(_0504_),
    .X(_0534_));
 sky130_fd_sc_hd__and2b_1 _0992_ (.A_N(_0500_),
    .B(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__mux4_1 _0993_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(\po_0.regf_0.rf[13][2] ),
    .A2(\po_0.regf_0.rf[14][2] ),
    .A3(\po_0.regf_0.rf[15][2] ),
    .S0(_0507_),
    .S1(_0508_),
    .X(_0536_));
 sky130_fd_sc_hd__a21bo_1 _0994_ (.A1(_0536_),
    .A2(_0511_),
    .B1_N(_0512_),
    .X(_0537_));
 sky130_fd_sc_hd__mux4_1 _0995_ (.A0(\po_0.regf_0.rf[0][2] ),
    .A1(\po_0.regf_0.rf[1][2] ),
    .A2(\po_0.regf_0.rf[2][2] ),
    .A3(\po_0.regf_0.rf[3][2] ),
    .S0(_0515_),
    .S1(_0516_),
    .X(_0538_));
 sky130_fd_sc_hd__and2b_1 _0996_ (.A_N(_0514_),
    .B(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__mux4_1 _0997_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(\po_0.regf_0.rf[5][2] ),
    .A2(\po_0.regf_0.rf[6][2] ),
    .A3(\po_0.regf_0.rf[7][2] ),
    .S0(_0507_),
    .S1(_0508_),
    .X(_0540_));
 sky130_fd_sc_hd__a21o_1 _0998_ (.A1(_0540_),
    .A2(_0511_),
    .B1(_0520_),
    .X(_0541_));
 sky130_fd_sc_hd__o22a_1 _0999_ (.A1(_0535_),
    .A2(_0537_),
    .B1(_0539_),
    .B2(_0541_),
    .X(\po_0.regf_0._5_[2] ));
 sky130_fd_sc_hd__mux4_1 _1000_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(\po_0.regf_0.rf[13][3] ),
    .A2(\po_0.regf_0.rf[14][3] ),
    .A3(\po_0.regf_0.rf[15][3] ),
    .S0(_0522_),
    .S1(_0523_),
    .X(_0542_));
 sky130_fd_sc_hd__a21bo_1 _1001_ (.A1(_0542_),
    .A2(_0525_),
    .B1_N(_0007_),
    .X(_0543_));
 sky130_fd_sc_hd__mux4_1 _1002_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(\po_0.regf_0.rf[9][3] ),
    .A2(\po_0.regf_0.rf[10][3] ),
    .A3(\po_0.regf_0.rf[11][3] ),
    .S0(_0515_),
    .S1(_0516_),
    .X(_0544_));
 sky130_fd_sc_hd__and2b_1 _1003_ (.A_N(_0514_),
    .B(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__mux4_1 _1004_ (.A0(\po_0.regf_0.rf[0][3] ),
    .A1(\po_0.regf_0.rf[1][3] ),
    .A2(\po_0.regf_0.rf[2][3] ),
    .A3(\po_0.regf_0.rf[3][3] ),
    .S0(_0529_),
    .S1(_0530_),
    .X(_0546_));
 sky130_fd_sc_hd__mux4_1 _1005_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(\po_0.regf_0.rf[5][3] ),
    .A2(\po_0.regf_0.rf[6][3] ),
    .A3(\po_0.regf_0.rf[7][3] ),
    .S0(_0529_),
    .S1(_0530_),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _1006_ (.A0(_0546_),
    .A1(_0547_),
    .S(_0510_),
    .X(_0548_));
 sky130_fd_sc_hd__o22a_1 _1007_ (.A1(_0543_),
    .A2(_0545_),
    .B1(_0520_),
    .B2(_0548_),
    .X(\po_0.regf_0._5_[3] ));
 sky130_fd_sc_hd__mux4_1 _1008_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(\po_0.regf_0.rf[9][4] ),
    .A2(\po_0.regf_0.rf[10][4] ),
    .A3(\po_0.regf_0.rf[11][4] ),
    .S0(_0502_),
    .S1(_0504_),
    .X(_0549_));
 sky130_fd_sc_hd__and2b_1 _1009_ (.A_N(_0500_),
    .B(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__mux4_1 _1010_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(\po_0.regf_0.rf[13][4] ),
    .A2(\po_0.regf_0.rf[14][4] ),
    .A3(\po_0.regf_0.rf[15][4] ),
    .S0(_0522_),
    .S1(_0523_),
    .X(_0551_));
 sky130_fd_sc_hd__a21bo_1 _1011_ (.A1(_0551_),
    .A2(_0525_),
    .B1_N(_0512_),
    .X(_0552_));
 sky130_fd_sc_hd__mux4_1 _1012_ (.A0(\po_0.regf_0.rf[0][4] ),
    .A1(\po_0.regf_0.rf[1][4] ),
    .A2(\po_0.regf_0.rf[2][4] ),
    .A3(\po_0.regf_0.rf[3][4] ),
    .S0(_0515_),
    .S1(_0516_),
    .X(_0553_));
 sky130_fd_sc_hd__and2b_1 _1013_ (.A_N(_0514_),
    .B(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__mux4_1 _1014_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(\po_0.regf_0.rf[5][4] ),
    .A2(\po_0.regf_0.rf[6][4] ),
    .A3(\po_0.regf_0.rf[7][4] ),
    .S0(_0507_),
    .S1(_0508_),
    .X(_0555_));
 sky130_fd_sc_hd__a21o_1 _1015_ (.A1(_0555_),
    .A2(_0511_),
    .B1(_0512_),
    .X(_0556_));
 sky130_fd_sc_hd__o22a_1 _1016_ (.A1(_0550_),
    .A2(_0552_),
    .B1(_0554_),
    .B2(_0556_),
    .X(\po_0.regf_0._5_[4] ));
 sky130_fd_sc_hd__mux4_1 _1017_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(\po_0.regf_0.rf[13][5] ),
    .A2(\po_0.regf_0.rf[14][5] ),
    .A3(\po_0.regf_0.rf[15][5] ),
    .S0(_0522_),
    .S1(_0523_),
    .X(_0557_));
 sky130_fd_sc_hd__a21bo_1 _1018_ (.A1(_0557_),
    .A2(_0525_),
    .B1_N(_0007_),
    .X(_0558_));
 sky130_fd_sc_hd__mux4_1 _1019_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(\po_0.regf_0.rf[9][5] ),
    .A2(\po_0.regf_0.rf[10][5] ),
    .A3(\po_0.regf_0.rf[11][5] ),
    .S0(_0502_),
    .S1(_0504_),
    .X(_0559_));
 sky130_fd_sc_hd__and2b_1 _1020_ (.A_N(_0500_),
    .B(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__mux4_1 _1021_ (.A0(\po_0.regf_0.rf[0][5] ),
    .A1(\po_0.regf_0.rf[1][5] ),
    .A2(\po_0.regf_0.rf[2][5] ),
    .A3(\po_0.regf_0.rf[3][5] ),
    .S0(_0529_),
    .S1(_0530_),
    .X(_0561_));
 sky130_fd_sc_hd__mux4_1 _1022_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(\po_0.regf_0.rf[5][5] ),
    .A2(\po_0.regf_0.rf[6][5] ),
    .A3(\po_0.regf_0.rf[7][5] ),
    .S0(_0501_),
    .S1(_0503_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _1023_ (.A0(_0561_),
    .A1(_0562_),
    .S(_0510_),
    .X(_0563_));
 sky130_fd_sc_hd__o22a_1 _1024_ (.A1(_0558_),
    .A2(_0560_),
    .B1(_0520_),
    .B2(_0563_),
    .X(\po_0.regf_0._5_[5] ));
 sky130_fd_sc_hd__mux4_1 _1025_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(\po_0.regf_0.rf[9][6] ),
    .A2(\po_0.regf_0.rf[10][6] ),
    .A3(\po_0.regf_0.rf[11][6] ),
    .S0(_0502_),
    .S1(_0504_),
    .X(_0564_));
 sky130_fd_sc_hd__and2b_1 _1026_ (.A_N(_0500_),
    .B(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__mux4_1 _1027_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(\po_0.regf_0.rf[13][6] ),
    .A2(\po_0.regf_0.rf[14][6] ),
    .A3(\po_0.regf_0.rf[15][6] ),
    .S0(_0522_),
    .S1(_0523_),
    .X(_0566_));
 sky130_fd_sc_hd__a21bo_1 _1028_ (.A1(_0566_),
    .A2(_0525_),
    .B1_N(_0512_),
    .X(_0567_));
 sky130_fd_sc_hd__mux4_1 _1029_ (.A0(\po_0.regf_0.rf[0][6] ),
    .A1(\po_0.regf_0.rf[1][6] ),
    .A2(\po_0.regf_0.rf[2][6] ),
    .A3(\po_0.regf_0.rf[3][6] ),
    .S0(_0515_),
    .S1(_0516_),
    .X(_0568_));
 sky130_fd_sc_hd__and2b_1 _1030_ (.A_N(_0514_),
    .B(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__mux4_1 _1031_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(\po_0.regf_0.rf[5][6] ),
    .A2(\po_0.regf_0.rf[6][6] ),
    .A3(\po_0.regf_0.rf[7][6] ),
    .S0(_0507_),
    .S1(_0508_),
    .X(_0570_));
 sky130_fd_sc_hd__a21o_1 _1032_ (.A1(_0570_),
    .A2(_0511_),
    .B1(_0512_),
    .X(_0571_));
 sky130_fd_sc_hd__o22a_1 _1033_ (.A1(_0565_),
    .A2(_0567_),
    .B1(_0569_),
    .B2(_0571_),
    .X(\po_0.regf_0._5_[6] ));
 sky130_fd_sc_hd__mux4_1 _1034_ (.A0(\po_0.regf_0.rf[12][7] ),
    .A1(\po_0.regf_0.rf[13][7] ),
    .A2(\po_0.regf_0.rf[14][7] ),
    .A3(\po_0.regf_0.rf[15][7] ),
    .S0(_0522_),
    .S1(_0523_),
    .X(_0572_));
 sky130_fd_sc_hd__a21bo_1 _1035_ (.A1(_0572_),
    .A2(_0525_),
    .B1_N(_0007_),
    .X(_0573_));
 sky130_fd_sc_hd__mux4_1 _1036_ (.A0(\po_0.regf_0.rf[8][7] ),
    .A1(\po_0.regf_0.rf[9][7] ),
    .A2(\po_0.regf_0.rf[10][7] ),
    .A3(\po_0.regf_0.rf[11][7] ),
    .S0(_0502_),
    .S1(_0504_),
    .X(_0574_));
 sky130_fd_sc_hd__and2b_1 _1037_ (.A_N(_0500_),
    .B(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__mux4_1 _1038_ (.A0(\po_0.regf_0.rf[0][7] ),
    .A1(\po_0.regf_0.rf[1][7] ),
    .A2(\po_0.regf_0.rf[2][7] ),
    .A3(\po_0.regf_0.rf[3][7] ),
    .S0(_0529_),
    .S1(_0530_),
    .X(_0576_));
 sky130_fd_sc_hd__mux4_1 _1039_ (.A0(\po_0.regf_0.rf[4][7] ),
    .A1(\po_0.regf_0.rf[5][7] ),
    .A2(\po_0.regf_0.rf[6][7] ),
    .A3(\po_0.regf_0.rf[7][7] ),
    .S0(_0501_),
    .S1(_0503_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _1040_ (.A0(_0576_),
    .A1(_0577_),
    .S(_0510_),
    .X(_0578_));
 sky130_fd_sc_hd__o22a_1 _1041_ (.A1(_0573_),
    .A2(_0575_),
    .B1(_0520_),
    .B2(_0578_),
    .X(\po_0.regf_0._5_[7] ));
 sky130_fd_sc_hd__buf_2 _1042_ (.A(_0000_),
    .X(_0579_));
 sky130_fd_sc_hd__clkbuf_4 _1043_ (.A(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__clkbuf_2 _1044_ (.A(_0001_),
    .X(_0581_));
 sky130_fd_sc_hd__buf_2 _1045_ (.A(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__mux4_1 _1046_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(\po_0.regf_0.rf[13][0] ),
    .A2(\po_0.regf_0.rf[14][0] ),
    .A3(\po_0.regf_0.rf[15][0] ),
    .S0(_0580_),
    .S1(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__clkbuf_2 _1047_ (.A(_0002_),
    .X(_0584_));
 sky130_fd_sc_hd__clkbuf_2 _1048_ (.A(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__clkbuf_2 _1049_ (.A(_0003_),
    .X(_0586_));
 sky130_fd_sc_hd__a21bo_1 _1050_ (.A1(_0583_),
    .A2(_0585_),
    .B1_N(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_2 _1051_ (.A(_0584_),
    .X(_0588_));
 sky130_fd_sc_hd__clkbuf_4 _1052_ (.A(_0579_),
    .X(_0589_));
 sky130_fd_sc_hd__buf_2 _1053_ (.A(_0581_),
    .X(_0590_));
 sky130_fd_sc_hd__mux4_1 _1054_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(\po_0.regf_0.rf[9][0] ),
    .A2(\po_0.regf_0.rf[10][0] ),
    .A3(\po_0.regf_0.rf[11][0] ),
    .S0(_0589_),
    .S1(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__and2b_1 _1055_ (.A_N(_0588_),
    .B(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__buf_2 _1056_ (.A(_0003_),
    .X(_0593_));
 sky130_fd_sc_hd__clkbuf_4 _1057_ (.A(_0579_),
    .X(_0594_));
 sky130_fd_sc_hd__buf_2 _1058_ (.A(_0581_),
    .X(_0595_));
 sky130_fd_sc_hd__mux4_1 _1059_ (.A0(\po_0.regf_0.rf[0][0] ),
    .A1(\po_0.regf_0.rf[1][0] ),
    .A2(\po_0.regf_0.rf[2][0] ),
    .A3(\po_0.regf_0.rf[3][0] ),
    .S0(_0594_),
    .S1(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__clkbuf_4 _1060_ (.A(_0000_),
    .X(_0597_));
 sky130_fd_sc_hd__buf_2 _1061_ (.A(_0001_),
    .X(_0598_));
 sky130_fd_sc_hd__mux4_1 _1062_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(\po_0.regf_0.rf[5][0] ),
    .A2(\po_0.regf_0.rf[6][0] ),
    .A3(\po_0.regf_0.rf[7][0] ),
    .S0(_0597_),
    .S1(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__clkbuf_2 _1063_ (.A(_0002_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _1064_ (.A0(_0596_),
    .A1(_0599_),
    .S(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__o22a_1 _1065_ (.A1(_0587_),
    .A2(_0592_),
    .B1(_0593_),
    .B2(_0601_),
    .X(\po_0.regf_0._3_[0] ));
 sky130_fd_sc_hd__mux4_1 _1066_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(\po_0.regf_0.rf[13][1] ),
    .A2(\po_0.regf_0.rf[14][1] ),
    .A3(\po_0.regf_0.rf[15][1] ),
    .S0(_0580_),
    .S1(_0582_),
    .X(_0602_));
 sky130_fd_sc_hd__a21bo_1 _1067_ (.A1(_0602_),
    .A2(_0585_),
    .B1_N(_0003_),
    .X(_0603_));
 sky130_fd_sc_hd__mux4_1 _1068_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(\po_0.regf_0.rf[9][1] ),
    .A2(\po_0.regf_0.rf[10][1] ),
    .A3(\po_0.regf_0.rf[11][1] ),
    .S0(_0589_),
    .S1(_0590_),
    .X(_0604_));
 sky130_fd_sc_hd__and2b_1 _1069_ (.A_N(_0588_),
    .B(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__mux4_1 _1070_ (.A0(\po_0.regf_0.rf[0][1] ),
    .A1(\po_0.regf_0.rf[1][1] ),
    .A2(\po_0.regf_0.rf[2][1] ),
    .A3(\po_0.regf_0.rf[3][1] ),
    .S0(_0594_),
    .S1(_0595_),
    .X(_0606_));
 sky130_fd_sc_hd__mux4_1 _1071_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(\po_0.regf_0.rf[5][1] ),
    .A2(\po_0.regf_0.rf[6][1] ),
    .A3(\po_0.regf_0.rf[7][1] ),
    .S0(_0597_),
    .S1(_0598_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _1072_ (.A0(_0606_),
    .A1(_0607_),
    .S(_0600_),
    .X(_0608_));
 sky130_fd_sc_hd__o22a_1 _1073_ (.A1(_0603_),
    .A2(_0605_),
    .B1(_0593_),
    .B2(_0608_),
    .X(\po_0.regf_0._3_[1] ));
 sky130_fd_sc_hd__mux4_1 _1074_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(\po_0.regf_0.rf[13][2] ),
    .A2(\po_0.regf_0.rf[14][2] ),
    .A3(\po_0.regf_0.rf[15][2] ),
    .S0(_0580_),
    .S1(_0582_),
    .X(_0609_));
 sky130_fd_sc_hd__a21bo_1 _1075_ (.A1(_0609_),
    .A2(_0585_),
    .B1_N(_0003_),
    .X(_0610_));
 sky130_fd_sc_hd__mux4_1 _1076_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(\po_0.regf_0.rf[9][2] ),
    .A2(\po_0.regf_0.rf[10][2] ),
    .A3(\po_0.regf_0.rf[11][2] ),
    .S0(_0589_),
    .S1(_0590_),
    .X(_0611_));
 sky130_fd_sc_hd__and2b_1 _1077_ (.A_N(_0588_),
    .B(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__mux4_1 _1078_ (.A0(\po_0.regf_0.rf[0][2] ),
    .A1(\po_0.regf_0.rf[1][2] ),
    .A2(\po_0.regf_0.rf[2][2] ),
    .A3(\po_0.regf_0.rf[3][2] ),
    .S0(_0597_),
    .S1(_0598_),
    .X(_0613_));
 sky130_fd_sc_hd__mux4_1 _1079_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(\po_0.regf_0.rf[5][2] ),
    .A2(\po_0.regf_0.rf[6][2] ),
    .A3(\po_0.regf_0.rf[7][2] ),
    .S0(_0597_),
    .S1(_0598_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _1080_ (.A0(_0613_),
    .A1(_0614_),
    .S(_0584_),
    .X(_0615_));
 sky130_fd_sc_hd__o22a_1 _1081_ (.A1(_0610_),
    .A2(_0612_),
    .B1(_0593_),
    .B2(_0615_),
    .X(\po_0.regf_0._3_[2] ));
 sky130_fd_sc_hd__clkbuf_4 _1082_ (.A(_0579_),
    .X(_0616_));
 sky130_fd_sc_hd__buf_2 _1083_ (.A(_0581_),
    .X(_0617_));
 sky130_fd_sc_hd__mux4_1 _1084_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(\po_0.regf_0.rf[5][3] ),
    .A2(\po_0.regf_0.rf[6][3] ),
    .A3(\po_0.regf_0.rf[7][3] ),
    .S0(_0616_),
    .S1(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__a21o_1 _1085_ (.A1(_0618_),
    .A2(_0585_),
    .B1(_0586_),
    .X(_0619_));
 sky130_fd_sc_hd__mux4_1 _1086_ (.A0(\po_0.regf_0.rf[0][3] ),
    .A1(\po_0.regf_0.rf[1][3] ),
    .A2(\po_0.regf_0.rf[2][3] ),
    .A3(\po_0.regf_0.rf[3][3] ),
    .S0(_0589_),
    .S1(_0590_),
    .X(_0620_));
 sky130_fd_sc_hd__and2b_1 _1087_ (.A_N(_0588_),
    .B(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__mux4_1 _1088_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(\po_0.regf_0.rf[13][3] ),
    .A2(\po_0.regf_0.rf[14][3] ),
    .A3(\po_0.regf_0.rf[15][3] ),
    .S0(_0616_),
    .S1(_0617_),
    .X(_0622_));
 sky130_fd_sc_hd__clkbuf_2 _1089_ (.A(_0584_),
    .X(_0623_));
 sky130_fd_sc_hd__a21bo_1 _1090_ (.A1(_0622_),
    .A2(_0623_),
    .B1_N(_0586_),
    .X(_0624_));
 sky130_fd_sc_hd__mux4_1 _1091_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(\po_0.regf_0.rf[9][3] ),
    .A2(\po_0.regf_0.rf[10][3] ),
    .A3(\po_0.regf_0.rf[11][3] ),
    .S0(_0580_),
    .S1(_0582_),
    .X(_0625_));
 sky130_fd_sc_hd__and2b_1 _1092_ (.A_N(_0623_),
    .B(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__o22a_1 _1093_ (.A1(_0619_),
    .A2(_0621_),
    .B1(_0624_),
    .B2(_0626_),
    .X(\po_0.regf_0._3_[3] ));
 sky130_fd_sc_hd__mux4_1 _1094_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(\po_0.regf_0.rf[13][4] ),
    .A2(\po_0.regf_0.rf[14][4] ),
    .A3(\po_0.regf_0.rf[15][4] ),
    .S0(_0580_),
    .S1(_0582_),
    .X(_0627_));
 sky130_fd_sc_hd__a21bo_1 _1095_ (.A1(_0627_),
    .A2(_0585_),
    .B1_N(_0003_),
    .X(_0628_));
 sky130_fd_sc_hd__mux4_1 _1096_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(\po_0.regf_0.rf[9][4] ),
    .A2(\po_0.regf_0.rf[10][4] ),
    .A3(\po_0.regf_0.rf[11][4] ),
    .S0(_0594_),
    .S1(_0595_),
    .X(_0629_));
 sky130_fd_sc_hd__and2b_1 _1097_ (.A_N(_0600_),
    .B(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__mux4_1 _1098_ (.A0(\po_0.regf_0.rf[0][4] ),
    .A1(\po_0.regf_0.rf[1][4] ),
    .A2(\po_0.regf_0.rf[2][4] ),
    .A3(\po_0.regf_0.rf[3][4] ),
    .S0(_0597_),
    .S1(_0598_),
    .X(_0631_));
 sky130_fd_sc_hd__mux4_1 _1099_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(\po_0.regf_0.rf[5][4] ),
    .A2(\po_0.regf_0.rf[6][4] ),
    .A3(\po_0.regf_0.rf[7][4] ),
    .S0(_0579_),
    .S1(_0581_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _1100_ (.A0(_0631_),
    .A1(_0632_),
    .S(_0584_),
    .X(_0633_));
 sky130_fd_sc_hd__o22a_1 _1101_ (.A1(_0628_),
    .A2(_0630_),
    .B1(_0593_),
    .B2(_0633_),
    .X(\po_0.regf_0._3_[4] ));
 sky130_fd_sc_hd__mux4_1 _1102_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(\po_0.regf_0.rf[13][5] ),
    .A2(\po_0.regf_0.rf[14][5] ),
    .A3(\po_0.regf_0.rf[15][5] ),
    .S0(_0580_),
    .S1(_0582_),
    .X(_0634_));
 sky130_fd_sc_hd__a21bo_1 _1103_ (.A1(_0634_),
    .A2(_0585_),
    .B1_N(_0003_),
    .X(_0635_));
 sky130_fd_sc_hd__mux4_1 _1104_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(\po_0.regf_0.rf[9][5] ),
    .A2(\po_0.regf_0.rf[10][5] ),
    .A3(\po_0.regf_0.rf[11][5] ),
    .S0(_0594_),
    .S1(_0595_),
    .X(_0636_));
 sky130_fd_sc_hd__and2b_1 _1105_ (.A_N(_0600_),
    .B(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__mux4_1 _1106_ (.A0(\po_0.regf_0.rf[0][5] ),
    .A1(\po_0.regf_0.rf[1][5] ),
    .A2(\po_0.regf_0.rf[2][5] ),
    .A3(\po_0.regf_0.rf[3][5] ),
    .S0(_0597_),
    .S1(_0598_),
    .X(_0638_));
 sky130_fd_sc_hd__mux4_1 _1107_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(\po_0.regf_0.rf[5][5] ),
    .A2(\po_0.regf_0.rf[6][5] ),
    .A3(\po_0.regf_0.rf[7][5] ),
    .S0(_0579_),
    .S1(_0581_),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _1108_ (.A0(_0638_),
    .A1(_0639_),
    .S(_0584_),
    .X(_0640_));
 sky130_fd_sc_hd__o22a_1 _1109_ (.A1(_0635_),
    .A2(_0637_),
    .B1(_0593_),
    .B2(_0640_),
    .X(\po_0.regf_0._3_[5] ));
 sky130_fd_sc_hd__mux4_1 _1110_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(\po_0.regf_0.rf[9][6] ),
    .A2(\po_0.regf_0.rf[10][6] ),
    .A3(\po_0.regf_0.rf[11][6] ),
    .S0(_0594_),
    .S1(_0595_),
    .X(_0641_));
 sky130_fd_sc_hd__and2b_1 _1111_ (.A_N(_0600_),
    .B(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__mux4_1 _1112_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(\po_0.regf_0.rf[13][6] ),
    .A2(\po_0.regf_0.rf[14][6] ),
    .A3(\po_0.regf_0.rf[15][6] ),
    .S0(_0616_),
    .S1(_0617_),
    .X(_0643_));
 sky130_fd_sc_hd__a21bo_1 _1113_ (.A1(_0643_),
    .A2(_0623_),
    .B1_N(_0586_),
    .X(_0644_));
 sky130_fd_sc_hd__mux4_1 _1114_ (.A0(\po_0.regf_0.rf[0][6] ),
    .A1(\po_0.regf_0.rf[1][6] ),
    .A2(\po_0.regf_0.rf[2][6] ),
    .A3(\po_0.regf_0.rf[3][6] ),
    .S0(_0589_),
    .S1(_0590_),
    .X(_0645_));
 sky130_fd_sc_hd__and2b_1 _1115_ (.A_N(_0588_),
    .B(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__mux4_1 _1116_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(\po_0.regf_0.rf[5][6] ),
    .A2(\po_0.regf_0.rf[6][6] ),
    .A3(\po_0.regf_0.rf[7][6] ),
    .S0(_0616_),
    .S1(_0617_),
    .X(_0647_));
 sky130_fd_sc_hd__a21o_1 _1117_ (.A1(_0647_),
    .A2(_0623_),
    .B1(_0593_),
    .X(_0648_));
 sky130_fd_sc_hd__o22a_1 _1118_ (.A1(_0642_),
    .A2(_0644_),
    .B1(_0646_),
    .B2(_0648_),
    .X(\po_0.regf_0._3_[6] ));
 sky130_fd_sc_hd__mux4_1 _1119_ (.A0(\po_0.regf_0.rf[8][7] ),
    .A1(\po_0.regf_0.rf[9][7] ),
    .A2(\po_0.regf_0.rf[10][7] ),
    .A3(\po_0.regf_0.rf[11][7] ),
    .S0(_0594_),
    .S1(_0595_),
    .X(_0649_));
 sky130_fd_sc_hd__and2b_1 _1120_ (.A_N(_0600_),
    .B(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__mux4_1 _1121_ (.A0(\po_0.regf_0.rf[12][7] ),
    .A1(\po_0.regf_0.rf[13][7] ),
    .A2(\po_0.regf_0.rf[14][7] ),
    .A3(\po_0.regf_0.rf[15][7] ),
    .S0(_0616_),
    .S1(_0617_),
    .X(_0651_));
 sky130_fd_sc_hd__a21bo_1 _1122_ (.A1(_0651_),
    .A2(_0623_),
    .B1_N(_0586_),
    .X(_0652_));
 sky130_fd_sc_hd__mux4_1 _1123_ (.A0(\po_0.regf_0.rf[0][7] ),
    .A1(\po_0.regf_0.rf[1][7] ),
    .A2(\po_0.regf_0.rf[2][7] ),
    .A3(\po_0.regf_0.rf[3][7] ),
    .S0(_0589_),
    .S1(_0590_),
    .X(_0653_));
 sky130_fd_sc_hd__and2b_1 _1124_ (.A_N(_0588_),
    .B(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__mux4_1 _1125_ (.A0(\po_0.regf_0.rf[4][7] ),
    .A1(\po_0.regf_0.rf[5][7] ),
    .A2(\po_0.regf_0.rf[6][7] ),
    .A3(\po_0.regf_0.rf[7][7] ),
    .S0(_0616_),
    .S1(_0617_),
    .X(_0655_));
 sky130_fd_sc_hd__a21o_1 _1126_ (.A1(_0655_),
    .A2(_0623_),
    .B1(_0586_),
    .X(_0656_));
 sky130_fd_sc_hd__o22a_1 _1127_ (.A1(_0650_),
    .A2(_0652_),
    .B1(_0654_),
    .B2(_0656_),
    .X(\po_0.regf_0._3_[7] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1128_ (.A(_0486_),
    .X(_0657_));
 sky130_fd_sc_hd__and3_2 _1129_ (.A(_0657_),
    .B(_0492_),
    .C(\uc_0.bc_0._85_[3] ),
    .X(_0658_));
 sky130_fd_sc_hd__buf_2 _1130_ (.A(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__buf_2 _1131_ (.A(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _1132_ (.A0(\po_0.regf_0.rq_addr[0] ),
    .A1(\po_0.muxf_0.rf_w_data[4] ),
    .S(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__clkbuf_1 _1133_ (.A(_0661_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _1134_ (.A0(\po_0.regf_0.rq_addr[1] ),
    .A1(\po_0.muxf_0.rf_w_data[5] ),
    .S(_0660_),
    .X(_0662_));
 sky130_fd_sc_hd__clkbuf_1 _1135_ (.A(_0662_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _1136_ (.A0(\po_0.regf_0.rq_addr[2] ),
    .A1(\po_0.muxf_0.rf_w_data[6] ),
    .S(_0660_),
    .X(_0663_));
 sky130_fd_sc_hd__clkbuf_1 _1137_ (.A(_0663_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _1138_ (.A0(\po_0.regf_0.rq_addr[3] ),
    .A1(\po_0.muxf_0.rf_w_data[7] ),
    .S(_0660_),
    .X(_0664_));
 sky130_fd_sc_hd__clkbuf_1 _1139_ (.A(_0664_),
    .X(_0015_));
 sky130_fd_sc_hd__a221o_2 _1140_ (.A1(_0463_),
    .A2(_0465_),
    .B1(_0467_),
    .B2(_0469_),
    .C1(_0472_),
    .X(_0665_));
 sky130_fd_sc_hd__nand3_4 _1141_ (.A(\uc_0.bc_0._85_[2] ),
    .B(_0496_),
    .C(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__nor3_2 _1142_ (.A(net60),
    .B(_0665_),
    .C(_0492_),
    .Y(_0667_));
 sky130_fd_sc_hd__or3b_1 _1143_ (.A(net60),
    .B(_0496_),
    .C_N(_0486_),
    .X(_0668_));
 sky130_fd_sc_hd__o32ai_4 _1144_ (.A1(_0487_),
    .A2(_0493_),
    .A3(_0666_),
    .B1(_0667_),
    .B2(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__buf_2 _1145_ (.A(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _1146_ (.A0(\po_0.regf_0.rp_addr[0] ),
    .A1(\uc_0.bc_0._14_[0] ),
    .S(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__clkbuf_1 _1147_ (.A(_0671_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _1148_ (.A0(\po_0.regf_0.rp_addr[1] ),
    .A1(\uc_0.bc_0._14_[1] ),
    .S(_0670_),
    .X(_0672_));
 sky130_fd_sc_hd__clkbuf_1 _1149_ (.A(_0672_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _1150_ (.A0(\po_0.regf_0.rp_addr[2] ),
    .A1(\uc_0.bc_0._14_[2] ),
    .S(_0670_),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_1 _1151_ (.A(_0673_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _1152_ (.A0(\po_0.regf_0.rp_addr[3] ),
    .A1(\uc_0.bc_0._14_[3] ),
    .S(_0670_),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_1 _1153_ (.A(_0674_),
    .X(_0011_));
 sky130_fd_sc_hd__clkbuf_2 _1154_ (.A(\uc_0._21_[0] ),
    .X(_0675_));
 sky130_fd_sc_hd__buf_2 _1155_ (.A(_0488_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _1156_ (.A0(\po_0.muxf_0.rf_w_data[0] ),
    .A1(_0675_),
    .S(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__clkbuf_1 _1157_ (.A(_0677_),
    .X(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[0] ));
 sky130_fd_sc_hd__mux2_1 _1158_ (.A0(\po_0.muxf_0.rf_w_data[1] ),
    .A1(\uc_0._21_[1] ),
    .S(_0676_),
    .X(_0678_));
 sky130_fd_sc_hd__clkbuf_1 _1159_ (.A(_0678_),
    .X(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[1] ));
 sky130_fd_sc_hd__clkbuf_2 _1160_ (.A(\uc_0._21_[2] ),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _1161_ (.A0(\po_0.muxf_0.rf_w_data[2] ),
    .A1(_0679_),
    .S(_0676_),
    .X(_0680_));
 sky130_fd_sc_hd__clkbuf_1 _1162_ (.A(_0680_),
    .X(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[2] ));
 sky130_fd_sc_hd__mux2_1 _1163_ (.A0(\po_0.muxf_0.rf_w_data[3] ),
    .A1(\uc_0._21_[3] ),
    .S(_0676_),
    .X(_0681_));
 sky130_fd_sc_hd__clkbuf_1 _1164_ (.A(_0681_),
    .X(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[3] ));
 sky130_fd_sc_hd__mux2_1 _1165_ (.A0(\po_0.muxf_0.rf_w_data[4] ),
    .A1(\uc_0._21_[4] ),
    .S(_0676_),
    .X(_0682_));
 sky130_fd_sc_hd__clkbuf_1 _1166_ (.A(_0682_),
    .X(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[4] ));
 sky130_fd_sc_hd__clkbuf_2 _1167_ (.A(\uc_0._21_[5] ),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _1168_ (.A0(\po_0.muxf_0.rf_w_data[5] ),
    .A1(_0683_),
    .S(_0488_),
    .X(_0684_));
 sky130_fd_sc_hd__clkbuf_1 _1169_ (.A(_0684_),
    .X(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[5] ));
 sky130_fd_sc_hd__clkbuf_2 _1170_ (.A(\uc_0._21_[6] ),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _1171_ (.A0(\po_0.muxf_0.rf_w_data[6] ),
    .A1(_0685_),
    .S(_0488_),
    .X(_0686_));
 sky130_fd_sc_hd__clkbuf_1 _1172_ (.A(_0686_),
    .X(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[6] ));
 sky130_fd_sc_hd__mux2_1 _1173_ (.A0(\po_0.muxf_0.rf_w_data[7] ),
    .A1(\uc_0._21_[7] ),
    .S(_0488_),
    .X(_0687_));
 sky130_fd_sc_hd__clkbuf_1 _1174_ (.A(_0687_),
    .X(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[7] ));
 sky130_fd_sc_hd__buf_2 _1175_ (.A(_0472_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _1176_ (.A0(\uc_0.bc_0._14_[0] ),
    .A1(_0675_),
    .S(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__clkbuf_1 _1177_ (.A(_0689_),
    .X(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[0] ));
 sky130_fd_sc_hd__mux2_1 _1178_ (.A0(\uc_0.bc_0._14_[1] ),
    .A1(\uc_0._21_[1] ),
    .S(_0688_),
    .X(_0690_));
 sky130_fd_sc_hd__clkbuf_1 _1179_ (.A(_0690_),
    .X(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[1] ));
 sky130_fd_sc_hd__mux2_1 _1180_ (.A0(\uc_0.bc_0._14_[2] ),
    .A1(_0679_),
    .S(_0688_),
    .X(_0691_));
 sky130_fd_sc_hd__clkbuf_1 _1181_ (.A(_0691_),
    .X(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[2] ));
 sky130_fd_sc_hd__mux2_1 _1182_ (.A0(\uc_0.bc_0._14_[3] ),
    .A1(\uc_0._21_[3] ),
    .S(_0688_),
    .X(_0692_));
 sky130_fd_sc_hd__clkbuf_1 _1183_ (.A(_0692_),
    .X(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[3] ));
 sky130_fd_sc_hd__mux2_1 _1184_ (.A0(\uc_0.bc_0._14_[4] ),
    .A1(\uc_0._21_[4] ),
    .S(_0688_),
    .X(_0693_));
 sky130_fd_sc_hd__clkbuf_1 _1185_ (.A(_0693_),
    .X(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[4] ));
 sky130_fd_sc_hd__mux2_1 _1186_ (.A0(_0464_),
    .A1(_0683_),
    .S(_0472_),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_1 _1187_ (.A(_0694_),
    .X(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[5] ));
 sky130_fd_sc_hd__mux2_1 _1188_ (.A0(\uc_0.bc_0._14_[6] ),
    .A1(_0685_),
    .S(_0472_),
    .X(_0695_));
 sky130_fd_sc_hd__clkbuf_1 _1189_ (.A(_0695_),
    .X(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[6] ));
 sky130_fd_sc_hd__mux2_1 _1190_ (.A0(\uc_0.bc_0._14_[7] ),
    .A1(\uc_0._21_[7] ),
    .S(_0472_),
    .X(_0696_));
 sky130_fd_sc_hd__clkbuf_1 _1191_ (.A(_0696_),
    .X(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[7] ));
 sky130_fd_sc_hd__a21bo_1 _1192_ (.A1(_0462_),
    .A2(_0466_),
    .B1_N(_0470_),
    .X(_0697_));
 sky130_fd_sc_hd__clkbuf_2 _1193_ (.A(_0697_),
    .X(net46));
 sky130_fd_sc_hd__a21o_1 _1194_ (.A1(net46),
    .A2(_0468_),
    .B1(_0469_),
    .X(net47));
 sky130_fd_sc_hd__and4b_1 _1195_ (.A_N(_0462_),
    .B(_0466_),
    .C(_0470_),
    .D(_0468_),
    .X(_0698_));
 sky130_fd_sc_hd__a21oi_1 _1196_ (.A1(_0470_),
    .A2(_0468_),
    .B1(_0466_),
    .Y(_0699_));
 sky130_fd_sc_hd__nor2_1 _1197_ (.A(_0698_),
    .B(_0699_),
    .Y(net48));
 sky130_fd_sc_hd__a31o_2 _1198_ (.A1(_0470_),
    .A2(_0468_),
    .A3(_0466_),
    .B1(_0462_),
    .X(net49));
 sky130_fd_sc_hd__and2b_1 _1199_ (.A_N(_0479_),
    .B(\po_0._1_[0] ),
    .X(_0700_));
 sky130_fd_sc_hd__or2b_1 _1200_ (.A(\po_0._1_[1] ),
    .B_N(net20),
    .X(_0701_));
 sky130_fd_sc_hd__or2b_1 _1201_ (.A(net20),
    .B_N(\po_0._1_[1] ),
    .X(_0702_));
 sky130_fd_sc_hd__nand2_1 _1202_ (.A(_0701_),
    .B(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__xor2_1 _1203_ (.A(_0700_),
    .B(_0703_),
    .X(\po_0.alu_0._10_[1] ));
 sky130_fd_sc_hd__and2b_1 _1204_ (.A_N(_0478_),
    .B(\po_0._1_[1] ),
    .X(_0704_));
 sky130_fd_sc_hd__o21ai_1 _1205_ (.A1(_0700_),
    .A2(_0704_),
    .B1(_0701_),
    .Y(_0705_));
 sky130_fd_sc_hd__nand2_1 _1206_ (.A(_0480_),
    .B(\po_0._1_[2] ),
    .Y(_0706_));
 sky130_fd_sc_hd__or2_1 _1207_ (.A(net21),
    .B(\po_0._1_[2] ),
    .X(_0707_));
 sky130_fd_sc_hd__nand2_2 _1208_ (.A(_0706_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__xor2_1 _1209_ (.A(_0705_),
    .B(_0708_),
    .X(\po_0.alu_0._10_[2] ));
 sky130_fd_sc_hd__nand2_1 _1210_ (.A(net51),
    .B(\po_0._1_[3] ),
    .Y(_0709_));
 sky130_fd_sc_hd__or2_1 _1211_ (.A(net51),
    .B(\po_0._1_[3] ),
    .X(_0710_));
 sky130_fd_sc_hd__and2_1 _1212_ (.A(_0709_),
    .B(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1213_ (.A(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__and2b_1 _1214_ (.A_N(\po_0._1_[2] ),
    .B(_0480_),
    .X(_0713_));
 sky130_fd_sc_hd__a21oi_1 _1215_ (.A1(_0705_),
    .A2(_0708_),
    .B1(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__xor2_1 _1216_ (.A(_0712_),
    .B(_0714_),
    .X(\po_0.alu_0._10_[3] ));
 sky130_fd_sc_hd__and2_1 _1217_ (.A(net50),
    .B(\po_0._1_[4] ),
    .X(_0715_));
 sky130_fd_sc_hd__nor2_1 _1218_ (.A(net50),
    .B(\po_0._1_[4] ),
    .Y(_0716_));
 sky130_fd_sc_hd__or2b_1 _1219_ (.A(\po_0._1_[3] ),
    .B_N(net51),
    .X(_0717_));
 sky130_fd_sc_hd__o21ai_1 _1220_ (.A1(_0712_),
    .A2(_0714_),
    .B1(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__o21ai_1 _1221_ (.A1(_0715_),
    .A2(_0716_),
    .B1(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__or3_1 _1222_ (.A(_0715_),
    .B(_0716_),
    .C(_0718_),
    .X(_0720_));
 sky130_fd_sc_hd__and2_1 _1223_ (.A(_0719_),
    .B(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__clkbuf_1 _1224_ (.A(_0721_),
    .X(\po_0.alu_0._10_[4] ));
 sky130_fd_sc_hd__or2b_1 _1225_ (.A(\po_0._1_[4] ),
    .B_N(net50),
    .X(_0722_));
 sky130_fd_sc_hd__and2_1 _1226_ (.A(net24),
    .B(\po_0._1_[5] ),
    .X(_0723_));
 sky130_fd_sc_hd__nor2_1 _1227_ (.A(net24),
    .B(\po_0._1_[5] ),
    .Y(_0724_));
 sky130_fd_sc_hd__nor2_1 _1228_ (.A(_0723_),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__a21oi_1 _1229_ (.A1(_0719_),
    .A2(_0722_),
    .B1(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__nand3_1 _1230_ (.A(_0719_),
    .B(_0725_),
    .C(_0722_),
    .Y(_0727_));
 sky130_fd_sc_hd__and2b_1 _1231_ (.A_N(_0726_),
    .B(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__clkbuf_1 _1232_ (.A(_0728_),
    .X(\po_0.alu_0._10_[5] ));
 sky130_fd_sc_hd__and2_1 _1233_ (.A(net25),
    .B(\po_0._1_[6] ),
    .X(_0729_));
 sky130_fd_sc_hd__nor2_1 _1234_ (.A(net25),
    .B(\po_0._1_[6] ),
    .Y(_0730_));
 sky130_fd_sc_hd__or2_1 _1235_ (.A(_0729_),
    .B(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__clkbuf_2 _1236_ (.A(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__and2b_1 _1237_ (.A_N(\po_0._1_[5] ),
    .B(net24),
    .X(_0733_));
 sky130_fd_sc_hd__nor2_1 _1238_ (.A(_0726_),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__xnor2_1 _1239_ (.A(_0732_),
    .B(_0734_),
    .Y(\po_0.alu_0._10_[6] ));
 sky130_fd_sc_hd__o21ai_1 _1240_ (.A1(_0726_),
    .A2(_0733_),
    .B1(_0732_),
    .Y(_0735_));
 sky130_fd_sc_hd__xnor2_2 _1241_ (.A(net26),
    .B(\po_0._1_[7] ),
    .Y(_0736_));
 sky130_fd_sc_hd__or2b_1 _1242_ (.A(\po_0._1_[6] ),
    .B_N(net25),
    .X(_0737_));
 sky130_fd_sc_hd__nand3_1 _1243_ (.A(_0735_),
    .B(_0736_),
    .C(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__a21o_1 _1244_ (.A1(_0735_),
    .A2(_0737_),
    .B1(_0736_),
    .X(_0739_));
 sky130_fd_sc_hd__nand2_1 _1245_ (.A(_0738_),
    .B(_0739_),
    .Y(\po_0.alu_0._10_[7] ));
 sky130_fd_sc_hd__and2b_1 _1246_ (.A_N(\po_0.muxf_0.s1 ),
    .B(\po_0.muxf_0.s0 ),
    .X(_0740_));
 sky130_fd_sc_hd__clkbuf_2 _1247_ (.A(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__and2b_1 _1248_ (.A_N(\po_0.muxf_0.s0 ),
    .B(\po_0.muxf_0.s1 ),
    .X(_0742_));
 sky130_fd_sc_hd__clkbuf_2 _1249_ (.A(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__nor2_2 _1250_ (.A(_0450_),
    .B(_0447_),
    .Y(_0744_));
 sky130_fd_sc_hd__nand2b_2 _1251_ (.A_N(\po_0.alu_0.s1 ),
    .B(\po_0.alu_0.s0 ),
    .Y(_0745_));
 sky130_fd_sc_hd__mux2_1 _1252_ (.A0(\po_0.alu_0._10_[0] ),
    .A1(\po_0.alu_0._11_[0] ),
    .S(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__or3_1 _1253_ (.A(_0479_),
    .B(_0450_),
    .C(_0447_),
    .X(_0747_));
 sky130_fd_sc_hd__nor2_2 _1254_ (.A(_0740_),
    .B(_0742_),
    .Y(_0748_));
 sky130_fd_sc_hd__o211a_1 _1255_ (.A1(_0744_),
    .A2(_0746_),
    .B1(_0747_),
    .C1(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__a221o_2 _1256_ (.A1(net1),
    .A2(_0741_),
    .B1(_0743_),
    .B2(\po_0.muxf_0.rf_w_data[0] ),
    .C1(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__clkbuf_2 _1257_ (.A(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1258_ (.A(\po_0.regf_0.w_addr[1] ),
    .X(_0752_));
 sky130_fd_sc_hd__buf_2 _1259_ (.A(\po_0.regf_0.w_wr ),
    .X(_0753_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1260_ (.A(\po_0.regf_0.w_addr[3] ),
    .X(_0754_));
 sky130_fd_sc_hd__and2b_1 _1261_ (.A_N(_0754_),
    .B(\po_0.regf_0.w_addr[2] ),
    .X(_0755_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1262_ (.A(\po_0.regf_0.w_addr[0] ),
    .X(_0756_));
 sky130_fd_sc_hd__and4b_2 _1263_ (.A_N(_0752_),
    .B(_0753_),
    .C(_0755_),
    .D(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__clkbuf_2 _1264_ (.A(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_1 _1265_ (.A0(\po_0.regf_0.rf[5][0] ),
    .A1(_0751_),
    .S(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__clkbuf_1 _1266_ (.A(_0759_),
    .X(_0016_));
 sky130_fd_sc_hd__and2b_1 _1267_ (.A_N(\po_0._1_[1] ),
    .B(_0478_),
    .X(_0760_));
 sky130_fd_sc_hd__a211o_1 _1268_ (.A1(_0479_),
    .A2(\po_0._1_[0] ),
    .B1(_0760_),
    .C1(_0704_),
    .X(_0761_));
 sky130_fd_sc_hd__and2b_1 _1269_ (.A_N(\po_0.alu_0.s1 ),
    .B(_0447_),
    .X(_0762_));
 sky130_fd_sc_hd__o21bai_1 _1270_ (.A1(_0760_),
    .A2(_0704_),
    .B1_N(_0498_),
    .Y(_0763_));
 sky130_fd_sc_hd__a22o_1 _1271_ (.A1(_0450_),
    .A2(\po_0.alu_0._11_[1] ),
    .B1(_0744_),
    .B2(_0478_),
    .X(_0764_));
 sky130_fd_sc_hd__a31o_1 _1272_ (.A1(_0761_),
    .A2(_0762_),
    .A3(_0763_),
    .B1(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__a22o_1 _1273_ (.A1(net2),
    .A2(_0740_),
    .B1(_0742_),
    .B2(\po_0.muxf_0.rf_w_data[1] ),
    .X(_0766_));
 sky130_fd_sc_hd__a21o_2 _1274_ (.A1(_0765_),
    .A2(_0748_),
    .B1(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__clkbuf_2 _1275_ (.A(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__mux2_1 _1276_ (.A0(\po_0.regf_0.rf[5][1] ),
    .A1(_0768_),
    .S(_0758_),
    .X(_0769_));
 sky130_fd_sc_hd__clkbuf_1 _1277_ (.A(_0769_),
    .X(_0017_));
 sky130_fd_sc_hd__a22o_1 _1278_ (.A1(_0450_),
    .A2(\po_0.alu_0._11_[2] ),
    .B1(_0744_),
    .B2(_0480_),
    .X(_0770_));
 sky130_fd_sc_hd__and2_1 _1279_ (.A(_0478_),
    .B(\po_0._1_[1] ),
    .X(_0771_));
 sky130_fd_sc_hd__a31oi_2 _1280_ (.A1(_0703_),
    .A2(\po_0._1_[0] ),
    .A3(_0479_),
    .B1(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__o21ai_1 _1281_ (.A1(_0708_),
    .A2(_0772_),
    .B1(_0762_),
    .Y(_0773_));
 sky130_fd_sc_hd__a21oi_1 _1282_ (.A1(_0708_),
    .A2(_0772_),
    .B1(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__o21a_1 _1283_ (.A1(_0770_),
    .A2(_0774_),
    .B1(_0748_),
    .X(_0775_));
 sky130_fd_sc_hd__a221o_2 _1284_ (.A1(net3),
    .A2(_0741_),
    .B1(_0743_),
    .B2(\po_0.muxf_0.rf_w_data[2] ),
    .C1(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__clkbuf_2 _1285_ (.A(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _1286_ (.A0(\po_0.regf_0.rf[5][2] ),
    .A1(_0777_),
    .S(_0758_),
    .X(_0778_));
 sky130_fd_sc_hd__clkbuf_1 _1287_ (.A(_0778_),
    .X(_0018_));
 sky130_fd_sc_hd__o21ai_1 _1288_ (.A1(_0708_),
    .A2(_0772_),
    .B1(_0706_),
    .Y(_0779_));
 sky130_fd_sc_hd__a21oi_1 _1289_ (.A1(_0779_),
    .A2(_0712_),
    .B1(_0745_),
    .Y(_0780_));
 sky130_fd_sc_hd__o21ai_1 _1290_ (.A1(_0712_),
    .A2(_0779_),
    .B1(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__nand2_1 _1291_ (.A(_0745_),
    .B(\po_0.alu_0._11_[3] ),
    .Y(_0782_));
 sky130_fd_sc_hd__o211ai_1 _1292_ (.A1(_0452_),
    .A2(_0448_),
    .B1(_0781_),
    .C1(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__or3_1 _1293_ (.A(net51),
    .B(_0451_),
    .C(_0447_),
    .X(_0784_));
 sky130_fd_sc_hd__a22o_1 _1294_ (.A1(net4),
    .A2(_0740_),
    .B1(_0742_),
    .B2(\po_0.muxf_0.rf_w_data[3] ),
    .X(_0785_));
 sky130_fd_sc_hd__a31o_2 _1295_ (.A1(_0783_),
    .A2(_0784_),
    .A3(_0748_),
    .B1(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__clkbuf_2 _1296_ (.A(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__mux2_1 _1297_ (.A0(\po_0.regf_0.rf[5][3] ),
    .A1(_0787_),
    .S(_0758_),
    .X(_0788_));
 sky130_fd_sc_hd__clkbuf_1 _1298_ (.A(_0788_),
    .X(_0019_));
 sky130_fd_sc_hd__nand2_1 _1299_ (.A(_0478_),
    .B(\po_0._1_[1] ),
    .Y(_0789_));
 sky130_fd_sc_hd__nand4_1 _1300_ (.A(_0706_),
    .B(_0707_),
    .C(_0709_),
    .D(_0710_),
    .Y(_0790_));
 sky130_fd_sc_hd__a21oi_1 _1301_ (.A1(_0763_),
    .A2(_0789_),
    .B1(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__and2_1 _1302_ (.A(net51),
    .B(\po_0._1_[3] ),
    .X(_0792_));
 sky130_fd_sc_hd__nor2_1 _1303_ (.A(_0715_),
    .B(_0716_),
    .Y(_0793_));
 sky130_fd_sc_hd__a311o_1 _1304_ (.A1(_0480_),
    .A2(_0710_),
    .A3(\po_0._1_[2] ),
    .B1(_0792_),
    .C1(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__a31o_1 _1305_ (.A1(_0710_),
    .A2(\po_0._1_[2] ),
    .A3(_0480_),
    .B1(_0792_),
    .X(_0795_));
 sky130_fd_sc_hd__o21ai_1 _1306_ (.A1(_0795_),
    .A2(_0791_),
    .B1(_0793_),
    .Y(_0796_));
 sky130_fd_sc_hd__o211ai_1 _1307_ (.A1(_0791_),
    .A2(_0794_),
    .B1(_0762_),
    .C1(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__a22oi_1 _1308_ (.A1(_0451_),
    .A2(\po_0.alu_0._11_[4] ),
    .B1(_0744_),
    .B2(net50),
    .Y(_0798_));
 sky130_fd_sc_hd__or2_1 _1309_ (.A(_0740_),
    .B(_0742_),
    .X(_0799_));
 sky130_fd_sc_hd__a21oi_1 _1310_ (.A1(_0797_),
    .A2(_0798_),
    .B1(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__a221o_2 _1311_ (.A1(net5),
    .A2(_0741_),
    .B1(_0743_),
    .B2(\po_0.muxf_0.rf_w_data[4] ),
    .C1(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__clkbuf_2 _1312_ (.A(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _1313_ (.A0(\po_0.regf_0.rf[5][4] ),
    .A1(_0802_),
    .S(_0757_),
    .X(_0803_));
 sky130_fd_sc_hd__clkbuf_1 _1314_ (.A(_0803_),
    .X(_0020_));
 sky130_fd_sc_hd__nand2_1 _1315_ (.A(net50),
    .B(\po_0._1_[4] ),
    .Y(_0804_));
 sky130_fd_sc_hd__a2bb2o_1 _1316_ (.A1_N(_0723_),
    .A2_N(_0724_),
    .B1(_0796_),
    .B2(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__a31oi_1 _1317_ (.A1(_0804_),
    .A2(_0796_),
    .A3(_0725_),
    .B1(_0745_),
    .Y(_0806_));
 sky130_fd_sc_hd__nand2_1 _1318_ (.A(_0805_),
    .B(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__or2b_1 _1319_ (.A(\po_0.alu_0._11_[5] ),
    .B_N(_0450_),
    .X(_0808_));
 sky130_fd_sc_hd__o311a_1 _1320_ (.A1(net24),
    .A2(_0451_),
    .A3(_0447_),
    .B1(_0808_),
    .C1(_0748_),
    .X(_0809_));
 sky130_fd_sc_hd__nand2_1 _1321_ (.A(_0807_),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__a22oi_1 _1322_ (.A1(net6),
    .A2(_0741_),
    .B1(_0743_),
    .B2(\po_0.muxf_0.rf_w_data[5] ),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_2 _1323_ (.A(_0810_),
    .B(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__clkbuf_2 _1324_ (.A(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _1325_ (.A0(\po_0.regf_0.rf[5][5] ),
    .A1(_0813_),
    .S(_0757_),
    .X(_0814_));
 sky130_fd_sc_hd__clkbuf_1 _1326_ (.A(_0814_),
    .X(_0021_));
 sky130_fd_sc_hd__nor4_1 _1327_ (.A(_0715_),
    .B(_0716_),
    .C(_0723_),
    .D(_0724_),
    .Y(_0815_));
 sky130_fd_sc_hd__o21ai_1 _1328_ (.A1(_0795_),
    .A2(_0791_),
    .B1(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__o21ba_1 _1329_ (.A1(_0804_),
    .A2(_0724_),
    .B1_N(_0723_),
    .X(_0817_));
 sky130_fd_sc_hd__a31oi_1 _1330_ (.A1(_0732_),
    .A2(_0816_),
    .A3(_0817_),
    .B1(_0745_),
    .Y(_0818_));
 sky130_fd_sc_hd__a21o_1 _1331_ (.A1(_0816_),
    .A2(_0817_),
    .B1(_0732_),
    .X(_0819_));
 sky130_fd_sc_hd__a22o_1 _1332_ (.A1(_0451_),
    .A2(\po_0.alu_0._11_[6] ),
    .B1(_0744_),
    .B2(net25),
    .X(_0820_));
 sky130_fd_sc_hd__a21oi_2 _1333_ (.A1(_0818_),
    .A2(_0819_),
    .B1(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__a22oi_2 _1334_ (.A1(net7),
    .A2(_0741_),
    .B1(_0743_),
    .B2(\po_0.muxf_0.rf_w_data[6] ),
    .Y(_0822_));
 sky130_fd_sc_hd__o21ai_4 _1335_ (.A1(_0799_),
    .A2(_0821_),
    .B1(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__clkbuf_2 _1336_ (.A(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _1337_ (.A0(\po_0.regf_0.rf[5][6] ),
    .A1(_0824_),
    .S(_0757_),
    .X(_0825_));
 sky130_fd_sc_hd__clkbuf_1 _1338_ (.A(_0825_),
    .X(_0022_));
 sky130_fd_sc_hd__inv_2 _1339_ (.A(_0736_),
    .Y(_0826_));
 sky130_fd_sc_hd__nand3b_1 _1340_ (.A_N(_0729_),
    .B(_0826_),
    .C(_0819_),
    .Y(_0827_));
 sky130_fd_sc_hd__a21oi_1 _1341_ (.A1(_0816_),
    .A2(_0817_),
    .B1(_0732_),
    .Y(_0828_));
 sky130_fd_sc_hd__o21ai_1 _1342_ (.A1(_0729_),
    .A2(_0828_),
    .B1(_0736_),
    .Y(_0829_));
 sky130_fd_sc_hd__nand3_1 _1343_ (.A(_0827_),
    .B(_0762_),
    .C(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__or2b_1 _1344_ (.A(\po_0.alu_0._11_[7] ),
    .B_N(_0451_),
    .X(_0831_));
 sky130_fd_sc_hd__o311a_1 _1345_ (.A1(net26),
    .A2(_0452_),
    .A3(_0448_),
    .B1(_0831_),
    .C1(_0748_),
    .X(_0832_));
 sky130_fd_sc_hd__a22o_1 _1346_ (.A1(net8),
    .A2(_0741_),
    .B1(_0743_),
    .B2(\po_0.muxf_0.rf_w_data[7] ),
    .X(_0833_));
 sky130_fd_sc_hd__a21oi_4 _1347_ (.A1(_0830_),
    .A2(_0832_),
    .B1(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__clkbuf_2 _1348_ (.A(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__nor2_1 _1349_ (.A(\po_0.regf_0.rf[5][7] ),
    .B(_0758_),
    .Y(_0836_));
 sky130_fd_sc_hd__a21oi_1 _1350_ (.A1(_0758_),
    .A2(_0835_),
    .B1(_0836_),
    .Y(_0023_));
 sky130_fd_sc_hd__clkbuf_2 _1351_ (.A(_0750_),
    .X(_0837_));
 sky130_fd_sc_hd__clkbuf_2 _1352_ (.A(\po_0.regf_0.w_addr[1] ),
    .X(_0838_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1353_ (.A(\po_0.regf_0.w_wr ),
    .X(_0839_));
 sky130_fd_sc_hd__and4b_2 _1354_ (.A_N(_0756_),
    .B(_0838_),
    .C(_0839_),
    .D(_0755_),
    .X(_0840_));
 sky130_fd_sc_hd__buf_2 _1355_ (.A(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _1356_ (.A0(\po_0.regf_0.rf[6][0] ),
    .A1(_0837_),
    .S(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__clkbuf_1 _1357_ (.A(_0842_),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_2 _1358_ (.A(_0767_),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _1359_ (.A0(\po_0.regf_0.rf[6][1] ),
    .A1(_0843_),
    .S(_0841_),
    .X(_0844_));
 sky130_fd_sc_hd__clkbuf_1 _1360_ (.A(_0844_),
    .X(_0025_));
 sky130_fd_sc_hd__clkbuf_2 _1361_ (.A(_0776_),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_1 _1362_ (.A0(\po_0.regf_0.rf[6][2] ),
    .A1(_0845_),
    .S(_0841_),
    .X(_0846_));
 sky130_fd_sc_hd__clkbuf_1 _1363_ (.A(_0846_),
    .X(_0026_));
 sky130_fd_sc_hd__clkbuf_2 _1364_ (.A(_0786_),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_1 _1365_ (.A0(\po_0.regf_0.rf[6][3] ),
    .A1(_0847_),
    .S(_0841_),
    .X(_0848_));
 sky130_fd_sc_hd__clkbuf_1 _1366_ (.A(_0848_),
    .X(_0027_));
 sky130_fd_sc_hd__clkbuf_2 _1367_ (.A(_0801_),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _1368_ (.A0(\po_0.regf_0.rf[6][4] ),
    .A1(_0849_),
    .S(_0840_),
    .X(_0850_));
 sky130_fd_sc_hd__clkbuf_1 _1369_ (.A(_0850_),
    .X(_0028_));
 sky130_fd_sc_hd__clkbuf_2 _1370_ (.A(_0812_),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_1 _1371_ (.A0(\po_0.regf_0.rf[6][5] ),
    .A1(_0851_),
    .S(_0840_),
    .X(_0852_));
 sky130_fd_sc_hd__clkbuf_1 _1372_ (.A(_0852_),
    .X(_0029_));
 sky130_fd_sc_hd__clkbuf_2 _1373_ (.A(_0823_),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_1 _1374_ (.A0(\po_0.regf_0.rf[6][6] ),
    .A1(_0853_),
    .S(_0840_),
    .X(_0854_));
 sky130_fd_sc_hd__clkbuf_1 _1375_ (.A(_0854_),
    .X(_0030_));
 sky130_fd_sc_hd__clkbuf_2 _1376_ (.A(_0834_),
    .X(_0855_));
 sky130_fd_sc_hd__nor2_1 _1377_ (.A(\po_0.regf_0.rf[6][7] ),
    .B(_0841_),
    .Y(_0856_));
 sky130_fd_sc_hd__a21oi_1 _1378_ (.A1(_0855_),
    .A2(_0841_),
    .B1(_0856_),
    .Y(_0031_));
 sky130_fd_sc_hd__nand3_1 _1379_ (.A(\po_0.regf_0.w_addr[0] ),
    .B(\po_0.regf_0.w_addr[1] ),
    .C(\po_0.regf_0.w_wr ),
    .Y(_0857_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1380_ (.A(\po_0.regf_0.w_addr[2] ),
    .X(_0858_));
 sky130_fd_sc_hd__or3b_2 _1381_ (.A(_0754_),
    .B(_0857_),
    .C_N(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__buf_2 _1382_ (.A(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _1383_ (.A0(_0751_),
    .A1(\po_0.regf_0.rf[7][0] ),
    .S(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__clkbuf_1 _1384_ (.A(_0861_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _1385_ (.A0(_0768_),
    .A1(\po_0.regf_0.rf[7][1] ),
    .S(_0860_),
    .X(_0862_));
 sky130_fd_sc_hd__clkbuf_1 _1386_ (.A(_0862_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _1387_ (.A0(_0777_),
    .A1(\po_0.regf_0.rf[7][2] ),
    .S(_0860_),
    .X(_0863_));
 sky130_fd_sc_hd__clkbuf_1 _1388_ (.A(_0863_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _1389_ (.A0(_0787_),
    .A1(\po_0.regf_0.rf[7][3] ),
    .S(_0860_),
    .X(_0864_));
 sky130_fd_sc_hd__clkbuf_1 _1390_ (.A(_0864_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _1391_ (.A0(_0802_),
    .A1(\po_0.regf_0.rf[7][4] ),
    .S(_0859_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_1 _1392_ (.A(_0865_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _1393_ (.A0(_0813_),
    .A1(\po_0.regf_0.rf[7][5] ),
    .S(_0859_),
    .X(_0866_));
 sky130_fd_sc_hd__clkbuf_1 _1394_ (.A(_0866_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _1395_ (.A0(_0824_),
    .A1(\po_0.regf_0.rf[7][6] ),
    .S(_0859_),
    .X(_0867_));
 sky130_fd_sc_hd__clkbuf_1 _1396_ (.A(_0867_),
    .X(_0038_));
 sky130_fd_sc_hd__nand2_1 _1397_ (.A(_0860_),
    .B(\po_0.regf_0.rf[7][7] ),
    .Y(_0868_));
 sky130_fd_sc_hd__o21ai_1 _1398_ (.A1(_0860_),
    .A2(_0835_),
    .B1(_0868_),
    .Y(_0039_));
 sky130_fd_sc_hd__buf_2 _1399_ (.A(\po_0.regf_0.w_addr[0] ),
    .X(_0869_));
 sky130_fd_sc_hd__and2b_1 _1400_ (.A_N(_0858_),
    .B(\po_0.regf_0.w_addr[3] ),
    .X(_0870_));
 sky130_fd_sc_hd__and4bb_2 _1401_ (.A_N(_0869_),
    .B_N(_0752_),
    .C(_0839_),
    .D(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__buf_2 _1402_ (.A(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _1403_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(_0837_),
    .S(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__clkbuf_1 _1404_ (.A(_0873_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _1405_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(_0843_),
    .S(_0872_),
    .X(_0874_));
 sky130_fd_sc_hd__clkbuf_1 _1406_ (.A(_0874_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _1407_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(_0845_),
    .S(_0872_),
    .X(_0875_));
 sky130_fd_sc_hd__clkbuf_1 _1408_ (.A(_0875_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _1409_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(_0847_),
    .S(_0872_),
    .X(_0876_));
 sky130_fd_sc_hd__clkbuf_1 _1410_ (.A(_0876_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _1411_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(_0849_),
    .S(_0871_),
    .X(_0877_));
 sky130_fd_sc_hd__clkbuf_1 _1412_ (.A(_0877_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _1413_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(_0851_),
    .S(_0871_),
    .X(_0878_));
 sky130_fd_sc_hd__clkbuf_1 _1414_ (.A(_0878_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _1415_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(_0853_),
    .S(_0871_),
    .X(_0879_));
 sky130_fd_sc_hd__clkbuf_1 _1416_ (.A(_0879_),
    .X(_0046_));
 sky130_fd_sc_hd__nor2_1 _1417_ (.A(\po_0.regf_0.rf[8][7] ),
    .B(_0872_),
    .Y(_0880_));
 sky130_fd_sc_hd__a21oi_1 _1418_ (.A1(_0855_),
    .A2(_0872_),
    .B1(_0880_),
    .Y(_0047_));
 sky130_fd_sc_hd__and4b_2 _1419_ (.A_N(_0752_),
    .B(_0753_),
    .C(_0870_),
    .D(_0756_),
    .X(_0184_));
 sky130_fd_sc_hd__buf_2 _1420_ (.A(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _1421_ (.A0(\po_0.regf_0.rf[9][0] ),
    .A1(_0837_),
    .S(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _1422_ (.A(_0186_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _1423_ (.A0(\po_0.regf_0.rf[9][1] ),
    .A1(_0843_),
    .S(_0185_),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_1 _1424_ (.A(_0187_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _1425_ (.A0(\po_0.regf_0.rf[9][2] ),
    .A1(_0845_),
    .S(_0185_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_1 _1426_ (.A(_0188_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _1427_ (.A0(\po_0.regf_0.rf[9][3] ),
    .A1(_0847_),
    .S(_0185_),
    .X(_0189_));
 sky130_fd_sc_hd__clkbuf_1 _1428_ (.A(_0189_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _1429_ (.A0(\po_0.regf_0.rf[9][4] ),
    .A1(_0849_),
    .S(_0184_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_1 _1430_ (.A(_0190_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1431_ (.A0(\po_0.regf_0.rf[9][5] ),
    .A1(_0851_),
    .S(_0184_),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_1 _1432_ (.A(_0191_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _1433_ (.A0(\po_0.regf_0.rf[9][6] ),
    .A1(_0853_),
    .S(_0184_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _1434_ (.A(_0192_),
    .X(_0054_));
 sky130_fd_sc_hd__nor2_1 _1435_ (.A(\po_0.regf_0.rf[9][7] ),
    .B(_0185_),
    .Y(_0193_));
 sky130_fd_sc_hd__a21oi_1 _1436_ (.A1(_0855_),
    .A2(_0185_),
    .B1(_0193_),
    .Y(_0055_));
 sky130_fd_sc_hd__nor2_1 _1437_ (.A(_0858_),
    .B(_0754_),
    .Y(_0194_));
 sky130_fd_sc_hd__and4b_2 _1438_ (.A_N(_0752_),
    .B(_0839_),
    .C(_0194_),
    .D(_0756_),
    .X(_0195_));
 sky130_fd_sc_hd__buf_2 _1439_ (.A(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _1440_ (.A0(\po_0.regf_0.rf[1][0] ),
    .A1(_0837_),
    .S(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_1 _1441_ (.A(_0197_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _1442_ (.A0(\po_0.regf_0.rf[1][1] ),
    .A1(_0843_),
    .S(_0196_),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_1 _1443_ (.A(_0198_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(\po_0.regf_0.rf[1][2] ),
    .A1(_0845_),
    .S(_0196_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_1 _1445_ (.A(_0199_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _1446_ (.A0(\po_0.regf_0.rf[1][3] ),
    .A1(_0847_),
    .S(_0196_),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_1 _1447_ (.A(_0200_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _1448_ (.A0(\po_0.regf_0.rf[1][4] ),
    .A1(_0849_),
    .S(_0195_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_1 _1449_ (.A(_0201_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1450_ (.A0(\po_0.regf_0.rf[1][5] ),
    .A1(_0851_),
    .S(_0195_),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_1 _1451_ (.A(_0202_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1452_ (.A0(\po_0.regf_0.rf[1][6] ),
    .A1(_0853_),
    .S(_0195_),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_1 _1453_ (.A(_0203_),
    .X(_0062_));
 sky130_fd_sc_hd__nor2_1 _1454_ (.A(\po_0.regf_0.rf[1][7] ),
    .B(_0196_),
    .Y(_0204_));
 sky130_fd_sc_hd__a21oi_1 _1455_ (.A1(_0855_),
    .A2(_0196_),
    .B1(_0204_),
    .Y(_0063_));
 sky130_fd_sc_hd__and2_2 _1456_ (.A(_0858_),
    .B(_0754_),
    .X(_0205_));
 sky130_fd_sc_hd__nand4_4 _1457_ (.A(_0869_),
    .B(_0838_),
    .C(_0753_),
    .D(_0205_),
    .Y(_0206_));
 sky130_fd_sc_hd__buf_2 _1458_ (.A(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _1459_ (.A0(_0751_),
    .A1(\po_0.regf_0.rf[15][0] ),
    .S(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_1 _1460_ (.A(_0208_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1461_ (.A0(_0768_),
    .A1(\po_0.regf_0.rf[15][1] ),
    .S(_0207_),
    .X(_0209_));
 sky130_fd_sc_hd__clkbuf_1 _1462_ (.A(_0209_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1463_ (.A0(_0777_),
    .A1(\po_0.regf_0.rf[15][2] ),
    .S(_0207_),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_1 _1464_ (.A(_0210_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1465_ (.A0(_0787_),
    .A1(\po_0.regf_0.rf[15][3] ),
    .S(_0207_),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_1 _1466_ (.A(_0211_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(_0802_),
    .A1(\po_0.regf_0.rf[15][4] ),
    .S(_0206_),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_1 _1468_ (.A(_0212_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1469_ (.A0(_0813_),
    .A1(\po_0.regf_0.rf[15][5] ),
    .S(_0206_),
    .X(_0213_));
 sky130_fd_sc_hd__clkbuf_1 _1470_ (.A(_0213_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1471_ (.A0(_0824_),
    .A1(\po_0.regf_0.rf[15][6] ),
    .S(_0206_),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_1 _1472_ (.A(_0214_),
    .X(_0070_));
 sky130_fd_sc_hd__nand2_1 _1473_ (.A(_0207_),
    .B(\po_0.regf_0.rf[15][7] ),
    .Y(_0215_));
 sky130_fd_sc_hd__o21ai_1 _1474_ (.A1(_0207_),
    .A2(_0835_),
    .B1(_0215_),
    .Y(_0071_));
 sky130_fd_sc_hd__and4b_2 _1475_ (.A_N(_0756_),
    .B(_0838_),
    .C(_0839_),
    .D(_0205_),
    .X(_0216_));
 sky130_fd_sc_hd__buf_2 _1476_ (.A(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _1477_ (.A0(\po_0.regf_0.rf[14][0] ),
    .A1(_0837_),
    .S(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__clkbuf_1 _1478_ (.A(_0218_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1479_ (.A0(\po_0.regf_0.rf[14][1] ),
    .A1(_0843_),
    .S(_0217_),
    .X(_0219_));
 sky130_fd_sc_hd__clkbuf_1 _1480_ (.A(_0219_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1481_ (.A0(\po_0.regf_0.rf[14][2] ),
    .A1(_0845_),
    .S(_0217_),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_1 _1482_ (.A(_0220_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1483_ (.A0(\po_0.regf_0.rf[14][3] ),
    .A1(_0847_),
    .S(_0217_),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_1 _1484_ (.A(_0221_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _1485_ (.A0(\po_0.regf_0.rf[14][4] ),
    .A1(_0849_),
    .S(_0216_),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_1 _1486_ (.A(_0222_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1487_ (.A0(\po_0.regf_0.rf[14][5] ),
    .A1(_0851_),
    .S(_0216_),
    .X(_0223_));
 sky130_fd_sc_hd__clkbuf_1 _1488_ (.A(_0223_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1489_ (.A0(\po_0.regf_0.rf[14][6] ),
    .A1(_0853_),
    .S(_0216_),
    .X(_0224_));
 sky130_fd_sc_hd__clkbuf_1 _1490_ (.A(_0224_),
    .X(_0078_));
 sky130_fd_sc_hd__nor2_1 _1491_ (.A(\po_0.regf_0.rf[14][7] ),
    .B(_0217_),
    .Y(_0225_));
 sky130_fd_sc_hd__a21oi_1 _1492_ (.A1(_0855_),
    .A2(_0217_),
    .B1(_0225_),
    .Y(_0079_));
 sky130_fd_sc_hd__nand4b_4 _1493_ (.A_N(_0838_),
    .B(_0753_),
    .C(_0205_),
    .D(_0869_),
    .Y(_0226_));
 sky130_fd_sc_hd__buf_2 _1494_ (.A(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(_0751_),
    .A1(\po_0.regf_0.rf[13][0] ),
    .S(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_1 _1496_ (.A(_0228_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _1497_ (.A0(_0768_),
    .A1(\po_0.regf_0.rf[13][1] ),
    .S(_0227_),
    .X(_0229_));
 sky130_fd_sc_hd__clkbuf_1 _1498_ (.A(_0229_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _1499_ (.A0(_0777_),
    .A1(\po_0.regf_0.rf[13][2] ),
    .S(_0227_),
    .X(_0230_));
 sky130_fd_sc_hd__clkbuf_1 _1500_ (.A(_0230_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _1501_ (.A0(_0787_),
    .A1(\po_0.regf_0.rf[13][3] ),
    .S(_0227_),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_1 _1502_ (.A(_0231_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _1503_ (.A0(_0802_),
    .A1(\po_0.regf_0.rf[13][4] ),
    .S(_0226_),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_1 _1504_ (.A(_0232_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _1505_ (.A0(_0813_),
    .A1(\po_0.regf_0.rf[13][5] ),
    .S(_0226_),
    .X(_0233_));
 sky130_fd_sc_hd__clkbuf_1 _1506_ (.A(_0233_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _1507_ (.A0(_0824_),
    .A1(\po_0.regf_0.rf[13][6] ),
    .S(_0226_),
    .X(_0234_));
 sky130_fd_sc_hd__clkbuf_1 _1508_ (.A(_0234_),
    .X(_0086_));
 sky130_fd_sc_hd__nand2_1 _1509_ (.A(_0227_),
    .B(\po_0.regf_0.rf[13][7] ),
    .Y(_0235_));
 sky130_fd_sc_hd__o21ai_1 _1510_ (.A1(_0227_),
    .A2(_0835_),
    .B1(_0235_),
    .Y(_0087_));
 sky130_fd_sc_hd__and4bb_2 _1511_ (.A_N(_0869_),
    .B_N(\po_0.regf_0.w_addr[1] ),
    .C(_0839_),
    .D(_0205_),
    .X(_0236_));
 sky130_fd_sc_hd__buf_2 _1512_ (.A(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _1513_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(_0837_),
    .S(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__clkbuf_1 _1514_ (.A(_0238_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _1515_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(_0843_),
    .S(_0237_),
    .X(_0239_));
 sky130_fd_sc_hd__clkbuf_1 _1516_ (.A(_0239_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1517_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(_0845_),
    .S(_0237_),
    .X(_0240_));
 sky130_fd_sc_hd__clkbuf_1 _1518_ (.A(_0240_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _1519_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(_0847_),
    .S(_0237_),
    .X(_0241_));
 sky130_fd_sc_hd__clkbuf_1 _1520_ (.A(_0241_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _1521_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(_0849_),
    .S(_0236_),
    .X(_0242_));
 sky130_fd_sc_hd__clkbuf_1 _1522_ (.A(_0242_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _1523_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(_0851_),
    .S(_0236_),
    .X(_0243_));
 sky130_fd_sc_hd__clkbuf_1 _1524_ (.A(_0243_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _1525_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(_0853_),
    .S(_0236_),
    .X(_0244_));
 sky130_fd_sc_hd__clkbuf_1 _1526_ (.A(_0244_),
    .X(_0094_));
 sky130_fd_sc_hd__nor2_1 _1527_ (.A(\po_0.regf_0.rf[12][7] ),
    .B(_0237_),
    .Y(_0245_));
 sky130_fd_sc_hd__a21oi_1 _1528_ (.A1(_0855_),
    .A2(_0237_),
    .B1(_0245_),
    .Y(_0095_));
 sky130_fd_sc_hd__clkbuf_2 _1529_ (.A(\uc_0._00_ ),
    .X(_0246_));
 sky130_fd_sc_hd__clkbuf_2 _1530_ (.A(\uc_0._02_ ),
    .X(_0247_));
 sky130_fd_sc_hd__nor2_2 _1531_ (.A(_0246_),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__clkbuf_2 _1532_ (.A(net37),
    .X(_0249_));
 sky130_fd_sc_hd__clkbuf_2 _1533_ (.A(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__xnor2_1 _1534_ (.A(_0250_),
    .B(_0675_),
    .Y(_0251_));
 sky130_fd_sc_hd__clkbuf_2 _1535_ (.A(_0247_),
    .X(_0252_));
 sky130_fd_sc_hd__nor3_2 _1536_ (.A(\uc_0._01_ ),
    .B(\uc_0._00_ ),
    .C(\uc_0._02_ ),
    .Y(_0253_));
 sky130_fd_sc_hd__mux2_1 _1537_ (.A0(_0252_),
    .A1(_0253_),
    .S(_0250_),
    .X(_0254_));
 sky130_fd_sc_hd__a31o_1 _1538_ (.A1(\uc_0._01_ ),
    .A2(_0248_),
    .A3(_0251_),
    .B1(_0254_),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_2 _1539_ (.A(net38),
    .X(_0255_));
 sky130_fd_sc_hd__or3_1 _1540_ (.A(\uc_0._01_ ),
    .B(_0246_),
    .C(\uc_0._02_ ),
    .X(_0256_));
 sky130_fd_sc_hd__clkbuf_2 _1541_ (.A(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__and2_1 _1542_ (.A(net38),
    .B(\uc_0._21_[1] ),
    .X(_0258_));
 sky130_fd_sc_hd__nor2_2 _1543_ (.A(net38),
    .B(\uc_0._21_[1] ),
    .Y(_0259_));
 sky130_fd_sc_hd__or4_1 _1544_ (.A(_0249_),
    .B(_0675_),
    .C(_0258_),
    .D(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__o22ai_2 _1545_ (.A1(net37),
    .A2(\uc_0._21_[0] ),
    .B1(_0258_),
    .B2(_0259_),
    .Y(_0261_));
 sky130_fd_sc_hd__o21ai_1 _1546_ (.A1(_0249_),
    .A2(_0255_),
    .B1(_0247_),
    .Y(_0262_));
 sky130_fd_sc_hd__a21oi_1 _1547_ (.A1(_0250_),
    .A2(_0255_),
    .B1(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__clkbuf_2 _1548_ (.A(_0253_),
    .X(_0264_));
 sky130_fd_sc_hd__a311o_1 _1549_ (.A1(_0260_),
    .A2(_0248_),
    .A3(_0261_),
    .B1(_0263_),
    .C1(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__o21a_1 _1550_ (.A1(_0255_),
    .A2(_0257_),
    .B1(_0265_),
    .X(_0097_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1551_ (.A(net57),
    .X(_0266_));
 sky130_fd_sc_hd__inv_2 _1552_ (.A(_0247_),
    .Y(_0267_));
 sky130_fd_sc_hd__a21oi_1 _1553_ (.A1(_0250_),
    .A2(_0255_),
    .B1(_0266_),
    .Y(_0268_));
 sky130_fd_sc_hd__and3_1 _1554_ (.A(_0249_),
    .B(_0255_),
    .C(_0266_),
    .X(_0269_));
 sky130_fd_sc_hd__o31ai_1 _1555_ (.A1(_0267_),
    .A2(_0268_),
    .A3(_0269_),
    .B1(_0257_),
    .Y(_0270_));
 sky130_fd_sc_hd__nor2_2 _1556_ (.A(\uc_0._21_[2] ),
    .B(net57),
    .Y(_0271_));
 sky130_fd_sc_hd__nand2_1 _1557_ (.A(_0679_),
    .B(net57),
    .Y(_0272_));
 sky130_fd_sc_hd__nand3b_1 _1558_ (.A_N(_0271_),
    .B(_0272_),
    .C(_0259_),
    .Y(_0273_));
 sky130_fd_sc_hd__o221a_1 _1559_ (.A1(_0250_),
    .A2(_0675_),
    .B1(_0258_),
    .B2(_0259_),
    .C1(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__and2_1 _1560_ (.A(\uc_0._21_[2] ),
    .B(net57),
    .X(_0275_));
 sky130_fd_sc_hd__o22ai_4 _1561_ (.A1(net38),
    .A2(\uc_0._21_[1] ),
    .B1(_0271_),
    .B2(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__a21boi_1 _1562_ (.A1(_0276_),
    .A2(_0273_),
    .B1_N(_0261_),
    .Y(_0277_));
 sky130_fd_sc_hd__a2111oi_1 _1563_ (.A1(_0274_),
    .A2(_0276_),
    .B1(_0252_),
    .C1(_0246_),
    .D1(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__o22a_1 _1564_ (.A1(_0266_),
    .A2(_0257_),
    .B1(_0270_),
    .B2(_0278_),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_2 _1565_ (.A(net40),
    .X(_0279_));
 sky130_fd_sc_hd__o21ai_1 _1566_ (.A1(_0279_),
    .A2(_0269_),
    .B1(_0247_),
    .Y(_0280_));
 sky130_fd_sc_hd__and4_1 _1567_ (.A(_0249_),
    .B(net38),
    .C(_0266_),
    .D(_0279_),
    .X(_0281_));
 sky130_fd_sc_hd__o221ai_2 _1568_ (.A1(_0249_),
    .A2(_0675_),
    .B1(_0258_),
    .B2(_0259_),
    .C1(_0273_),
    .Y(_0282_));
 sky130_fd_sc_hd__and2_1 _1569_ (.A(\uc_0._21_[3] ),
    .B(net40),
    .X(_0283_));
 sky130_fd_sc_hd__o21ai_1 _1570_ (.A1(\uc_0._21_[3] ),
    .A2(net40),
    .B1(_0271_),
    .Y(_0284_));
 sky130_fd_sc_hd__nor2_2 _1571_ (.A(\uc_0._21_[3] ),
    .B(net40),
    .Y(_0285_));
 sky130_fd_sc_hd__o22ai_1 _1572_ (.A1(_0679_),
    .A2(net57),
    .B1(_0285_),
    .B2(_0283_),
    .Y(_0286_));
 sky130_fd_sc_hd__o21ai_1 _1573_ (.A1(_0283_),
    .A2(_0284_),
    .B1(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__a21oi_1 _1574_ (.A1(_0276_),
    .A2(_0282_),
    .B1(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__a311o_1 _1575_ (.A1(_0276_),
    .A2(_0282_),
    .A3(_0287_),
    .B1(\uc_0._02_ ),
    .C1(_0246_),
    .X(_0289_));
 sky130_fd_sc_hd__o22ai_1 _1576_ (.A1(_0280_),
    .A2(_0281_),
    .B1(_0288_),
    .B2(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__mux2_1 _1577_ (.A0(_0290_),
    .A1(_0279_),
    .S(_0253_),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _1578_ (.A(_0291_),
    .X(_0099_));
 sky130_fd_sc_hd__clkbuf_2 _1579_ (.A(net41),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_2 _1580_ (.A(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__nand2_1 _1581_ (.A(_0293_),
    .B(_0281_),
    .Y(_0294_));
 sky130_fd_sc_hd__a41o_1 _1582_ (.A1(_0250_),
    .A2(_0255_),
    .A3(_0266_),
    .A4(_0279_),
    .B1(_0293_),
    .X(_0295_));
 sky130_fd_sc_hd__a31o_1 _1583_ (.A1(_0294_),
    .A2(_0252_),
    .A3(_0295_),
    .B1(_0264_),
    .X(_0296_));
 sky130_fd_sc_hd__and2b_1 _1584_ (.A_N(net41),
    .B(\uc_0._21_[4] ),
    .X(_0297_));
 sky130_fd_sc_hd__and2b_1 _1585_ (.A_N(\uc_0._21_[4] ),
    .B(_0292_),
    .X(_0298_));
 sky130_fd_sc_hd__or3_1 _1586_ (.A(_0285_),
    .B(_0297_),
    .C(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__o21ai_1 _1587_ (.A1(_0297_),
    .A2(_0298_),
    .B1(_0285_),
    .Y(_0300_));
 sky130_fd_sc_hd__o21ai_1 _1588_ (.A1(_0679_),
    .A2(net39),
    .B1(_0259_),
    .Y(_0301_));
 sky130_fd_sc_hd__nor2_1 _1589_ (.A(_0275_),
    .B(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__o21ai_1 _1590_ (.A1(_0261_),
    .A2(_0302_),
    .B1(_0276_),
    .Y(_0303_));
 sky130_fd_sc_hd__o21a_1 _1591_ (.A1(_0283_),
    .A2(_0284_),
    .B1(_0286_),
    .X(_0304_));
 sky130_fd_sc_hd__o22a_1 _1592_ (.A1(_0679_),
    .A2(_0266_),
    .B1(_0285_),
    .B2(_0283_),
    .X(_0305_));
 sky130_fd_sc_hd__a221o_1 _1593_ (.A1(_0299_),
    .A2(_0300_),
    .B1(_0303_),
    .B2(_0304_),
    .C1(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__nand2_1 _1594_ (.A(_0299_),
    .B(_0300_),
    .Y(_0307_));
 sky130_fd_sc_hd__o21bai_1 _1595_ (.A1(_0305_),
    .A2(_0288_),
    .B1_N(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__and3_1 _1596_ (.A(_0306_),
    .B(_0248_),
    .C(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__o22a_1 _1597_ (.A1(_0293_),
    .A2(_0257_),
    .B1(_0296_),
    .B2(_0309_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_2 _1598_ (.A(net56),
    .X(_0310_));
 sky130_fd_sc_hd__a31o_1 _1599_ (.A1(_0279_),
    .A2(_0293_),
    .A3(_0269_),
    .B1(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__nand4_1 _1600_ (.A(_0279_),
    .B(_0293_),
    .C(_0310_),
    .D(_0269_),
    .Y(_0312_));
 sky130_fd_sc_hd__a31o_1 _1601_ (.A1(_0311_),
    .A2(_0252_),
    .A3(_0312_),
    .B1(_0264_),
    .X(_0313_));
 sky130_fd_sc_hd__nor2_1 _1602_ (.A(net56),
    .B(_0683_),
    .Y(_0314_));
 sky130_fd_sc_hd__and2_1 _1603_ (.A(net56),
    .B(\uc_0._21_[5] ),
    .X(_0315_));
 sky130_fd_sc_hd__nor4_1 _1604_ (.A(_0292_),
    .B(\uc_0._21_[4] ),
    .C(_0314_),
    .D(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__o22a_1 _1605_ (.A1(_0292_),
    .A2(\uc_0._21_[4] ),
    .B1(_0314_),
    .B2(_0315_),
    .X(_0317_));
 sky130_fd_sc_hd__or2_1 _1606_ (.A(_0316_),
    .B(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__inv_2 _1607_ (.A(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__a21oi_1 _1608_ (.A1(_0303_),
    .A2(_0304_),
    .B1(_0305_),
    .Y(_0320_));
 sky130_fd_sc_hd__o32ai_4 _1609_ (.A1(_0285_),
    .A2(_0297_),
    .A3(_0298_),
    .B1(_0307_),
    .B2(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__a311o_1 _1610_ (.A1(_0299_),
    .A2(_0308_),
    .A3(_0318_),
    .B1(_0247_),
    .C1(_0246_),
    .X(_0322_));
 sky130_fd_sc_hd__a21oi_1 _1611_ (.A1(_0319_),
    .A2(_0321_),
    .B1(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__o22a_1 _1612_ (.A1(_0310_),
    .A2(_0257_),
    .B1(_0313_),
    .B2(_0323_),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_2 _1613_ (.A(net43),
    .X(_0324_));
 sky130_fd_sc_hd__a31o_1 _1614_ (.A1(_0293_),
    .A2(_0310_),
    .A3(_0281_),
    .B1(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__nand4_1 _1615_ (.A(_0292_),
    .B(_0310_),
    .C(net43),
    .D(_0281_),
    .Y(_0326_));
 sky130_fd_sc_hd__a31oi_1 _1616_ (.A1(_0325_),
    .A2(_0326_),
    .A3(_0252_),
    .B1(_0264_),
    .Y(_0327_));
 sky130_fd_sc_hd__a21oi_1 _1617_ (.A1(_0299_),
    .A2(_0308_),
    .B1(_0318_),
    .Y(_0328_));
 sky130_fd_sc_hd__xnor2_1 _1618_ (.A(\uc_0._21_[6] ),
    .B(net43),
    .Y(_0329_));
 sky130_fd_sc_hd__o21ai_2 _1619_ (.A1(net56),
    .A2(_0683_),
    .B1(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__or3_1 _1620_ (.A(net56),
    .B(_0683_),
    .C(_0329_),
    .X(_0331_));
 sky130_fd_sc_hd__o211ai_1 _1621_ (.A1(_0317_),
    .A2(_0328_),
    .B1(_0330_),
    .C1(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__a221o_1 _1622_ (.A1(_0330_),
    .A2(_0331_),
    .B1(_0321_),
    .B2(_0319_),
    .C1(_0317_),
    .X(_0333_));
 sky130_fd_sc_hd__nand3_1 _1623_ (.A(_0332_),
    .B(_0248_),
    .C(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__o2bb2a_1 _1624_ (.A1_N(_0327_),
    .A2_N(_0334_),
    .B1(_0257_),
    .B2(_0324_),
    .X(_0102_));
 sky130_fd_sc_hd__inv_2 _1625_ (.A(net44),
    .Y(_0335_));
 sky130_fd_sc_hd__xnor2_1 _1626_ (.A(\uc_0._21_[7] ),
    .B(net44),
    .Y(_0336_));
 sky130_fd_sc_hd__o21ba_1 _1627_ (.A1(_0685_),
    .A2(_0324_),
    .B1_N(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__nor3b_1 _1628_ (.A(_0685_),
    .B(_0324_),
    .C_N(_0336_),
    .Y(_0338_));
 sky130_fd_sc_hd__nand2_1 _1629_ (.A(_0330_),
    .B(_0331_),
    .Y(_0339_));
 sky130_fd_sc_hd__a21oi_1 _1630_ (.A1(_0321_),
    .A2(_0319_),
    .B1(_0317_),
    .Y(_0340_));
 sky130_fd_sc_hd__o21a_1 _1631_ (.A1(net56),
    .A2(_0683_),
    .B1(_0329_),
    .X(_0341_));
 sky130_fd_sc_hd__o21bai_1 _1632_ (.A1(_0339_),
    .A2(_0340_),
    .B1_N(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__o21ai_1 _1633_ (.A1(_0337_),
    .A2(_0338_),
    .B1(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__o21a_1 _1634_ (.A1(_0685_),
    .A2(net43),
    .B1(_0336_),
    .X(_0344_));
 sky130_fd_sc_hd__nor3_1 _1635_ (.A(_0685_),
    .B(_0324_),
    .C(_0336_),
    .Y(_0345_));
 sky130_fd_sc_hd__o221ai_1 _1636_ (.A1(_0344_),
    .A2(_0345_),
    .B1(_0339_),
    .B2(_0340_),
    .C1(_0330_),
    .Y(_0346_));
 sky130_fd_sc_hd__nand3_1 _1637_ (.A(_0343_),
    .B(_0248_),
    .C(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__or2_1 _1638_ (.A(_0335_),
    .B(_0326_),
    .X(_0348_));
 sky130_fd_sc_hd__a41o_1 _1639_ (.A1(_0292_),
    .A2(_0310_),
    .A3(_0324_),
    .A4(_0281_),
    .B1(net44),
    .X(_0349_));
 sky130_fd_sc_hd__a31oi_1 _1640_ (.A1(_0348_),
    .A2(_0349_),
    .A3(_0252_),
    .B1(_0264_),
    .Y(_0350_));
 sky130_fd_sc_hd__a22oi_1 _1641_ (.A1(_0335_),
    .A2(_0264_),
    .B1(_0347_),
    .B2(_0350_),
    .Y(_0103_));
 sky130_fd_sc_hd__and4bb_2 _1642_ (.A_N(_0756_),
    .B_N(\po_0.regf_0.w_addr[1] ),
    .C(_0839_),
    .D(_0755_),
    .X(_0351_));
 sky130_fd_sc_hd__buf_2 _1643_ (.A(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _1644_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(_0750_),
    .S(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_1 _1645_ (.A(_0353_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _1646_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(_0767_),
    .S(_0352_),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _1647_ (.A(_0354_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1648_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(_0776_),
    .S(_0352_),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _1649_ (.A(_0355_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _1650_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(_0786_),
    .S(_0352_),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_1 _1651_ (.A(_0356_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1652_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(_0801_),
    .S(_0351_),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _1653_ (.A(_0357_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _1654_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(_0812_),
    .S(_0351_),
    .X(_0358_));
 sky130_fd_sc_hd__clkbuf_1 _1655_ (.A(_0358_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1656_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(_0823_),
    .S(_0351_),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _1657_ (.A(_0359_),
    .X(_0110_));
 sky130_fd_sc_hd__nor2_1 _1658_ (.A(\po_0.regf_0.rf[4][7] ),
    .B(_0352_),
    .Y(_0360_));
 sky130_fd_sc_hd__a21oi_1 _1659_ (.A1(_0834_),
    .A2(_0352_),
    .B1(_0360_),
    .Y(_0111_));
 sky130_fd_sc_hd__or4b_1 _1660_ (.A(_0665_),
    .B(\uc_0.bc_0._85_[2] ),
    .C(\uc_0.bc_0._85_[3] ),
    .D_N(\uc_0.bc_0._85_[0] ),
    .X(_0361_));
 sky130_fd_sc_hd__buf_2 _1661_ (.A(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__o21a_1 _1662_ (.A1(_0487_),
    .A2(_0246_),
    .B1(_0362_),
    .X(_0112_));
 sky130_fd_sc_hd__and4_2 _1663_ (.A(_0869_),
    .B(_0838_),
    .C(_0753_),
    .D(_0194_),
    .X(_0363_));
 sky130_fd_sc_hd__buf_2 _1664_ (.A(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _1665_ (.A0(\po_0.regf_0.rf[3][0] ),
    .A1(_0750_),
    .S(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _1666_ (.A(_0365_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1667_ (.A0(\po_0.regf_0.rf[3][1] ),
    .A1(_0767_),
    .S(_0364_),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _1668_ (.A(_0366_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _1669_ (.A0(\po_0.regf_0.rf[3][2] ),
    .A1(_0776_),
    .S(_0364_),
    .X(_0367_));
 sky130_fd_sc_hd__clkbuf_1 _1670_ (.A(_0367_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _1671_ (.A0(\po_0.regf_0.rf[3][3] ),
    .A1(_0786_),
    .S(_0364_),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_1 _1672_ (.A(_0368_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _1673_ (.A0(\po_0.regf_0.rf[3][4] ),
    .A1(_0801_),
    .S(_0363_),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _1674_ (.A(_0369_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _1675_ (.A0(\po_0.regf_0.rf[3][5] ),
    .A1(_0812_),
    .S(_0363_),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_1 _1676_ (.A(_0370_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _1677_ (.A0(\po_0.regf_0.rf[3][6] ),
    .A1(_0823_),
    .S(_0363_),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_1 _1678_ (.A(_0371_),
    .X(_0119_));
 sky130_fd_sc_hd__nor2_1 _1679_ (.A(\po_0.regf_0.rf[3][7] ),
    .B(_0364_),
    .Y(_0372_));
 sky130_fd_sc_hd__a21oi_1 _1680_ (.A1(_0834_),
    .A2(_0364_),
    .B1(_0372_),
    .Y(_0120_));
 sky130_fd_sc_hd__and4b_2 _1681_ (.A_N(\po_0.regf_0.w_addr[0] ),
    .B(_0752_),
    .C(\po_0.regf_0.w_wr ),
    .D(_0870_),
    .X(_0373_));
 sky130_fd_sc_hd__buf_2 _1682_ (.A(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _1683_ (.A0(\po_0.regf_0.rf[10][0] ),
    .A1(_0750_),
    .S(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _1684_ (.A(_0375_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _1685_ (.A0(\po_0.regf_0.rf[10][1] ),
    .A1(_0767_),
    .S(_0374_),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _1686_ (.A(_0376_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _1687_ (.A0(\po_0.regf_0.rf[10][2] ),
    .A1(_0776_),
    .S(_0374_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _1688_ (.A(_0377_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1689_ (.A0(\po_0.regf_0.rf[10][3] ),
    .A1(_0786_),
    .S(_0374_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _1690_ (.A(_0378_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _1691_ (.A0(\po_0.regf_0.rf[10][4] ),
    .A1(_0801_),
    .S(_0373_),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_1 _1692_ (.A(_0379_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _1693_ (.A0(\po_0.regf_0.rf[10][5] ),
    .A1(_0812_),
    .S(_0373_),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _1694_ (.A(_0380_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1695_ (.A0(\po_0.regf_0.rf[10][6] ),
    .A1(_0823_),
    .S(_0373_),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_1 _1696_ (.A(_0381_),
    .X(_0127_));
 sky130_fd_sc_hd__nor2_1 _1697_ (.A(\po_0.regf_0.rf[10][7] ),
    .B(_0374_),
    .Y(_0382_));
 sky130_fd_sc_hd__a21oi_1 _1698_ (.A1(_0834_),
    .A2(_0374_),
    .B1(_0382_),
    .Y(_0128_));
 sky130_fd_sc_hd__and4b_2 _1699_ (.A_N(\po_0.regf_0.w_addr[0] ),
    .B(_0752_),
    .C(\po_0.regf_0.w_wr ),
    .D(_0194_),
    .X(_0383_));
 sky130_fd_sc_hd__buf_2 _1700_ (.A(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _1701_ (.A0(\po_0.regf_0.rf[2][0] ),
    .A1(_0750_),
    .S(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_1 _1702_ (.A(_0385_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _1703_ (.A0(\po_0.regf_0.rf[2][1] ),
    .A1(_0767_),
    .S(_0384_),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_1 _1704_ (.A(_0386_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _1705_ (.A0(\po_0.regf_0.rf[2][2] ),
    .A1(_0776_),
    .S(_0384_),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_1 _1706_ (.A(_0387_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _1707_ (.A0(\po_0.regf_0.rf[2][3] ),
    .A1(_0786_),
    .S(_0384_),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_1 _1708_ (.A(_0388_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _1709_ (.A0(\po_0.regf_0.rf[2][4] ),
    .A1(_0801_),
    .S(_0383_),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_1 _1710_ (.A(_0389_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _1711_ (.A0(\po_0.regf_0.rf[2][5] ),
    .A1(_0812_),
    .S(_0383_),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _1712_ (.A(_0390_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _1713_ (.A0(\po_0.regf_0.rf[2][6] ),
    .A1(_0823_),
    .S(_0383_),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_1 _1714_ (.A(_0391_),
    .X(_0135_));
 sky130_fd_sc_hd__nor2_1 _1715_ (.A(\po_0.regf_0.rf[2][7] ),
    .B(_0384_),
    .Y(_0392_));
 sky130_fd_sc_hd__a21oi_1 _1716_ (.A1(_0834_),
    .A2(_0384_),
    .B1(_0392_),
    .Y(_0136_));
 sky130_fd_sc_hd__or4bb_4 _1717_ (.A(\po_0.regf_0.w_addr[0] ),
    .B(\po_0.regf_0.w_addr[1] ),
    .C_N(\po_0.regf_0.w_wr ),
    .D_N(_0194_),
    .X(_0393_));
 sky130_fd_sc_hd__buf_2 _1718_ (.A(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _1719_ (.A0(_0751_),
    .A1(\po_0.regf_0.rf[0][0] ),
    .S(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _1720_ (.A(_0395_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _1721_ (.A0(_0768_),
    .A1(\po_0.regf_0.rf[0][1] ),
    .S(_0394_),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _1722_ (.A(_0396_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _1723_ (.A0(_0777_),
    .A1(\po_0.regf_0.rf[0][2] ),
    .S(_0394_),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_1 _1724_ (.A(_0397_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _1725_ (.A0(_0787_),
    .A1(\po_0.regf_0.rf[0][3] ),
    .S(_0394_),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_1 _1726_ (.A(_0398_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _1727_ (.A0(_0802_),
    .A1(\po_0.regf_0.rf[0][4] ),
    .S(_0393_),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _1728_ (.A(_0399_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _1729_ (.A0(_0813_),
    .A1(\po_0.regf_0.rf[0][5] ),
    .S(_0393_),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_1 _1730_ (.A(_0400_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _1731_ (.A0(_0824_),
    .A1(\po_0.regf_0.rf[0][6] ),
    .S(_0393_),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _1732_ (.A(_0401_),
    .X(_0143_));
 sky130_fd_sc_hd__nand2_1 _1733_ (.A(_0394_),
    .B(\po_0.regf_0.rf[0][7] ),
    .Y(_0402_));
 sky130_fd_sc_hd__o21ai_1 _1734_ (.A1(_0394_),
    .A2(_0835_),
    .B1(_0402_),
    .Y(_0144_));
 sky130_fd_sc_hd__and2_1 _1735_ (.A(_0657_),
    .B(\uc_0.bc_0._85_[3] ),
    .X(_0403_));
 sky130_fd_sc_hd__a21oi_1 _1736_ (.A1(_0403_),
    .A2(_0667_),
    .B1(\po_0.muxf_0.s1 ),
    .Y(_0404_));
 sky130_fd_sc_hd__and4b_1 _1737_ (.A_N(_0657_),
    .B(_0493_),
    .C(_0496_),
    .D(\uc_0.bc_0._85_[1] ),
    .X(_0405_));
 sky130_fd_sc_hd__a211oi_1 _1738_ (.A1(_0493_),
    .A2(_0403_),
    .B1(_0404_),
    .C1(_0405_),
    .Y(_0145_));
 sky130_fd_sc_hd__a31o_1 _1739_ (.A1(_0657_),
    .A2(\uc_0.bc_0._85_[3] ),
    .A3(_0667_),
    .B1(_0660_),
    .X(_0406_));
 sky130_fd_sc_hd__o21ba_1 _1740_ (.A1(\po_0.muxf_0.s0 ),
    .A2(_0405_),
    .B1_N(_0406_),
    .X(_0146_));
 sky130_fd_sc_hd__or3_1 _1741_ (.A(_0487_),
    .B(_0657_),
    .C(_0496_),
    .X(_0407_));
 sky130_fd_sc_hd__a21bo_1 _1742_ (.A1(_0362_),
    .A2(\uc_0._01_ ),
    .B1_N(_0407_),
    .X(_0147_));
 sky130_fd_sc_hd__a2111oi_1 _1743_ (.A1(_0489_),
    .A2(_0267_),
    .B1(_0487_),
    .C1(_0688_),
    .D1(_0676_),
    .Y(_0148_));
 sky130_fd_sc_hd__or3b_4 _1744_ (.A(_0857_),
    .B(_0858_),
    .C_N(_0754_),
    .X(_0408_));
 sky130_fd_sc_hd__buf_2 _1745_ (.A(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _1746_ (.A0(_0751_),
    .A1(\po_0.regf_0.rf[11][0] ),
    .S(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_1 _1747_ (.A(_0410_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _1748_ (.A0(_0768_),
    .A1(\po_0.regf_0.rf[11][1] ),
    .S(_0409_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _1749_ (.A(_0411_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _1750_ (.A0(_0777_),
    .A1(\po_0.regf_0.rf[11][2] ),
    .S(_0409_),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_1 _1751_ (.A(_0412_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _1752_ (.A0(_0787_),
    .A1(\po_0.regf_0.rf[11][3] ),
    .S(_0409_),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_1 _1753_ (.A(_0413_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _1754_ (.A0(_0802_),
    .A1(\po_0.regf_0.rf[11][4] ),
    .S(_0408_),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _1755_ (.A(_0414_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _1756_ (.A0(_0813_),
    .A1(\po_0.regf_0.rf[11][5] ),
    .S(_0408_),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _1757_ (.A(_0415_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _1758_ (.A0(_0824_),
    .A1(\po_0.regf_0.rf[11][6] ),
    .S(_0408_),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _1759_ (.A(_0416_),
    .X(_0155_));
 sky130_fd_sc_hd__nand2_1 _1760_ (.A(_0409_),
    .B(\po_0.regf_0.rf[11][7] ),
    .Y(_0417_));
 sky130_fd_sc_hd__o21ai_1 _1761_ (.A1(_0409_),
    .A2(_0835_),
    .B1(_0417_),
    .Y(_0156_));
 sky130_fd_sc_hd__clkbuf_4 _1762_ (.A(_0666_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _1763_ (.A0(\po_0.muxf_0.rf_w_data[0] ),
    .A1(net27),
    .S(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _1764_ (.A(_0419_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _1765_ (.A0(\po_0.muxf_0.rf_w_data[1] ),
    .A1(net28),
    .S(_0418_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_1 _1766_ (.A(_0420_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _1767_ (.A0(\po_0.muxf_0.rf_w_data[2] ),
    .A1(net29),
    .S(_0418_),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _1768_ (.A(_0421_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _1769_ (.A0(\po_0.muxf_0.rf_w_data[3] ),
    .A1(net30),
    .S(_0418_),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _1770_ (.A(_0422_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _1771_ (.A0(\po_0.muxf_0.rf_w_data[4] ),
    .A1(net31),
    .S(_0418_),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _1772_ (.A(_0423_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _1773_ (.A0(\po_0.muxf_0.rf_w_data[5] ),
    .A1(net32),
    .S(_0418_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_1 _1774_ (.A(_0424_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _1775_ (.A0(\po_0.muxf_0.rf_w_data[6] ),
    .A1(net33),
    .S(_0666_),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_1 _1776_ (.A(_0425_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _1777_ (.A0(\po_0.muxf_0.rf_w_data[7] ),
    .A1(net34),
    .S(_0666_),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_1 _1778_ (.A(_0426_),
    .X(_0164_));
 sky130_fd_sc_hd__a21o_1 _1779_ (.A1(_0362_),
    .A2(net35),
    .B1(_0405_),
    .X(_0165_));
 sky130_fd_sc_hd__or3_1 _1780_ (.A(_0487_),
    .B(_0493_),
    .C(_0666_),
    .X(_0427_));
 sky130_fd_sc_hd__a21bo_1 _1781_ (.A1(_0362_),
    .A2(net36),
    .B1_N(_0427_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _1782_ (.A0(_0452_),
    .A1(\uc_0.bc_0._85_[1] ),
    .S(_0660_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_1 _1783_ (.A(_0428_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _1784_ (.A0(_0448_),
    .A1(_0464_),
    .S(_0659_),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_1 _1785_ (.A(_0429_),
    .X(_0168_));
 sky130_fd_sc_hd__a32o_1 _1786_ (.A1(_0657_),
    .A2(_0493_),
    .A3(\uc_0.bc_0._85_[3] ),
    .B1(_0361_),
    .B2(net55),
    .X(_0169_));
 sky130_fd_sc_hd__a21o_1 _1787_ (.A1(_0362_),
    .A2(net52),
    .B1(_0670_),
    .X(_0170_));
 sky130_fd_sc_hd__a211o_2 _1788_ (.A1(_0403_),
    .A2(_0667_),
    .B1(_0405_),
    .C1(_0658_),
    .X(_0430_));
 sky130_fd_sc_hd__a21o_1 _1789_ (.A1(_0362_),
    .A2(_0753_),
    .B1(_0430_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _1790_ (.A0(\po_0.regf_0.rq_addr[0] ),
    .A1(\po_0.muxf_0.rf_w_data[4] ),
    .S(_0659_),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _1791_ (.A(_0431_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _1792_ (.A0(\po_0.regf_0.rq_addr[1] ),
    .A1(\po_0.muxf_0.rf_w_data[5] ),
    .S(_0659_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _1793_ (.A(_0432_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _1794_ (.A0(\po_0.regf_0.rq_addr[2] ),
    .A1(\po_0.muxf_0.rf_w_data[6] ),
    .S(_0659_),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _1795_ (.A(_0433_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _1796_ (.A0(\po_0.regf_0.rq_addr[3] ),
    .A1(\po_0.muxf_0.rf_w_data[7] ),
    .S(_0659_),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_1 _1797_ (.A(_0434_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _1798_ (.A0(\po_0.regf_0.rp_addr[0] ),
    .A1(\uc_0.bc_0._14_[0] ),
    .S(_0670_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_1 _1799_ (.A(_0435_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _1800_ (.A0(\po_0.regf_0.rp_addr[1] ),
    .A1(\uc_0.bc_0._14_[1] ),
    .S(_0669_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _1801_ (.A(_0436_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _1802_ (.A0(\po_0.regf_0.rp_addr[2] ),
    .A1(\uc_0.bc_0._14_[2] ),
    .S(_0669_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _1803_ (.A(_0437_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _1804_ (.A0(\po_0.regf_0.rp_addr[3] ),
    .A1(\uc_0.bc_0._14_[3] ),
    .S(_0669_),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _1805_ (.A(_0438_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _1806_ (.A0(\uc_0.bc_0._14_[0] ),
    .A1(\po_0.muxf_0.rf_w_data[0] ),
    .S(_0658_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _1807_ (.A0(_0869_),
    .A1(_0439_),
    .S(_0430_),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_1 _1808_ (.A(_0440_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _1809_ (.A0(\uc_0.bc_0._14_[1] ),
    .A1(\po_0.muxf_0.rf_w_data[1] ),
    .S(_0658_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _1810_ (.A0(_0838_),
    .A1(_0441_),
    .S(_0430_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _1811_ (.A(_0442_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _1812_ (.A0(\uc_0.bc_0._14_[2] ),
    .A1(\po_0.muxf_0.rf_w_data[2] ),
    .S(_0658_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _1813_ (.A0(_0858_),
    .A1(_0443_),
    .S(_0430_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_1 _1814_ (.A(_0444_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _1815_ (.A0(\uc_0.bc_0._14_[3] ),
    .A1(\po_0.muxf_0.rf_w_data[3] ),
    .S(_0658_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _1816_ (.A0(_0754_),
    .A1(_0445_),
    .S(_0430_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _1817_ (.A(_0446_),
    .X(_0183_));
 sky130_fd_sc_hd__dfxtp_1 _1818_ (.CLK(net92),
    .D(_0016_),
    .Q(\po_0.regf_0.rf[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1819_ (.CLK(net88),
    .D(_0017_),
    .Q(\po_0.regf_0.rf[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1820_ (.CLK(net92),
    .D(_0018_),
    .Q(\po_0.regf_0.rf[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1821_ (.CLK(net88),
    .D(_0019_),
    .Q(\po_0.regf_0.rf[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1822_ (.CLK(net105),
    .D(_0020_),
    .Q(\po_0.regf_0.rf[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1823_ (.CLK(net104),
    .D(_0021_),
    .Q(\po_0.regf_0.rf[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1824_ (.CLK(net104),
    .D(_0022_),
    .Q(\po_0.regf_0.rf[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1825_ (.CLK(net92),
    .D(_0023_),
    .Q(\po_0.regf_0.rf[5][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1826_ (.D(\po_0.regf_0._5_[0] ),
    .GATE(net55),
    .Q(\po_0._1_[0] ));
 sky130_fd_sc_hd__dlxtp_1 _1827_ (.D(\po_0.regf_0._5_[1] ),
    .GATE(net54),
    .Q(\po_0._1_[1] ));
 sky130_fd_sc_hd__dlxtp_1 _1828_ (.D(\po_0.regf_0._5_[2] ),
    .GATE(net55),
    .Q(\po_0._1_[2] ));
 sky130_fd_sc_hd__dlxtp_1 _1829_ (.D(\po_0.regf_0._5_[3] ),
    .GATE(net54),
    .Q(\po_0._1_[3] ));
 sky130_fd_sc_hd__dlxtp_1 _1830_ (.D(\po_0.regf_0._5_[4] ),
    .GATE(net54),
    .Q(\po_0._1_[4] ));
 sky130_fd_sc_hd__dlxtp_1 _1831_ (.D(\po_0.regf_0._5_[5] ),
    .GATE(net54),
    .Q(\po_0._1_[5] ));
 sky130_fd_sc_hd__dlxtp_1 _1832_ (.D(\po_0.regf_0._5_[6] ),
    .GATE(net54),
    .Q(\po_0._1_[6] ));
 sky130_fd_sc_hd__dlxtp_1 _1833_ (.D(\po_0.regf_0._5_[7] ),
    .GATE(net54),
    .Q(\po_0._1_[7] ));
 sky130_fd_sc_hd__dlxtp_1 _1834_ (.D(\po_0.regf_0._3_[0] ),
    .GATE(net52),
    .Q(net19));
 sky130_fd_sc_hd__dlxtp_1 _1835_ (.D(\po_0.regf_0._3_[1] ),
    .GATE(net52),
    .Q(net20));
 sky130_fd_sc_hd__dlxtp_1 _1836_ (.D(\po_0.regf_0._3_[2] ),
    .GATE(net53),
    .Q(net21));
 sky130_fd_sc_hd__dlxtp_1 _1837_ (.D(\po_0.regf_0._3_[3] ),
    .GATE(net52),
    .Q(net22));
 sky130_fd_sc_hd__dlxtp_1 _1838_ (.D(\po_0.regf_0._3_[4] ),
    .GATE(net53),
    .Q(net23));
 sky130_fd_sc_hd__dlxtp_1 _1839_ (.D(\po_0.regf_0._3_[5] ),
    .GATE(net52),
    .Q(net24));
 sky130_fd_sc_hd__dlxtp_1 _1840_ (.D(\po_0.regf_0._3_[6] ),
    .GATE(net53),
    .Q(net25));
 sky130_fd_sc_hd__dlxtp_1 _1841_ (.D(\po_0.regf_0._3_[7] ),
    .GATE(net52),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _1842_ (.CLK(net92),
    .D(_0024_),
    .Q(\po_0.regf_0.rf[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1843_ (.CLK(net83),
    .D(_0025_),
    .Q(\po_0.regf_0.rf[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1844_ (.CLK(net85),
    .D(_0026_),
    .Q(\po_0.regf_0.rf[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1845_ (.CLK(net88),
    .D(_0027_),
    .Q(\po_0.regf_0.rf[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1846_ (.CLK(net105),
    .D(_0028_),
    .Q(\po_0.regf_0.rf[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1847_ (.CLK(net104),
    .D(_0029_),
    .Q(\po_0.regf_0.rf[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1848_ (.CLK(net104),
    .D(_0030_),
    .Q(\po_0.regf_0.rf[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1849_ (.CLK(net89),
    .D(_0031_),
    .Q(\po_0.regf_0.rf[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1850_ (.CLK(net92),
    .D(_0032_),
    .Q(\po_0.regf_0.rf[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1851_ (.CLK(net89),
    .D(_0033_),
    .Q(\po_0.regf_0.rf[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1852_ (.CLK(net95),
    .D(_0034_),
    .Q(\po_0.regf_0.rf[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1853_ (.CLK(net88),
    .D(_0035_),
    .Q(\po_0.regf_0.rf[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1854_ (.CLK(net106),
    .D(_0036_),
    .Q(\po_0.regf_0.rf[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1855_ (.CLK(net104),
    .D(_0037_),
    .Q(\po_0.regf_0.rf[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1856_ (.CLK(net104),
    .D(_0038_),
    .Q(\po_0.regf_0.rf[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1857_ (.CLK(net89),
    .D(_0039_),
    .Q(\po_0.regf_0.rf[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1858_ (.CLK(net86),
    .D(_0040_),
    .Q(\po_0.regf_0.rf[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1859_ (.CLK(net82),
    .D(_0041_),
    .Q(\po_0.regf_0.rf[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1860_ (.CLK(net86),
    .D(_0042_),
    .Q(\po_0.regf_0.rf[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1861_ (.CLK(net82),
    .D(_0043_),
    .Q(\po_0.regf_0.rf[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1862_ (.CLK(net99),
    .D(_0044_),
    .Q(\po_0.regf_0.rf[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1863_ (.CLK(net97),
    .D(_0045_),
    .Q(\po_0.regf_0.rf[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1864_ (.CLK(net97),
    .D(_0046_),
    .Q(\po_0.regf_0.rf[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1865_ (.CLK(net84),
    .D(_0047_),
    .Q(\po_0.regf_0.rf[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1866_ (.CLK(net78),
    .D(_0008_),
    .Q(_0000_));
 sky130_fd_sc_hd__dfxtp_1 _1867_ (.CLK(net78),
    .D(_0009_),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_1 _1868_ (.CLK(net78),
    .D(_0010_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_2 _1869_ (.CLK(net75),
    .D(_0011_),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_1 _1870_ (.CLK(net85),
    .D(_0048_),
    .Q(\po_0.regf_0.rf[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1871_ (.CLK(net82),
    .D(_0049_),
    .Q(\po_0.regf_0.rf[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1872_ (.CLK(net86),
    .D(_0050_),
    .Q(\po_0.regf_0.rf[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1873_ (.CLK(net83),
    .D(_0051_),
    .Q(\po_0.regf_0.rf[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1874_ (.CLK(net100),
    .D(_0052_),
    .Q(\po_0.regf_0.rf[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1875_ (.CLK(net98),
    .D(_0053_),
    .Q(\po_0.regf_0.rf[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1876_ (.CLK(net98),
    .D(_0054_),
    .Q(\po_0.regf_0.rf[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1877_ (.CLK(net83),
    .D(_0055_),
    .Q(\po_0.regf_0.rf[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1878_ (.CLK(net68),
    .D(_0056_),
    .Q(\po_0.regf_0.rf[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1879_ (.CLK(net65),
    .D(_0057_),
    .Q(\po_0.regf_0.rf[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1880_ (.CLK(net68),
    .D(_0058_),
    .Q(\po_0.regf_0.rf[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1881_ (.CLK(net65),
    .D(_0059_),
    .Q(\po_0.regf_0.rf[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1882_ (.CLK(net99),
    .D(_0060_),
    .Q(\po_0.regf_0.rf[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1883_ (.CLK(net97),
    .D(_0061_),
    .Q(\po_0.regf_0.rf[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1884_ (.CLK(net97),
    .D(_0062_),
    .Q(\po_0.regf_0.rf[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1885_ (.CLK(net65),
    .D(_0063_),
    .Q(\po_0.regf_0.rf[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1886_ (.CLK(net93),
    .D(_0064_),
    .Q(\po_0.regf_0.rf[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1887_ (.CLK(net90),
    .D(_0065_),
    .Q(\po_0.regf_0.rf[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1888_ (.CLK(net93),
    .D(_0066_),
    .Q(\po_0.regf_0.rf[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1889_ (.CLK(net90),
    .D(_0067_),
    .Q(\po_0.regf_0.rf[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1890_ (.CLK(net105),
    .D(_0068_),
    .Q(\po_0.regf_0.rf[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1891_ (.CLK(net103),
    .D(_0069_),
    .Q(\po_0.regf_0.rf[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1892_ (.CLK(net102),
    .D(_0070_),
    .Q(\po_0.regf_0.rf[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1893_ (.CLK(net90),
    .D(_0071_),
    .Q(\po_0.regf_0.rf[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1894_ (.CLK(net92),
    .D(_0072_),
    .Q(\po_0.regf_0.rf[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1895_ (.CLK(net90),
    .D(_0073_),
    .Q(\po_0.regf_0.rf[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1896_ (.CLK(net95),
    .D(_0074_),
    .Q(\po_0.regf_0.rf[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1897_ (.CLK(net88),
    .D(_0075_),
    .Q(\po_0.regf_0.rf[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1898_ (.CLK(net105),
    .D(_0076_),
    .Q(\po_0.regf_0.rf[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1899_ (.CLK(net103),
    .D(_0077_),
    .Q(\po_0.regf_0.rf[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1900_ (.CLK(net102),
    .D(_0078_),
    .Q(\po_0.regf_0.rf[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1901_ (.CLK(net89),
    .D(_0079_),
    .Q(\po_0.regf_0.rf[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1902_ (.CLK(net93),
    .D(_0080_),
    .Q(\po_0.regf_0.rf[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1903_ (.CLK(net91),
    .D(_0081_),
    .Q(\po_0.regf_0.rf[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1904_ (.CLK(net93),
    .D(_0082_),
    .Q(\po_0.regf_0.rf[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1905_ (.CLK(net90),
    .D(_0083_),
    .Q(\po_0.regf_0.rf[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1906_ (.CLK(net105),
    .D(_0084_),
    .Q(\po_0.regf_0.rf[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1907_ (.CLK(net103),
    .D(_0085_),
    .Q(\po_0.regf_0.rf[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1908_ (.CLK(net102),
    .D(_0086_),
    .Q(\po_0.regf_0.rf[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1909_ (.CLK(net93),
    .D(_0087_),
    .Q(\po_0.regf_0.rf[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1910_ (.CLK(net93),
    .D(_0088_),
    .Q(\po_0.regf_0.rf[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1911_ (.CLK(net90),
    .D(_0089_),
    .Q(\po_0.regf_0.rf[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1912_ (.CLK(net94),
    .D(_0090_),
    .Q(\po_0.regf_0.rf[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1913_ (.CLK(net88),
    .D(_0091_),
    .Q(\po_0.regf_0.rf[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1914_ (.CLK(net105),
    .D(_0092_),
    .Q(\po_0.regf_0.rf[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1915_ (.CLK(net103),
    .D(_0093_),
    .Q(\po_0.regf_0.rf[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1916_ (.CLK(net102),
    .D(_0094_),
    .Q(\po_0.regf_0.rf[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1917_ (.CLK(net89),
    .D(_0095_),
    .Q(\po_0.regf_0.rf[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1918_ (.CLK(net73),
    .D(_0096_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_2 _1919_ (.CLK(net73),
    .D(_0097_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _1920_ (.CLK(net71),
    .D(_0098_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_2 _1921_ (.CLK(net71),
    .D(_0099_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _1922_ (.CLK(net72),
    .D(_0100_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _1923_ (.CLK(net71),
    .D(_0101_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_2 _1924_ (.CLK(net71),
    .D(_0102_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_2 _1925_ (.CLK(net71),
    .D(_0103_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _1926_ (.CLK(net85),
    .D(_0104_),
    .Q(\po_0.regf_0.rf[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1927_ (.CLK(net83),
    .D(_0105_),
    .Q(\po_0.regf_0.rf[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1928_ (.CLK(net85),
    .D(_0106_),
    .Q(\po_0.regf_0.rf[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1929_ (.CLK(net83),
    .D(_0107_),
    .Q(\po_0.regf_0.rf[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1930_ (.CLK(net100),
    .D(_0108_),
    .Q(\po_0.regf_0.rf[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1931_ (.CLK(net98),
    .D(_0109_),
    .Q(\po_0.regf_0.rf[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1932_ (.CLK(net98),
    .D(_0110_),
    .Q(\po_0.regf_0.rf[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1933_ (.CLK(net85),
    .D(_0111_),
    .Q(\po_0.regf_0.rf[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1934_ (.CLK(net71),
    .D(net9),
    .Q(\uc_0._21_[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1935_ (.CLK(net103),
    .D(net10),
    .Q(\uc_0._21_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1936_ (.CLK(net80),
    .D(net11),
    .Q(\uc_0._21_[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1937_ (.CLK(net64),
    .D(net12),
    .Q(\uc_0._21_[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1938_ (.CLK(net64),
    .D(net13),
    .Q(\uc_0._21_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1939_ (.CLK(net64),
    .D(net14),
    .Q(\uc_0._21_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1940_ (.CLK(net64),
    .D(net15),
    .Q(\uc_0._21_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1941_ (.CLK(net63),
    .D(net16),
    .Q(\uc_0._21_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1942_ (.CLK(net72),
    .D(_0112_),
    .Q(\uc_0._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _1943_ (.CLK(net74),
    .D(_0012_),
    .Q(_0004_));
 sky130_fd_sc_hd__dfxtp_1 _1944_ (.CLK(net75),
    .D(_0013_),
    .Q(_0005_));
 sky130_fd_sc_hd__dfxtp_1 _1945_ (.CLK(net75),
    .D(_0014_),
    .Q(_0006_));
 sky130_fd_sc_hd__dfxtp_2 _1946_ (.CLK(net69),
    .D(_0015_),
    .Q(_0007_));
 sky130_fd_sc_hd__dfxtp_1 _1947_ (.CLK(net68),
    .D(_0113_),
    .Q(\po_0.regf_0.rf[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1948_ (.CLK(net67),
    .D(_0114_),
    .Q(\po_0.regf_0.rf[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1949_ (.CLK(net69),
    .D(_0115_),
    .Q(\po_0.regf_0.rf[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1950_ (.CLK(net67),
    .D(_0116_),
    .Q(\po_0.regf_0.rf[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1951_ (.CLK(net78),
    .D(_0117_),
    .Q(\po_0.regf_0.rf[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1952_ (.CLK(net76),
    .D(_0118_),
    .Q(\po_0.regf_0.rf[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1953_ (.CLK(net75),
    .D(_0119_),
    .Q(\po_0.regf_0.rf[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1954_ (.CLK(net66),
    .D(_0120_),
    .Q(\po_0.regf_0.rf[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1955_ (.CLK(net86),
    .D(_0121_),
    .Q(\po_0.regf_0.rf[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1956_ (.CLK(net82),
    .D(_0122_),
    .Q(\po_0.regf_0.rf[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1957_ (.CLK(net86),
    .D(_0123_),
    .Q(\po_0.regf_0.rf[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1958_ (.CLK(net82),
    .D(_0124_),
    .Q(\po_0.regf_0.rf[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1959_ (.CLK(net99),
    .D(_0125_),
    .Q(\po_0.regf_0.rf[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1960_ (.CLK(net97),
    .D(_0126_),
    .Q(\po_0.regf_0.rf[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1961_ (.CLK(net97),
    .D(_0127_),
    .Q(\po_0.regf_0.rf[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1962_ (.CLK(net84),
    .D(_0128_),
    .Q(\po_0.regf_0.rf[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1963_ (.CLK(net68),
    .D(_0129_),
    .Q(\po_0.regf_0.rf[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1964_ (.CLK(net65),
    .D(_0130_),
    .Q(\po_0.regf_0.rf[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1965_ (.CLK(net68),
    .D(_0131_),
    .Q(\po_0.regf_0.rf[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1966_ (.CLK(net65),
    .D(_0132_),
    .Q(\po_0.regf_0.rf[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1967_ (.CLK(net76),
    .D(_0133_),
    .Q(\po_0.regf_0.rf[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1968_ (.CLK(net76),
    .D(_0134_),
    .Q(\po_0.regf_0.rf[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1969_ (.CLK(net75),
    .D(_0135_),
    .Q(\po_0.regf_0.rf[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1970_ (.CLK(net66),
    .D(_0136_),
    .Q(\po_0.regf_0.rf[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1971_ (.CLK(net68),
    .D(_0137_),
    .Q(\po_0.regf_0.rf[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1972_ (.CLK(net66),
    .D(_0138_),
    .Q(\po_0.regf_0.rf[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1973_ (.CLK(net69),
    .D(_0139_),
    .Q(\po_0.regf_0.rf[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1974_ (.CLK(net65),
    .D(_0140_),
    .Q(\po_0.regf_0.rf[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1975_ (.CLK(net78),
    .D(_0141_),
    .Q(\po_0.regf_0.rf[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1976_ (.CLK(net76),
    .D(_0142_),
    .Q(\po_0.regf_0.rf[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1977_ (.CLK(net75),
    .D(_0143_),
    .Q(\po_0.regf_0.rf[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1978_ (.CLK(net66),
    .D(_0144_),
    .Q(\po_0.regf_0.rf[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1979_ (.CLK(net74),
    .D(_0145_),
    .Q(\po_0.muxf_0.s1 ));
 sky130_fd_sc_hd__dfxtp_1 _1980_ (.CLK(net74),
    .D(_0146_),
    .Q(\po_0.muxf_0.s0 ));
 sky130_fd_sc_hd__dfxtp_1 _1981_ (.CLK(net63),
    .D(\uc_0.bc_0._85_[0] ),
    .Q(\uc_0.bc_0._12_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1982_ (.CLK(net63),
    .D(\uc_0.bc_0._85_[1] ),
    .Q(\uc_0.bc_0._12_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1983_ (.CLK(net72),
    .D(\uc_0.bc_0._85_[2] ),
    .Q(\uc_0.bc_0._12_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1984_ (.CLK(net63),
    .D(\uc_0.bc_0._85_[3] ),
    .Q(\uc_0.bc_0._12_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1985_ (.CLK(net72),
    .D(_0147_),
    .Q(\uc_0._01_ ));
 sky130_fd_sc_hd__dfxtp_1 _1986_ (.CLK(net72),
    .D(_0148_),
    .Q(\uc_0._02_ ));
 sky130_fd_sc_hd__dfxtp_1 _1987_ (.CLK(net85),
    .D(_0149_),
    .Q(\po_0.regf_0.rf[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1988_ (.CLK(net82),
    .D(_0150_),
    .Q(\po_0.regf_0.rf[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1989_ (.CLK(net87),
    .D(_0151_),
    .Q(\po_0.regf_0.rf[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1990_ (.CLK(net83),
    .D(_0152_),
    .Q(\po_0.regf_0.rf[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1991_ (.CLK(net100),
    .D(_0153_),
    .Q(\po_0.regf_0.rf[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1992_ (.CLK(net98),
    .D(_0154_),
    .Q(\po_0.regf_0.rf[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1993_ (.CLK(net98),
    .D(_0155_),
    .Q(\po_0.regf_0.rf[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1994_ (.CLK(net84),
    .D(_0156_),
    .Q(\po_0.regf_0.rf[11][7] ));
 sky130_fd_sc_hd__dlxtn_1 _1995_ (.D(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[0] ),
    .GATE_N(net61),
    .Q(\po_0.muxf_0.rf_w_data[0] ));
 sky130_fd_sc_hd__dlxtn_2 _1996_ (.D(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[1] ),
    .GATE_N(net61),
    .Q(\po_0.muxf_0.rf_w_data[1] ));
 sky130_fd_sc_hd__dlxtn_2 _1997_ (.D(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[2] ),
    .GATE_N(net61),
    .Q(\po_0.muxf_0.rf_w_data[2] ));
 sky130_fd_sc_hd__dlxtn_2 _1998_ (.D(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[3] ),
    .GATE_N(net61),
    .Q(\po_0.muxf_0.rf_w_data[3] ));
 sky130_fd_sc_hd__dlxtn_2 _1999_ (.D(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[4] ),
    .GATE_N(net59),
    .Q(\po_0.muxf_0.rf_w_data[4] ));
 sky130_fd_sc_hd__dlxtn_2 _2000_ (.D(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[5] ),
    .GATE_N(net58),
    .Q(\po_0.muxf_0.rf_w_data[5] ));
 sky130_fd_sc_hd__dlxtn_1 _2001_ (.D(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[6] ),
    .GATE_N(net59),
    .Q(\po_0.muxf_0.rf_w_data[6] ));
 sky130_fd_sc_hd__dlxtn_1 _2002_ (.D(\uc_0.bc_0.359$func$/openlane/designs/vahid6i/src/vahid6i.v:987$36.$result[7] ),
    .GATE_N(net58),
    .Q(\po_0.muxf_0.rf_w_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2003_ (.CLK(net80),
    .D(_0157_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _2004_ (.CLK(net106),
    .D(_0158_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _2005_ (.CLK(net94),
    .D(_0159_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _2006_ (.CLK(net94),
    .D(_0160_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _2007_ (.CLK(net102),
    .D(_0161_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _2008_ (.CLK(net102),
    .D(_0162_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _2009_ (.CLK(net74),
    .D(_0163_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _2010_ (.CLK(net63),
    .D(_0164_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _2011_ (.CLK(net80),
    .D(_0165_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _2012_ (.CLK(net79),
    .D(_0166_),
    .Q(net36));
 sky130_fd_sc_hd__dlxtn_1 _2013_ (.D(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[0] ),
    .GATE_N(net62),
    .Q(\uc_0.bc_0._14_[0] ));
 sky130_fd_sc_hd__dlxtn_1 _2014_ (.D(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[1] ),
    .GATE_N(net61),
    .Q(\uc_0.bc_0._14_[1] ));
 sky130_fd_sc_hd__dlxtn_1 _2015_ (.D(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[2] ),
    .GATE_N(net62),
    .Q(\uc_0.bc_0._14_[2] ));
 sky130_fd_sc_hd__dlxtn_1 _2016_ (.D(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[3] ),
    .GATE_N(net61),
    .Q(\uc_0.bc_0._14_[3] ));
 sky130_fd_sc_hd__dlxtn_1 _2017_ (.D(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[4] ),
    .GATE_N(net59),
    .Q(\uc_0.bc_0._14_[4] ));
 sky130_fd_sc_hd__dlxtn_1 _2018_ (.D(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[5] ),
    .GATE_N(net59),
    .Q(\uc_0.bc_0._14_[5] ));
 sky130_fd_sc_hd__dlxtn_1 _2019_ (.D(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[6] ),
    .GATE_N(net58),
    .Q(\uc_0.bc_0._14_[6] ));
 sky130_fd_sc_hd__dlxtn_1 _2020_ (.D(\uc_0.bc_0.358$func$/openlane/designs/vahid6i/src/vahid6i.v:960$35.$result[7] ),
    .GATE_N(net58),
    .Q(\uc_0.bc_0._14_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2021_ (.CLK(net70),
    .D(_0167_),
    .Q(\po_0.alu_0.s1 ));
 sky130_fd_sc_hd__dfxtp_1 _2022_ (.CLK(net63),
    .D(_0168_),
    .Q(\po_0.alu_0.s0 ));
 sky130_fd_sc_hd__dfxtp_1 _2023_ (.CLK(net72),
    .D(_0169_),
    .Q(\po_0.regf_0.rq_rd ));
 sky130_fd_sc_hd__dfxtp_1 _2024_ (.CLK(net77),
    .D(_0170_),
    .Q(\po_0.regf_0.rp_rd ));
 sky130_fd_sc_hd__dfxtp_1 _2025_ (.CLK(net99),
    .D(_0171_),
    .Q(\po_0.regf_0.w_wr ));
 sky130_fd_sc_hd__dfxtp_1 _2026_ (.CLK(net74),
    .D(_0172_),
    .Q(\po_0.regf_0.rq_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2027_ (.CLK(net69),
    .D(_0173_),
    .Q(\po_0.regf_0.rq_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2028_ (.CLK(net74),
    .D(_0174_),
    .Q(\po_0.regf_0.rq_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2029_ (.CLK(net64),
    .D(_0175_),
    .Q(\po_0.regf_0.rq_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2030_ (.CLK(net79),
    .D(_0176_),
    .Q(\po_0.regf_0.rp_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2031_ (.CLK(net78),
    .D(_0177_),
    .Q(\po_0.regf_0.rp_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2032_ (.CLK(net79),
    .D(_0178_),
    .Q(\po_0.regf_0.rp_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2033_ (.CLK(net77),
    .D(_0179_),
    .Q(\po_0.regf_0.rp_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2034_ (.CLK(net99),
    .D(_0180_),
    .Q(\po_0.regf_0.w_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2035_ (.CLK(net79),
    .D(_0181_),
    .Q(\po_0.regf_0.w_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2036_ (.CLK(net100),
    .D(_0182_),
    .Q(\po_0.regf_0.w_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2037_ (.CLK(net99),
    .D(_0183_),
    .Q(\po_0.regf_0.w_addr[3] ));
 sky130_fd_sc_hd__clkbuf_1 _2039_ (.A(net91),
    .X(net45));
 sky130_fd_sc_hd__ebufn_1 _2040_ (.A(\po_0.alu_0._10_[0] ),
    .TE_B(_0881_),
    .Z(\po_0.alu_0._11_[0] ));
 sky130_fd_sc_hd__ebufn_1 _2041_ (.A(\po_0.alu_0._10_[1] ),
    .TE_B(_0882_),
    .Z(\po_0.alu_0._11_[1] ));
 sky130_fd_sc_hd__ebufn_1 _2042_ (.A(\po_0.alu_0._10_[2] ),
    .TE_B(_0883_),
    .Z(\po_0.alu_0._11_[2] ));
 sky130_fd_sc_hd__ebufn_1 _2043_ (.A(\po_0.alu_0._10_[3] ),
    .TE_B(_0884_),
    .Z(\po_0.alu_0._11_[3] ));
 sky130_fd_sc_hd__ebufn_1 _2044_ (.A(\po_0.alu_0._10_[4] ),
    .TE_B(_0885_),
    .Z(\po_0.alu_0._11_[4] ));
 sky130_fd_sc_hd__ebufn_1 _2045_ (.A(\po_0.alu_0._10_[5] ),
    .TE_B(_0886_),
    .Z(\po_0.alu_0._11_[5] ));
 sky130_fd_sc_hd__ebufn_1 _2046_ (.A(\po_0.alu_0._10_[6] ),
    .TE_B(_0887_),
    .Z(\po_0.alu_0._11_[6] ));
 sky130_fd_sc_hd__ebufn_1 _2047_ (.A(\po_0.alu_0._10_[7] ),
    .TE_B(_0888_),
    .Z(\po_0.alu_0._11_[7] ));
 sky130_fd_sc_hd__clkbuf_1 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout101 (.A(net108),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(net107),
    .X(net102));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout103 (.A(net107),
    .X(net103));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout104 (.A(net107),
    .X(net104));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 fanout109 (.A(net17),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(net23),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout51 (.A(net22),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(\po_0.regf_0.rp_rd ),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 fanout53 (.A(\po_0.regf_0.rp_rd ),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout54 (.A(\po_0.regf_0.rq_rd ),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 fanout55 (.A(\po_0.regf_0.rq_rd ),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 fanout56 (.A(net42),
    .X(net56));
 sky130_fd_sc_hd__buf_2 fanout57 (.A(net39),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout58 (.A(net60),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout60 (.A(net18),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 fanout62 (.A(net18),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 fanout63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 fanout64 (.A(net70),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(net67),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout67 (.A(net70),
    .X(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout70 (.A(net109),
    .X(net70));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout71 (.A(net73),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 fanout72 (.A(net81),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 fanout73 (.A(net81),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 fanout74 (.A(net77),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(net77),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout77 (.A(net81),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 fanout78 (.A(net80),
    .X(net78));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 fanout81 (.A(net109),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 fanout82 (.A(net84),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout84 (.A(net87),
    .X(net84));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 fanout87 (.A(net96),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout88 (.A(net91),
    .X(net88));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout91 (.A(net96),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 fanout92 (.A(net95),
    .X(net92));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout93 (.A(net95),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout96 (.A(net108),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 fanout97 (.A(net101),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 fanout98 (.A(net101),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 fanout99 (.A(net101),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(D_R_data[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(I_data[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(I_data[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(I_data[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(I_data[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(I_data[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(I_data[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(I_data[7]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(clock),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(reset),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(D_R_data[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(D_R_data[2]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(D_R_data[3]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(D_R_data[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(D_R_data[5]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(D_R_data[6]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(D_R_data[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(I_data[0]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(D_W_data[0]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(D_W_data[1]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(D_W_data[2]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(D_W_data[3]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(D_W_data[4]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(D_W_data[5]));
 sky130_fd_sc_hd__clkbuf_4 output25 (.A(net25),
    .X(D_W_data[6]));
 sky130_fd_sc_hd__clkbuf_4 output26 (.A(net26),
    .X(D_W_data[7]));
 sky130_fd_sc_hd__clkbuf_4 output27 (.A(net27),
    .X(D_addr[0]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(D_addr[1]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(D_addr[2]));
 sky130_fd_sc_hd__clkbuf_4 output30 (.A(net30),
    .X(D_addr[3]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(D_addr[4]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(D_addr[5]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(D_addr[6]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(D_addr[7]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(D_rd));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(D_wr));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net37),
    .X(I_addr[0]));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net38),
    .X(I_addr[1]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net57),
    .X(I_addr[2]));
 sky130_fd_sc_hd__clkbuf_4 output40 (.A(net40),
    .X(I_addr[3]));
 sky130_fd_sc_hd__clkbuf_4 output41 (.A(net41),
    .X(I_addr[4]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(I_addr[5]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(I_addr[6]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(I_addr[7]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(led_clock));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(leds[0]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(leds[1]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(leds[2]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(leds[3]));
 sky130_fd_sc_hd__conb_1 vahid6i_110 (.HI(net110));
 assign I_rd = net110;
endmodule
