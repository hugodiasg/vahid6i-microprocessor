magic
tech sky130A
magscale 1 2
timestamp 1680791366
<< viali >>
rect 1777 37417 1811 37451
rect 22569 37417 22603 37451
rect 31769 37349 31803 37383
rect 4629 37281 4663 37315
rect 17693 37281 17727 37315
rect 19257 37281 19291 37315
rect 28457 37281 28491 37315
rect 1685 37213 1719 37247
rect 4905 37213 4939 37247
rect 7205 37213 7239 37247
rect 10425 37213 10459 37247
rect 13645 37213 13679 37247
rect 16221 37213 16255 37247
rect 17969 37213 18003 37247
rect 19533 37213 19567 37247
rect 20361 37213 20395 37247
rect 22753 37213 22787 37247
rect 25881 37213 25915 37247
rect 28733 37213 28767 37247
rect 35081 37213 35115 37247
rect 36185 37213 36219 37247
rect 2237 37145 2271 37179
rect 22477 37145 22511 37179
rect 31585 37145 31619 37179
rect 35909 37145 35943 37179
rect 2329 37077 2363 37111
rect 7389 37077 7423 37111
rect 10609 37077 10643 37111
rect 13829 37077 13863 37111
rect 16405 37077 16439 37111
rect 20177 37077 20211 37111
rect 22937 37077 22971 37111
rect 26065 37077 26099 37111
rect 34897 37077 34931 37111
rect 36369 37077 36403 37111
rect 6837 36873 6871 36907
rect 17141 36873 17175 36907
rect 18981 36873 19015 36907
rect 20637 36873 20671 36907
rect 22293 36873 22327 36907
rect 17662 36805 17696 36839
rect 19502 36805 19536 36839
rect 22998 36805 23032 36839
rect 30113 36805 30147 36839
rect 7021 36737 7055 36771
rect 7113 36737 7147 36771
rect 16497 36737 16531 36771
rect 17325 36737 17359 36771
rect 19165 36737 19199 36771
rect 21649 36737 21683 36771
rect 22201 36737 22235 36771
rect 22753 36737 22787 36771
rect 7389 36669 7423 36703
rect 17417 36669 17451 36703
rect 19257 36669 19291 36703
rect 22477 36669 22511 36703
rect 21833 36601 21867 36635
rect 30297 36601 30331 36635
rect 16313 36533 16347 36567
rect 18797 36533 18831 36567
rect 21465 36533 21499 36567
rect 24133 36533 24167 36567
rect 17233 36329 17267 36363
rect 17969 36329 18003 36363
rect 19533 36329 19567 36363
rect 22661 36329 22695 36363
rect 18613 36193 18647 36227
rect 19993 36193 20027 36227
rect 20085 36193 20119 36227
rect 21281 36193 21315 36227
rect 30205 36193 30239 36227
rect 31125 36193 31159 36227
rect 5825 36125 5859 36159
rect 15853 36125 15887 36159
rect 16120 36125 16154 36159
rect 17693 36125 17727 36159
rect 18337 36125 18371 36159
rect 21548 36125 21582 36159
rect 29929 36125 29963 36159
rect 30849 36125 30883 36159
rect 6092 36057 6126 36091
rect 7205 35989 7239 36023
rect 17509 35989 17543 36023
rect 18429 35989 18463 36023
rect 19901 35989 19935 36023
rect 6377 35785 6411 35819
rect 16681 35785 16715 35819
rect 17141 35785 17175 35819
rect 29377 35785 29411 35819
rect 31033 35785 31067 35819
rect 29898 35717 29932 35751
rect 6561 35649 6595 35683
rect 17049 35649 17083 35683
rect 19441 35649 19475 35683
rect 19708 35649 19742 35683
rect 29285 35649 29319 35683
rect 29561 35649 29595 35683
rect 17325 35581 17359 35615
rect 29653 35581 29687 35615
rect 20821 35445 20855 35479
rect 29101 35445 29135 35479
rect 6193 35241 6227 35275
rect 9045 35241 9079 35275
rect 19717 35241 19751 35275
rect 29745 35241 29779 35275
rect 6745 35105 6779 35139
rect 9229 35105 9263 35139
rect 9689 35105 9723 35139
rect 14657 35105 14691 35139
rect 20637 35105 20671 35139
rect 25053 35105 25087 35139
rect 30205 35105 30239 35139
rect 30297 35105 30331 35139
rect 1409 35037 1443 35071
rect 6653 35037 6687 35071
rect 8953 35037 8987 35071
rect 9597 35037 9631 35071
rect 9781 35037 9815 35071
rect 17233 35037 17267 35071
rect 19901 35037 19935 35071
rect 20453 35037 20487 35071
rect 21097 35037 21131 35071
rect 21189 35037 21223 35071
rect 22845 35037 22879 35071
rect 24593 35037 24627 35071
rect 24961 35037 24995 35071
rect 6561 34969 6595 35003
rect 14473 34969 14507 35003
rect 17478 34969 17512 35003
rect 21434 34969 21468 35003
rect 23112 34969 23146 35003
rect 25298 34969 25332 35003
rect 1593 34901 1627 34935
rect 9229 34901 9263 34935
rect 14105 34901 14139 34935
rect 14565 34901 14599 34935
rect 18613 34901 18647 34935
rect 19993 34901 20027 34935
rect 20361 34901 20395 34935
rect 20913 34901 20947 34935
rect 22569 34901 22603 34935
rect 24225 34901 24259 34935
rect 24409 34901 24443 34935
rect 24777 34901 24811 34935
rect 26433 34901 26467 34935
rect 30113 34901 30147 34935
rect 5181 34697 5215 34731
rect 5733 34697 5767 34731
rect 6653 34697 6687 34731
rect 9873 34697 9907 34731
rect 11345 34697 11379 34731
rect 14841 34697 14875 34731
rect 16681 34697 16715 34731
rect 17049 34697 17083 34731
rect 18245 34697 18279 34731
rect 19993 34697 20027 34731
rect 21833 34697 21867 34731
rect 23857 34697 23891 34731
rect 24317 34697 24351 34731
rect 26065 34697 26099 34731
rect 7174 34629 7208 34663
rect 8760 34629 8794 34663
rect 15384 34629 15418 34663
rect 18705 34629 18739 34663
rect 22201 34629 22235 34663
rect 4068 34561 4102 34595
rect 5641 34561 5675 34595
rect 6837 34561 6871 34595
rect 8493 34561 8527 34595
rect 9965 34561 9999 34595
rect 10232 34561 10266 34595
rect 11529 34561 11563 34595
rect 11713 34561 11747 34595
rect 11897 34561 11931 34595
rect 12164 34561 12198 34595
rect 13461 34561 13495 34595
rect 13728 34561 13762 34595
rect 15117 34561 15151 34595
rect 16865 34561 16899 34595
rect 17233 34561 17267 34595
rect 18613 34561 18647 34595
rect 19073 34561 19107 34595
rect 19809 34561 19843 34595
rect 24225 34561 24259 34595
rect 26433 34561 26467 34595
rect 3801 34493 3835 34527
rect 5917 34493 5951 34527
rect 6929 34493 6963 34527
rect 17325 34493 17359 34527
rect 17601 34493 17635 34527
rect 18797 34493 18831 34527
rect 22293 34493 22327 34527
rect 22477 34493 22511 34527
rect 24501 34493 24535 34527
rect 25145 34493 25179 34527
rect 25421 34493 25455 34527
rect 26525 34493 26559 34527
rect 26709 34493 26743 34527
rect 5273 34425 5307 34459
rect 19257 34425 19291 34459
rect 8309 34357 8343 34391
rect 11621 34357 11655 34391
rect 13277 34357 13311 34391
rect 16497 34357 16531 34391
rect 4261 34153 4295 34187
rect 7113 34153 7147 34187
rect 9137 34153 9171 34187
rect 10425 34153 10459 34187
rect 12265 34153 12299 34187
rect 13645 34153 13679 34187
rect 16221 34153 16255 34187
rect 10333 34085 10367 34119
rect 12541 34085 12575 34119
rect 4813 34017 4847 34051
rect 6929 34017 6963 34051
rect 7573 34017 7607 34051
rect 7757 34017 7791 34051
rect 10517 34017 10551 34051
rect 13001 34017 13035 34051
rect 13185 34017 13219 34051
rect 16681 34017 16715 34051
rect 16865 34017 16899 34051
rect 4445 33949 4479 33983
rect 6653 33949 6687 33983
rect 10241 33949 10275 33983
rect 12449 33949 12483 33983
rect 12909 33949 12943 33983
rect 13829 33949 13863 33983
rect 14105 33949 14139 33983
rect 5080 33881 5114 33915
rect 6745 33881 6779 33915
rect 9045 33881 9079 33915
rect 14372 33881 14406 33915
rect 16589 33881 16623 33915
rect 6193 33813 6227 33847
rect 6285 33813 6319 33847
rect 7481 33813 7515 33847
rect 15485 33813 15519 33847
rect 5181 33609 5215 33643
rect 14289 33609 14323 33643
rect 17141 33609 17175 33643
rect 26525 33609 26559 33643
rect 17662 33541 17696 33575
rect 27230 33541 27264 33575
rect 5365 33473 5399 33507
rect 14473 33473 14507 33507
rect 17325 33473 17359 33507
rect 17417 33473 17451 33507
rect 19421 33473 19455 33507
rect 21925 33473 21959 33507
rect 22192 33473 22226 33507
rect 24041 33473 24075 33507
rect 26709 33473 26743 33507
rect 36185 33473 36219 33507
rect 19165 33405 19199 33439
rect 24133 33405 24167 33439
rect 24317 33405 24351 33439
rect 26985 33405 27019 33439
rect 36369 33337 36403 33371
rect 18797 33269 18831 33303
rect 20545 33269 20579 33303
rect 23305 33269 23339 33303
rect 23673 33269 23707 33303
rect 28365 33269 28399 33303
rect 3065 33065 3099 33099
rect 14289 33065 14323 33099
rect 17509 33065 17543 33099
rect 18889 33065 18923 33099
rect 23949 33065 23983 33099
rect 26433 33065 26467 33099
rect 19349 32997 19383 33031
rect 3801 32929 3835 32963
rect 6653 32929 6687 32963
rect 7297 32929 7331 32963
rect 7573 32929 7607 32963
rect 7849 32929 7883 32963
rect 10701 32929 10735 32963
rect 11253 32929 11287 32963
rect 14841 32929 14875 32963
rect 18061 32929 18095 32963
rect 19993 32929 20027 32963
rect 20177 32929 20211 32963
rect 20821 32929 20855 32963
rect 21214 32929 21248 32963
rect 22109 32929 22143 32963
rect 22293 32929 22327 32963
rect 22753 32929 22787 32963
rect 23146 32929 23180 32963
rect 23305 32929 23339 32963
rect 24685 32929 24719 32963
rect 25145 32929 25179 32963
rect 26893 32929 26927 32963
rect 27077 32929 27111 32963
rect 1685 32861 1719 32895
rect 3617 32861 3651 32895
rect 6837 32861 6871 32895
rect 7690 32861 7724 32895
rect 10057 32861 10091 32895
rect 10241 32861 10275 32895
rect 10977 32861 11011 32895
rect 11094 32861 11128 32895
rect 12449 32861 12483 32895
rect 14657 32861 14691 32895
rect 15485 32861 15519 32895
rect 17877 32861 17911 32895
rect 19073 32861 19107 32895
rect 19717 32861 19751 32895
rect 20361 32861 20395 32895
rect 21097 32861 21131 32895
rect 21373 32861 21407 32895
rect 23029 32861 23063 32895
rect 24225 32861 24259 32895
rect 24501 32861 24535 32895
rect 25421 32861 25455 32895
rect 25538 32861 25572 32895
rect 25697 32861 25731 32895
rect 26801 32861 26835 32895
rect 1952 32793 1986 32827
rect 4046 32793 4080 32827
rect 14749 32793 14783 32827
rect 15752 32793 15786 32827
rect 3433 32725 3467 32759
rect 5181 32725 5215 32759
rect 8493 32725 8527 32759
rect 11897 32725 11931 32759
rect 12265 32725 12299 32759
rect 16865 32725 16899 32759
rect 17969 32725 18003 32759
rect 19809 32725 19843 32759
rect 22017 32725 22051 32759
rect 24041 32725 24075 32759
rect 26341 32725 26375 32759
rect 1961 32521 1995 32555
rect 2697 32521 2731 32555
rect 3893 32521 3927 32555
rect 4261 32521 4295 32555
rect 16129 32521 16163 32555
rect 19441 32521 19475 32555
rect 22385 32521 22419 32555
rect 22845 32521 22879 32555
rect 27721 32521 27755 32555
rect 2789 32453 2823 32487
rect 4353 32453 4387 32487
rect 12164 32453 12198 32487
rect 16221 32453 16255 32487
rect 18889 32453 18923 32487
rect 23388 32453 23422 32487
rect 28242 32453 28276 32487
rect 1409 32385 1443 32419
rect 2145 32385 2179 32419
rect 6469 32385 6503 32419
rect 6653 32385 6687 32419
rect 7527 32385 7561 32419
rect 8657 32385 8691 32419
rect 9873 32385 9907 32419
rect 11897 32385 11931 32419
rect 13921 32385 13955 32419
rect 14774 32385 14808 32419
rect 17049 32385 17083 32419
rect 17233 32385 17267 32419
rect 17969 32385 18003 32419
rect 19257 32385 19291 32419
rect 19625 32385 19659 32419
rect 22477 32385 22511 32419
rect 23029 32385 23063 32419
rect 24593 32385 24627 32419
rect 24777 32385 24811 32419
rect 25630 32385 25664 32419
rect 27905 32385 27939 32419
rect 2973 32317 3007 32351
rect 4537 32317 4571 32351
rect 7389 32317 7423 32351
rect 7665 32317 7699 32351
rect 8401 32317 8435 32351
rect 10149 32317 10183 32351
rect 13737 32317 13771 32351
rect 14657 32317 14691 32351
rect 14933 32317 14967 32351
rect 16405 32317 16439 32351
rect 18086 32317 18120 32351
rect 18245 32317 18279 32351
rect 22661 32317 22695 32351
rect 23121 32317 23155 32351
rect 25513 32317 25547 32351
rect 25789 32317 25823 32351
rect 27997 32317 28031 32351
rect 2329 32249 2363 32283
rect 7113 32249 7147 32283
rect 14381 32249 14415 32283
rect 17693 32249 17727 32283
rect 22017 32249 22051 32283
rect 24501 32249 24535 32283
rect 25237 32249 25271 32283
rect 1593 32181 1627 32215
rect 8309 32181 8343 32215
rect 9781 32181 9815 32215
rect 13277 32181 13311 32215
rect 15577 32181 15611 32215
rect 15761 32181 15795 32215
rect 19809 32181 19843 32215
rect 26433 32181 26467 32215
rect 29377 32181 29411 32215
rect 8401 31977 8435 32011
rect 11897 31977 11931 32011
rect 12449 31977 12483 32011
rect 28549 31977 28583 32011
rect 9321 31909 9355 31943
rect 10701 31909 10735 31943
rect 15945 31909 15979 31943
rect 17693 31909 17727 31943
rect 30757 31909 30791 31943
rect 4537 31841 4571 31875
rect 6101 31841 6135 31875
rect 9045 31841 9079 31875
rect 9873 31841 9907 31875
rect 10057 31841 10091 31875
rect 10977 31841 11011 31875
rect 11094 31841 11128 31875
rect 11253 31841 11287 31875
rect 12909 31841 12943 31875
rect 13001 31841 13035 31875
rect 14105 31841 14139 31875
rect 14289 31841 14323 31875
rect 14749 31841 14783 31875
rect 15142 31841 15176 31875
rect 17049 31841 17083 31875
rect 17233 31841 17267 31875
rect 17969 31841 18003 31875
rect 18086 31841 18120 31875
rect 18889 31841 18923 31875
rect 29193 31841 29227 31875
rect 31401 31841 31435 31875
rect 5457 31773 5491 31807
rect 5641 31773 5675 31807
rect 6377 31773 6411 31807
rect 6494 31773 6528 31807
rect 6653 31773 6687 31807
rect 7297 31773 7331 31807
rect 8401 31773 8435 31807
rect 8677 31773 8711 31807
rect 8953 31773 8987 31807
rect 9137 31773 9171 31807
rect 9321 31773 9355 31807
rect 9597 31773 9631 31807
rect 9781 31773 9815 31807
rect 9965 31773 9999 31807
rect 10241 31773 10275 31807
rect 15025 31773 15059 31807
rect 15301 31773 15335 31807
rect 16221 31773 16255 31807
rect 18245 31773 18279 31807
rect 27077 31773 27111 31807
rect 29009 31773 29043 31807
rect 29837 31773 29871 31807
rect 31217 31773 31251 31807
rect 4353 31705 4387 31739
rect 27344 31705 27378 31739
rect 28917 31705 28951 31739
rect 3893 31637 3927 31671
rect 4261 31637 4295 31671
rect 8585 31637 8619 31671
rect 9505 31637 9539 31671
rect 12817 31637 12851 31671
rect 16037 31637 16071 31671
rect 28457 31637 28491 31671
rect 29653 31637 29687 31671
rect 31125 31637 31159 31671
rect 3249 31433 3283 31467
rect 10701 31433 10735 31467
rect 24501 31433 24535 31467
rect 27261 31433 27295 31467
rect 27905 31433 27939 31467
rect 3770 31365 3804 31399
rect 9566 31365 9600 31399
rect 27997 31365 28031 31399
rect 29644 31365 29678 31399
rect 1593 31297 1627 31331
rect 1860 31297 1894 31331
rect 3433 31297 3467 31331
rect 7389 31297 7423 31331
rect 7481 31297 7515 31331
rect 19901 31297 19935 31331
rect 23121 31297 23155 31331
rect 23857 31297 23891 31331
rect 24317 31297 24351 31331
rect 25145 31297 25179 31331
rect 26157 31297 26191 31331
rect 27445 31297 27479 31331
rect 29377 31297 29411 31331
rect 31125 31297 31159 31331
rect 31953 31297 31987 31331
rect 3525 31229 3559 31263
rect 7573 31229 7607 31263
rect 9321 31229 9355 31263
rect 24961 31229 24995 31263
rect 25881 31229 25915 31263
rect 26019 31229 26053 31263
rect 28181 31229 28215 31263
rect 30849 31229 30883 31263
rect 4905 31161 4939 31195
rect 23305 31161 23339 31195
rect 24133 31161 24167 31195
rect 25605 31161 25639 31195
rect 27537 31161 27571 31195
rect 2973 31093 3007 31127
rect 7021 31093 7055 31127
rect 19717 31093 19751 31127
rect 26801 31093 26835 31127
rect 30757 31093 30791 31127
rect 31769 31093 31803 31127
rect 1961 30889 1995 30923
rect 8585 30889 8619 30923
rect 29745 30889 29779 30923
rect 2329 30821 2363 30855
rect 2881 30753 2915 30787
rect 5273 30753 5307 30787
rect 5457 30753 5491 30787
rect 5917 30753 5951 30787
rect 6193 30753 6227 30787
rect 6331 30753 6365 30787
rect 6469 30753 6503 30787
rect 21281 30753 21315 30787
rect 25329 30753 25363 30787
rect 25789 30753 25823 30787
rect 26341 30753 26375 30787
rect 30205 30753 30239 30787
rect 30297 30753 30331 30787
rect 2145 30685 2179 30719
rect 2697 30685 2731 30719
rect 2789 30685 2823 30719
rect 5181 30685 5215 30719
rect 7205 30685 7239 30719
rect 11989 30685 12023 30719
rect 14289 30685 14323 30719
rect 17325 30685 17359 30719
rect 19441 30685 19475 30719
rect 19708 30685 19742 30719
rect 21189 30685 21223 30719
rect 22845 30685 22879 30719
rect 24593 30685 24627 30719
rect 25145 30685 25179 30719
rect 26065 30685 26099 30719
rect 26182 30685 26216 30719
rect 30757 30685 30791 30719
rect 31024 30685 31058 30719
rect 7472 30617 7506 30651
rect 12256 30617 12290 30651
rect 21526 30617 21560 30651
rect 23112 30617 23146 30651
rect 4997 30549 5031 30583
rect 7113 30549 7147 30583
rect 13369 30549 13403 30583
rect 14105 30549 14139 30583
rect 17417 30549 17451 30583
rect 20821 30549 20855 30583
rect 21005 30549 21039 30583
rect 22661 30549 22695 30583
rect 24225 30549 24259 30583
rect 24409 30549 24443 30583
rect 26985 30549 27019 30583
rect 30113 30549 30147 30583
rect 32137 30549 32171 30583
rect 7849 30345 7883 30379
rect 12357 30345 12391 30379
rect 13093 30345 13127 30379
rect 16957 30345 16991 30379
rect 19901 30345 19935 30379
rect 20361 30345 20395 30379
rect 21833 30345 21867 30379
rect 22201 30345 22235 30379
rect 23765 30345 23799 30379
rect 13912 30277 13946 30311
rect 17478 30277 17512 30311
rect 22293 30277 22327 30311
rect 4629 30209 4663 30243
rect 4896 30209 4930 30243
rect 6929 30209 6963 30243
rect 8033 30209 8067 30243
rect 8760 30209 8794 30243
rect 9965 30209 9999 30243
rect 10232 30209 10266 30243
rect 11529 30209 11563 30243
rect 11713 30209 11747 30243
rect 12541 30209 12575 30243
rect 13001 30209 13035 30243
rect 13645 30209 13679 30243
rect 15384 30209 15418 30243
rect 16865 30209 16899 30243
rect 17141 30209 17175 30243
rect 18797 30209 18831 30243
rect 19533 30209 19567 30243
rect 20269 30209 20303 30243
rect 23213 30209 23247 30243
rect 24133 30209 24167 30243
rect 24225 30209 24259 30243
rect 25053 30209 25087 30243
rect 27353 30209 27387 30243
rect 27813 30209 27847 30243
rect 27905 30209 27939 30243
rect 36185 30209 36219 30243
rect 7205 30141 7239 30175
rect 8493 30141 8527 30175
rect 13277 30141 13311 30175
rect 15117 30141 15151 30175
rect 17233 30141 17267 30175
rect 20545 30141 20579 30175
rect 22477 30141 22511 30175
rect 24317 30141 24351 30175
rect 25329 30141 25363 30175
rect 27997 30141 28031 30175
rect 12633 30073 12667 30107
rect 16681 30073 16715 30107
rect 23397 30073 23431 30107
rect 27445 30073 27479 30107
rect 6009 30005 6043 30039
rect 9873 30005 9907 30039
rect 11345 30005 11379 30039
rect 11529 30005 11563 30039
rect 15025 30005 15059 30039
rect 16497 30005 16531 30039
rect 18613 30005 18647 30039
rect 18889 30005 18923 30039
rect 19717 30005 19751 30039
rect 27169 30005 27203 30039
rect 36369 30005 36403 30039
rect 5273 29801 5307 29835
rect 9137 29801 9171 29835
rect 10333 29801 10367 29835
rect 14105 29801 14139 29835
rect 16129 29801 16163 29835
rect 17417 29801 17451 29835
rect 28273 29801 28307 29835
rect 5181 29733 5215 29767
rect 3801 29665 3835 29699
rect 5733 29665 5767 29699
rect 5825 29665 5859 29699
rect 7297 29665 7331 29699
rect 9229 29665 9263 29699
rect 9689 29665 9723 29699
rect 14657 29665 14691 29699
rect 16589 29665 16623 29699
rect 16773 29665 16807 29699
rect 17969 29665 18003 29699
rect 24961 29665 24995 29699
rect 26893 29665 26927 29699
rect 3617 29597 3651 29631
rect 5641 29597 5675 29631
rect 7113 29597 7147 29631
rect 8953 29597 8987 29631
rect 9045 29597 9079 29631
rect 9597 29597 9631 29631
rect 9781 29597 9815 29631
rect 10333 29597 10367 29631
rect 10609 29597 10643 29631
rect 14473 29597 14507 29631
rect 24869 29597 24903 29631
rect 27160 29597 27194 29631
rect 29377 29597 29411 29631
rect 29561 29597 29595 29631
rect 31217 29597 31251 29631
rect 4046 29529 4080 29563
rect 17785 29529 17819 29563
rect 25206 29529 25240 29563
rect 29806 29529 29840 29563
rect 3433 29461 3467 29495
rect 6745 29461 6779 29495
rect 7205 29461 7239 29495
rect 10517 29461 10551 29495
rect 14565 29461 14599 29495
rect 16497 29461 16531 29495
rect 17877 29461 17911 29495
rect 24685 29461 24719 29495
rect 26341 29461 26375 29495
rect 29193 29461 29227 29495
rect 30941 29461 30975 29495
rect 31033 29461 31067 29495
rect 4261 29257 4295 29291
rect 4629 29257 4663 29291
rect 6009 29257 6043 29291
rect 7849 29257 7883 29291
rect 25145 29257 25179 29291
rect 25513 29257 25547 29291
rect 29561 29257 29595 29291
rect 29929 29257 29963 29291
rect 6714 29189 6748 29223
rect 30840 29189 30874 29223
rect 1593 29121 1627 29155
rect 1777 29121 1811 29155
rect 2044 29121 2078 29155
rect 4721 29121 4755 29155
rect 6193 29121 6227 29155
rect 6469 29121 6503 29155
rect 12541 29121 12575 29155
rect 18337 29121 18371 29155
rect 18604 29121 18638 29155
rect 19809 29121 19843 29155
rect 21005 29121 21039 29155
rect 22661 29121 22695 29155
rect 22928 29121 22962 29155
rect 27261 29121 27295 29155
rect 28181 29121 28215 29155
rect 28298 29121 28332 29155
rect 28457 29121 28491 29155
rect 30573 29121 30607 29155
rect 4905 29053 4939 29087
rect 19993 29053 20027 29087
rect 20729 29053 20763 29087
rect 20846 29053 20880 29087
rect 21649 29053 21683 29087
rect 25605 29053 25639 29087
rect 25789 29053 25823 29087
rect 27445 29053 27479 29087
rect 30021 29053 30055 29087
rect 30205 29053 30239 29087
rect 1409 28985 1443 29019
rect 12357 28985 12391 29019
rect 20453 28985 20487 29019
rect 27905 28985 27939 29019
rect 29101 28985 29135 29019
rect 3157 28917 3191 28951
rect 19717 28917 19751 28951
rect 24041 28917 24075 28951
rect 31953 28917 31987 28951
rect 2053 28713 2087 28747
rect 19257 28713 19291 28747
rect 23029 28713 23063 28747
rect 25421 28713 25455 28747
rect 30757 28713 30791 28747
rect 2421 28645 2455 28679
rect 5825 28645 5859 28679
rect 8953 28645 8987 28679
rect 13553 28645 13587 28679
rect 14749 28645 14783 28679
rect 3065 28577 3099 28611
rect 5181 28577 5215 28611
rect 6101 28577 6135 28611
rect 6377 28577 6411 28611
rect 10885 28577 10919 28611
rect 11278 28577 11312 28611
rect 11437 28577 11471 28611
rect 12173 28577 12207 28611
rect 14105 28577 14139 28611
rect 15142 28577 15176 28611
rect 15301 28577 15335 28611
rect 16957 28577 16991 28611
rect 17601 28577 17635 28611
rect 17877 28577 17911 28611
rect 19993 28577 20027 28611
rect 20177 28577 20211 28611
rect 21189 28577 21223 28611
rect 21465 28577 21499 28611
rect 21582 28577 21616 28611
rect 23949 28577 23983 28611
rect 27445 28577 27479 28611
rect 28089 28577 28123 28611
rect 28365 28577 28399 28611
rect 28482 28577 28516 28611
rect 31217 28577 31251 28611
rect 31309 28577 31343 28611
rect 2237 28509 2271 28543
rect 5365 28509 5399 28543
rect 6218 28509 6252 28543
rect 9229 28509 9263 28543
rect 9321 28509 9355 28543
rect 9505 28509 9539 28543
rect 10241 28509 10275 28543
rect 10425 28509 10459 28543
rect 11161 28509 11195 28543
rect 12440 28509 12474 28543
rect 14289 28509 14323 28543
rect 15025 28509 15059 28543
rect 17141 28509 17175 28543
rect 17994 28509 18028 28543
rect 18153 28509 18187 28543
rect 19441 28509 19475 28543
rect 19901 28509 19935 28543
rect 20545 28509 20579 28543
rect 20729 28509 20763 28543
rect 21741 28509 21775 28543
rect 23213 28509 23247 28543
rect 23765 28509 23799 28543
rect 25237 28509 25271 28543
rect 27629 28509 27663 28543
rect 28641 28509 28675 28543
rect 2789 28441 2823 28475
rect 8953 28441 8987 28475
rect 9413 28441 9447 28475
rect 23673 28441 23707 28475
rect 25881 28441 25915 28475
rect 2881 28373 2915 28407
rect 7021 28373 7055 28407
rect 9137 28373 9171 28407
rect 12081 28373 12115 28407
rect 15945 28373 15979 28407
rect 18797 28373 18831 28407
rect 19533 28373 19567 28407
rect 22385 28373 22419 28407
rect 23305 28373 23339 28407
rect 25973 28373 26007 28407
rect 29285 28373 29319 28407
rect 31125 28373 31159 28407
rect 4997 28169 5031 28203
rect 9781 28169 9815 28203
rect 12541 28169 12575 28203
rect 12909 28169 12943 28203
rect 16221 28169 16255 28203
rect 19717 28169 19751 28203
rect 20453 28169 20487 28203
rect 21005 28169 21039 28203
rect 27169 28169 27203 28203
rect 8668 28101 8702 28135
rect 22078 28101 22112 28135
rect 27077 28101 27111 28135
rect 28733 28101 28767 28135
rect 3884 28033 3918 28067
rect 8401 28033 8435 28067
rect 13001 28033 13035 28067
rect 13369 28033 13403 28067
rect 14289 28033 14323 28067
rect 14406 28033 14440 28067
rect 15669 28033 15703 28067
rect 16129 28033 16163 28067
rect 16865 28033 16899 28067
rect 17785 28033 17819 28067
rect 17902 28033 17936 28067
rect 18061 28033 18095 28067
rect 18889 28033 18923 28067
rect 19349 28033 19383 28067
rect 19533 28033 19567 28067
rect 20361 28033 20395 28067
rect 20821 28033 20855 28067
rect 21557 28033 21591 28067
rect 23489 28033 23523 28067
rect 24409 28033 24443 28067
rect 24547 28033 24581 28067
rect 25688 28033 25722 28067
rect 3617 27965 3651 27999
rect 13185 27965 13219 27999
rect 13553 27965 13587 27999
rect 14565 27965 14599 27999
rect 16405 27965 16439 27999
rect 17049 27965 17083 27999
rect 17509 27965 17543 27999
rect 21833 27965 21867 27999
rect 23673 27965 23707 27999
rect 24685 27965 24719 27999
rect 25421 27965 25455 27999
rect 28825 27965 28859 27999
rect 28917 27965 28951 27999
rect 14013 27897 14047 27931
rect 15761 27897 15795 27931
rect 19165 27897 19199 27931
rect 21373 27897 21407 27931
rect 24133 27897 24167 27931
rect 15209 27829 15243 27863
rect 15485 27829 15519 27863
rect 18705 27829 18739 27863
rect 18981 27829 19015 27863
rect 23213 27829 23247 27863
rect 25329 27829 25363 27863
rect 26801 27829 26835 27863
rect 28365 27829 28399 27863
rect 3893 27625 3927 27659
rect 21189 27625 21223 27659
rect 4169 27557 4203 27591
rect 5641 27557 5675 27591
rect 18705 27557 18739 27591
rect 29377 27557 29411 27591
rect 31033 27557 31067 27591
rect 31861 27557 31895 27591
rect 3525 27489 3559 27523
rect 4813 27489 4847 27523
rect 5181 27489 5215 27523
rect 5917 27489 5951 27523
rect 6055 27489 6089 27523
rect 6929 27489 6963 27523
rect 7573 27489 7607 27523
rect 10057 27489 10091 27523
rect 10241 27489 10275 27523
rect 10701 27489 10735 27523
rect 11094 27489 11128 27523
rect 21833 27489 21867 27523
rect 24593 27489 24627 27523
rect 25053 27489 25087 27523
rect 25467 27489 25501 27523
rect 25605 27489 25639 27523
rect 26893 27489 26927 27523
rect 30389 27489 30423 27523
rect 31217 27489 31251 27523
rect 1409 27421 1443 27455
rect 3341 27421 3375 27455
rect 4077 27421 4111 27455
rect 4537 27421 4571 27455
rect 4997 27421 5031 27455
rect 6193 27421 6227 27455
rect 7113 27421 7147 27455
rect 7849 27421 7883 27455
rect 7966 27421 8000 27455
rect 8125 27421 8159 27455
rect 10977 27421 11011 27455
rect 11253 27421 11287 27455
rect 14289 27421 14323 27455
rect 15209 27421 15243 27455
rect 15476 27421 15510 27455
rect 17325 27421 17359 27455
rect 19257 27421 19291 27455
rect 24409 27421 24443 27455
rect 25329 27421 25363 27455
rect 26709 27421 26743 27455
rect 27905 27421 27939 27455
rect 27997 27421 28031 27455
rect 31585 27421 31619 27455
rect 36185 27421 36219 27455
rect 1676 27353 1710 27387
rect 17592 27353 17626 27387
rect 21557 27353 21591 27387
rect 28242 27353 28276 27387
rect 30849 27353 30883 27387
rect 31677 27353 31711 27387
rect 2789 27285 2823 27319
rect 2881 27285 2915 27319
rect 3249 27285 3283 27319
rect 4629 27285 4663 27319
rect 6837 27285 6871 27319
rect 8769 27285 8803 27319
rect 11897 27285 11931 27319
rect 14105 27285 14139 27319
rect 16589 27285 16623 27319
rect 19441 27285 19475 27319
rect 21649 27285 21683 27319
rect 26249 27285 26283 27319
rect 26341 27285 26375 27319
rect 26801 27285 26835 27319
rect 27721 27285 27755 27319
rect 30665 27285 30699 27319
rect 30757 27285 30791 27319
rect 31493 27285 31527 27319
rect 36369 27285 36403 27319
rect 1777 27081 1811 27115
rect 2789 27081 2823 27115
rect 11345 27081 11379 27115
rect 15025 27081 15059 27115
rect 18613 27081 18647 27115
rect 25973 27081 26007 27115
rect 26433 27081 26467 27115
rect 30665 27081 30699 27115
rect 31125 27081 31159 27115
rect 3310 27013 3344 27047
rect 13912 27013 13946 27047
rect 20545 27013 20579 27047
rect 21005 27013 21039 27047
rect 32597 27013 32631 27047
rect 1961 26945 1995 26979
rect 2973 26945 3007 26979
rect 6837 26945 6871 26979
rect 7573 26945 7607 26979
rect 7690 26945 7724 26979
rect 9413 26945 9447 26979
rect 10232 26945 10266 26979
rect 11529 26945 11563 26979
rect 11713 26945 11747 26979
rect 12449 26945 12483 26979
rect 17325 26945 17359 26979
rect 17601 26945 17635 26979
rect 19901 26945 19935 26979
rect 20729 26945 20763 26979
rect 22937 26945 22971 26979
rect 23121 26945 23155 26979
rect 23213 26945 23247 26979
rect 25053 26945 25087 26979
rect 26157 26945 26191 26979
rect 26341 26945 26375 26979
rect 28365 26945 28399 26979
rect 29653 26945 29687 26979
rect 31033 26945 31067 26979
rect 31217 26945 31251 26979
rect 32137 26945 32171 26979
rect 32689 26945 32723 26979
rect 33333 26945 33367 26979
rect 33517 26945 33551 26979
rect 3065 26877 3099 26911
rect 6653 26877 6687 26911
rect 7849 26877 7883 26911
rect 9965 26877 9999 26911
rect 13645 26877 13679 26911
rect 18705 26877 18739 26911
rect 18797 26877 18831 26911
rect 30481 26877 30515 26911
rect 4445 26809 4479 26843
rect 7297 26809 7331 26843
rect 29837 26809 29871 26843
rect 8493 26741 8527 26775
rect 9505 26741 9539 26775
rect 11529 26741 11563 26775
rect 12265 26741 12299 26775
rect 18245 26741 18279 26775
rect 19717 26741 19751 26775
rect 21097 26741 21131 26775
rect 22753 26741 22787 26775
rect 25145 26741 25179 26775
rect 28457 26741 28491 26775
rect 4169 26537 4203 26571
rect 10149 26537 10183 26571
rect 13645 26537 13679 26571
rect 14105 26537 14139 26571
rect 17417 26537 17451 26571
rect 17601 26537 17635 26571
rect 32413 26537 32447 26571
rect 22753 26469 22787 26503
rect 4813 26401 4847 26435
rect 8769 26401 8803 26435
rect 8953 26401 8987 26435
rect 14657 26401 14691 26435
rect 17141 26401 17175 26435
rect 21465 26401 21499 26435
rect 21833 26401 21867 26435
rect 23857 26401 23891 26435
rect 30297 26401 30331 26435
rect 4537 26333 4571 26367
rect 9229 26333 9263 26367
rect 10149 26333 10183 26367
rect 10425 26333 10459 26367
rect 11897 26333 11931 26367
rect 12164 26333 12198 26367
rect 14473 26333 14507 26367
rect 17785 26333 17819 26367
rect 19349 26333 19383 26367
rect 19616 26333 19650 26367
rect 21097 26333 21131 26367
rect 21373 26333 21407 26367
rect 21925 26333 21959 26367
rect 23397 26333 23431 26367
rect 23765 26333 23799 26367
rect 24593 26333 24627 26367
rect 30481 26333 30515 26367
rect 30941 26333 30975 26367
rect 31493 26333 31527 26367
rect 31861 26333 31895 26367
rect 31953 26333 31987 26367
rect 32689 26333 32723 26367
rect 4629 26265 4663 26299
rect 8585 26265 8619 26299
rect 13553 26265 13587 26299
rect 14565 26265 14599 26299
rect 16957 26265 16991 26299
rect 17325 26265 17359 26299
rect 20913 26265 20947 26299
rect 22109 26265 22143 26299
rect 22569 26265 22603 26299
rect 24041 26265 24075 26299
rect 30849 26265 30883 26299
rect 31033 26265 31067 26299
rect 10333 26197 10367 26231
rect 13277 26197 13311 26231
rect 20729 26197 20763 26231
rect 21281 26197 21315 26231
rect 24409 26197 24443 26231
rect 2237 25993 2271 26027
rect 6837 25993 6871 26027
rect 12449 25993 12483 26027
rect 12817 25993 12851 26027
rect 17049 25993 17083 26027
rect 18981 25993 19015 26027
rect 19901 25993 19935 26027
rect 20361 25993 20395 26027
rect 22937 25993 22971 26027
rect 26985 25993 27019 26027
rect 33333 25993 33367 26027
rect 2697 25925 2731 25959
rect 8493 25925 8527 25959
rect 22845 25925 22879 25959
rect 24400 25925 24434 25959
rect 2053 25857 2087 25891
rect 2605 25857 2639 25891
rect 6745 25857 6779 25891
rect 7941 25857 7975 25891
rect 8309 25857 8343 25891
rect 9128 25857 9162 25891
rect 10333 25857 10367 25891
rect 10517 25857 10551 25891
rect 11897 25857 11931 25891
rect 13461 25857 13495 25891
rect 15117 25857 15151 25891
rect 15384 25857 15418 25891
rect 17509 25857 17543 25891
rect 18245 25857 18279 25891
rect 18797 25857 18831 25891
rect 19073 25857 19107 25891
rect 20269 25857 20303 25891
rect 22661 25857 22695 25891
rect 23305 25857 23339 25891
rect 24133 25857 24167 25891
rect 26341 25857 26375 25891
rect 27353 25857 27387 25891
rect 28089 25857 28123 25891
rect 31401 25857 31435 25891
rect 32137 25857 32171 25891
rect 33149 25857 33183 25891
rect 33517 25857 33551 25891
rect 2789 25789 2823 25823
rect 7021 25789 7055 25823
rect 7481 25789 7515 25823
rect 7849 25789 7883 25823
rect 8861 25789 8895 25823
rect 11529 25789 11563 25823
rect 11989 25789 12023 25823
rect 12909 25789 12943 25823
rect 13093 25789 13127 25823
rect 14381 25789 14415 25823
rect 14749 25789 14783 25823
rect 14841 25789 14875 25823
rect 17141 25789 17175 25823
rect 17325 25789 17359 25823
rect 17877 25789 17911 25823
rect 18337 25789 18371 25823
rect 20545 25789 20579 25823
rect 23397 25789 23431 25823
rect 27445 25789 27479 25823
rect 27537 25789 27571 25823
rect 32321 25789 32355 25823
rect 32597 25789 32631 25823
rect 32689 25789 32723 25823
rect 32965 25789 32999 25823
rect 16497 25721 16531 25755
rect 17693 25721 17727 25755
rect 33885 25721 33919 25755
rect 1869 25653 1903 25687
rect 6377 25653 6411 25687
rect 8125 25653 8159 25687
rect 10241 25653 10275 25687
rect 10425 25653 10459 25687
rect 12173 25653 12207 25687
rect 13553 25653 13587 25687
rect 15025 25653 15059 25687
rect 16681 25653 16715 25687
rect 18521 25653 18555 25687
rect 18613 25653 18647 25687
rect 23581 25653 23615 25687
rect 25513 25653 25547 25687
rect 26157 25653 26191 25687
rect 27905 25653 27939 25687
rect 31493 25653 31527 25687
rect 33977 25653 34011 25687
rect 2881 25449 2915 25483
rect 9321 25449 9355 25483
rect 24501 25449 24535 25483
rect 27353 25449 27387 25483
rect 31677 25449 31711 25483
rect 32321 25449 32355 25483
rect 10793 25381 10827 25415
rect 4721 25313 4755 25347
rect 5549 25313 5583 25347
rect 5825 25313 5859 25347
rect 6101 25313 6135 25347
rect 7481 25313 7515 25347
rect 7573 25313 7607 25347
rect 9413 25313 9447 25347
rect 10609 25313 10643 25347
rect 11437 25313 11471 25347
rect 25145 25313 25179 25347
rect 27629 25313 27663 25347
rect 31401 25313 31435 25347
rect 31861 25313 31895 25347
rect 32781 25313 32815 25347
rect 33977 25313 34011 25347
rect 1501 25245 1535 25279
rect 1768 25245 1802 25279
rect 3985 25245 4019 25279
rect 4905 25245 4939 25279
rect 5089 25245 5123 25279
rect 5942 25245 5976 25279
rect 7113 25245 7147 25279
rect 7941 25245 7975 25279
rect 9137 25245 9171 25279
rect 9229 25245 9263 25279
rect 10333 25245 10367 25279
rect 10425 25245 10459 25279
rect 10701 25245 10735 25279
rect 14841 25245 14875 25279
rect 15117 25245 15151 25279
rect 16129 25245 16163 25279
rect 19073 25245 19107 25279
rect 19257 25245 19291 25279
rect 24961 25245 24995 25279
rect 25973 25245 26007 25279
rect 26240 25245 26274 25279
rect 27896 25245 27930 25279
rect 29377 25245 29411 25279
rect 29561 25245 29595 25279
rect 31493 25245 31527 25279
rect 32229 25245 32263 25279
rect 33057 25245 33091 25279
rect 33701 25245 33735 25279
rect 4445 25177 4479 25211
rect 8125 25177 8159 25211
rect 11253 25177 11287 25211
rect 15025 25177 15059 25211
rect 19502 25177 19536 25211
rect 29806 25177 29840 25211
rect 31033 25177 31067 25211
rect 3801 25109 3835 25143
rect 4077 25109 4111 25143
rect 4537 25109 4571 25143
rect 6745 25109 6779 25143
rect 7757 25109 7791 25143
rect 10149 25109 10183 25143
rect 11161 25109 11195 25143
rect 14657 25109 14691 25143
rect 15945 25109 15979 25143
rect 18889 25109 18923 25143
rect 20637 25109 20671 25143
rect 24869 25109 24903 25143
rect 29009 25109 29043 25143
rect 29193 25109 29227 25143
rect 30941 25109 30975 25143
rect 31309 25109 31343 25143
rect 32045 25109 32079 25143
rect 4721 24905 4755 24939
rect 19625 24905 19659 24939
rect 19993 24905 20027 24939
rect 20085 24905 20119 24939
rect 23673 24905 23707 24939
rect 24133 24905 24167 24939
rect 27905 24905 27939 24939
rect 28273 24905 28307 24939
rect 29469 24905 29503 24939
rect 29837 24905 29871 24939
rect 30573 24905 30607 24939
rect 33885 24905 33919 24939
rect 3608 24837 3642 24871
rect 7573 24837 7607 24871
rect 24041 24837 24075 24871
rect 1409 24769 1443 24803
rect 6561 24769 6595 24803
rect 6653 24769 6687 24803
rect 6929 24769 6963 24803
rect 7665 24769 7699 24803
rect 12081 24769 12115 24803
rect 12348 24769 12382 24803
rect 13645 24769 13679 24803
rect 14381 24769 14415 24803
rect 14473 24769 14507 24803
rect 14749 24769 14783 24803
rect 17601 24769 17635 24803
rect 17693 24769 17727 24803
rect 17969 24769 18003 24803
rect 18061 24769 18095 24803
rect 21097 24769 21131 24803
rect 21189 24769 21223 24803
rect 21465 24769 21499 24803
rect 22569 24769 22603 24803
rect 22661 24769 22695 24803
rect 22937 24769 22971 24803
rect 29929 24769 29963 24803
rect 31033 24769 31067 24803
rect 32413 24769 32447 24803
rect 32761 24769 32795 24803
rect 1685 24701 1719 24735
rect 3341 24701 3375 24735
rect 7849 24701 7883 24735
rect 14105 24701 14139 24735
rect 14657 24701 14691 24735
rect 14841 24701 14875 24735
rect 15301 24701 15335 24735
rect 17877 24701 17911 24735
rect 20269 24701 20303 24735
rect 21373 24701 21407 24735
rect 23029 24701 23063 24735
rect 24225 24701 24259 24735
rect 28365 24701 28399 24735
rect 28457 24701 28491 24735
rect 30021 24701 30055 24735
rect 30297 24701 30331 24735
rect 30665 24701 30699 24735
rect 30757 24701 30791 24735
rect 31125 24701 31159 24735
rect 31401 24701 31435 24735
rect 32505 24701 32539 24735
rect 6837 24633 6871 24667
rect 14013 24633 14047 24667
rect 15117 24633 15151 24667
rect 23397 24633 23431 24667
rect 23489 24633 23523 24667
rect 6377 24565 6411 24599
rect 7205 24565 7239 24599
rect 13461 24565 13495 24599
rect 14197 24565 14231 24599
rect 17417 24565 17451 24599
rect 18245 24565 18279 24599
rect 20913 24565 20947 24599
rect 22385 24565 22419 24599
rect 22845 24565 22879 24599
rect 32229 24565 32263 24599
rect 11529 24361 11563 24395
rect 12357 24361 12391 24395
rect 18061 24361 18095 24395
rect 18613 24361 18647 24395
rect 21281 24361 21315 24395
rect 21833 24361 21867 24395
rect 22109 24361 22143 24395
rect 23673 24361 23707 24395
rect 28457 24361 28491 24395
rect 32413 24361 32447 24395
rect 2789 24293 2823 24327
rect 5457 24293 5491 24327
rect 11437 24293 11471 24327
rect 12633 24293 12667 24327
rect 17877 24293 17911 24327
rect 18521 24293 18555 24327
rect 21189 24293 21223 24327
rect 21649 24293 21683 24327
rect 25329 24293 25363 24327
rect 4997 24225 5031 24259
rect 5733 24225 5767 24259
rect 7297 24225 7331 24259
rect 8769 24225 8803 24259
rect 8953 24225 8987 24259
rect 11069 24225 11103 24259
rect 13093 24225 13127 24259
rect 13277 24225 13311 24259
rect 17601 24225 17635 24259
rect 24685 24225 24719 24259
rect 27261 24225 27295 24259
rect 27537 24225 27571 24259
rect 27675 24225 27709 24259
rect 1409 24157 1443 24191
rect 4813 24157 4847 24191
rect 5850 24157 5884 24191
rect 6009 24157 6043 24191
rect 7021 24157 7055 24191
rect 7113 24157 7147 24191
rect 7389 24157 7423 24191
rect 8585 24157 8619 24191
rect 12541 24157 12575 24191
rect 13001 24157 13035 24191
rect 21373 24157 21407 24191
rect 21925 24157 21959 24191
rect 22293 24157 22327 24191
rect 22569 24157 22603 24191
rect 23397 24157 23431 24191
rect 23489 24157 23523 24191
rect 23765 24157 23799 24191
rect 24869 24157 24903 24191
rect 25605 24157 25639 24191
rect 25722 24157 25756 24191
rect 25881 24157 25915 24191
rect 26617 24157 26651 24191
rect 26801 24157 26835 24191
rect 27813 24157 27847 24191
rect 32597 24157 32631 24191
rect 36185 24157 36219 24191
rect 1676 24089 1710 24123
rect 9198 24089 9232 24123
rect 18153 24089 18187 24123
rect 20821 24089 20855 24123
rect 6653 24021 6687 24055
rect 6837 24021 6871 24055
rect 10333 24021 10367 24055
rect 23213 24021 23247 24055
rect 26525 24021 26559 24055
rect 36369 24021 36403 24055
rect 1777 23817 1811 23851
rect 2145 23817 2179 23851
rect 2513 23817 2547 23851
rect 7021 23817 7055 23851
rect 7573 23817 7607 23851
rect 8499 23817 8533 23851
rect 11713 23817 11747 23851
rect 14473 23817 14507 23851
rect 18521 23817 18555 23851
rect 21649 23817 21683 23851
rect 22385 23817 22419 23851
rect 23581 23817 23615 23851
rect 30297 23817 30331 23851
rect 33425 23817 33459 23851
rect 8401 23749 8435 23783
rect 23121 23749 23155 23783
rect 23673 23749 23707 23783
rect 33333 23749 33367 23783
rect 1961 23681 1995 23715
rect 2605 23681 2639 23715
rect 2973 23681 3007 23715
rect 3240 23681 3274 23715
rect 6561 23681 6595 23715
rect 8585 23681 8619 23715
rect 8677 23681 8711 23715
rect 9045 23681 9079 23715
rect 9137 23681 9171 23715
rect 9229 23681 9263 23715
rect 9505 23681 9539 23715
rect 11621 23681 11655 23715
rect 11897 23681 11931 23715
rect 12633 23681 12667 23715
rect 13829 23681 13863 23715
rect 15117 23681 15151 23715
rect 15384 23681 15418 23715
rect 17601 23681 17635 23715
rect 17877 23681 17911 23715
rect 19349 23681 19383 23715
rect 19441 23681 19475 23715
rect 19809 23681 19843 23715
rect 20729 23681 20763 23715
rect 22293 23681 22327 23715
rect 24685 23681 24719 23715
rect 24869 23681 24903 23715
rect 25605 23681 25639 23715
rect 25722 23681 25756 23715
rect 26985 23681 27019 23715
rect 27169 23681 27203 23715
rect 27905 23681 27939 23715
rect 28022 23681 28056 23715
rect 28917 23681 28951 23715
rect 29184 23681 29218 23715
rect 2697 23613 2731 23647
rect 7113 23613 7147 23647
rect 9689 23613 9723 23647
rect 10425 23613 10459 23647
rect 10563 23613 10597 23647
rect 10701 23613 10735 23647
rect 12817 23613 12851 23647
rect 13553 23613 13587 23647
rect 13670 23613 13704 23647
rect 16681 23613 16715 23647
rect 16865 23613 16899 23647
rect 17718 23613 17752 23647
rect 19625 23613 19659 23647
rect 19993 23613 20027 23647
rect 20846 23613 20880 23647
rect 21005 23613 21039 23647
rect 24133 23613 24167 23647
rect 25881 23613 25915 23647
rect 28181 23613 28215 23647
rect 6837 23545 6871 23579
rect 7389 23545 7423 23579
rect 10149 23545 10183 23579
rect 13277 23545 13311 23579
rect 17325 23545 17359 23579
rect 20453 23545 20487 23579
rect 23397 23545 23431 23579
rect 24041 23545 24075 23579
rect 25329 23545 25363 23579
rect 27629 23545 27663 23579
rect 4353 23477 4387 23511
rect 11345 23477 11379 23511
rect 12081 23477 12115 23511
rect 16497 23477 16531 23511
rect 18981 23477 19015 23511
rect 26525 23477 26559 23511
rect 28825 23477 28859 23511
rect 3801 23273 3835 23307
rect 11713 23273 11747 23307
rect 15669 23273 15703 23307
rect 29193 23273 29227 23307
rect 34529 23273 34563 23307
rect 2881 23205 2915 23239
rect 5089 23205 5123 23239
rect 20453 23205 20487 23239
rect 32781 23205 32815 23239
rect 3341 23137 3375 23171
rect 3525 23137 3559 23171
rect 5641 23137 5675 23171
rect 9873 23137 9907 23171
rect 10057 23137 10091 23171
rect 10517 23137 10551 23171
rect 10910 23137 10944 23171
rect 16405 23137 16439 23171
rect 16497 23137 16531 23171
rect 19809 23137 19843 23171
rect 19993 23137 20027 23171
rect 20729 23137 20763 23171
rect 20846 23137 20880 23171
rect 24961 23137 24995 23171
rect 26341 23137 26375 23171
rect 26525 23137 26559 23171
rect 30113 23137 30147 23171
rect 30389 23137 30423 23171
rect 32045 23137 32079 23171
rect 32413 23137 32447 23171
rect 3985 23069 4019 23103
rect 5549 23069 5583 23103
rect 10793 23069 10827 23103
rect 11069 23069 11103 23103
rect 14473 23069 14507 23103
rect 15853 23069 15887 23103
rect 18981 23069 19015 23103
rect 19257 23069 19291 23103
rect 21005 23069 21039 23103
rect 23949 23069 23983 23103
rect 24777 23069 24811 23103
rect 27629 23069 27663 23103
rect 27721 23069 27755 23103
rect 29377 23069 29411 23103
rect 29929 23069 29963 23103
rect 31033 23069 31067 23103
rect 31769 23069 31803 23103
rect 33149 23069 33183 23103
rect 3249 23001 3283 23035
rect 4813 23001 4847 23035
rect 27966 23001 28000 23035
rect 31125 23001 31159 23035
rect 31309 23001 31343 23035
rect 33416 23001 33450 23035
rect 4905 22933 4939 22967
rect 5457 22933 5491 22967
rect 14289 22933 14323 22967
rect 15945 22933 15979 22967
rect 16313 22933 16347 22967
rect 18797 22933 18831 22967
rect 19441 22933 19475 22967
rect 21649 22933 21683 22967
rect 23765 22933 23799 22967
rect 24409 22933 24443 22967
rect 24869 22933 24903 22967
rect 25881 22933 25915 22967
rect 26249 22933 26283 22967
rect 27445 22933 27479 22967
rect 29101 22933 29135 22967
rect 29561 22933 29595 22967
rect 30021 22933 30055 22967
rect 30573 22933 30607 22967
rect 30941 22933 30975 22967
rect 31585 22933 31619 22967
rect 31677 22933 31711 22967
rect 32873 22933 32907 22967
rect 5457 22729 5491 22763
rect 19901 22729 19935 22763
rect 24777 22729 24811 22763
rect 27997 22729 28031 22763
rect 32321 22729 32355 22763
rect 33793 22729 33827 22763
rect 14718 22661 14752 22695
rect 18788 22661 18822 22695
rect 23664 22661 23698 22695
rect 28365 22661 28399 22695
rect 1409 22593 1443 22627
rect 4077 22593 4111 22627
rect 4344 22593 4378 22627
rect 7573 22593 7607 22627
rect 7840 22593 7874 22627
rect 9045 22593 9079 22627
rect 9229 22593 9263 22627
rect 12541 22593 12575 22627
rect 13461 22593 13495 22627
rect 13599 22593 13633 22627
rect 14473 22593 14507 22627
rect 18153 22593 18187 22627
rect 25697 22593 25731 22627
rect 31033 22593 31067 22627
rect 31677 22593 31711 22627
rect 31861 22593 31895 22627
rect 32137 22593 32171 22627
rect 32321 22593 32355 22627
rect 32413 22593 32447 22627
rect 32873 22593 32907 22627
rect 33977 22593 34011 22627
rect 12725 22525 12759 22559
rect 13737 22525 13771 22559
rect 18521 22525 18555 22559
rect 23397 22525 23431 22559
rect 28457 22525 28491 22559
rect 28641 22525 28675 22559
rect 30757 22525 30791 22559
rect 33149 22525 33183 22559
rect 1593 22457 1627 22491
rect 8953 22457 8987 22491
rect 13185 22457 13219 22491
rect 9045 22389 9079 22423
rect 14381 22389 14415 22423
rect 15853 22389 15887 22423
rect 18337 22389 18371 22423
rect 25789 22389 25823 22423
rect 31677 22389 31711 22423
rect 4629 22185 4663 22219
rect 7941 22185 7975 22219
rect 10609 22185 10643 22219
rect 14197 22185 14231 22219
rect 26985 22185 27019 22219
rect 6929 22117 6963 22151
rect 12817 22117 12851 22151
rect 9229 22049 9263 22083
rect 13553 22049 13587 22083
rect 14749 22049 14783 22083
rect 16221 22049 16255 22083
rect 16405 22049 16439 22083
rect 16865 22049 16899 22083
rect 17141 22049 17175 22083
rect 17258 22049 17292 22083
rect 17417 22049 17451 22083
rect 21373 22049 21407 22083
rect 25605 22049 25639 22083
rect 30665 22049 30699 22083
rect 31309 22049 31343 22083
rect 32781 22049 32815 22083
rect 33517 22049 33551 22083
rect 1593 21981 1627 22015
rect 4813 21981 4847 22015
rect 8217 21981 8251 22015
rect 10701 21981 10735 22015
rect 10885 21981 10919 22015
rect 11437 21981 11471 22015
rect 13277 21981 13311 22015
rect 14565 21981 14599 22015
rect 21281 21981 21315 22015
rect 25513 21981 25547 22015
rect 30481 21981 30515 22015
rect 31033 21981 31067 22015
rect 32505 21981 32539 22015
rect 33333 21981 33367 22015
rect 1860 21913 1894 21947
rect 6653 21913 6687 21947
rect 7941 21913 7975 21947
rect 9474 21913 9508 21947
rect 11704 21913 11738 21947
rect 14657 21913 14691 21947
rect 21618 21913 21652 21947
rect 25850 21913 25884 21947
rect 30205 21913 30239 21947
rect 2973 21845 3007 21879
rect 7113 21845 7147 21879
rect 8125 21845 8159 21879
rect 10793 21845 10827 21879
rect 12909 21845 12943 21879
rect 13369 21845 13403 21879
rect 18061 21845 18095 21879
rect 21097 21845 21131 21879
rect 22753 21845 22787 21879
rect 25329 21845 25363 21879
rect 30573 21845 30607 21879
rect 30849 21845 30883 21879
rect 32137 21845 32171 21879
rect 32597 21845 32631 21879
rect 32965 21845 32999 21879
rect 33425 21845 33459 21879
rect 1961 21641 1995 21675
rect 2237 21641 2271 21675
rect 2697 21641 2731 21675
rect 6193 21641 6227 21675
rect 7941 21641 7975 21675
rect 11805 21641 11839 21675
rect 16773 21641 16807 21675
rect 18429 21641 18463 21675
rect 21833 21641 21867 21675
rect 22201 21641 22235 21675
rect 22293 21641 22327 21675
rect 25053 21641 25087 21675
rect 28733 21641 28767 21675
rect 9321 21573 9355 21607
rect 17294 21573 17328 21607
rect 2145 21505 2179 21539
rect 2605 21505 2639 21539
rect 4537 21505 4571 21539
rect 5273 21505 5307 21539
rect 7205 21505 7239 21539
rect 7297 21505 7331 21539
rect 7757 21505 7791 21539
rect 8033 21505 8067 21539
rect 9505 21505 9539 21539
rect 9597 21505 9631 21539
rect 11989 21505 12023 21539
rect 15945 21505 15979 21539
rect 16957 21505 16991 21539
rect 17049 21505 17083 21539
rect 20637 21505 20671 21539
rect 23121 21505 23155 21539
rect 23388 21505 23422 21539
rect 24961 21505 24995 21539
rect 28641 21505 28675 21539
rect 33333 21505 33367 21539
rect 2881 21437 2915 21471
rect 4353 21437 4387 21471
rect 5411 21437 5445 21471
rect 5549 21437 5583 21471
rect 6837 21437 6871 21471
rect 16037 21437 16071 21471
rect 16221 21437 16255 21471
rect 20269 21437 20303 21471
rect 20729 21437 20763 21471
rect 21005 21437 21039 21471
rect 22477 21437 22511 21471
rect 25145 21437 25179 21471
rect 28825 21437 28859 21471
rect 4997 21369 5031 21403
rect 9321 21369 9355 21403
rect 21373 21369 21407 21403
rect 7481 21301 7515 21335
rect 7573 21301 7607 21335
rect 15577 21301 15611 21335
rect 20913 21301 20947 21335
rect 21465 21301 21499 21335
rect 24501 21301 24535 21335
rect 24593 21301 24627 21335
rect 28273 21301 28307 21335
rect 33149 21301 33183 21335
rect 9873 21097 9907 21131
rect 16313 21097 16347 21131
rect 17325 21097 17359 21131
rect 19717 21097 19751 21131
rect 20361 21097 20395 21131
rect 23397 21097 23431 21131
rect 27261 21097 27295 21131
rect 27905 21097 27939 21131
rect 29377 21097 29411 21131
rect 32321 21097 32355 21131
rect 6469 21029 6503 21063
rect 7665 21029 7699 21063
rect 10885 21029 10919 21063
rect 13737 21029 13771 21063
rect 17141 21029 17175 21063
rect 25145 21029 25179 21063
rect 27721 21029 27755 21063
rect 30849 21029 30883 21063
rect 31401 21029 31435 21063
rect 32873 21029 32907 21063
rect 2789 20961 2823 20995
rect 4353 20961 4387 20995
rect 4629 20961 4663 20995
rect 5273 20961 5307 20995
rect 5549 20961 5583 20995
rect 5666 20961 5700 20995
rect 7205 20961 7239 20995
rect 9321 20961 9355 20995
rect 10977 20961 11011 20995
rect 11437 20961 11471 20995
rect 11529 20961 11563 20995
rect 14197 20961 14231 20995
rect 14565 20961 14599 20995
rect 17785 20961 17819 20995
rect 17877 20961 17911 20995
rect 18521 20961 18555 20995
rect 20545 20961 20579 20995
rect 24777 20961 24811 20995
rect 25697 20961 25731 20995
rect 25789 20961 25823 20995
rect 26433 20961 26467 20995
rect 26709 20961 26743 20995
rect 27997 20961 28031 20995
rect 30389 20961 30423 20995
rect 30941 20961 30975 20995
rect 33149 20961 33183 20995
rect 2605 20893 2639 20927
rect 3617 20893 3651 20927
rect 4813 20893 4847 20927
rect 5825 20893 5859 20927
rect 6929 20893 6963 20927
rect 7021 20893 7055 20927
rect 7297 20893 7331 20927
rect 9413 20893 9447 20927
rect 11069 20893 11103 20927
rect 11989 20893 12023 20927
rect 12173 20893 12207 20927
rect 12265 20893 12299 20927
rect 14657 20893 14691 20927
rect 14933 20893 14967 20927
rect 16773 20893 16807 20927
rect 17693 20893 17727 20927
rect 18613 20893 18647 20927
rect 19901 20893 19935 20927
rect 20085 20893 20119 20927
rect 20177 20893 20211 20927
rect 20453 20893 20487 20927
rect 20729 20893 20763 20927
rect 20913 20893 20947 20927
rect 21005 20893 21039 20927
rect 23581 20893 23615 20927
rect 26525 20893 26559 20927
rect 26985 20893 27019 20927
rect 27077 20893 27111 20927
rect 27353 20893 27387 20927
rect 29745 20893 29779 20927
rect 30481 20893 30515 20927
rect 31769 20893 31803 20927
rect 32137 20893 32171 20927
rect 32689 20893 32723 20927
rect 33405 20893 33439 20927
rect 2697 20825 2731 20859
rect 4169 20825 4203 20859
rect 7389 20825 7423 20859
rect 8953 20825 8987 20859
rect 9781 20825 9815 20859
rect 10517 20825 10551 20859
rect 13461 20825 13495 20859
rect 15200 20825 15234 20859
rect 18797 20825 18831 20859
rect 19625 20825 19659 20859
rect 25973 20825 26007 20859
rect 27445 20825 27479 20859
rect 28264 20825 28298 20859
rect 31677 20825 31711 20859
rect 36093 20825 36127 20859
rect 2237 20757 2271 20791
rect 3433 20757 3467 20791
rect 3801 20757 3835 20791
rect 4261 20757 4295 20791
rect 6745 20757 6779 20791
rect 7849 20757 7883 20791
rect 9597 20757 9631 20791
rect 11713 20757 11747 20791
rect 11805 20757 11839 20791
rect 13921 20757 13955 20791
rect 14841 20757 14875 20791
rect 17233 20757 17267 20791
rect 18153 20757 18187 20791
rect 25237 20757 25271 20791
rect 25329 20757 25363 20791
rect 26065 20757 26099 20791
rect 26801 20757 26835 20791
rect 29561 20757 29595 20791
rect 31217 20757 31251 20791
rect 31585 20757 31619 20791
rect 31953 20757 31987 20791
rect 34529 20757 34563 20791
rect 36369 20757 36403 20791
rect 2881 20553 2915 20587
rect 4445 20553 4479 20587
rect 8125 20553 8159 20587
rect 8769 20553 8803 20587
rect 14473 20553 14507 20587
rect 15301 20553 15335 20587
rect 18337 20553 18371 20587
rect 19441 20553 19475 20587
rect 20637 20553 20671 20587
rect 22293 20553 22327 20587
rect 25237 20553 25271 20587
rect 27721 20553 27755 20587
rect 28089 20553 28123 20587
rect 28549 20553 28583 20587
rect 30665 20553 30699 20587
rect 33517 20553 33551 20587
rect 3332 20485 3366 20519
rect 20177 20485 20211 20519
rect 22201 20485 22235 20519
rect 25145 20485 25179 20519
rect 26341 20485 26375 20519
rect 28457 20485 28491 20519
rect 30849 20485 30883 20519
rect 31493 20485 31527 20519
rect 32382 20485 32416 20519
rect 1501 20417 1535 20451
rect 1768 20417 1802 20451
rect 3065 20417 3099 20451
rect 7389 20417 7423 20451
rect 8677 20417 8711 20451
rect 9321 20417 9355 20451
rect 10885 20417 10919 20451
rect 10977 20417 11011 20451
rect 11253 20417 11287 20451
rect 12725 20417 12759 20451
rect 13001 20417 13035 20451
rect 14381 20417 14415 20451
rect 15485 20417 15519 20451
rect 17417 20417 17451 20451
rect 17509 20417 17543 20451
rect 17785 20417 17819 20451
rect 18245 20417 18279 20451
rect 19349 20417 19383 20451
rect 23121 20417 23155 20451
rect 24317 20417 24351 20451
rect 24409 20417 24443 20451
rect 24685 20417 24719 20451
rect 26157 20417 26191 20451
rect 27629 20417 27663 20451
rect 29009 20417 29043 20451
rect 31677 20417 31711 20451
rect 31861 20417 31895 20451
rect 31953 20417 31987 20451
rect 32137 20417 32171 20451
rect 7113 20349 7147 20383
rect 8953 20349 8987 20383
rect 11161 20349 11195 20383
rect 14657 20349 14691 20383
rect 18521 20349 18555 20383
rect 22385 20349 22419 20383
rect 25329 20349 25363 20383
rect 28641 20349 28675 20383
rect 29193 20349 29227 20383
rect 30389 20349 30423 20383
rect 30757 20349 30791 20383
rect 20545 20281 20579 20315
rect 23305 20281 23339 20315
rect 24777 20281 24811 20315
rect 8309 20213 8343 20247
rect 9505 20213 9539 20247
rect 10701 20213 10735 20247
rect 13737 20213 13771 20247
rect 14013 20213 14047 20247
rect 17233 20213 17267 20247
rect 17693 20213 17727 20247
rect 17877 20213 17911 20247
rect 21833 20213 21867 20247
rect 24133 20213 24167 20247
rect 24593 20213 24627 20247
rect 31033 20213 31067 20247
rect 1869 20009 1903 20043
rect 6837 20009 6871 20043
rect 8493 20009 8527 20043
rect 10977 20009 11011 20043
rect 13369 20009 13403 20043
rect 13829 20009 13863 20043
rect 23581 20009 23615 20043
rect 32689 20009 32723 20043
rect 6653 19941 6687 19975
rect 10793 19941 10827 19975
rect 16957 19941 16991 19975
rect 10517 19873 10551 19907
rect 15025 19873 15059 19907
rect 16589 19873 16623 19907
rect 21465 19873 21499 19907
rect 33241 19873 33275 19907
rect 2053 19805 2087 19839
rect 6377 19805 6411 19839
rect 8217 19805 8251 19839
rect 8309 19805 8343 19839
rect 8585 19805 8619 19839
rect 13553 19805 13587 19839
rect 13645 19805 13679 19839
rect 13921 19805 13955 19839
rect 15301 19805 15335 19839
rect 16405 19805 16439 19839
rect 16773 19805 16807 19839
rect 21373 19805 21407 19839
rect 22937 19805 22971 19839
rect 23397 19805 23431 19839
rect 27997 19805 28031 19839
rect 29929 19805 29963 19839
rect 33057 19805 33091 19839
rect 34345 19805 34379 19839
rect 19993 19737 20027 19771
rect 21710 19737 21744 19771
rect 34529 19737 34563 19771
rect 34805 19737 34839 19771
rect 8033 19669 8067 19703
rect 15945 19669 15979 19703
rect 16313 19669 16347 19703
rect 20085 19669 20119 19703
rect 21189 19669 21223 19703
rect 22845 19669 22879 19703
rect 23121 19669 23155 19703
rect 28181 19669 28215 19703
rect 29745 19669 29779 19703
rect 33149 19669 33183 19703
rect 34897 19669 34931 19703
rect 12541 19465 12575 19499
rect 14749 19465 14783 19499
rect 19257 19465 19291 19499
rect 22017 19465 22051 19499
rect 25329 19465 25363 19499
rect 26065 19465 26099 19499
rect 35541 19465 35575 19499
rect 1501 19397 1535 19431
rect 2973 19397 3007 19431
rect 4169 19397 4203 19431
rect 26341 19397 26375 19431
rect 29736 19397 29770 19431
rect 33241 19397 33275 19431
rect 2421 19329 2455 19363
rect 2881 19329 2915 19363
rect 3985 19329 4019 19363
rect 4353 19329 4387 19363
rect 4721 19329 4755 19363
rect 8300 19329 8334 19363
rect 12449 19329 12483 19363
rect 12909 19329 12943 19363
rect 15301 19329 15335 19363
rect 16957 19329 16991 19363
rect 18245 19329 18279 19363
rect 18521 19329 18555 19363
rect 19993 19329 20027 19363
rect 21833 19329 21867 19363
rect 23397 19329 23431 19363
rect 25421 19329 25455 19363
rect 25881 19329 25915 19363
rect 26985 19329 27019 19363
rect 29469 19329 29503 19363
rect 34161 19329 34195 19363
rect 34428 19329 34462 19363
rect 3157 19261 3191 19295
rect 8033 19261 8067 19295
rect 12725 19261 12759 19295
rect 13093 19261 13127 19295
rect 13553 19261 13587 19295
rect 13829 19261 13863 19295
rect 13946 19261 13980 19295
rect 14105 19261 14139 19295
rect 15025 19261 15059 19295
rect 16681 19261 16715 19295
rect 25605 19261 25639 19295
rect 27169 19261 27203 19295
rect 27905 19261 27939 19295
rect 28043 19261 28077 19295
rect 28191 19261 28225 19295
rect 28825 19261 28859 19295
rect 33425 19261 33459 19295
rect 2513 19193 2547 19227
rect 4537 19193 4571 19227
rect 27629 19193 27663 19227
rect 1593 19125 1627 19159
rect 2237 19125 2271 19159
rect 4813 19125 4847 19159
rect 9413 19125 9447 19159
rect 12081 19125 12115 19159
rect 20177 19125 20211 19159
rect 23673 19125 23707 19159
rect 24961 19125 24995 19159
rect 26433 19125 26467 19159
rect 30849 19125 30883 19159
rect 3249 18921 3283 18955
rect 6193 18921 6227 18955
rect 8125 18921 8159 18955
rect 8953 18921 8987 18955
rect 11253 18921 11287 18955
rect 12909 18921 12943 18955
rect 16221 18921 16255 18955
rect 18245 18921 18279 18955
rect 21465 18921 21499 18955
rect 22017 18921 22051 18955
rect 26249 18921 26283 18955
rect 29193 18921 29227 18955
rect 29837 18921 29871 18955
rect 33793 18921 33827 18955
rect 20269 18853 20303 18887
rect 27169 18853 27203 18887
rect 4353 18785 4387 18819
rect 4997 18785 5031 18819
rect 9413 18785 9447 18819
rect 9597 18785 9631 18819
rect 10057 18785 10091 18819
rect 14841 18785 14875 18819
rect 16405 18785 16439 18819
rect 17049 18785 17083 18819
rect 20662 18785 20696 18819
rect 20821 18785 20855 18819
rect 25053 18785 25087 18819
rect 25446 18785 25480 18819
rect 25605 18785 25639 18819
rect 27997 18785 28031 18819
rect 28549 18785 28583 18819
rect 30389 18785 30423 18819
rect 32413 18785 32447 18819
rect 34989 18785 35023 18819
rect 1869 18717 1903 18751
rect 2136 18717 2170 18751
rect 4537 18717 4571 18751
rect 5273 18717 5307 18751
rect 5411 18717 5445 18751
rect 5549 18717 5583 18751
rect 9137 18717 9171 18751
rect 9229 18717 9263 18751
rect 10333 18717 10367 18751
rect 10471 18717 10505 18751
rect 10609 18717 10643 18751
rect 11529 18717 11563 18751
rect 16589 18717 16623 18751
rect 17325 18717 17359 18751
rect 17442 18717 17476 18751
rect 17601 18717 17635 18751
rect 19625 18717 19659 18751
rect 19809 18717 19843 18751
rect 20545 18717 20579 18751
rect 21833 18717 21867 18751
rect 24409 18717 24443 18751
rect 24593 18717 24627 18751
rect 25329 18717 25363 18751
rect 26985 18717 27019 18751
rect 27353 18717 27387 18751
rect 27537 18717 27571 18751
rect 28273 18717 28307 18751
rect 28390 18717 28424 18751
rect 30205 18717 30239 18751
rect 30297 18717 30331 18751
rect 30941 18717 30975 18751
rect 34713 18717 34747 18751
rect 8033 18649 8067 18683
rect 8953 18649 8987 18683
rect 11796 18649 11830 18683
rect 15108 18649 15142 18683
rect 31208 18649 31242 18683
rect 32658 18649 32692 18683
rect 32321 18581 32355 18615
rect 6193 18377 6227 18411
rect 8217 18377 8251 18411
rect 9045 18377 9079 18411
rect 11345 18377 11379 18411
rect 11897 18377 11931 18411
rect 14749 18377 14783 18411
rect 15209 18377 15243 18411
rect 18521 18377 18555 18411
rect 21189 18377 21223 18411
rect 22201 18377 22235 18411
rect 24869 18377 24903 18411
rect 26341 18377 26375 18411
rect 28641 18377 28675 18411
rect 31217 18377 31251 18411
rect 32229 18377 32263 18411
rect 35357 18377 35391 18411
rect 2697 18309 2731 18343
rect 27997 18309 28031 18343
rect 28549 18309 28583 18343
rect 30757 18309 30791 18343
rect 4353 18241 4387 18275
rect 4537 18241 4571 18275
rect 8953 18241 8987 18275
rect 9137 18241 9171 18275
rect 9505 18241 9539 18275
rect 10425 18241 10459 18275
rect 10542 18241 10576 18275
rect 10701 18241 10735 18275
rect 12081 18241 12115 18275
rect 12909 18241 12943 18275
rect 13093 18241 13127 18275
rect 13829 18241 13863 18275
rect 13946 18241 13980 18275
rect 15393 18241 15427 18275
rect 16681 18241 16715 18275
rect 17601 18241 17635 18275
rect 17877 18241 17911 18275
rect 18613 18241 18647 18275
rect 19349 18241 19383 18275
rect 20269 18241 20303 18275
rect 20545 18241 20579 18275
rect 22937 18241 22971 18275
rect 23213 18241 23247 18275
rect 23949 18241 23983 18275
rect 24225 18241 24259 18275
rect 25217 18241 25251 18275
rect 27261 18241 27295 18275
rect 31401 18241 31435 18275
rect 32413 18241 32447 18275
rect 33057 18241 33091 18275
rect 33324 18241 33358 18275
rect 35173 18241 35207 18275
rect 2789 18173 2823 18207
rect 2973 18173 3007 18207
rect 5273 18173 5307 18207
rect 5411 18173 5445 18207
rect 5549 18173 5583 18207
rect 6377 18173 6411 18207
rect 6561 18173 6595 18207
rect 7297 18173 7331 18207
rect 7414 18173 7448 18207
rect 7573 18173 7607 18207
rect 9689 18173 9723 18207
rect 14105 18173 14139 18207
rect 16865 18173 16899 18207
rect 17718 18173 17752 18207
rect 19533 18173 19567 18207
rect 20386 18173 20420 18207
rect 22293 18173 22327 18207
rect 22477 18173 22511 18207
rect 23029 18173 23063 18207
rect 23673 18173 23707 18207
rect 24066 18173 24100 18207
rect 24961 18173 24995 18207
rect 26985 18173 27019 18207
rect 30849 18173 30883 18207
rect 30941 18173 30975 18207
rect 34713 18173 34747 18207
rect 35081 18173 35115 18207
rect 4997 18105 5031 18139
rect 7021 18105 7055 18139
rect 10149 18105 10183 18139
rect 13553 18105 13587 18139
rect 17325 18105 17359 18139
rect 19993 18105 20027 18139
rect 28181 18105 28215 18139
rect 30389 18105 30423 18139
rect 2329 18037 2363 18071
rect 18797 18037 18831 18071
rect 21833 18037 21867 18071
rect 22753 18037 22787 18071
rect 34437 18037 34471 18071
rect 5181 17833 5215 17867
rect 7849 17833 7883 17867
rect 9689 17833 9723 17867
rect 10195 17833 10229 17867
rect 22109 17833 22143 17867
rect 23857 17833 23891 17867
rect 24961 17833 24995 17867
rect 30941 17833 30975 17867
rect 33517 17833 33551 17867
rect 6653 17765 6687 17799
rect 27353 17765 27387 17799
rect 6009 17697 6043 17731
rect 6929 17697 6963 17731
rect 9873 17697 9907 17731
rect 10977 17697 11011 17731
rect 14565 17697 14599 17731
rect 14657 17697 14691 17731
rect 17601 17697 17635 17731
rect 28089 17697 28123 17731
rect 29561 17697 29595 17731
rect 1409 17629 1443 17663
rect 3801 17629 3835 17663
rect 6193 17629 6227 17663
rect 7046 17629 7080 17663
rect 7205 17629 7239 17663
rect 9505 17629 9539 17663
rect 9597 17629 9631 17663
rect 9965 17629 9999 17663
rect 10885 17629 10919 17663
rect 11069 17629 11103 17663
rect 17417 17629 17451 17663
rect 18981 17629 19015 17663
rect 19257 17629 19291 17663
rect 20729 17629 20763 17663
rect 22477 17629 22511 17663
rect 22744 17629 22778 17663
rect 25145 17629 25179 17663
rect 25881 17629 25915 17663
rect 25973 17629 26007 17663
rect 27813 17629 27847 17663
rect 33701 17629 33735 17663
rect 1676 17561 1710 17595
rect 4068 17561 4102 17595
rect 14473 17561 14507 17595
rect 19502 17561 19536 17595
rect 20996 17561 21030 17595
rect 26240 17561 26274 17595
rect 29806 17561 29840 17595
rect 2789 17493 2823 17527
rect 9321 17493 9355 17527
rect 9873 17493 9907 17527
rect 14105 17493 14139 17527
rect 17049 17493 17083 17527
rect 17509 17493 17543 17527
rect 18797 17493 18831 17527
rect 20637 17493 20671 17527
rect 25697 17493 25731 17527
rect 27445 17493 27479 17527
rect 27905 17493 27939 17527
rect 1869 17289 1903 17323
rect 3985 17289 4019 17323
rect 4445 17289 4479 17323
rect 4813 17289 4847 17323
rect 4905 17289 4939 17323
rect 6101 17289 6135 17323
rect 6837 17289 6871 17323
rect 11069 17289 11103 17323
rect 12909 17289 12943 17323
rect 13277 17289 13311 17323
rect 14933 17289 14967 17323
rect 18061 17289 18095 17323
rect 18889 17289 18923 17323
rect 19257 17289 19291 17323
rect 21005 17289 21039 17323
rect 22845 17289 22879 17323
rect 23213 17289 23247 17323
rect 26249 17289 26283 17323
rect 27077 17289 27111 17323
rect 28733 17289 28767 17323
rect 29469 17289 29503 17323
rect 32137 17289 32171 17323
rect 33609 17289 33643 17323
rect 13798 17221 13832 17255
rect 23305 17221 23339 17255
rect 27598 17221 27632 17255
rect 2053 17153 2087 17187
rect 4169 17153 4203 17187
rect 6009 17153 6043 17187
rect 9956 17153 9990 17187
rect 11529 17153 11563 17187
rect 11796 17153 11830 17187
rect 13461 17153 13495 17187
rect 13553 17153 13587 17187
rect 16221 17153 16255 17187
rect 16681 17153 16715 17187
rect 16948 17153 16982 17187
rect 21189 17153 21223 17187
rect 26433 17153 26467 17187
rect 27261 17153 27295 17187
rect 29653 17153 29687 17187
rect 32505 17153 32539 17187
rect 33977 17153 34011 17187
rect 36461 17153 36495 17187
rect 5089 17085 5123 17119
rect 6929 17085 6963 17119
rect 7021 17085 7055 17119
rect 9689 17085 9723 17119
rect 19349 17085 19383 17119
rect 19441 17085 19475 17119
rect 23397 17085 23431 17119
rect 27353 17085 27387 17119
rect 32597 17085 32631 17119
rect 32781 17085 32815 17119
rect 34069 17085 34103 17119
rect 34253 17085 34287 17119
rect 6469 16949 6503 16983
rect 16405 16949 16439 16983
rect 36277 16949 36311 16983
rect 11805 16745 11839 16779
rect 17233 16745 17267 16779
rect 27721 16745 27755 16779
rect 29745 16745 29779 16779
rect 32965 16745 32999 16779
rect 34529 16745 34563 16779
rect 8769 16677 8803 16711
rect 4261 16609 4295 16643
rect 4445 16609 4479 16643
rect 5917 16609 5951 16643
rect 7389 16609 7423 16643
rect 12725 16609 12759 16643
rect 14933 16609 14967 16643
rect 16957 16609 16991 16643
rect 23765 16609 23799 16643
rect 23949 16609 23983 16643
rect 28181 16609 28215 16643
rect 28365 16609 28399 16643
rect 30297 16609 30331 16643
rect 31033 16609 31067 16643
rect 31125 16609 31159 16643
rect 31585 16609 31619 16643
rect 33149 16609 33183 16643
rect 4813 16541 4847 16575
rect 8953 16541 8987 16575
rect 9137 16541 9171 16575
rect 11989 16541 12023 16575
rect 12449 16541 12483 16575
rect 17417 16541 17451 16575
rect 24869 16541 24903 16575
rect 28089 16541 28123 16575
rect 34897 16541 34931 16575
rect 6184 16473 6218 16507
rect 7656 16473 7690 16507
rect 15200 16473 15234 16507
rect 16773 16473 16807 16507
rect 23673 16473 23707 16507
rect 25136 16473 25170 16507
rect 30205 16473 30239 16507
rect 30941 16473 30975 16507
rect 31852 16473 31886 16507
rect 33416 16473 33450 16507
rect 3801 16405 3835 16439
rect 4169 16405 4203 16439
rect 4629 16405 4663 16439
rect 7297 16405 7331 16439
rect 9045 16405 9079 16439
rect 12081 16405 12115 16439
rect 12541 16405 12575 16439
rect 16313 16405 16347 16439
rect 16405 16405 16439 16439
rect 16865 16405 16899 16439
rect 23305 16405 23339 16439
rect 26249 16405 26283 16439
rect 30113 16405 30147 16439
rect 30573 16405 30607 16439
rect 34713 16405 34747 16439
rect 3801 16201 3835 16235
rect 6377 16201 6411 16235
rect 8217 16201 8251 16235
rect 10241 16201 10275 16235
rect 12265 16201 12299 16235
rect 13921 16201 13955 16235
rect 15301 16201 15335 16235
rect 19809 16201 19843 16235
rect 21557 16201 21591 16235
rect 22661 16201 22695 16235
rect 24317 16201 24351 16235
rect 25789 16201 25823 16235
rect 26341 16201 26375 16235
rect 28917 16201 28951 16235
rect 30573 16201 30607 16235
rect 31769 16201 31803 16235
rect 32137 16201 32171 16235
rect 32505 16201 32539 16235
rect 32965 16201 32999 16235
rect 33793 16201 33827 16235
rect 34161 16201 34195 16235
rect 4620 16133 4654 16167
rect 8033 16133 8067 16167
rect 12786 16133 12820 16167
rect 23182 16133 23216 16167
rect 25697 16133 25731 16167
rect 29438 16133 29472 16167
rect 33425 16133 33459 16167
rect 34253 16133 34287 16167
rect 1409 16065 1443 16099
rect 2421 16065 2455 16099
rect 2688 16065 2722 16099
rect 4353 16065 4387 16099
rect 6561 16065 6595 16099
rect 8309 16065 8343 16099
rect 8861 16065 8895 16099
rect 9128 16065 9162 16099
rect 10333 16065 10367 16099
rect 10517 16065 10551 16099
rect 12449 16065 12483 16099
rect 12541 16065 12575 16099
rect 15485 16065 15519 16099
rect 17601 16065 17635 16099
rect 18429 16065 18463 16099
rect 18696 16065 18730 16099
rect 20433 16065 20467 16099
rect 22845 16065 22879 16099
rect 25973 16065 26007 16099
rect 26525 16065 26559 16099
rect 29101 16065 29135 16099
rect 31953 16065 31987 16099
rect 33333 16065 33367 16099
rect 20177 15997 20211 16031
rect 22937 15997 22971 16031
rect 29193 15997 29227 16031
rect 32597 15997 32631 16031
rect 32689 15997 32723 16031
rect 33609 15997 33643 16031
rect 34345 15997 34379 16031
rect 8033 15929 8067 15963
rect 1593 15861 1627 15895
rect 5733 15861 5767 15895
rect 10333 15861 10367 15895
rect 17785 15861 17819 15895
rect 26157 15861 26191 15895
rect 2881 15657 2915 15691
rect 4813 15657 4847 15691
rect 9045 15657 9079 15691
rect 12909 15657 12943 15691
rect 18705 15657 18739 15691
rect 20085 15657 20119 15691
rect 22109 15657 22143 15691
rect 23673 15657 23707 15691
rect 26985 15657 27019 15691
rect 28825 15657 28859 15691
rect 29745 15657 29779 15691
rect 16129 15589 16163 15623
rect 27813 15589 27847 15623
rect 5365 15521 5399 15555
rect 13553 15521 13587 15555
rect 16773 15521 16807 15555
rect 19809 15521 19843 15555
rect 27537 15521 27571 15555
rect 28457 15521 28491 15555
rect 30205 15521 30239 15555
rect 30297 15521 30331 15555
rect 3065 15453 3099 15487
rect 5181 15453 5215 15487
rect 9045 15453 9079 15487
rect 9321 15453 9355 15487
rect 10517 15453 10551 15487
rect 10793 15453 10827 15487
rect 13277 15453 13311 15487
rect 18889 15453 18923 15487
rect 19625 15453 19659 15487
rect 20269 15453 20303 15487
rect 20637 15453 20671 15487
rect 20729 15453 20763 15487
rect 22293 15453 22327 15487
rect 24593 15453 24627 15487
rect 27353 15453 27387 15487
rect 28641 15453 28675 15487
rect 30113 15453 30147 15487
rect 13369 15385 13403 15419
rect 19717 15385 19751 15419
rect 20974 15385 21008 15419
rect 22538 15385 22572 15419
rect 24860 15385 24894 15419
rect 5273 15317 5307 15351
rect 9229 15317 9263 15351
rect 11529 15317 11563 15351
rect 16497 15317 16531 15351
rect 16589 15317 16623 15351
rect 19257 15317 19291 15351
rect 20453 15317 20487 15351
rect 25973 15317 26007 15351
rect 27445 15317 27479 15351
rect 28181 15317 28215 15351
rect 28273 15317 28307 15351
rect 6377 15113 6411 15147
rect 6745 15113 6779 15147
rect 16497 15113 16531 15147
rect 16681 15113 16715 15147
rect 25145 15113 25179 15147
rect 33609 15113 33643 15147
rect 4445 15045 4479 15079
rect 15384 15045 15418 15079
rect 25513 15045 25547 15079
rect 4537 14977 4571 15011
rect 5549 14977 5583 15011
rect 7849 14977 7883 15011
rect 8125 14977 8159 15011
rect 13829 14977 13863 15011
rect 14105 14977 14139 15011
rect 15117 14977 15151 15011
rect 16865 14977 16899 15011
rect 17601 14977 17635 15011
rect 22569 14977 22603 15011
rect 25329 14977 25363 15011
rect 25605 14977 25639 15011
rect 27445 14977 27479 15011
rect 31861 14977 31895 15011
rect 34253 14977 34287 15011
rect 4721 14909 4755 14943
rect 6837 14909 6871 14943
rect 6929 14909 6963 14943
rect 17325 14909 17359 14943
rect 27537 14909 27571 14943
rect 27629 14909 27663 14943
rect 33701 14909 33735 14943
rect 33793 14909 33827 14943
rect 4077 14773 4111 14807
rect 5365 14773 5399 14807
rect 8861 14773 8895 14807
rect 14841 14773 14875 14807
rect 18337 14773 18371 14807
rect 22385 14773 22419 14807
rect 27077 14773 27111 14807
rect 31677 14773 31711 14807
rect 33241 14773 33275 14807
rect 34069 14773 34103 14807
rect 6469 14569 6503 14603
rect 9873 14569 9907 14603
rect 19257 14569 19291 14603
rect 22293 14569 22327 14603
rect 27905 14569 27939 14603
rect 11713 14501 11747 14535
rect 30573 14501 30607 14535
rect 30757 14501 30791 14535
rect 34345 14501 34379 14535
rect 10241 14433 10275 14467
rect 19717 14433 19751 14467
rect 19809 14433 19843 14467
rect 21005 14433 21039 14467
rect 22937 14433 22971 14467
rect 26525 14433 26559 14467
rect 29561 14433 29595 14467
rect 31309 14433 31343 14467
rect 33333 14433 33367 14467
rect 3985 14365 4019 14399
rect 5089 14365 5123 14399
rect 5356 14365 5390 14399
rect 7113 14365 7147 14399
rect 7389 14365 7423 14399
rect 9781 14365 9815 14399
rect 10517 14365 10551 14399
rect 10701 14365 10735 14399
rect 12081 14365 12115 14399
rect 12173 14365 12207 14399
rect 13645 14365 13679 14399
rect 14105 14365 14139 14399
rect 15485 14365 15519 14399
rect 15761 14365 15795 14399
rect 18521 14365 18555 14399
rect 25421 14365 25455 14399
rect 25697 14365 25731 14399
rect 29377 14365 29411 14399
rect 29837 14365 29871 14399
rect 31585 14365 31619 14399
rect 31861 14365 31895 14399
rect 33241 14365 33275 14399
rect 33609 14365 33643 14399
rect 36185 14365 36219 14399
rect 11437 14297 11471 14331
rect 14289 14297 14323 14331
rect 22753 14297 22787 14331
rect 24501 14297 24535 14331
rect 26792 14297 26826 14331
rect 31125 14297 31159 14331
rect 3801 14229 3835 14263
rect 8125 14229 8159 14263
rect 10701 14229 10735 14263
rect 11897 14229 11931 14263
rect 12357 14229 12391 14263
rect 13737 14229 13771 14263
rect 14473 14229 14507 14263
rect 16497 14229 16531 14263
rect 18337 14229 18371 14263
rect 19625 14229 19659 14263
rect 20453 14229 20487 14263
rect 20821 14229 20855 14263
rect 20913 14229 20947 14263
rect 22661 14229 22695 14263
rect 24593 14229 24627 14263
rect 26433 14229 26467 14263
rect 29193 14229 29227 14263
rect 31217 14229 31251 14263
rect 32597 14229 32631 14263
rect 33057 14229 33091 14263
rect 36369 14229 36403 14263
rect 4537 14025 4571 14059
rect 7941 14025 7975 14059
rect 10609 14025 10643 14059
rect 11161 14025 11195 14059
rect 19349 14025 19383 14059
rect 21373 14025 21407 14059
rect 23397 14025 23431 14059
rect 23857 14025 23891 14059
rect 25697 14025 25731 14059
rect 26985 14025 27019 14059
rect 29561 14025 29595 14059
rect 29929 14025 29963 14059
rect 30573 14025 30607 14059
rect 33149 14025 33183 14059
rect 33517 14025 33551 14059
rect 3424 13957 3458 13991
rect 12541 13957 12575 13991
rect 13185 13957 13219 13991
rect 22284 13957 22318 13991
rect 24378 13957 24412 13991
rect 3157 13889 3191 13923
rect 6929 13889 6963 13923
rect 7205 13889 7239 13923
rect 8401 13889 8435 13923
rect 8585 13889 8619 13923
rect 9321 13889 9355 13923
rect 10149 13889 10183 13923
rect 10701 13889 10735 13923
rect 12173 13889 12207 13923
rect 12357 13889 12391 13923
rect 13093 13889 13127 13923
rect 13277 13889 13311 13923
rect 13553 13889 13587 13923
rect 13718 13889 13752 13923
rect 13829 13889 13863 13923
rect 13921 13889 13955 13923
rect 14013 13889 14047 13923
rect 14289 13889 14323 13923
rect 14473 13889 14507 13923
rect 14565 13889 14599 13923
rect 14749 13889 14783 13923
rect 17969 13889 18003 13923
rect 18236 13889 18270 13923
rect 19993 13889 20027 13923
rect 20260 13889 20294 13923
rect 21649 13889 21683 13923
rect 24041 13889 24075 13923
rect 24133 13889 24167 13923
rect 25881 13889 25915 13923
rect 27169 13889 27203 13923
rect 28457 13889 28491 13923
rect 29285 13889 29319 13923
rect 30757 13889 30791 13923
rect 31125 13889 31159 13923
rect 31953 13889 31987 13923
rect 9505 13821 9539 13855
rect 11529 13821 11563 13855
rect 11713 13821 11747 13855
rect 11897 13821 11931 13855
rect 13001 13821 13035 13855
rect 14933 13821 14967 13855
rect 22017 13821 22051 13855
rect 28181 13821 28215 13855
rect 30021 13821 30055 13855
rect 30113 13821 30147 13855
rect 30849 13821 30883 13855
rect 33609 13821 33643 13855
rect 33701 13821 33735 13855
rect 10977 13753 11011 13787
rect 12817 13753 12851 13787
rect 25513 13753 25547 13787
rect 8493 13685 8527 13719
rect 10241 13685 10275 13719
rect 13369 13685 13403 13719
rect 14289 13685 14323 13719
rect 21465 13685 21499 13719
rect 16405 13481 16439 13515
rect 17877 13481 17911 13515
rect 19257 13481 19291 13515
rect 20269 13481 20303 13515
rect 20729 13481 20763 13515
rect 22293 13481 22327 13515
rect 24409 13481 24443 13515
rect 28917 13481 28951 13515
rect 30941 13481 30975 13515
rect 8125 13413 8159 13447
rect 10333 13413 10367 13447
rect 28089 13413 28123 13447
rect 10517 13345 10551 13379
rect 11713 13345 11747 13379
rect 11989 13345 12023 13379
rect 15393 13345 15427 13379
rect 16497 13345 16531 13379
rect 18429 13345 18463 13379
rect 19717 13345 19751 13379
rect 19809 13345 19843 13379
rect 21189 13345 21223 13379
rect 21373 13345 21407 13379
rect 22937 13345 22971 13379
rect 24961 13345 24995 13379
rect 26341 13345 26375 13379
rect 28641 13345 28675 13379
rect 31493 13345 31527 13379
rect 33333 13345 33367 13379
rect 4445 13277 4479 13311
rect 4721 13277 4755 13311
rect 6009 13277 6043 13311
rect 6285 13277 6319 13311
rect 8401 13277 8435 13311
rect 10241 13277 10275 13311
rect 11621 13277 11655 13311
rect 15669 13277 15703 13311
rect 19625 13277 19659 13311
rect 20453 13277 20487 13311
rect 21097 13277 21131 13311
rect 22661 13277 22695 13311
rect 22753 13277 22787 13311
rect 24869 13277 24903 13311
rect 27169 13277 27203 13311
rect 29101 13277 29135 13311
rect 33057 13277 33091 13311
rect 8125 13209 8159 13243
rect 16764 13209 16798 13243
rect 18153 13209 18187 13243
rect 30573 13209 30607 13243
rect 31309 13209 31343 13243
rect 5457 13141 5491 13175
rect 7021 13141 7055 13175
rect 8309 13141 8343 13175
rect 10517 13141 10551 13175
rect 24777 13141 24811 13175
rect 25789 13141 25823 13175
rect 26157 13141 26191 13175
rect 26249 13141 26283 13175
rect 26985 13141 27019 13175
rect 28457 13141 28491 13175
rect 28549 13141 28583 13175
rect 31401 13141 31435 13175
rect 7573 12937 7607 12971
rect 8677 12937 8711 12971
rect 8769 12937 8803 12971
rect 8861 12937 8895 12971
rect 13645 12937 13679 12971
rect 13829 12937 13863 12971
rect 16681 12937 16715 12971
rect 25421 12937 25455 12971
rect 30297 12937 30331 12971
rect 32781 12937 32815 12971
rect 34069 12937 34103 12971
rect 36001 12937 36035 12971
rect 9781 12869 9815 12903
rect 15117 12869 15151 12903
rect 15853 12869 15887 12903
rect 1501 12801 1535 12835
rect 4997 12801 5031 12835
rect 5273 12801 5307 12835
rect 6653 12801 6687 12835
rect 7389 12801 7423 12835
rect 7573 12801 7607 12835
rect 8585 12801 8619 12835
rect 9413 12801 9447 12835
rect 9597 12801 9631 12835
rect 13277 12801 13311 12835
rect 13461 12801 13495 12835
rect 13737 12801 13771 12835
rect 14197 12801 14231 12835
rect 14933 12801 14967 12835
rect 15209 12801 15243 12835
rect 15301 12801 15335 12835
rect 15577 12801 15611 12835
rect 15761 12801 15795 12835
rect 15945 12801 15979 12835
rect 16865 12801 16899 12835
rect 25605 12801 25639 12835
rect 25973 12801 26007 12835
rect 26801 12801 26835 12835
rect 27261 12801 27295 12835
rect 29184 12801 29218 12835
rect 32965 12801 32999 12835
rect 33057 12801 33091 12835
rect 33333 12801 33367 12835
rect 34877 12801 34911 12835
rect 5641 12733 5675 12767
rect 6377 12733 6411 12767
rect 7665 12733 7699 12767
rect 7941 12733 7975 12767
rect 8953 12733 8987 12767
rect 14013 12733 14047 12767
rect 14105 12733 14139 12767
rect 14289 12733 14323 12767
rect 18245 12733 18279 12767
rect 25697 12733 25731 12767
rect 26985 12733 27019 12767
rect 28917 12733 28951 12767
rect 34621 12733 34655 12767
rect 15485 12665 15519 12699
rect 18613 12665 18647 12699
rect 1593 12597 1627 12631
rect 16129 12597 16163 12631
rect 18705 12597 18739 12631
rect 27997 12597 28031 12631
rect 9229 12393 9263 12427
rect 9505 12393 9539 12427
rect 11621 12393 11655 12427
rect 12541 12393 12575 12427
rect 18889 12393 18923 12427
rect 22937 12393 22971 12427
rect 25789 12393 25823 12427
rect 27077 12393 27111 12427
rect 29193 12393 29227 12427
rect 32965 12393 32999 12427
rect 34713 12393 34747 12427
rect 9597 12325 9631 12359
rect 11161 12325 11195 12359
rect 7757 12257 7791 12291
rect 9689 12257 9723 12291
rect 10149 12257 10183 12291
rect 10241 12257 10275 12291
rect 11805 12257 11839 12291
rect 12173 12257 12207 12291
rect 21281 12257 21315 12291
rect 23673 12257 23707 12291
rect 24409 12257 24443 12291
rect 27721 12257 27755 12291
rect 30021 12257 30055 12291
rect 30113 12257 30147 12291
rect 31493 12227 31527 12261
rect 33425 12257 33459 12291
rect 33517 12257 33551 12291
rect 4629 12189 4663 12223
rect 5733 12189 5767 12223
rect 6009 12189 6043 12223
rect 7113 12189 7147 12223
rect 7481 12189 7515 12223
rect 7941 12189 7975 12223
rect 9137 12189 9171 12223
rect 9321 12189 9355 12223
rect 9413 12189 9447 12223
rect 9781 12189 9815 12223
rect 9965 12189 9999 12223
rect 10517 12189 10551 12223
rect 11437 12189 11471 12223
rect 11529 12189 11563 12223
rect 12403 12189 12437 12223
rect 12633 12189 12667 12223
rect 15117 12189 15151 12223
rect 15301 12189 15335 12223
rect 15761 12189 15795 12223
rect 18245 12189 18279 12223
rect 18338 12189 18372 12223
rect 18710 12189 18744 12223
rect 19533 12189 19567 12223
rect 19681 12189 19715 12223
rect 19998 12189 20032 12223
rect 22753 12189 22787 12223
rect 23857 12189 23891 12223
rect 23949 12189 23983 12223
rect 24133 12189 24167 12223
rect 24225 12189 24259 12223
rect 27445 12189 27479 12223
rect 29377 12189 29411 12223
rect 31217 12189 31251 12223
rect 31309 12189 31343 12223
rect 31953 12189 31987 12223
rect 32137 12189 32171 12223
rect 34897 12189 34931 12223
rect 35173 12189 35207 12223
rect 7297 12121 7331 12155
rect 11161 12121 11195 12155
rect 11805 12121 11839 12155
rect 15945 12121 15979 12155
rect 17969 12121 18003 12155
rect 18153 12121 18187 12155
rect 18521 12121 18555 12155
rect 18613 12121 18647 12155
rect 19809 12121 19843 12155
rect 19901 12121 19935 12155
rect 21548 12121 21582 12155
rect 24654 12121 24688 12155
rect 33333 12121 33367 12155
rect 4997 12053 5031 12087
rect 8125 12053 8159 12087
rect 11345 12053 11379 12087
rect 15117 12053 15151 12087
rect 16129 12053 16163 12087
rect 20177 12053 20211 12087
rect 22661 12053 22695 12087
rect 27537 12053 27571 12087
rect 29561 12053 29595 12087
rect 29929 12053 29963 12087
rect 31493 12053 31527 12087
rect 32045 12053 32079 12087
rect 35081 12053 35115 12087
rect 7205 11849 7239 11883
rect 11805 11849 11839 11883
rect 12725 11849 12759 11883
rect 14381 11849 14415 11883
rect 18981 11849 19015 11883
rect 20085 11849 20119 11883
rect 21833 11849 21867 11883
rect 24501 11849 24535 11883
rect 7573 11781 7607 11815
rect 7665 11781 7699 11815
rect 9321 11781 9355 11815
rect 12081 11781 12115 11815
rect 15301 11781 15335 11815
rect 18153 11781 18187 11815
rect 18889 11781 18923 11815
rect 24225 11781 24259 11815
rect 3893 11713 3927 11747
rect 4169 11713 4203 11747
rect 6929 11713 6963 11747
rect 7021 11713 7055 11747
rect 7481 11713 7515 11747
rect 7849 11713 7883 11747
rect 7941 11713 7975 11747
rect 8493 11713 8527 11747
rect 10425 11713 10459 11747
rect 11713 11713 11747 11747
rect 12173 11713 12207 11747
rect 12357 11713 12391 11747
rect 12449 11713 12483 11747
rect 12541 11713 12575 11747
rect 13093 11713 13127 11747
rect 13829 11713 13863 11747
rect 14013 11713 14047 11747
rect 14105 11713 14139 11747
rect 14197 11713 14231 11747
rect 15485 11713 15519 11747
rect 15577 11713 15611 11747
rect 17049 11713 17083 11747
rect 17417 11713 17451 11747
rect 17969 11713 18003 11747
rect 19441 11713 19475 11747
rect 19589 11713 19623 11747
rect 19717 11713 19751 11747
rect 19809 11713 19843 11747
rect 19947 11713 19981 11747
rect 22017 11713 22051 11747
rect 22293 11713 22327 11747
rect 22477 11713 22511 11747
rect 23029 11713 23063 11747
rect 23765 11713 23799 11747
rect 23857 11713 23891 11747
rect 24317 11713 24351 11747
rect 24593 11713 24627 11747
rect 30297 11713 30331 11747
rect 30481 11713 30515 11747
rect 30941 11713 30975 11747
rect 31585 11713 31619 11747
rect 32229 11713 32263 11747
rect 33149 11713 33183 11747
rect 33241 11713 33275 11747
rect 33701 11713 33735 11747
rect 34989 11713 35023 11747
rect 35256 11713 35290 11747
rect 8217 11645 8251 11679
rect 8309 11645 8343 11679
rect 8401 11645 8435 11679
rect 10333 11645 10367 11679
rect 13277 11645 13311 11679
rect 18245 11645 18279 11679
rect 22569 11645 22603 11679
rect 22753 11645 22787 11679
rect 22845 11645 22879 11679
rect 22937 11645 22971 11679
rect 24133 11645 24167 11679
rect 31217 11645 31251 11679
rect 31769 11645 31803 11679
rect 33517 11645 33551 11679
rect 9689 11577 9723 11611
rect 11897 11577 11931 11611
rect 13737 11577 13771 11611
rect 18521 11577 18555 11611
rect 24041 11577 24075 11611
rect 24317 11577 24351 11611
rect 31677 11577 31711 11611
rect 33333 11577 33367 11611
rect 4905 11509 4939 11543
rect 7297 11509 7331 11543
rect 8033 11509 8067 11543
rect 9781 11509 9815 11543
rect 10793 11509 10827 11543
rect 11989 11509 12023 11543
rect 15301 11509 15335 11543
rect 18705 11509 18739 11543
rect 30297 11509 30331 11543
rect 32321 11509 32355 11543
rect 33885 11509 33919 11543
rect 36369 11509 36403 11543
rect 7205 11305 7239 11339
rect 7573 11305 7607 11339
rect 12265 11305 12299 11339
rect 16773 11305 16807 11339
rect 19809 11305 19843 11339
rect 22293 11305 22327 11339
rect 22477 11305 22511 11339
rect 23489 11305 23523 11339
rect 31309 11305 31343 11339
rect 36277 11305 36311 11339
rect 9413 11237 9447 11271
rect 14289 11237 14323 11271
rect 7389 11169 7423 11203
rect 11621 11169 11655 11203
rect 17417 11169 17451 11203
rect 19533 11169 19567 11203
rect 21097 11169 21131 11203
rect 28825 11169 28859 11203
rect 7113 11101 7147 11135
rect 7481 11101 7515 11135
rect 9413 11101 9447 11135
rect 9689 11101 9723 11135
rect 11805 11101 11839 11135
rect 14565 11101 14599 11135
rect 14657 11101 14691 11135
rect 14749 11101 14783 11135
rect 14933 11101 14967 11135
rect 15209 11101 15243 11135
rect 18521 11101 18555 11135
rect 18705 11101 18739 11135
rect 18797 11101 18831 11135
rect 18889 11101 18923 11135
rect 19441 11101 19475 11135
rect 19630 11079 19664 11113
rect 19901 11101 19935 11135
rect 19993 11101 20027 11135
rect 20269 11101 20303 11135
rect 20453 11101 20487 11135
rect 20729 11101 20763 11135
rect 20913 11101 20947 11135
rect 23121 11101 23155 11135
rect 23305 11101 23339 11135
rect 26341 11101 26375 11135
rect 28089 11101 28123 11135
rect 28273 11101 28307 11135
rect 28549 11101 28583 11135
rect 28641 11101 28675 11135
rect 31033 11101 31067 11135
rect 31125 11101 31159 11135
rect 31861 11101 31895 11135
rect 31953 11101 31987 11135
rect 32045 11101 32079 11135
rect 32229 11101 32263 11135
rect 35265 11101 35299 11135
rect 36461 11101 36495 11135
rect 9597 11033 9631 11067
rect 19257 11033 19291 11067
rect 19533 11033 19567 11067
rect 22109 11033 22143 11067
rect 26525 11033 26559 11067
rect 15025 10965 15059 10999
rect 17141 10965 17175 10999
rect 17233 10965 17267 10999
rect 19073 10965 19107 10999
rect 22293 10965 22327 10999
rect 28457 10965 28491 10999
rect 28825 10965 28859 10999
rect 35081 10965 35115 10999
rect 7481 10761 7515 10795
rect 10241 10761 10275 10795
rect 14105 10761 14139 10795
rect 14473 10761 14507 10795
rect 14841 10761 14875 10795
rect 16313 10761 16347 10795
rect 18061 10761 18095 10795
rect 24777 10761 24811 10795
rect 28641 10761 28675 10795
rect 31493 10761 31527 10795
rect 36369 10761 36403 10795
rect 6009 10693 6043 10727
rect 16926 10693 16960 10727
rect 24869 10693 24903 10727
rect 25666 10693 25700 10727
rect 29285 10693 29319 10727
rect 34529 10693 34563 10727
rect 4997 10625 5031 10659
rect 5089 10625 5123 10659
rect 5181 10625 5215 10659
rect 5549 10625 5583 10659
rect 5733 10625 5767 10659
rect 5825 10625 5859 10659
rect 5917 10625 5951 10659
rect 7205 10625 7239 10659
rect 7297 10625 7331 10659
rect 10333 10625 10367 10659
rect 10701 10625 10735 10659
rect 13737 10625 13771 10659
rect 16497 10625 16531 10659
rect 21557 10625 21591 10659
rect 21925 10625 21959 10659
rect 24409 10625 24443 10659
rect 25053 10625 25087 10659
rect 25237 10625 25271 10659
rect 27629 10625 27663 10659
rect 27905 10625 27939 10659
rect 28273 10625 28307 10659
rect 28457 10625 28491 10659
rect 28825 10625 28859 10659
rect 28917 10625 28951 10659
rect 29193 10625 29227 10659
rect 29653 10625 29687 10659
rect 31309 10625 31343 10659
rect 31401 10625 31435 10659
rect 31677 10625 31711 10659
rect 32229 10625 32263 10659
rect 32689 10625 32723 10659
rect 33057 10625 33091 10659
rect 33609 10625 33643 10659
rect 33793 10625 33827 10659
rect 34069 10625 34103 10659
rect 34253 10625 34287 10659
rect 35245 10625 35279 10659
rect 5365 10557 5399 10591
rect 7481 10557 7515 10591
rect 10977 10557 11011 10591
rect 13829 10557 13863 10591
rect 14933 10557 14967 10591
rect 15025 10557 15059 10591
rect 16681 10557 16715 10591
rect 24501 10557 24535 10591
rect 25329 10557 25363 10591
rect 25421 10557 25455 10591
rect 28549 10557 28583 10591
rect 29469 10557 29503 10591
rect 31769 10557 31803 10591
rect 31953 10557 31987 10591
rect 32781 10557 32815 10591
rect 32965 10557 32999 10591
rect 33885 10557 33919 10591
rect 34989 10557 35023 10591
rect 5825 10489 5859 10523
rect 27905 10489 27939 10523
rect 29561 10489 29595 10523
rect 32321 10489 32355 10523
rect 13737 10421 13771 10455
rect 21373 10421 21407 10455
rect 22017 10421 22051 10455
rect 24593 10421 24627 10455
rect 26801 10421 26835 10455
rect 28089 10421 28123 10455
rect 29101 10421 29135 10455
rect 29469 10421 29503 10455
rect 31861 10421 31895 10455
rect 34621 10421 34655 10455
rect 6929 10217 6963 10251
rect 7941 10217 7975 10251
rect 12541 10217 12575 10251
rect 14105 10217 14139 10251
rect 15117 10217 15151 10251
rect 16773 10217 16807 10251
rect 17877 10217 17911 10251
rect 27813 10217 27847 10251
rect 28733 10217 28767 10251
rect 33241 10217 33275 10251
rect 6469 10149 6503 10183
rect 7665 10149 7699 10183
rect 22753 10149 22787 10183
rect 26157 10149 26191 10183
rect 29837 10149 29871 10183
rect 34437 10149 34471 10183
rect 5917 10081 5951 10115
rect 7113 10081 7147 10115
rect 8953 10081 8987 10115
rect 11713 10081 11747 10115
rect 14749 10081 14783 10115
rect 17325 10081 17359 10115
rect 19257 10081 19291 10115
rect 21557 10081 21591 10115
rect 21833 10081 21867 10115
rect 21925 10081 21959 10115
rect 24777 10081 24811 10115
rect 28917 10081 28951 10115
rect 30481 10081 30515 10115
rect 31493 10081 31527 10115
rect 33425 10081 33459 10115
rect 33517 10081 33551 10115
rect 33977 10081 34011 10115
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 4077 10013 4111 10047
rect 4261 10013 4295 10047
rect 4445 10013 4479 10047
rect 4721 10013 4755 10047
rect 6101 10013 6135 10047
rect 6377 10013 6411 10047
rect 6745 10013 6779 10047
rect 6837 10013 6871 10047
rect 7205 10013 7239 10047
rect 7389 10013 7423 10047
rect 7757 10013 7791 10047
rect 7849 10013 7883 10047
rect 12357 10013 12391 10047
rect 12449 10013 12483 10047
rect 13553 10013 13587 10047
rect 13645 10013 13679 10047
rect 14289 10013 14323 10047
rect 14933 10013 14967 10047
rect 17141 10013 17175 10047
rect 18153 10013 18187 10047
rect 20913 10013 20947 10047
rect 21097 10013 21131 10047
rect 21373 10013 21407 10047
rect 22569 10013 22603 10047
rect 22753 10013 22787 10047
rect 22937 10013 22971 10047
rect 23121 10013 23155 10047
rect 23213 10013 23247 10047
rect 23489 10013 23523 10047
rect 24409 10013 24443 10047
rect 26985 10013 27019 10047
rect 27169 10013 27203 10047
rect 27353 10013 27387 10047
rect 27537 10013 27571 10047
rect 28641 10013 28675 10047
rect 30113 10013 30147 10047
rect 30205 10013 30239 10047
rect 31125 10013 31159 10047
rect 31953 10013 31987 10047
rect 32413 10013 32447 10047
rect 32597 10013 32631 10047
rect 32689 10013 32723 10047
rect 32781 10013 32815 10047
rect 32965 10013 32999 10047
rect 33609 10013 33643 10047
rect 33701 10013 33735 10047
rect 34069 10013 34103 10047
rect 34805 10013 34839 10047
rect 1501 9945 1535 9979
rect 3893 9945 3927 9979
rect 4537 9945 4571 9979
rect 4905 9945 4939 9979
rect 5089 9945 5123 9979
rect 5273 9945 5307 9979
rect 6469 9945 6503 9979
rect 11897 9945 11931 9979
rect 12265 9945 12299 9979
rect 17785 9945 17819 9979
rect 19524 9945 19558 9979
rect 20729 9945 20763 9979
rect 21005 9945 21039 9979
rect 21235 9945 21269 9979
rect 22042 9945 22076 9979
rect 25044 9945 25078 9979
rect 27721 9945 27755 9979
rect 28917 9945 28951 9979
rect 29837 9945 29871 9979
rect 1593 9877 1627 9911
rect 6285 9877 6319 9911
rect 6653 9877 6687 9911
rect 7113 9877 7147 9911
rect 8309 9877 8343 9911
rect 9183 9877 9217 9911
rect 11989 9877 12023 9911
rect 12081 9877 12115 9911
rect 12725 9877 12759 9911
rect 13553 9877 13587 9911
rect 17233 9877 17267 9911
rect 18245 9877 18279 9911
rect 20637 9877 20671 9911
rect 22201 9877 22235 9911
rect 23029 9877 23063 9911
rect 24593 9877 24627 9911
rect 30021 9877 30055 9911
rect 31309 9877 31343 9911
rect 31769 9877 31803 9911
rect 31861 9877 31895 9911
rect 33149 9877 33183 9911
rect 34897 9877 34931 9911
rect 6469 9673 6503 9707
rect 11989 9673 12023 9707
rect 15117 9673 15151 9707
rect 19349 9673 19383 9707
rect 21557 9673 21591 9707
rect 26157 9673 26191 9707
rect 32689 9673 32723 9707
rect 33793 9673 33827 9707
rect 5365 9605 5399 9639
rect 10057 9605 10091 9639
rect 12909 9605 12943 9639
rect 30113 9605 30147 9639
rect 30205 9605 30239 9639
rect 33241 9605 33275 9639
rect 5089 9537 5123 9571
rect 5181 9537 5215 9571
rect 6377 9537 6411 9571
rect 6745 9537 6779 9571
rect 8309 9537 8343 9571
rect 8953 9537 8987 9571
rect 9413 9537 9447 9571
rect 9597 9537 9631 9571
rect 9689 9537 9723 9571
rect 9781 9537 9815 9571
rect 10517 9537 10551 9571
rect 10701 9537 10735 9571
rect 10793 9537 10827 9571
rect 10885 9537 10919 9571
rect 11529 9537 11563 9571
rect 11805 9537 11839 9571
rect 12633 9537 12667 9571
rect 12817 9537 12851 9571
rect 13006 9537 13040 9571
rect 15301 9537 15335 9571
rect 16681 9537 16715 9571
rect 18236 9537 18270 9571
rect 20913 9537 20947 9571
rect 21373 9537 21407 9571
rect 23581 9537 23615 9571
rect 23949 9537 23983 9571
rect 24225 9537 24259 9571
rect 24685 9537 24719 9571
rect 25145 9537 25179 9571
rect 25881 9537 25915 9571
rect 25973 9537 26007 9571
rect 30021 9537 30055 9571
rect 30389 9537 30423 9571
rect 30481 9537 30515 9571
rect 30573 9537 30607 9571
rect 30757 9537 30791 9571
rect 32321 9537 32355 9571
rect 32597 9537 32631 9571
rect 33517 9537 33551 9571
rect 34161 9537 34195 9571
rect 5365 9469 5399 9503
rect 6561 9469 6595 9503
rect 8585 9469 8619 9503
rect 9045 9469 9079 9503
rect 10057 9469 10091 9503
rect 11897 9469 11931 9503
rect 12909 9469 12943 9503
rect 17969 9469 18003 9503
rect 21189 9469 21223 9503
rect 22385 9469 22419 9503
rect 22661 9469 22695 9503
rect 25513 9469 25547 9503
rect 33333 9469 33367 9503
rect 34253 9469 34287 9503
rect 34345 9469 34379 9503
rect 6745 9401 6779 9435
rect 8401 9401 8435 9435
rect 9413 9401 9447 9435
rect 9873 9401 9907 9435
rect 16865 9401 16899 9435
rect 23765 9401 23799 9435
rect 32413 9401 32447 9435
rect 8493 9333 8527 9367
rect 9321 9333 9355 9367
rect 11069 9333 11103 9367
rect 11621 9333 11655 9367
rect 21097 9333 21131 9367
rect 29837 9333 29871 9367
rect 30573 9333 30607 9367
rect 30941 9333 30975 9367
rect 32137 9333 32171 9367
rect 32505 9333 32539 9367
rect 33425 9333 33459 9367
rect 33701 9333 33735 9367
rect 4629 9129 4663 9163
rect 10977 9129 11011 9163
rect 13001 9129 13035 9163
rect 13369 9129 13403 9163
rect 14473 9129 14507 9163
rect 14841 9129 14875 9163
rect 23121 9129 23155 9163
rect 23581 9129 23615 9163
rect 23673 9129 23707 9163
rect 24041 9129 24075 9163
rect 10517 9061 10551 9095
rect 16497 9061 16531 9095
rect 27537 9061 27571 9095
rect 11253 8993 11287 9027
rect 16129 8993 16163 9027
rect 21373 8993 21407 9027
rect 22753 8993 22787 9027
rect 22937 8993 22971 9027
rect 4445 8925 4479 8959
rect 10425 8925 10459 8959
rect 10609 8925 10643 8959
rect 11161 8925 11195 8959
rect 11345 8925 11379 8959
rect 11437 8925 11471 8959
rect 11621 8925 11655 8959
rect 12909 8925 12943 8959
rect 14381 8925 14415 8959
rect 15853 8925 15887 8959
rect 16589 8925 16623 8959
rect 16865 8925 16899 8959
rect 17325 8925 17359 8959
rect 17592 8925 17626 8959
rect 21649 8925 21683 8959
rect 22385 8925 22419 8959
rect 22569 8925 22603 8959
rect 23029 8925 23063 8959
rect 23397 8925 23431 8959
rect 23673 8925 23707 8959
rect 23857 8925 23891 8959
rect 27813 8925 27847 8959
rect 27905 8925 27939 8959
rect 27998 8925 28032 8959
rect 28370 8925 28404 8959
rect 30389 8925 30423 8959
rect 16313 8857 16347 8891
rect 16681 8857 16715 8891
rect 17049 8857 17083 8891
rect 27537 8857 27571 8891
rect 27721 8857 27755 8891
rect 28181 8857 28215 8891
rect 28273 8857 28307 8891
rect 4905 8789 4939 8823
rect 15485 8789 15519 8823
rect 15945 8789 15979 8823
rect 16405 8789 16439 8823
rect 18705 8789 18739 8823
rect 28549 8789 28583 8823
rect 30481 8789 30515 8823
rect 10425 8585 10459 8619
rect 13829 8585 13863 8619
rect 15945 8585 15979 8619
rect 23949 8585 23983 8619
rect 26801 8585 26835 8619
rect 29393 8585 29427 8619
rect 32337 8585 32371 8619
rect 34161 8585 34195 8619
rect 17141 8517 17175 8551
rect 29193 8517 29227 8551
rect 32137 8517 32171 8551
rect 32597 8517 32631 8551
rect 34069 8517 34103 8551
rect 34437 8517 34471 8551
rect 7113 8449 7147 8483
rect 7297 8449 7331 8483
rect 9781 8449 9815 8483
rect 12541 8449 12575 8483
rect 12817 8449 12851 8483
rect 13005 8471 13039 8505
rect 13369 8449 13403 8483
rect 14013 8449 14047 8483
rect 14832 8449 14866 8483
rect 16957 8449 16991 8483
rect 17233 8449 17267 8483
rect 21097 8449 21131 8483
rect 21281 8449 21315 8483
rect 21833 8449 21867 8483
rect 22201 8449 22235 8483
rect 22569 8449 22603 8483
rect 23857 8449 23891 8483
rect 24409 8449 24443 8483
rect 26525 8449 26559 8483
rect 27353 8449 27387 8483
rect 27721 8449 27755 8483
rect 27905 8449 27939 8483
rect 28365 8449 28399 8483
rect 28825 8449 28859 8483
rect 32781 8449 32815 8483
rect 32873 8449 32907 8483
rect 9965 8381 9999 8415
rect 14289 8381 14323 8415
rect 14381 8381 14415 8415
rect 14565 8381 14599 8415
rect 24133 8381 24167 8415
rect 26801 8381 26835 8415
rect 12633 8313 12667 8347
rect 12725 8313 12759 8347
rect 13645 8313 13679 8347
rect 17233 8313 17267 8347
rect 21097 8313 21131 8347
rect 21925 8313 21959 8347
rect 26617 8313 26651 8347
rect 27445 8313 27479 8347
rect 32597 8313 32631 8347
rect 34621 8313 34655 8347
rect 7113 8245 7147 8279
rect 12357 8245 12391 8279
rect 29377 8245 29411 8279
rect 29561 8245 29595 8279
rect 32321 8245 32355 8279
rect 32505 8245 32539 8279
rect 6193 8041 6227 8075
rect 10517 8041 10551 8075
rect 10977 8041 11011 8075
rect 11345 8041 11379 8075
rect 13829 8041 13863 8075
rect 15117 8041 15151 8075
rect 17877 8041 17911 8075
rect 18889 8041 18923 8075
rect 19073 8041 19107 8075
rect 25881 8041 25915 8075
rect 26617 8041 26651 8075
rect 27629 8041 27663 8075
rect 30205 8041 30239 8075
rect 33517 8041 33551 8075
rect 8033 7973 8067 8007
rect 21465 7973 21499 8007
rect 26433 7973 26467 8007
rect 27353 7973 27387 8007
rect 28089 7973 28123 8007
rect 30849 7973 30883 8007
rect 32781 7973 32815 8007
rect 4721 7905 4755 7939
rect 7113 7905 7147 7939
rect 7573 7905 7607 7939
rect 7849 7905 7883 7939
rect 8217 7905 8251 7939
rect 12173 7905 12207 7939
rect 17509 7905 17543 7939
rect 20913 7905 20947 7939
rect 21097 7905 21131 7939
rect 27629 7905 27663 7939
rect 30389 7905 30423 7939
rect 30573 7905 30607 7939
rect 30665 7905 30699 7939
rect 31033 7905 31067 7939
rect 31493 7905 31527 7939
rect 33149 7905 33183 7939
rect 4445 7837 4479 7871
rect 4629 7837 4663 7871
rect 4905 7837 4939 7871
rect 5089 7837 5123 7871
rect 5181 7837 5215 7871
rect 5273 7837 5307 7871
rect 5549 7837 5583 7871
rect 5825 7837 5859 7871
rect 5917 7837 5951 7871
rect 6101 7837 6135 7871
rect 6377 7837 6411 7871
rect 6653 7837 6687 7871
rect 6837 7837 6871 7871
rect 7205 7837 7239 7871
rect 7665 7837 7699 7871
rect 7757 7837 7791 7871
rect 8033 7837 8067 7871
rect 8125 7837 8159 7871
rect 8309 7837 8343 7871
rect 8401 7837 8435 7871
rect 8585 7837 8619 7871
rect 9873 7837 9907 7871
rect 10057 7837 10091 7871
rect 10885 7837 10919 7871
rect 11897 7837 11931 7871
rect 12081 7837 12115 7871
rect 13737 7837 13771 7871
rect 14105 7837 14139 7871
rect 14381 7837 14415 7871
rect 15301 7837 15335 7871
rect 17233 7837 17267 7871
rect 18429 7837 18463 7871
rect 18521 7837 18555 7871
rect 18889 7837 18923 7871
rect 19257 7837 19291 7871
rect 20821 7837 20855 7871
rect 21465 7837 21499 7871
rect 21649 7837 21683 7871
rect 21833 7837 21867 7871
rect 22753 7837 22787 7871
rect 22845 7837 22879 7871
rect 23121 7837 23155 7871
rect 23949 7837 23983 7871
rect 24501 7837 24535 7871
rect 27261 7837 27295 7871
rect 27445 7837 27479 7871
rect 27537 7837 27571 7871
rect 28365 7837 28399 7871
rect 28549 7837 28583 7871
rect 29929 7837 29963 7871
rect 30021 7837 30055 7871
rect 30297 7837 30331 7871
rect 30757 7837 30791 7871
rect 31125 7837 31159 7871
rect 31217 7837 31251 7871
rect 31309 7837 31343 7871
rect 31677 7837 31711 7871
rect 31769 7837 31803 7871
rect 32045 7837 32079 7871
rect 32137 7837 32171 7871
rect 32597 7837 32631 7871
rect 33333 7837 33367 7871
rect 33609 7837 33643 7871
rect 34713 7837 34747 7871
rect 34969 7837 35003 7871
rect 36461 7837 36495 7871
rect 5457 7769 5491 7803
rect 7481 7769 7515 7803
rect 11989 7769 12023 7803
rect 17718 7769 17752 7803
rect 19524 7769 19558 7803
rect 24746 7769 24780 7803
rect 26157 7769 26191 7803
rect 29193 7769 29227 7803
rect 30459 7769 30493 7803
rect 32229 7769 32263 7803
rect 32505 7769 32539 7803
rect 33793 7769 33827 7803
rect 4629 7701 4663 7735
rect 5365 7701 5399 7735
rect 6929 7701 6963 7735
rect 8493 7701 8527 7735
rect 12403 7701 12437 7735
rect 17601 7701 17635 7735
rect 20637 7701 20671 7735
rect 21741 7701 21775 7735
rect 22569 7701 22603 7735
rect 27905 7701 27939 7735
rect 28273 7701 28307 7735
rect 29285 7701 29319 7735
rect 29745 7701 29779 7735
rect 31953 7701 31987 7735
rect 32413 7701 32447 7735
rect 33885 7701 33919 7735
rect 36093 7701 36127 7735
rect 36277 7701 36311 7735
rect 7205 7497 7239 7531
rect 7849 7497 7883 7531
rect 10057 7497 10091 7531
rect 10333 7497 10367 7531
rect 11805 7497 11839 7531
rect 13737 7497 13771 7531
rect 19993 7497 20027 7531
rect 21005 7497 21039 7531
rect 23121 7497 23155 7531
rect 23489 7497 23523 7531
rect 24133 7497 24167 7531
rect 27445 7497 27479 7531
rect 29929 7497 29963 7531
rect 30757 7497 30791 7531
rect 33517 7497 33551 7531
rect 6009 7429 6043 7463
rect 7481 7429 7515 7463
rect 16948 7429 16982 7463
rect 21925 7429 21959 7463
rect 23581 7429 23615 7463
rect 25228 7429 25262 7463
rect 30021 7429 30055 7463
rect 31861 7429 31895 7463
rect 33885 7429 33919 7463
rect 34253 7429 34287 7463
rect 34897 7429 34931 7463
rect 5917 7361 5951 7395
rect 6101 7361 6135 7395
rect 7113 7361 7147 7395
rect 7389 7361 7423 7395
rect 7757 7361 7791 7395
rect 7941 7361 7975 7395
rect 10241 7361 10275 7395
rect 10517 7361 10551 7395
rect 11989 7361 12023 7395
rect 12357 7361 12391 7395
rect 12633 7361 12667 7395
rect 13277 7361 13311 7395
rect 14381 7361 14415 7395
rect 19901 7361 19935 7395
rect 20085 7361 20119 7395
rect 21189 7361 21223 7395
rect 21373 7361 21407 7395
rect 21465 7361 21499 7395
rect 21649 7361 21683 7395
rect 22109 7361 22143 7395
rect 22201 7361 22235 7395
rect 22293 7361 22327 7395
rect 22385 7361 22419 7395
rect 24133 7361 24167 7395
rect 24409 7361 24443 7395
rect 24593 7361 24627 7395
rect 29101 7361 29135 7395
rect 30481 7361 30515 7395
rect 31033 7361 31067 7395
rect 31217 7361 31251 7395
rect 31493 7361 31527 7395
rect 31953 7361 31987 7395
rect 32321 7361 32355 7395
rect 32413 7361 32447 7395
rect 32689 7361 32723 7395
rect 33701 7361 33735 7395
rect 33793 7361 33827 7395
rect 34069 7361 34103 7395
rect 34161 7361 34195 7395
rect 34437 7361 34471 7395
rect 34529 7361 34563 7395
rect 34621 7361 34655 7395
rect 7297 7293 7331 7327
rect 14105 7293 14139 7327
rect 16681 7293 16715 7327
rect 23765 7293 23799 7327
rect 24225 7293 24259 7327
rect 24961 7293 24995 7327
rect 26985 7293 27019 7327
rect 30113 7293 30147 7327
rect 30757 7293 30791 7327
rect 31631 7293 31665 7327
rect 32597 7293 32631 7327
rect 34713 7293 34747 7327
rect 34897 7293 34931 7327
rect 21281 7225 21315 7259
rect 27261 7225 27295 7259
rect 29193 7225 29227 7259
rect 31769 7225 31803 7259
rect 34253 7225 34287 7259
rect 13369 7157 13403 7191
rect 18061 7157 18095 7191
rect 24317 7157 24351 7191
rect 26341 7157 26375 7191
rect 29561 7157 29595 7191
rect 30573 7157 30607 7191
rect 31125 7157 31159 7191
rect 32137 7157 32171 7191
rect 10149 6953 10183 6987
rect 10425 6953 10459 6987
rect 11253 6953 11287 6987
rect 11437 6953 11471 6987
rect 23581 6953 23615 6987
rect 5733 6885 5767 6919
rect 5365 6817 5399 6851
rect 11529 6817 11563 6851
rect 15025 6817 15059 6851
rect 15209 6817 15243 6851
rect 18429 6817 18463 6851
rect 18777 6817 18811 6851
rect 21465 6817 21499 6851
rect 22385 6817 22419 6851
rect 31309 6817 31343 6851
rect 9965 6749 9999 6783
rect 10977 6749 11011 6783
rect 11805 6749 11839 6783
rect 14289 6749 14323 6783
rect 14933 6749 14967 6783
rect 18337 6749 18371 6783
rect 18521 6749 18555 6783
rect 18981 6749 19015 6783
rect 21649 6749 21683 6783
rect 21925 6749 21959 6783
rect 23397 6749 23431 6783
rect 25973 6749 26007 6783
rect 28917 6749 28951 6783
rect 29101 6749 29135 6783
rect 31401 6749 31435 6783
rect 31493 6749 31527 6783
rect 31585 6749 31619 6783
rect 33885 6749 33919 6783
rect 18153 6681 18187 6715
rect 18705 6681 18739 6715
rect 22017 6681 22051 6715
rect 22201 6681 22235 6715
rect 26157 6681 26191 6715
rect 5825 6613 5859 6647
rect 14105 6613 14139 6647
rect 14565 6613 14599 6647
rect 18889 6613 18923 6647
rect 21833 6613 21867 6647
rect 29101 6613 29135 6647
rect 31125 6613 31159 6647
rect 33977 6613 34011 6647
rect 5457 6409 5491 6443
rect 7573 6409 7607 6443
rect 10425 6409 10459 6443
rect 14565 6409 14599 6443
rect 15393 6409 15427 6443
rect 15485 6409 15519 6443
rect 17325 6409 17359 6443
rect 22661 6409 22695 6443
rect 23581 6409 23615 6443
rect 27813 6409 27847 6443
rect 1676 6341 1710 6375
rect 13452 6341 13486 6375
rect 15117 6341 15151 6375
rect 18521 6341 18555 6375
rect 19257 6341 19291 6375
rect 28365 6341 28399 6375
rect 1409 6273 1443 6307
rect 5181 6273 5215 6307
rect 5273 6273 5307 6307
rect 5733 6273 5767 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 7481 6273 7515 6307
rect 7665 6273 7699 6307
rect 7849 6273 7883 6307
rect 7941 6273 7975 6307
rect 8125 6273 8159 6307
rect 8217 6273 8251 6307
rect 8677 6273 8711 6307
rect 9965 6273 9999 6307
rect 11529 6273 11563 6307
rect 15301 6273 15335 6307
rect 15669 6273 15703 6307
rect 17233 6273 17267 6307
rect 17417 6273 17451 6307
rect 17601 6273 17635 6307
rect 18889 6273 18923 6307
rect 18981 6273 19015 6307
rect 20637 6273 20671 6307
rect 20821 6273 20855 6307
rect 22017 6273 22051 6307
rect 22109 6273 22143 6307
rect 22293 6273 22327 6307
rect 22385 6273 22419 6307
rect 22569 6273 22603 6307
rect 23397 6273 23431 6307
rect 23949 6273 23983 6307
rect 25329 6273 25363 6307
rect 25513 6273 25547 6307
rect 27629 6273 27663 6307
rect 27905 6273 27939 6307
rect 28181 6273 28215 6307
rect 28273 6273 28307 6307
rect 28549 6273 28583 6307
rect 28641 6273 28675 6307
rect 29469 6273 29503 6307
rect 31309 6273 31343 6307
rect 31401 6273 31435 6307
rect 31493 6273 31527 6307
rect 5457 6205 5491 6239
rect 5825 6205 5859 6239
rect 6469 6205 6503 6239
rect 8309 6205 8343 6239
rect 8953 6205 8987 6239
rect 11805 6205 11839 6239
rect 13185 6205 13219 6239
rect 17877 6205 17911 6239
rect 18705 6205 18739 6239
rect 18797 6205 18831 6239
rect 31217 6205 31251 6239
rect 6101 6137 6135 6171
rect 8585 6137 8619 6171
rect 8861 6137 8895 6171
rect 2789 6069 2823 6103
rect 8217 6069 8251 6103
rect 8769 6069 8803 6103
rect 10241 6069 10275 6103
rect 19349 6069 19383 6103
rect 20637 6069 20671 6103
rect 21833 6069 21867 6103
rect 23765 6069 23799 6103
rect 25329 6069 25363 6103
rect 27629 6069 27663 6103
rect 27997 6069 28031 6103
rect 29285 6069 29319 6103
rect 31033 6069 31067 6103
rect 1593 5865 1627 5899
rect 7573 5865 7607 5899
rect 8493 5865 8527 5899
rect 10701 5865 10735 5899
rect 11253 5865 11287 5899
rect 12173 5865 12207 5899
rect 12909 5865 12943 5899
rect 15853 5865 15887 5899
rect 21005 5865 21039 5899
rect 22937 5865 22971 5899
rect 24225 5865 24259 5899
rect 25697 5865 25731 5899
rect 27629 5865 27663 5899
rect 31585 5865 31619 5899
rect 31861 5865 31895 5899
rect 33609 5865 33643 5899
rect 8125 5797 8159 5831
rect 14749 5797 14783 5831
rect 17141 5797 17175 5831
rect 17877 5797 17911 5831
rect 24869 5797 24903 5831
rect 26525 5797 26559 5831
rect 10057 5729 10091 5763
rect 11437 5729 11471 5763
rect 17693 5729 17727 5763
rect 19441 5729 19475 5763
rect 26157 5729 26191 5763
rect 26617 5729 26651 5763
rect 27169 5729 27203 5763
rect 33701 5729 33735 5763
rect 1409 5661 1443 5695
rect 7297 5661 7331 5695
rect 7849 5661 7883 5695
rect 8677 5661 8711 5695
rect 8953 5661 8987 5695
rect 9137 5661 9171 5695
rect 9965 5661 9999 5695
rect 10241 5661 10275 5695
rect 10977 5661 11011 5695
rect 11529 5661 11563 5695
rect 11713 5661 11747 5695
rect 12265 5661 12299 5695
rect 12449 5661 12483 5695
rect 14933 5661 14967 5695
rect 15025 5661 15059 5695
rect 15117 5661 15151 5695
rect 15602 5661 15636 5695
rect 15853 5661 15887 5695
rect 16037 5661 16071 5695
rect 16773 5661 16807 5695
rect 18061 5661 18095 5695
rect 18245 5661 18279 5695
rect 19257 5661 19291 5695
rect 19717 5661 19751 5695
rect 19993 5661 20027 5695
rect 20177 5661 20211 5695
rect 20270 5661 20304 5695
rect 20545 5661 20579 5695
rect 20642 5661 20676 5695
rect 21189 5661 21223 5695
rect 21281 5661 21315 5695
rect 21465 5661 21499 5695
rect 21557 5661 21591 5695
rect 21833 5661 21867 5695
rect 21925 5661 21959 5695
rect 22199 5661 22233 5695
rect 23213 5661 23247 5695
rect 23489 5661 23523 5695
rect 24685 5661 24719 5695
rect 25881 5661 25915 5695
rect 25973 5661 26007 5695
rect 26249 5661 26283 5695
rect 26801 5661 26835 5695
rect 27629 5661 27663 5695
rect 27905 5661 27939 5695
rect 27997 5661 28031 5695
rect 29561 5661 29595 5695
rect 29817 5661 29851 5695
rect 31309 5661 31343 5695
rect 31401 5661 31435 5695
rect 31677 5661 31711 5695
rect 31769 5661 31803 5695
rect 32137 5661 32171 5695
rect 32229 5661 32263 5695
rect 32485 5661 32519 5695
rect 33977 5661 34011 5695
rect 8401 5593 8435 5627
rect 8585 5593 8619 5627
rect 14749 5593 14783 5627
rect 17141 5593 17175 5627
rect 17601 5593 17635 5627
rect 20453 5593 20487 5627
rect 26341 5593 26375 5627
rect 26709 5593 26743 5627
rect 26985 5593 27019 5627
rect 31861 5593 31895 5627
rect 7757 5525 7791 5559
rect 8309 5525 8343 5559
rect 9321 5525 9355 5559
rect 9781 5525 9815 5559
rect 15393 5525 15427 5559
rect 15485 5525 15519 5559
rect 15761 5525 15795 5559
rect 16865 5525 16899 5559
rect 19533 5525 19567 5559
rect 20821 5525 20855 5559
rect 21649 5525 21683 5559
rect 26433 5525 26467 5559
rect 27813 5525 27847 5559
rect 28089 5525 28123 5559
rect 30941 5525 30975 5559
rect 31125 5525 31159 5559
rect 31953 5525 31987 5559
rect 7665 5321 7699 5355
rect 9229 5321 9263 5355
rect 10517 5321 10551 5355
rect 12265 5321 12299 5355
rect 12541 5321 12575 5355
rect 17509 5321 17543 5355
rect 19993 5321 20027 5355
rect 22017 5321 22051 5355
rect 22385 5321 22419 5355
rect 23489 5321 23523 5355
rect 25421 5321 25455 5355
rect 27445 5321 27479 5355
rect 30849 5321 30883 5355
rect 34161 5321 34195 5355
rect 15117 5253 15151 5287
rect 20177 5253 20211 5287
rect 23857 5253 23891 5287
rect 27261 5253 27295 5287
rect 31769 5253 31803 5287
rect 7481 5185 7515 5219
rect 7757 5185 7791 5219
rect 9413 5185 9447 5219
rect 9873 5185 9907 5219
rect 10057 5185 10091 5219
rect 11529 5185 11563 5219
rect 12449 5185 12483 5219
rect 12725 5185 12759 5219
rect 14841 5185 14875 5219
rect 15761 5185 15795 5219
rect 16129 5185 16163 5219
rect 16221 5185 16255 5219
rect 16313 5185 16347 5219
rect 16405 5185 16439 5219
rect 16773 5185 16807 5219
rect 16957 5185 16991 5219
rect 17233 5185 17267 5219
rect 17417 5185 17451 5219
rect 19809 5185 19843 5219
rect 19901 5185 19935 5219
rect 20085 5185 20119 5219
rect 20269 5185 20303 5219
rect 20545 5185 20579 5219
rect 25237 5185 25271 5219
rect 27537 5185 27571 5219
rect 30757 5185 30791 5219
rect 32781 5185 32815 5219
rect 33037 5185 33071 5219
rect 36185 5185 36219 5219
rect 11989 5117 12023 5151
rect 15025 5117 15059 5151
rect 15485 5117 15519 5151
rect 15577 5117 15611 5151
rect 22477 5117 22511 5151
rect 22661 5117 22695 5151
rect 23949 5117 23983 5151
rect 24133 5117 24167 5151
rect 25053 5117 25087 5151
rect 7481 5049 7515 5083
rect 9689 5049 9723 5083
rect 20729 5049 20763 5083
rect 10333 4981 10367 5015
rect 11805 4981 11839 5015
rect 15945 4981 15979 5015
rect 27261 4981 27295 5015
rect 31861 4981 31895 5015
rect 36369 4981 36403 5015
rect 25513 4777 25547 4811
rect 28365 4777 28399 4811
rect 28733 4709 28767 4743
rect 31401 4709 31435 4743
rect 25145 4641 25179 4675
rect 25329 4641 25363 4675
rect 28641 4641 28675 4675
rect 16957 4573 16991 4607
rect 17233 4573 17267 4607
rect 25053 4573 25087 4607
rect 25513 4573 25547 4607
rect 25697 4573 25731 4607
rect 27537 4573 27571 4607
rect 27685 4573 27719 4607
rect 28002 4573 28036 4607
rect 28273 4573 28307 4607
rect 28549 4573 28583 4607
rect 29101 4573 29135 4607
rect 31217 4573 31251 4607
rect 16773 4505 16807 4539
rect 25421 4505 25455 4539
rect 27813 4505 27847 4539
rect 27905 4505 27939 4539
rect 28825 4505 28859 4539
rect 29009 4505 29043 4539
rect 17141 4437 17175 4471
rect 25881 4437 25915 4471
rect 28181 4437 28215 4471
rect 29101 4437 29135 4471
rect 19993 4233 20027 4267
rect 20085 4233 20119 4267
rect 22845 4233 22879 4267
rect 22753 4165 22787 4199
rect 6633 4097 6667 4131
rect 9577 4097 9611 4131
rect 18613 4097 18647 4131
rect 22017 4097 22051 4131
rect 25053 4097 25087 4131
rect 25237 4097 25271 4131
rect 25329 4097 25363 4131
rect 26249 4097 26283 4131
rect 26433 4097 26467 4131
rect 26525 4097 26559 4131
rect 26709 4097 26743 4131
rect 30297 4097 30331 4131
rect 30389 4097 30423 4131
rect 30481 4097 30515 4131
rect 30849 4097 30883 4131
rect 6377 4029 6411 4063
rect 9321 4029 9355 4063
rect 18705 4029 18739 4063
rect 18889 4029 18923 4063
rect 20269 4029 20303 4063
rect 22937 4029 22971 4063
rect 26617 4029 26651 4063
rect 30573 4029 30607 4063
rect 31033 4029 31067 4063
rect 10701 3961 10735 3995
rect 24869 3961 24903 3995
rect 25973 3961 26007 3995
rect 7757 3893 7791 3927
rect 18245 3893 18279 3927
rect 19625 3893 19659 3927
rect 21833 3893 21867 3927
rect 22385 3893 22419 3927
rect 26249 3893 26283 3927
rect 30113 3893 30147 3927
rect 22293 3689 22327 3723
rect 23489 3689 23523 3723
rect 34161 3689 34195 3723
rect 26893 3621 26927 3655
rect 28457 3621 28491 3655
rect 19257 3553 19291 3587
rect 20913 3553 20947 3587
rect 21097 3553 21131 3587
rect 22477 3553 22511 3587
rect 26157 3553 26191 3587
rect 26985 3553 27019 3587
rect 30113 3553 30147 3587
rect 31585 3553 31619 3587
rect 32321 3553 32355 3587
rect 15761 3485 15795 3519
rect 17693 3485 17727 3519
rect 17785 3485 17819 3519
rect 18061 3485 18095 3519
rect 19533 3485 19567 3519
rect 20361 3485 20395 3519
rect 21281 3485 21315 3519
rect 21557 3485 21591 3519
rect 22753 3485 22787 3519
rect 25881 3485 25915 3519
rect 25973 3485 26007 3519
rect 26525 3485 26559 3519
rect 26709 3485 26743 3519
rect 26801 3485 26835 3519
rect 27077 3485 27111 3519
rect 28181 3485 28215 3519
rect 28457 3485 28491 3519
rect 29742 3485 29776 3519
rect 30205 3485 30239 3519
rect 30849 3485 30883 3519
rect 30941 3485 30975 3519
rect 31309 3485 31343 3519
rect 31401 3485 31435 3519
rect 31493 3485 31527 3519
rect 31769 3485 31803 3519
rect 31861 3485 31895 3519
rect 31953 3485 31987 3519
rect 32413 3485 32447 3519
rect 32510 3463 32544 3497
rect 32781 3485 32815 3519
rect 33037 3485 33071 3519
rect 16028 3417 16062 3451
rect 26157 3417 26191 3451
rect 28365 3417 28399 3451
rect 32137 3417 32171 3451
rect 32321 3417 32355 3451
rect 17141 3349 17175 3383
rect 17509 3349 17543 3383
rect 18797 3349 18831 3383
rect 20453 3349 20487 3383
rect 20821 3349 20855 3383
rect 29561 3349 29595 3383
rect 29745 3349 29779 3383
rect 30665 3349 30699 3383
rect 31125 3349 31159 3383
rect 31217 3349 31251 3383
rect 31677 3349 31711 3383
rect 1409 3145 1443 3179
rect 16221 3145 16255 3179
rect 17049 3145 17083 3179
rect 18981 3145 19015 3179
rect 19441 3145 19475 3179
rect 19901 3145 19935 3179
rect 21189 3145 21223 3179
rect 21833 3145 21867 3179
rect 22201 3145 22235 3179
rect 22661 3145 22695 3179
rect 24777 3145 24811 3179
rect 25421 3145 25455 3179
rect 25697 3145 25731 3179
rect 26985 3145 27019 3179
rect 27537 3145 27571 3179
rect 30573 3145 30607 3179
rect 31401 3145 31435 3179
rect 31585 3145 31619 3179
rect 34161 3145 34195 3179
rect 3126 3077 3160 3111
rect 17141 3077 17175 3111
rect 28816 3077 28850 3111
rect 32137 3077 32171 3111
rect 32321 3077 32355 3111
rect 1593 3009 1627 3043
rect 2881 3009 2915 3043
rect 16405 3009 16439 3043
rect 17601 3009 17635 3043
rect 17868 3009 17902 3043
rect 19625 3009 19659 3043
rect 20085 3009 20119 3043
rect 20177 3009 20211 3043
rect 20453 3009 20487 3043
rect 22845 3009 22879 3043
rect 23949 3009 23983 3043
rect 24409 3009 24443 3043
rect 25053 3009 25087 3043
rect 25881 3009 25915 3043
rect 26157 3009 26191 3043
rect 26341 3009 26375 3043
rect 27169 3009 27203 3043
rect 27537 3009 27571 3043
rect 28549 3009 28583 3043
rect 30389 3009 30423 3043
rect 30481 3009 30515 3043
rect 30757 3009 30791 3043
rect 31309 3009 31343 3043
rect 31677 3009 31711 3043
rect 32781 3009 32815 3043
rect 33048 3009 33082 3043
rect 36093 3009 36127 3043
rect 17325 2941 17359 2975
rect 22293 2941 22327 2975
rect 22385 2941 22419 2975
rect 24317 2941 24351 2975
rect 25145 2941 25179 2975
rect 27445 2941 27479 2975
rect 27813 2941 27847 2975
rect 31493 2941 31527 2975
rect 32505 2941 32539 2975
rect 35633 2941 35667 2975
rect 4261 2873 4295 2907
rect 16681 2873 16715 2907
rect 24133 2873 24167 2907
rect 27629 2873 27663 2907
rect 30665 2873 30699 2907
rect 36277 2873 36311 2907
rect 27353 2805 27387 2839
rect 29929 2805 29963 2839
rect 5917 2601 5951 2635
rect 9137 2601 9171 2635
rect 18153 2601 18187 2635
rect 21373 2601 21407 2635
rect 25789 2601 25823 2635
rect 32965 2601 32999 2635
rect 3341 2533 3375 2567
rect 30389 2533 30423 2567
rect 25973 2465 26007 2499
rect 26157 2465 26191 2499
rect 35633 2465 35667 2499
rect 2881 2397 2915 2431
rect 6101 2397 6135 2431
rect 9321 2397 9355 2431
rect 11713 2397 11747 2431
rect 14933 2397 14967 2431
rect 18337 2397 18371 2431
rect 21557 2397 21591 2431
rect 23949 2397 23983 2431
rect 26065 2397 26099 2431
rect 27353 2397 27387 2431
rect 30573 2397 30607 2431
rect 33149 2397 33183 2431
rect 35909 2397 35943 2431
rect 1409 2329 1443 2363
rect 1777 2329 1811 2363
rect 30205 2329 30239 2363
rect 2237 2261 2271 2295
rect 2605 2261 2639 2295
rect 11897 2261 11931 2295
rect 15117 2261 15151 2295
rect 24133 2261 24167 2295
rect 27169 2261 27203 2295
rect 30665 2261 30699 2295
<< metal1 >>
rect 1104 37562 36800 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 36800 37562
rect 1104 37488 36800 37510
rect 934 37408 940 37460
rect 992 37448 998 37460
rect 1765 37451 1823 37457
rect 1765 37448 1777 37451
rect 992 37420 1777 37448
rect 992 37408 998 37420
rect 1765 37417 1777 37420
rect 1811 37417 1823 37451
rect 1765 37411 1823 37417
rect 21266 37408 21272 37460
rect 21324 37448 21330 37460
rect 22557 37451 22615 37457
rect 22557 37448 22569 37451
rect 21324 37420 22569 37448
rect 21324 37408 21330 37420
rect 22557 37417 22569 37420
rect 22603 37417 22615 37451
rect 22557 37411 22615 37417
rect 29914 37380 29920 37392
rect 26206 37352 29920 37380
rect 4614 37272 4620 37324
rect 4672 37272 4678 37324
rect 17034 37272 17040 37324
rect 17092 37312 17098 37324
rect 17681 37315 17739 37321
rect 17681 37312 17693 37315
rect 17092 37284 17693 37312
rect 17092 37272 17098 37284
rect 17681 37281 17693 37284
rect 17727 37312 17739 37315
rect 19245 37315 19303 37321
rect 17727 37284 18092 37312
rect 17727 37281 17739 37284
rect 17681 37275 17739 37281
rect 1673 37247 1731 37253
rect 1673 37213 1685 37247
rect 1719 37244 1731 37247
rect 4893 37247 4951 37253
rect 1719 37216 4292 37244
rect 1719 37213 1731 37216
rect 1673 37207 1731 37213
rect 1302 37136 1308 37188
rect 1360 37176 1366 37188
rect 2225 37179 2283 37185
rect 2225 37176 2237 37179
rect 1360 37148 2237 37176
rect 1360 37136 1366 37148
rect 2225 37145 2237 37148
rect 2271 37145 2283 37179
rect 4264 37176 4292 37216
rect 4893 37213 4905 37247
rect 4939 37244 4951 37247
rect 5442 37244 5448 37256
rect 4939 37216 5448 37244
rect 4939 37213 4951 37216
rect 4893 37207 4951 37213
rect 5442 37204 5448 37216
rect 5500 37204 5506 37256
rect 6822 37204 6828 37256
rect 6880 37244 6886 37256
rect 7193 37247 7251 37253
rect 7193 37244 7205 37247
rect 6880 37216 7205 37244
rect 6880 37204 6886 37216
rect 7193 37213 7205 37216
rect 7239 37213 7251 37247
rect 7193 37207 7251 37213
rect 10410 37204 10416 37256
rect 10468 37204 10474 37256
rect 12802 37204 12808 37256
rect 12860 37244 12866 37256
rect 13633 37247 13691 37253
rect 13633 37244 13645 37247
rect 12860 37216 13645 37244
rect 12860 37204 12866 37216
rect 13633 37213 13645 37216
rect 13679 37213 13691 37247
rect 13633 37207 13691 37213
rect 16209 37247 16267 37253
rect 16209 37213 16221 37247
rect 16255 37244 16267 37247
rect 16255 37216 17632 37244
rect 16255 37213 16267 37216
rect 16209 37207 16267 37213
rect 17218 37176 17224 37188
rect 4264 37148 17224 37176
rect 2225 37139 2283 37145
rect 17218 37136 17224 37148
rect 17276 37136 17282 37188
rect 17604 37176 17632 37216
rect 17862 37204 17868 37256
rect 17920 37244 17926 37256
rect 17957 37247 18015 37253
rect 17957 37244 17969 37247
rect 17920 37216 17969 37244
rect 17920 37204 17926 37216
rect 17957 37213 17969 37216
rect 18003 37213 18015 37247
rect 18064 37244 18092 37284
rect 19245 37281 19257 37315
rect 19291 37312 19303 37315
rect 26206 37312 26234 37352
rect 29914 37340 29920 37352
rect 29972 37340 29978 37392
rect 31754 37340 31760 37392
rect 31812 37340 31818 37392
rect 19291 37284 26234 37312
rect 19291 37281 19303 37284
rect 19245 37275 19303 37281
rect 28442 37272 28448 37324
rect 28500 37272 28506 37324
rect 19334 37244 19340 37256
rect 18064 37216 19340 37244
rect 17957 37207 18015 37213
rect 19334 37204 19340 37216
rect 19392 37244 19398 37256
rect 19521 37247 19579 37253
rect 19521 37244 19533 37247
rect 19392 37216 19533 37244
rect 19392 37204 19398 37216
rect 19521 37213 19533 37216
rect 19567 37213 19579 37247
rect 19521 37207 19579 37213
rect 19610 37204 19616 37256
rect 19668 37244 19674 37256
rect 20349 37247 20407 37253
rect 20349 37244 20361 37247
rect 19668 37216 20361 37244
rect 19668 37204 19674 37216
rect 20349 37213 20361 37216
rect 20395 37213 20407 37247
rect 20349 37207 20407 37213
rect 22278 37204 22284 37256
rect 22336 37244 22342 37256
rect 22741 37247 22799 37253
rect 22741 37244 22753 37247
rect 22336 37216 22753 37244
rect 22336 37204 22342 37216
rect 22741 37213 22753 37216
rect 22787 37213 22799 37247
rect 22741 37207 22799 37213
rect 25866 37204 25872 37256
rect 25924 37204 25930 37256
rect 28626 37204 28632 37256
rect 28684 37244 28690 37256
rect 28721 37247 28779 37253
rect 28721 37244 28733 37247
rect 28684 37216 28733 37244
rect 28684 37204 28690 37216
rect 28721 37213 28733 37216
rect 28767 37213 28779 37247
rect 28721 37207 28779 37213
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 35069 37247 35127 37253
rect 35069 37244 35081 37247
rect 34848 37216 35081 37244
rect 34848 37204 34854 37216
rect 35069 37213 35081 37216
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 36170 37204 36176 37256
rect 36228 37204 36234 37256
rect 20622 37176 20628 37188
rect 17604 37148 20628 37176
rect 20622 37136 20628 37148
rect 20680 37136 20686 37188
rect 22465 37179 22523 37185
rect 22465 37145 22477 37179
rect 22511 37176 22523 37179
rect 25130 37176 25136 37188
rect 22511 37148 25136 37176
rect 22511 37145 22523 37148
rect 22465 37139 22523 37145
rect 25130 37136 25136 37148
rect 25188 37136 25194 37188
rect 31478 37136 31484 37188
rect 31536 37176 31542 37188
rect 31573 37179 31631 37185
rect 31573 37176 31585 37179
rect 31536 37148 31585 37176
rect 31536 37136 31542 37148
rect 31573 37145 31585 37148
rect 31619 37145 31631 37179
rect 31573 37139 31631 37145
rect 35897 37179 35955 37185
rect 35897 37145 35909 37179
rect 35943 37176 35955 37179
rect 37366 37176 37372 37188
rect 35943 37148 37372 37176
rect 35943 37145 35955 37148
rect 35897 37139 35955 37145
rect 37366 37136 37372 37148
rect 37424 37136 37430 37188
rect 2314 37068 2320 37120
rect 2372 37068 2378 37120
rect 7374 37068 7380 37120
rect 7432 37068 7438 37120
rect 10594 37068 10600 37120
rect 10652 37068 10658 37120
rect 13538 37068 13544 37120
rect 13596 37108 13602 37120
rect 13817 37111 13875 37117
rect 13817 37108 13829 37111
rect 13596 37080 13829 37108
rect 13596 37068 13602 37080
rect 13817 37077 13829 37080
rect 13863 37077 13875 37111
rect 13817 37071 13875 37077
rect 16390 37068 16396 37120
rect 16448 37068 16454 37120
rect 20162 37068 20168 37120
rect 20220 37068 20226 37120
rect 22922 37068 22928 37120
rect 22980 37068 22986 37120
rect 26050 37068 26056 37120
rect 26108 37068 26114 37120
rect 30098 37068 30104 37120
rect 30156 37108 30162 37120
rect 34885 37111 34943 37117
rect 34885 37108 34897 37111
rect 30156 37080 34897 37108
rect 30156 37068 30162 37080
rect 34885 37077 34897 37080
rect 34931 37077 34943 37111
rect 34885 37071 34943 37077
rect 36354 37068 36360 37120
rect 36412 37068 36418 37120
rect 1104 37018 36800 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 36800 37018
rect 1104 36944 36800 36966
rect 6822 36864 6828 36916
rect 6880 36864 6886 36916
rect 17129 36907 17187 36913
rect 17129 36873 17141 36907
rect 17175 36873 17187 36907
rect 17129 36867 17187 36873
rect 18969 36907 19027 36913
rect 18969 36873 18981 36907
rect 19015 36873 19027 36907
rect 18969 36867 19027 36873
rect 17034 36836 17040 36848
rect 7116 36808 17040 36836
rect 6914 36728 6920 36780
rect 6972 36768 6978 36780
rect 7116 36777 7144 36808
rect 17034 36796 17040 36808
rect 17092 36796 17098 36848
rect 17144 36836 17172 36867
rect 17650 36839 17708 36845
rect 17650 36836 17662 36839
rect 17144 36808 17662 36836
rect 17650 36805 17662 36808
rect 17696 36805 17708 36839
rect 18984 36836 19012 36867
rect 20622 36864 20628 36916
rect 20680 36864 20686 36916
rect 22278 36864 22284 36916
rect 22336 36864 22342 36916
rect 19490 36839 19548 36845
rect 19490 36836 19502 36839
rect 18984 36808 19502 36836
rect 17650 36799 17708 36805
rect 19490 36805 19502 36808
rect 19536 36805 19548 36839
rect 19490 36799 19548 36805
rect 20162 36796 20168 36848
rect 20220 36836 20226 36848
rect 22986 36839 23044 36845
rect 22986 36836 22998 36839
rect 20220 36808 22998 36836
rect 20220 36796 20226 36808
rect 22986 36805 22998 36808
rect 23032 36805 23044 36839
rect 22986 36799 23044 36805
rect 30098 36796 30104 36848
rect 30156 36796 30162 36848
rect 7009 36771 7067 36777
rect 7009 36768 7021 36771
rect 6972 36740 7021 36768
rect 6972 36728 6978 36740
rect 7009 36737 7021 36740
rect 7055 36737 7067 36771
rect 7009 36731 7067 36737
rect 7101 36771 7159 36777
rect 7101 36737 7113 36771
rect 7147 36737 7159 36771
rect 7101 36731 7159 36737
rect 16485 36771 16543 36777
rect 16485 36737 16497 36771
rect 16531 36768 16543 36771
rect 16666 36768 16672 36780
rect 16531 36740 16672 36768
rect 16531 36737 16543 36740
rect 16485 36731 16543 36737
rect 7024 36700 7052 36731
rect 16666 36728 16672 36740
rect 16724 36728 16730 36780
rect 17313 36771 17371 36777
rect 17313 36737 17325 36771
rect 17359 36768 17371 36771
rect 17954 36768 17960 36780
rect 17359 36740 17960 36768
rect 17359 36737 17371 36740
rect 17313 36731 17371 36737
rect 17954 36728 17960 36740
rect 18012 36728 18018 36780
rect 19150 36728 19156 36780
rect 19208 36728 19214 36780
rect 21637 36771 21695 36777
rect 21637 36737 21649 36771
rect 21683 36768 21695 36771
rect 22189 36771 22247 36777
rect 21683 36740 21864 36768
rect 21683 36737 21695 36740
rect 21637 36731 21695 36737
rect 7377 36703 7435 36709
rect 7377 36700 7389 36703
rect 7024 36672 7389 36700
rect 7377 36669 7389 36672
rect 7423 36669 7435 36703
rect 7377 36663 7435 36669
rect 17402 36660 17408 36712
rect 17460 36660 17466 36712
rect 19242 36660 19248 36712
rect 19300 36660 19306 36712
rect 10410 36592 10416 36644
rect 10468 36632 10474 36644
rect 21836 36641 21864 36740
rect 22189 36737 22201 36771
rect 22235 36768 22247 36771
rect 22554 36768 22560 36780
rect 22235 36740 22560 36768
rect 22235 36737 22247 36740
rect 22189 36731 22247 36737
rect 22554 36728 22560 36740
rect 22612 36728 22618 36780
rect 22741 36771 22799 36777
rect 22741 36737 22753 36771
rect 22787 36768 22799 36771
rect 22830 36768 22836 36780
rect 22787 36740 22836 36768
rect 22787 36737 22799 36740
rect 22741 36731 22799 36737
rect 22830 36728 22836 36740
rect 22888 36728 22894 36780
rect 22465 36703 22523 36709
rect 22465 36669 22477 36703
rect 22511 36669 22523 36703
rect 22465 36663 22523 36669
rect 21821 36635 21879 36641
rect 10468 36604 16574 36632
rect 10468 36592 10474 36604
rect 16114 36524 16120 36576
rect 16172 36564 16178 36576
rect 16301 36567 16359 36573
rect 16301 36564 16313 36567
rect 16172 36536 16313 36564
rect 16172 36524 16178 36536
rect 16301 36533 16313 36536
rect 16347 36533 16359 36567
rect 16546 36564 16574 36604
rect 21821 36601 21833 36635
rect 21867 36601 21879 36635
rect 22480 36632 22508 36663
rect 22738 36632 22744 36644
rect 22480 36604 22744 36632
rect 21821 36595 21879 36601
rect 22738 36592 22744 36604
rect 22796 36592 22802 36644
rect 30285 36635 30343 36641
rect 30285 36601 30297 36635
rect 30331 36632 30343 36635
rect 30834 36632 30840 36644
rect 30331 36604 30840 36632
rect 30331 36601 30343 36604
rect 30285 36595 30343 36601
rect 30834 36592 30840 36604
rect 30892 36592 30898 36644
rect 18322 36564 18328 36576
rect 16546 36536 18328 36564
rect 16301 36527 16359 36533
rect 18322 36524 18328 36536
rect 18380 36564 18386 36576
rect 18785 36567 18843 36573
rect 18785 36564 18797 36567
rect 18380 36536 18797 36564
rect 18380 36524 18386 36536
rect 18785 36533 18797 36536
rect 18831 36533 18843 36567
rect 18785 36527 18843 36533
rect 21453 36567 21511 36573
rect 21453 36533 21465 36567
rect 21499 36564 21511 36567
rect 21542 36564 21548 36576
rect 21499 36536 21548 36564
rect 21499 36533 21511 36536
rect 21453 36527 21511 36533
rect 21542 36524 21548 36536
rect 21600 36524 21606 36576
rect 24118 36524 24124 36576
rect 24176 36524 24182 36576
rect 1104 36474 36800 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 36800 36474
rect 1104 36400 36800 36422
rect 17218 36320 17224 36372
rect 17276 36320 17282 36372
rect 17954 36320 17960 36372
rect 18012 36320 18018 36372
rect 19150 36320 19156 36372
rect 19208 36360 19214 36372
rect 19521 36363 19579 36369
rect 19521 36360 19533 36363
rect 19208 36332 19533 36360
rect 19208 36320 19214 36332
rect 19521 36329 19533 36332
rect 19567 36329 19579 36363
rect 19521 36323 19579 36329
rect 20732 36332 22232 36360
rect 20622 36292 20628 36304
rect 19996 36264 20628 36292
rect 18601 36227 18659 36233
rect 18601 36193 18613 36227
rect 18647 36224 18659 36227
rect 19058 36224 19064 36236
rect 18647 36196 19064 36224
rect 18647 36193 18659 36196
rect 18601 36187 18659 36193
rect 19058 36184 19064 36196
rect 19116 36184 19122 36236
rect 19996 36233 20024 36264
rect 20622 36252 20628 36264
rect 20680 36252 20686 36304
rect 19981 36227 20039 36233
rect 19981 36193 19993 36227
rect 20027 36193 20039 36227
rect 19981 36187 20039 36193
rect 20073 36227 20131 36233
rect 20073 36193 20085 36227
rect 20119 36224 20131 36227
rect 20732 36224 20760 36332
rect 22204 36292 22232 36332
rect 22278 36320 22284 36372
rect 22336 36360 22342 36372
rect 22649 36363 22707 36369
rect 22649 36360 22661 36363
rect 22336 36332 22661 36360
rect 22336 36320 22342 36332
rect 22649 36329 22661 36332
rect 22695 36329 22707 36363
rect 22649 36323 22707 36329
rect 22738 36320 22744 36372
rect 22796 36360 22802 36372
rect 30282 36360 30288 36372
rect 22796 36332 30288 36360
rect 22796 36320 22802 36332
rect 30282 36320 30288 36332
rect 30340 36320 30346 36372
rect 22756 36292 22784 36320
rect 22204 36264 22784 36292
rect 20119 36196 20760 36224
rect 20119 36193 20131 36196
rect 20073 36187 20131 36193
rect 3786 36116 3792 36168
rect 3844 36156 3850 36168
rect 5813 36159 5871 36165
rect 5813 36156 5825 36159
rect 3844 36128 5825 36156
rect 3844 36116 3850 36128
rect 5813 36125 5825 36128
rect 5859 36156 5871 36159
rect 8478 36156 8484 36168
rect 5859 36128 8484 36156
rect 5859 36125 5871 36128
rect 5813 36119 5871 36125
rect 8478 36116 8484 36128
rect 8536 36116 8542 36168
rect 16114 36165 16120 36168
rect 15841 36159 15899 36165
rect 15841 36125 15853 36159
rect 15887 36125 15899 36159
rect 16108 36156 16120 36165
rect 16075 36128 16120 36156
rect 15841 36119 15899 36125
rect 16108 36119 16120 36128
rect 6080 36091 6138 36097
rect 6080 36057 6092 36091
rect 6126 36088 6138 36091
rect 6362 36088 6368 36100
rect 6126 36060 6368 36088
rect 6126 36057 6138 36060
rect 6080 36051 6138 36057
rect 6362 36048 6368 36060
rect 6420 36048 6426 36100
rect 15856 36088 15884 36119
rect 16114 36116 16120 36119
rect 16172 36116 16178 36168
rect 17310 36116 17316 36168
rect 17368 36156 17374 36168
rect 17681 36159 17739 36165
rect 17681 36156 17693 36159
rect 17368 36128 17693 36156
rect 17368 36116 17374 36128
rect 17681 36125 17693 36128
rect 17727 36156 17739 36159
rect 17862 36156 17868 36168
rect 17727 36128 17868 36156
rect 17727 36125 17739 36128
rect 17681 36119 17739 36125
rect 17862 36116 17868 36128
rect 17920 36116 17926 36168
rect 18325 36159 18383 36165
rect 18325 36125 18337 36159
rect 18371 36156 18383 36159
rect 18414 36156 18420 36168
rect 18371 36128 18420 36156
rect 18371 36125 18383 36128
rect 18325 36119 18383 36125
rect 18414 36116 18420 36128
rect 18472 36116 18478 36168
rect 19076 36156 19104 36184
rect 20088 36156 20116 36187
rect 21266 36184 21272 36236
rect 21324 36184 21330 36236
rect 29270 36184 29276 36236
rect 29328 36224 29334 36236
rect 30193 36227 30251 36233
rect 30193 36224 30205 36227
rect 29328 36196 30205 36224
rect 29328 36184 29334 36196
rect 30193 36193 30205 36196
rect 30239 36193 30251 36227
rect 31113 36227 31171 36233
rect 31113 36224 31125 36227
rect 30193 36187 30251 36193
rect 30300 36196 31125 36224
rect 21542 36165 21548 36168
rect 21536 36156 21548 36165
rect 19076 36128 20116 36156
rect 21503 36128 21548 36156
rect 21536 36119 21548 36128
rect 21542 36116 21548 36119
rect 21600 36116 21606 36168
rect 29914 36116 29920 36168
rect 29972 36156 29978 36168
rect 30300 36156 30328 36196
rect 31113 36193 31125 36196
rect 31159 36224 31171 36227
rect 32766 36224 32772 36236
rect 31159 36196 32772 36224
rect 31159 36193 31171 36196
rect 31113 36187 31171 36193
rect 32766 36184 32772 36196
rect 32824 36184 32830 36236
rect 29972 36128 30328 36156
rect 29972 36116 29978 36128
rect 30834 36116 30840 36168
rect 30892 36116 30898 36168
rect 15856 36060 17448 36088
rect 17420 36032 17448 36060
rect 7190 35980 7196 36032
rect 7248 35980 7254 36032
rect 17402 35980 17408 36032
rect 17460 36020 17466 36032
rect 17497 36023 17555 36029
rect 17497 36020 17509 36023
rect 17460 35992 17509 36020
rect 17460 35980 17466 35992
rect 17497 35989 17509 35992
rect 17543 35989 17555 36023
rect 17497 35983 17555 35989
rect 18322 35980 18328 36032
rect 18380 36020 18386 36032
rect 18417 36023 18475 36029
rect 18417 36020 18429 36023
rect 18380 35992 18429 36020
rect 18380 35980 18386 35992
rect 18417 35989 18429 35992
rect 18463 35989 18475 36023
rect 18417 35983 18475 35989
rect 19518 35980 19524 36032
rect 19576 36020 19582 36032
rect 19889 36023 19947 36029
rect 19889 36020 19901 36023
rect 19576 35992 19901 36020
rect 19576 35980 19582 35992
rect 19889 35989 19901 35992
rect 19935 35989 19947 36023
rect 19889 35983 19947 35989
rect 1104 35930 36800 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 36800 35930
rect 1104 35856 36800 35878
rect 6362 35776 6368 35828
rect 6420 35776 6426 35828
rect 16666 35776 16672 35828
rect 16724 35776 16730 35828
rect 17129 35819 17187 35825
rect 17129 35785 17141 35819
rect 17175 35816 17187 35819
rect 17218 35816 17224 35828
rect 17175 35788 17224 35816
rect 17175 35785 17187 35788
rect 17129 35779 17187 35785
rect 17218 35776 17224 35788
rect 17276 35776 17282 35828
rect 29365 35819 29423 35825
rect 29365 35785 29377 35819
rect 29411 35785 29423 35819
rect 29365 35779 29423 35785
rect 19242 35708 19248 35760
rect 19300 35748 19306 35760
rect 21266 35748 21272 35760
rect 19300 35720 21272 35748
rect 19300 35708 19306 35720
rect 6178 35640 6184 35692
rect 6236 35680 6242 35692
rect 6549 35683 6607 35689
rect 6549 35680 6561 35683
rect 6236 35652 6561 35680
rect 6236 35640 6242 35652
rect 6549 35649 6561 35652
rect 6595 35649 6607 35683
rect 6549 35643 6607 35649
rect 16942 35640 16948 35692
rect 17000 35680 17006 35692
rect 19444 35689 19472 35720
rect 21266 35708 21272 35720
rect 21324 35708 21330 35760
rect 29380 35748 29408 35779
rect 30190 35776 30196 35828
rect 30248 35816 30254 35828
rect 31021 35819 31079 35825
rect 31021 35816 31033 35819
rect 30248 35788 31033 35816
rect 30248 35776 30254 35788
rect 31021 35785 31033 35788
rect 31067 35816 31079 35819
rect 36170 35816 36176 35828
rect 31067 35788 36176 35816
rect 31067 35785 31079 35788
rect 31021 35779 31079 35785
rect 36170 35776 36176 35788
rect 36228 35776 36234 35828
rect 29886 35751 29944 35757
rect 29886 35748 29898 35751
rect 29380 35720 29898 35748
rect 29886 35717 29898 35720
rect 29932 35717 29944 35751
rect 29886 35711 29944 35717
rect 19702 35689 19708 35692
rect 17037 35683 17095 35689
rect 17037 35680 17049 35683
rect 17000 35652 17049 35680
rect 17000 35640 17006 35652
rect 17037 35649 17049 35652
rect 17083 35649 17095 35683
rect 17037 35643 17095 35649
rect 19429 35683 19487 35689
rect 19429 35649 19441 35683
rect 19475 35649 19487 35683
rect 19429 35643 19487 35649
rect 19696 35643 19708 35689
rect 19702 35640 19708 35643
rect 19760 35640 19766 35692
rect 29270 35640 29276 35692
rect 29328 35640 29334 35692
rect 29549 35683 29607 35689
rect 29549 35649 29561 35683
rect 29595 35680 29607 35683
rect 29730 35680 29736 35692
rect 29595 35652 29736 35680
rect 29595 35649 29607 35652
rect 29549 35643 29607 35649
rect 29730 35640 29736 35652
rect 29788 35640 29794 35692
rect 17313 35615 17371 35621
rect 17313 35581 17325 35615
rect 17359 35612 17371 35615
rect 19058 35612 19064 35624
rect 17359 35584 19064 35612
rect 17359 35581 17371 35584
rect 17313 35575 17371 35581
rect 19058 35572 19064 35584
rect 19116 35572 19122 35624
rect 29641 35615 29699 35621
rect 29641 35581 29653 35615
rect 29687 35581 29699 35615
rect 29641 35575 29699 35581
rect 20809 35479 20867 35485
rect 20809 35445 20821 35479
rect 20855 35476 20867 35479
rect 20990 35476 20996 35488
rect 20855 35448 20996 35476
rect 20855 35445 20867 35448
rect 20809 35439 20867 35445
rect 20990 35436 20996 35448
rect 21048 35436 21054 35488
rect 29089 35479 29147 35485
rect 29089 35445 29101 35479
rect 29135 35476 29147 35479
rect 29656 35476 29684 35575
rect 30558 35476 30564 35488
rect 29135 35448 30564 35476
rect 29135 35445 29147 35448
rect 29089 35439 29147 35445
rect 30558 35436 30564 35448
rect 30616 35436 30622 35488
rect 1104 35386 36800 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 36800 35386
rect 1104 35312 36800 35334
rect 6178 35232 6184 35284
rect 6236 35232 6242 35284
rect 9033 35275 9091 35281
rect 9033 35241 9045 35275
rect 9079 35272 9091 35275
rect 10318 35272 10324 35284
rect 9079 35244 10324 35272
rect 9079 35241 9091 35244
rect 9033 35235 9091 35241
rect 10318 35232 10324 35244
rect 10376 35232 10382 35284
rect 19702 35232 19708 35284
rect 19760 35232 19766 35284
rect 24486 35272 24492 35284
rect 20640 35244 24492 35272
rect 9048 35176 9812 35204
rect 6730 35096 6736 35148
rect 6788 35136 6794 35148
rect 9048 35136 9076 35176
rect 6788 35108 9076 35136
rect 9217 35139 9275 35145
rect 6788 35096 6794 35108
rect 1397 35071 1455 35077
rect 1397 35037 1409 35071
rect 1443 35068 1455 35071
rect 2130 35068 2136 35080
rect 1443 35040 2136 35068
rect 1443 35037 1455 35040
rect 1397 35031 1455 35037
rect 2130 35028 2136 35040
rect 2188 35028 2194 35080
rect 6641 35071 6699 35077
rect 6641 35037 6653 35071
rect 6687 35068 6699 35071
rect 7190 35068 7196 35080
rect 6687 35040 7196 35068
rect 6687 35037 6699 35040
rect 6641 35031 6699 35037
rect 7190 35028 7196 35040
rect 7248 35028 7254 35080
rect 8956 35077 8984 35108
rect 9217 35105 9229 35139
rect 9263 35136 9275 35139
rect 9677 35139 9735 35145
rect 9677 35136 9689 35139
rect 9263 35108 9689 35136
rect 9263 35105 9275 35108
rect 9217 35099 9275 35105
rect 9677 35105 9689 35108
rect 9723 35105 9735 35139
rect 9677 35099 9735 35105
rect 9784 35077 9812 35176
rect 11698 35096 11704 35148
rect 11756 35136 11762 35148
rect 14645 35139 14703 35145
rect 14645 35136 14657 35139
rect 11756 35108 14657 35136
rect 11756 35096 11762 35108
rect 14645 35105 14657 35108
rect 14691 35136 14703 35139
rect 14691 35108 17356 35136
rect 14691 35105 14703 35108
rect 14645 35099 14703 35105
rect 8941 35071 8999 35077
rect 8941 35037 8953 35071
rect 8987 35037 8999 35071
rect 8941 35031 8999 35037
rect 9585 35071 9643 35077
rect 9585 35037 9597 35071
rect 9631 35037 9643 35071
rect 9585 35031 9643 35037
rect 9769 35071 9827 35077
rect 9769 35037 9781 35071
rect 9815 35068 9827 35071
rect 11054 35068 11060 35080
rect 9815 35040 11060 35068
rect 9815 35037 9827 35040
rect 9769 35031 9827 35037
rect 6549 35003 6607 35009
rect 6549 34969 6561 35003
rect 6595 35000 6607 35003
rect 7282 35000 7288 35012
rect 6595 34972 7288 35000
rect 6595 34969 6607 34972
rect 6549 34963 6607 34969
rect 7282 34960 7288 34972
rect 7340 34960 7346 35012
rect 9600 35000 9628 35031
rect 11054 35028 11060 35040
rect 11112 35028 11118 35080
rect 17126 35028 17132 35080
rect 17184 35068 17190 35080
rect 17221 35071 17279 35077
rect 17221 35068 17233 35071
rect 17184 35040 17233 35068
rect 17184 35028 17190 35040
rect 17221 35037 17233 35040
rect 17267 35037 17279 35071
rect 17328 35068 17356 35108
rect 19794 35096 19800 35148
rect 19852 35136 19858 35148
rect 20640 35145 20668 35244
rect 24486 35232 24492 35244
rect 24544 35232 24550 35284
rect 29730 35232 29736 35284
rect 29788 35232 29794 35284
rect 20625 35139 20683 35145
rect 20625 35136 20637 35139
rect 19852 35108 20637 35136
rect 19852 35096 19858 35108
rect 20625 35105 20637 35108
rect 20671 35105 20683 35139
rect 25041 35139 25099 35145
rect 25041 35136 25053 35139
rect 20625 35099 20683 35105
rect 23860 35108 25053 35136
rect 18782 35068 18788 35080
rect 17328 35040 18788 35068
rect 17221 35031 17279 35037
rect 18782 35028 18788 35040
rect 18840 35028 18846 35080
rect 19889 35071 19947 35077
rect 19889 35037 19901 35071
rect 19935 35068 19947 35071
rect 20441 35071 20499 35077
rect 19935 35040 20024 35068
rect 19935 35037 19947 35040
rect 19889 35031 19947 35037
rect 9858 35000 9864 35012
rect 9600 34972 9864 35000
rect 9858 34960 9864 34972
rect 9916 34960 9922 35012
rect 12894 34960 12900 35012
rect 12952 35000 12958 35012
rect 14461 35003 14519 35009
rect 14461 35000 14473 35003
rect 12952 34972 14473 35000
rect 12952 34960 12958 34972
rect 14461 34969 14473 34972
rect 14507 34969 14519 35003
rect 14461 34963 14519 34969
rect 17034 34960 17040 35012
rect 17092 35000 17098 35012
rect 17466 35003 17524 35009
rect 17466 35000 17478 35003
rect 17092 34972 17478 35000
rect 17092 34960 17098 34972
rect 17466 34969 17478 34972
rect 17512 34969 17524 35003
rect 17466 34963 17524 34969
rect 934 34892 940 34944
rect 992 34932 998 34944
rect 1581 34935 1639 34941
rect 1581 34932 1593 34935
rect 992 34904 1593 34932
rect 992 34892 998 34904
rect 1581 34901 1593 34904
rect 1627 34901 1639 34935
rect 1581 34895 1639 34901
rect 9214 34892 9220 34944
rect 9272 34892 9278 34944
rect 13814 34892 13820 34944
rect 13872 34932 13878 34944
rect 14093 34935 14151 34941
rect 14093 34932 14105 34935
rect 13872 34904 14105 34932
rect 13872 34892 13878 34904
rect 14093 34901 14105 34904
rect 14139 34901 14151 34935
rect 14093 34895 14151 34901
rect 14550 34892 14556 34944
rect 14608 34892 14614 34944
rect 15562 34892 15568 34944
rect 15620 34932 15626 34944
rect 17310 34932 17316 34944
rect 15620 34904 17316 34932
rect 15620 34892 15626 34904
rect 17310 34892 17316 34904
rect 17368 34892 17374 34944
rect 18601 34935 18659 34941
rect 18601 34901 18613 34935
rect 18647 34932 18659 34935
rect 18690 34932 18696 34944
rect 18647 34904 18696 34932
rect 18647 34901 18659 34904
rect 18601 34895 18659 34901
rect 18690 34892 18696 34904
rect 18748 34892 18754 34944
rect 19996 34941 20024 35040
rect 20441 35037 20453 35071
rect 20487 35068 20499 35071
rect 20990 35068 20996 35080
rect 20487 35040 20996 35068
rect 20487 35037 20499 35040
rect 20441 35031 20499 35037
rect 20990 35028 20996 35040
rect 21048 35028 21054 35080
rect 21082 35028 21088 35080
rect 21140 35028 21146 35080
rect 21177 35071 21235 35077
rect 21177 35037 21189 35071
rect 21223 35068 21235 35071
rect 21266 35068 21272 35080
rect 21223 35040 21272 35068
rect 21223 35037 21235 35040
rect 21177 35031 21235 35037
rect 21266 35028 21272 35040
rect 21324 35028 21330 35080
rect 22830 35028 22836 35080
rect 22888 35068 22894 35080
rect 23860 35068 23888 35108
rect 25041 35105 25053 35108
rect 25087 35105 25099 35139
rect 25041 35099 25099 35105
rect 22888 35040 23888 35068
rect 22888 35028 22894 35040
rect 23934 35028 23940 35080
rect 23992 35068 23998 35080
rect 24581 35071 24639 35077
rect 24581 35068 24593 35071
rect 23992 35040 24593 35068
rect 23992 35028 23998 35040
rect 24581 35037 24593 35040
rect 24627 35037 24639 35071
rect 24581 35031 24639 35037
rect 24946 35028 24952 35080
rect 25004 35028 25010 35080
rect 25056 35068 25084 35099
rect 30190 35096 30196 35148
rect 30248 35096 30254 35148
rect 30282 35096 30288 35148
rect 30340 35096 30346 35148
rect 25056 35040 25544 35068
rect 25516 35012 25544 35040
rect 21422 35003 21480 35009
rect 21422 35000 21434 35003
rect 20916 34972 21434 35000
rect 19981 34935 20039 34941
rect 19981 34901 19993 34935
rect 20027 34901 20039 34935
rect 19981 34895 20039 34901
rect 20346 34892 20352 34944
rect 20404 34892 20410 34944
rect 20916 34941 20944 34972
rect 21422 34969 21434 34972
rect 21468 34969 21480 35003
rect 21422 34963 21480 34969
rect 23100 35003 23158 35009
rect 23100 34969 23112 35003
rect 23146 35000 23158 35003
rect 25286 35003 25344 35009
rect 25286 35000 25298 35003
rect 23146 34972 24440 35000
rect 23146 34969 23158 34972
rect 23100 34963 23158 34969
rect 20901 34935 20959 34941
rect 20901 34901 20913 34935
rect 20947 34901 20959 34935
rect 20901 34895 20959 34901
rect 22094 34892 22100 34944
rect 22152 34932 22158 34944
rect 22557 34935 22615 34941
rect 22557 34932 22569 34935
rect 22152 34904 22569 34932
rect 22152 34892 22158 34904
rect 22557 34901 22569 34904
rect 22603 34901 22615 34935
rect 22557 34895 22615 34901
rect 24213 34935 24271 34941
rect 24213 34901 24225 34935
rect 24259 34932 24271 34935
rect 24302 34932 24308 34944
rect 24259 34904 24308 34932
rect 24259 34901 24271 34904
rect 24213 34895 24271 34901
rect 24302 34892 24308 34904
rect 24360 34892 24366 34944
rect 24412 34941 24440 34972
rect 24780 34972 25298 35000
rect 24780 34941 24808 34972
rect 25286 34969 25298 34972
rect 25332 34969 25344 35003
rect 25286 34963 25344 34969
rect 25498 34960 25504 35012
rect 25556 34960 25562 35012
rect 24397 34935 24455 34941
rect 24397 34901 24409 34935
rect 24443 34901 24455 34935
rect 24397 34895 24455 34901
rect 24765 34935 24823 34941
rect 24765 34901 24777 34935
rect 24811 34901 24823 34935
rect 24765 34895 24823 34901
rect 24854 34892 24860 34944
rect 24912 34932 24918 34944
rect 25590 34932 25596 34944
rect 24912 34904 25596 34932
rect 24912 34892 24918 34904
rect 25590 34892 25596 34904
rect 25648 34892 25654 34944
rect 26421 34935 26479 34941
rect 26421 34901 26433 34935
rect 26467 34932 26479 34935
rect 26510 34932 26516 34944
rect 26467 34904 26516 34932
rect 26467 34901 26479 34904
rect 26421 34895 26479 34901
rect 26510 34892 26516 34904
rect 26568 34892 26574 34944
rect 30098 34892 30104 34944
rect 30156 34892 30162 34944
rect 1104 34842 36800 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 36800 34842
rect 1104 34768 36800 34790
rect 5169 34731 5227 34737
rect 5169 34697 5181 34731
rect 5215 34728 5227 34731
rect 5721 34731 5779 34737
rect 5721 34728 5733 34731
rect 5215 34700 5733 34728
rect 5215 34697 5227 34700
rect 5169 34691 5227 34697
rect 5721 34697 5733 34700
rect 5767 34728 5779 34731
rect 6362 34728 6368 34740
rect 5767 34700 6368 34728
rect 5767 34697 5779 34700
rect 5721 34691 5779 34697
rect 6362 34688 6368 34700
rect 6420 34688 6426 34740
rect 6641 34731 6699 34737
rect 6641 34697 6653 34731
rect 6687 34728 6699 34731
rect 6687 34700 6914 34728
rect 6687 34697 6699 34700
rect 6641 34691 6699 34697
rect 6886 34660 6914 34700
rect 9858 34688 9864 34740
rect 9916 34688 9922 34740
rect 10042 34688 10048 34740
rect 10100 34728 10106 34740
rect 11333 34731 11391 34737
rect 11333 34728 11345 34731
rect 10100 34700 11345 34728
rect 10100 34688 10106 34700
rect 11333 34697 11345 34700
rect 11379 34697 11391 34731
rect 11333 34691 11391 34697
rect 7162 34663 7220 34669
rect 7162 34660 7174 34663
rect 6886 34632 7174 34660
rect 7162 34629 7174 34632
rect 7208 34629 7220 34663
rect 7162 34623 7220 34629
rect 8748 34663 8806 34669
rect 8748 34629 8760 34663
rect 8794 34660 8806 34663
rect 9214 34660 9220 34672
rect 8794 34632 9220 34660
rect 8794 34629 8806 34632
rect 8748 34623 8806 34629
rect 9214 34620 9220 34632
rect 9272 34620 9278 34672
rect 9968 34632 11284 34660
rect 4056 34595 4114 34601
rect 4056 34561 4068 34595
rect 4102 34592 4114 34595
rect 4614 34592 4620 34604
rect 4102 34564 4620 34592
rect 4102 34561 4114 34564
rect 4056 34555 4114 34561
rect 4614 34552 4620 34564
rect 4672 34552 4678 34604
rect 5626 34552 5632 34604
rect 5684 34552 5690 34604
rect 6825 34595 6883 34601
rect 6825 34561 6837 34595
rect 6871 34592 6883 34595
rect 7006 34592 7012 34604
rect 6871 34564 7012 34592
rect 6871 34561 6883 34564
rect 6825 34555 6883 34561
rect 7006 34552 7012 34564
rect 7064 34552 7070 34604
rect 8478 34552 8484 34604
rect 8536 34552 8542 34604
rect 9968 34601 9996 34632
rect 10226 34601 10232 34604
rect 9953 34595 10011 34601
rect 9953 34561 9965 34595
rect 9999 34561 10011 34595
rect 9953 34555 10011 34561
rect 10220 34555 10232 34601
rect 10226 34552 10232 34555
rect 10284 34552 10290 34604
rect 3786 34484 3792 34536
rect 3844 34484 3850 34536
rect 5905 34527 5963 34533
rect 5905 34493 5917 34527
rect 5951 34524 5963 34527
rect 6730 34524 6736 34536
rect 5951 34496 6736 34524
rect 5951 34493 5963 34496
rect 5905 34487 5963 34493
rect 6730 34484 6736 34496
rect 6788 34484 6794 34536
rect 6914 34484 6920 34536
rect 6972 34484 6978 34536
rect 11256 34524 11284 34632
rect 11348 34592 11376 34691
rect 13998 34688 14004 34740
rect 14056 34728 14062 34740
rect 14550 34728 14556 34740
rect 14056 34700 14556 34728
rect 14056 34688 14062 34700
rect 14550 34688 14556 34700
rect 14608 34728 14614 34740
rect 14829 34731 14887 34737
rect 14829 34728 14841 34731
rect 14608 34700 14841 34728
rect 14608 34688 14614 34700
rect 14829 34697 14841 34700
rect 14875 34697 14887 34731
rect 14829 34691 14887 34697
rect 16669 34731 16727 34737
rect 16669 34697 16681 34731
rect 16715 34697 16727 34731
rect 16669 34691 16727 34697
rect 14090 34660 14096 34672
rect 11900 34632 12434 34660
rect 11517 34595 11575 34601
rect 11517 34592 11529 34595
rect 11348 34564 11529 34592
rect 11517 34561 11529 34564
rect 11563 34561 11575 34595
rect 11517 34555 11575 34561
rect 11698 34552 11704 34604
rect 11756 34552 11762 34604
rect 11900 34601 11928 34632
rect 12158 34601 12164 34604
rect 11885 34595 11943 34601
rect 11885 34561 11897 34595
rect 11931 34561 11943 34595
rect 11885 34555 11943 34561
rect 12152 34555 12164 34601
rect 11900 34524 11928 34555
rect 12158 34552 12164 34555
rect 12216 34552 12222 34604
rect 12406 34592 12434 34632
rect 13464 34632 14096 34660
rect 13464 34601 13492 34632
rect 14090 34620 14096 34632
rect 14148 34620 14154 34672
rect 15372 34663 15430 34669
rect 15372 34629 15384 34663
rect 15418 34660 15430 34663
rect 16684 34660 16712 34691
rect 17034 34688 17040 34740
rect 17092 34688 17098 34740
rect 18233 34731 18291 34737
rect 18233 34697 18245 34731
rect 18279 34697 18291 34731
rect 18233 34691 18291 34697
rect 15418 34632 16712 34660
rect 15418 34629 15430 34632
rect 15372 34623 15430 34629
rect 13722 34601 13728 34604
rect 13449 34595 13507 34601
rect 13449 34592 13461 34595
rect 12406 34564 13461 34592
rect 13449 34561 13461 34564
rect 13495 34561 13507 34595
rect 13449 34555 13507 34561
rect 13716 34555 13728 34601
rect 13722 34552 13728 34555
rect 13780 34552 13786 34604
rect 14108 34592 14136 34620
rect 15105 34595 15163 34601
rect 15105 34592 15117 34595
rect 14108 34564 15117 34592
rect 15105 34561 15117 34564
rect 15151 34592 15163 34595
rect 15151 34564 16160 34592
rect 15151 34561 15163 34564
rect 15105 34555 15163 34561
rect 11256 34496 11928 34524
rect 16132 34524 16160 34564
rect 16850 34552 16856 34604
rect 16908 34552 16914 34604
rect 17221 34595 17279 34601
rect 17221 34561 17233 34595
rect 17267 34592 17279 34595
rect 18248 34592 18276 34691
rect 18322 34688 18328 34740
rect 18380 34728 18386 34740
rect 19981 34731 20039 34737
rect 19981 34728 19993 34731
rect 18380 34700 19993 34728
rect 18380 34688 18386 34700
rect 19981 34697 19993 34700
rect 20027 34697 20039 34731
rect 19981 34691 20039 34697
rect 21082 34688 21088 34740
rect 21140 34728 21146 34740
rect 21821 34731 21879 34737
rect 21821 34728 21833 34731
rect 21140 34700 21833 34728
rect 21140 34688 21146 34700
rect 21821 34697 21833 34700
rect 21867 34697 21879 34731
rect 21821 34691 21879 34697
rect 23845 34731 23903 34737
rect 23845 34697 23857 34731
rect 23891 34728 23903 34731
rect 23934 34728 23940 34740
rect 23891 34700 23940 34728
rect 23891 34697 23903 34700
rect 23845 34691 23903 34697
rect 23934 34688 23940 34700
rect 23992 34688 23998 34740
rect 24302 34688 24308 34740
rect 24360 34688 24366 34740
rect 24946 34688 24952 34740
rect 25004 34728 25010 34740
rect 26053 34731 26111 34737
rect 26053 34728 26065 34731
rect 25004 34700 26065 34728
rect 25004 34688 25010 34700
rect 26053 34697 26065 34700
rect 26099 34697 26111 34731
rect 26053 34691 26111 34697
rect 18690 34620 18696 34672
rect 18748 34620 18754 34672
rect 20346 34620 20352 34672
rect 20404 34660 20410 34672
rect 22189 34663 22247 34669
rect 22189 34660 22201 34663
rect 20404 34632 22201 34660
rect 20404 34620 20410 34632
rect 22189 34629 22201 34632
rect 22235 34629 22247 34663
rect 24320 34660 24348 34688
rect 25406 34660 25412 34672
rect 24320 34632 25412 34660
rect 22189 34623 22247 34629
rect 25406 34620 25412 34632
rect 25464 34620 25470 34672
rect 29270 34660 29276 34672
rect 25516 34632 29276 34660
rect 17267 34564 18276 34592
rect 18601 34595 18659 34601
rect 17267 34561 17279 34564
rect 17221 34555 17279 34561
rect 18601 34561 18613 34595
rect 18647 34561 18659 34595
rect 18601 34555 18659 34561
rect 19061 34595 19119 34601
rect 19061 34561 19073 34595
rect 19107 34561 19119 34595
rect 19061 34555 19119 34561
rect 17126 34524 17132 34536
rect 16132 34496 17132 34524
rect 17126 34484 17132 34496
rect 17184 34524 17190 34536
rect 17184 34496 17264 34524
rect 17184 34484 17190 34496
rect 5261 34459 5319 34465
rect 5261 34456 5273 34459
rect 4724 34428 5273 34456
rect 4724 34400 4752 34428
rect 5261 34425 5273 34428
rect 5307 34425 5319 34459
rect 5261 34419 5319 34425
rect 4706 34348 4712 34400
rect 4764 34348 4770 34400
rect 6932 34388 6960 34484
rect 17236 34456 17264 34496
rect 17310 34484 17316 34536
rect 17368 34484 17374 34536
rect 17589 34527 17647 34533
rect 17589 34524 17601 34527
rect 17420 34496 17601 34524
rect 17420 34456 17448 34496
rect 17589 34493 17601 34496
rect 17635 34493 17647 34527
rect 17589 34487 17647 34493
rect 17678 34484 17684 34536
rect 17736 34524 17742 34536
rect 18616 34524 18644 34555
rect 17736 34496 18644 34524
rect 17736 34484 17742 34496
rect 18782 34484 18788 34536
rect 18840 34484 18846 34536
rect 19076 34524 19104 34555
rect 19794 34552 19800 34604
rect 19852 34552 19858 34604
rect 23842 34552 23848 34604
rect 23900 34592 23906 34604
rect 24213 34595 24271 34601
rect 24213 34592 24225 34595
rect 23900 34564 24225 34592
rect 23900 34552 23906 34564
rect 24213 34561 24225 34564
rect 24259 34592 24271 34595
rect 24762 34592 24768 34604
rect 24259 34564 24768 34592
rect 24259 34561 24271 34564
rect 24213 34555 24271 34561
rect 24762 34552 24768 34564
rect 24820 34552 24826 34604
rect 25516 34592 25544 34632
rect 29270 34620 29276 34632
rect 29328 34620 29334 34672
rect 25148 34564 25544 34592
rect 19076 34496 20576 34524
rect 17236 34428 17448 34456
rect 18800 34456 18828 34484
rect 19245 34459 19303 34465
rect 19245 34456 19257 34459
rect 18800 34428 19257 34456
rect 19245 34425 19257 34428
rect 19291 34425 19303 34459
rect 20548 34456 20576 34496
rect 22094 34484 22100 34536
rect 22152 34524 22158 34536
rect 22281 34527 22339 34533
rect 22281 34524 22293 34527
rect 22152 34496 22293 34524
rect 22152 34484 22158 34496
rect 22281 34493 22293 34496
rect 22327 34493 22339 34527
rect 22281 34487 22339 34493
rect 22465 34527 22523 34533
rect 22465 34493 22477 34527
rect 22511 34493 22523 34527
rect 22465 34487 22523 34493
rect 22480 34456 22508 34487
rect 24486 34484 24492 34536
rect 24544 34484 24550 34536
rect 25038 34484 25044 34536
rect 25096 34524 25102 34536
rect 25148 34533 25176 34564
rect 25590 34552 25596 34604
rect 25648 34592 25654 34604
rect 26421 34595 26479 34601
rect 26421 34592 26433 34595
rect 25648 34564 26433 34592
rect 25648 34552 25654 34564
rect 26421 34561 26433 34564
rect 26467 34561 26479 34595
rect 26421 34555 26479 34561
rect 25133 34527 25191 34533
rect 25133 34524 25145 34527
rect 25096 34496 25145 34524
rect 25096 34484 25102 34496
rect 25133 34493 25145 34496
rect 25179 34493 25191 34527
rect 25133 34487 25191 34493
rect 25409 34527 25467 34533
rect 25409 34493 25421 34527
rect 25455 34524 25467 34527
rect 25498 34524 25504 34536
rect 25455 34496 25504 34524
rect 25455 34493 25467 34496
rect 25409 34487 25467 34493
rect 25498 34484 25504 34496
rect 25556 34524 25562 34536
rect 26326 34524 26332 34536
rect 25556 34496 26332 34524
rect 25556 34484 25562 34496
rect 26326 34484 26332 34496
rect 26384 34484 26390 34536
rect 26510 34484 26516 34536
rect 26568 34484 26574 34536
rect 26697 34527 26755 34533
rect 26697 34493 26709 34527
rect 26743 34493 26755 34527
rect 26697 34487 26755 34493
rect 24504 34456 24532 34484
rect 26602 34456 26608 34468
rect 20548 34428 22600 34456
rect 24504 34428 26608 34456
rect 19245 34419 19303 34425
rect 7098 34388 7104 34400
rect 6932 34360 7104 34388
rect 7098 34348 7104 34360
rect 7156 34348 7162 34400
rect 7558 34348 7564 34400
rect 7616 34388 7622 34400
rect 8297 34391 8355 34397
rect 8297 34388 8309 34391
rect 7616 34360 8309 34388
rect 7616 34348 7622 34360
rect 8297 34357 8309 34360
rect 8343 34357 8355 34391
rect 8297 34351 8355 34357
rect 11606 34348 11612 34400
rect 11664 34348 11670 34400
rect 12986 34348 12992 34400
rect 13044 34388 13050 34400
rect 13265 34391 13323 34397
rect 13265 34388 13277 34391
rect 13044 34360 13277 34388
rect 13044 34348 13050 34360
rect 13265 34357 13277 34360
rect 13311 34357 13323 34391
rect 13265 34351 13323 34357
rect 16485 34391 16543 34397
rect 16485 34357 16497 34391
rect 16531 34388 16543 34391
rect 16666 34388 16672 34400
rect 16531 34360 16672 34388
rect 16531 34357 16543 34360
rect 16485 34351 16543 34357
rect 16666 34348 16672 34360
rect 16724 34348 16730 34400
rect 22572 34388 22600 34428
rect 26602 34416 26608 34428
rect 26660 34416 26666 34468
rect 26712 34456 26740 34487
rect 28626 34456 28632 34468
rect 26712 34428 28632 34456
rect 26712 34388 26740 34428
rect 28626 34416 28632 34428
rect 28684 34416 28690 34468
rect 22572 34360 26740 34388
rect 1104 34298 36800 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 36800 34298
rect 1104 34224 36800 34246
rect 4249 34187 4307 34193
rect 4249 34153 4261 34187
rect 4295 34184 4307 34187
rect 4614 34184 4620 34196
rect 4295 34156 4620 34184
rect 4295 34153 4307 34156
rect 4249 34147 4307 34153
rect 4614 34144 4620 34156
rect 4672 34144 4678 34196
rect 7006 34144 7012 34196
rect 7064 34184 7070 34196
rect 7101 34187 7159 34193
rect 7101 34184 7113 34187
rect 7064 34156 7113 34184
rect 7064 34144 7070 34156
rect 7101 34153 7113 34156
rect 7147 34153 7159 34187
rect 7101 34147 7159 34153
rect 8478 34144 8484 34196
rect 8536 34184 8542 34196
rect 9125 34187 9183 34193
rect 9125 34184 9137 34187
rect 8536 34156 9137 34184
rect 8536 34144 8542 34156
rect 9125 34153 9137 34156
rect 9171 34153 9183 34187
rect 9125 34147 9183 34153
rect 10226 34144 10232 34196
rect 10284 34184 10290 34196
rect 10413 34187 10471 34193
rect 10413 34184 10425 34187
rect 10284 34156 10425 34184
rect 10284 34144 10290 34156
rect 10413 34153 10425 34156
rect 10459 34153 10471 34187
rect 10413 34147 10471 34153
rect 12158 34144 12164 34196
rect 12216 34184 12222 34196
rect 12253 34187 12311 34193
rect 12253 34184 12265 34187
rect 12216 34156 12265 34184
rect 12216 34144 12222 34156
rect 12253 34153 12265 34156
rect 12299 34153 12311 34187
rect 13633 34187 13691 34193
rect 12253 34147 12311 34153
rect 12406 34156 13216 34184
rect 10318 34076 10324 34128
rect 10376 34076 10382 34128
rect 11054 34076 11060 34128
rect 11112 34116 11118 34128
rect 12406 34116 12434 34156
rect 11112 34088 12434 34116
rect 12529 34119 12587 34125
rect 11112 34076 11118 34088
rect 12529 34085 12541 34119
rect 12575 34085 12587 34119
rect 12529 34079 12587 34085
rect 3786 34008 3792 34060
rect 3844 34048 3850 34060
rect 4801 34051 4859 34057
rect 4801 34048 4813 34051
rect 3844 34020 4813 34048
rect 3844 34008 3850 34020
rect 4801 34017 4813 34020
rect 4847 34017 4859 34051
rect 4801 34011 4859 34017
rect 6917 34051 6975 34057
rect 6917 34017 6929 34051
rect 6963 34017 6975 34051
rect 6917 34011 6975 34017
rect 4433 33983 4491 33989
rect 4433 33949 4445 33983
rect 4479 33980 4491 33983
rect 4706 33980 4712 33992
rect 4479 33952 4712 33980
rect 4479 33949 4491 33952
rect 4433 33943 4491 33949
rect 4706 33940 4712 33952
rect 4764 33940 4770 33992
rect 5626 33940 5632 33992
rect 5684 33980 5690 33992
rect 6641 33983 6699 33989
rect 6641 33980 6653 33983
rect 5684 33952 6653 33980
rect 5684 33940 5690 33952
rect 6641 33949 6653 33952
rect 6687 33949 6699 33983
rect 6932 33980 6960 34011
rect 7006 34008 7012 34060
rect 7064 34048 7070 34060
rect 7558 34048 7564 34060
rect 7064 34020 7564 34048
rect 7064 34008 7070 34020
rect 7558 34008 7564 34020
rect 7616 34008 7622 34060
rect 7745 34051 7803 34057
rect 7745 34017 7757 34051
rect 7791 34017 7803 34051
rect 7745 34011 7803 34017
rect 10505 34051 10563 34057
rect 10505 34017 10517 34051
rect 10551 34048 10563 34051
rect 11606 34048 11612 34060
rect 10551 34020 11612 34048
rect 10551 34017 10563 34020
rect 10505 34011 10563 34017
rect 7760 33980 7788 34011
rect 11606 34008 11612 34020
rect 11664 34008 11670 34060
rect 10229 33983 10287 33989
rect 10229 33980 10241 33983
rect 6932 33952 10241 33980
rect 6641 33943 6699 33949
rect 10229 33949 10241 33952
rect 10275 33949 10287 33983
rect 10229 33943 10287 33949
rect 12437 33983 12495 33989
rect 12437 33949 12449 33983
rect 12483 33980 12495 33983
rect 12544 33980 12572 34079
rect 12986 34008 12992 34060
rect 13044 34008 13050 34060
rect 13188 34057 13216 34156
rect 13633 34153 13645 34187
rect 13679 34184 13691 34187
rect 13722 34184 13728 34196
rect 13679 34156 13728 34184
rect 13679 34153 13691 34156
rect 13633 34147 13691 34153
rect 13722 34144 13728 34156
rect 13780 34144 13786 34196
rect 16209 34187 16267 34193
rect 16209 34153 16221 34187
rect 16255 34184 16267 34187
rect 16850 34184 16856 34196
rect 16255 34156 16856 34184
rect 16255 34153 16267 34156
rect 16209 34147 16267 34153
rect 16850 34144 16856 34156
rect 16908 34144 16914 34196
rect 26602 34144 26608 34196
rect 26660 34184 26666 34196
rect 30282 34184 30288 34196
rect 26660 34156 30288 34184
rect 26660 34144 26666 34156
rect 30282 34144 30288 34156
rect 30340 34144 30346 34196
rect 17862 34116 17868 34128
rect 16684 34088 17868 34116
rect 16684 34060 16712 34088
rect 17862 34076 17868 34088
rect 17920 34076 17926 34128
rect 13173 34051 13231 34057
rect 13173 34017 13185 34051
rect 13219 34048 13231 34051
rect 13219 34020 14228 34048
rect 13219 34017 13231 34020
rect 13173 34011 13231 34017
rect 12483 33952 12572 33980
rect 12483 33949 12495 33952
rect 12437 33943 12495 33949
rect 5068 33915 5126 33921
rect 5068 33881 5080 33915
rect 5114 33912 5126 33915
rect 5258 33912 5264 33924
rect 5114 33884 5264 33912
rect 5114 33881 5126 33884
rect 5068 33875 5126 33881
rect 5258 33872 5264 33884
rect 5316 33872 5322 33924
rect 6733 33915 6791 33921
rect 6733 33912 6745 33915
rect 6196 33884 6745 33912
rect 5350 33804 5356 33856
rect 5408 33844 5414 33856
rect 6196 33853 6224 33884
rect 6733 33881 6745 33884
rect 6779 33881 6791 33915
rect 6733 33875 6791 33881
rect 7098 33872 7104 33924
rect 7156 33912 7162 33924
rect 9033 33915 9091 33921
rect 9033 33912 9045 33915
rect 7156 33884 9045 33912
rect 7156 33872 7162 33884
rect 9033 33881 9045 33884
rect 9079 33912 9091 33915
rect 9766 33912 9772 33924
rect 9079 33884 9772 33912
rect 9079 33881 9091 33884
rect 9033 33875 9091 33881
rect 9766 33872 9772 33884
rect 9824 33872 9830 33924
rect 10244 33912 10272 33943
rect 12894 33940 12900 33992
rect 12952 33980 12958 33992
rect 13078 33980 13084 33992
rect 12952 33952 13084 33980
rect 12952 33940 12958 33952
rect 13078 33940 13084 33952
rect 13136 33940 13142 33992
rect 13814 33940 13820 33992
rect 13872 33940 13878 33992
rect 14090 33940 14096 33992
rect 14148 33940 14154 33992
rect 14200 33980 14228 34020
rect 16666 34008 16672 34060
rect 16724 34008 16730 34060
rect 16853 34051 16911 34057
rect 16853 34017 16865 34051
rect 16899 34048 16911 34051
rect 18322 34048 18328 34060
rect 16899 34020 18328 34048
rect 16899 34017 16911 34020
rect 16853 34011 16911 34017
rect 16868 33980 16896 34011
rect 18322 34008 18328 34020
rect 18380 34008 18386 34060
rect 14200 33952 16896 33980
rect 11698 33912 11704 33924
rect 10244 33884 11704 33912
rect 11698 33872 11704 33884
rect 11756 33872 11762 33924
rect 14366 33921 14372 33924
rect 14360 33875 14372 33921
rect 14366 33872 14372 33875
rect 14424 33872 14430 33924
rect 16577 33915 16635 33921
rect 16577 33881 16589 33915
rect 16623 33912 16635 33915
rect 17678 33912 17684 33924
rect 16623 33884 17684 33912
rect 16623 33881 16635 33884
rect 16577 33875 16635 33881
rect 17678 33872 17684 33884
rect 17736 33872 17742 33924
rect 6181 33847 6239 33853
rect 6181 33844 6193 33847
rect 5408 33816 6193 33844
rect 5408 33804 5414 33816
rect 6181 33813 6193 33816
rect 6227 33813 6239 33847
rect 6181 33807 6239 33813
rect 6270 33804 6276 33856
rect 6328 33804 6334 33856
rect 7282 33804 7288 33856
rect 7340 33844 7346 33856
rect 7469 33847 7527 33853
rect 7469 33844 7481 33847
rect 7340 33816 7481 33844
rect 7340 33804 7346 33816
rect 7469 33813 7481 33816
rect 7515 33813 7527 33847
rect 7469 33807 7527 33813
rect 15194 33804 15200 33856
rect 15252 33844 15258 33856
rect 15473 33847 15531 33853
rect 15473 33844 15485 33847
rect 15252 33816 15485 33844
rect 15252 33804 15258 33816
rect 15473 33813 15485 33816
rect 15519 33813 15531 33847
rect 15473 33807 15531 33813
rect 1104 33754 36800 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 36800 33754
rect 1104 33680 36800 33702
rect 5169 33643 5227 33649
rect 5169 33609 5181 33643
rect 5215 33640 5227 33643
rect 5258 33640 5264 33652
rect 5215 33612 5264 33640
rect 5215 33609 5227 33612
rect 5169 33603 5227 33609
rect 5258 33600 5264 33612
rect 5316 33600 5322 33652
rect 14277 33643 14335 33649
rect 14277 33609 14289 33643
rect 14323 33640 14335 33643
rect 14366 33640 14372 33652
rect 14323 33612 14372 33640
rect 14323 33609 14335 33612
rect 14277 33603 14335 33609
rect 14366 33600 14372 33612
rect 14424 33600 14430 33652
rect 17129 33643 17187 33649
rect 17129 33609 17141 33643
rect 17175 33609 17187 33643
rect 17129 33603 17187 33609
rect 26513 33643 26571 33649
rect 26513 33609 26525 33643
rect 26559 33609 26571 33643
rect 26513 33603 26571 33609
rect 17144 33572 17172 33603
rect 17650 33575 17708 33581
rect 17650 33572 17662 33575
rect 17144 33544 17662 33572
rect 17650 33541 17662 33544
rect 17696 33541 17708 33575
rect 26528 33572 26556 33603
rect 27218 33575 27276 33581
rect 27218 33572 27230 33575
rect 26528 33544 27230 33572
rect 17650 33535 17708 33541
rect 27218 33541 27230 33544
rect 27264 33541 27276 33575
rect 27218 33535 27276 33541
rect 5353 33507 5411 33513
rect 5353 33473 5365 33507
rect 5399 33504 5411 33507
rect 6270 33504 6276 33516
rect 5399 33476 6276 33504
rect 5399 33473 5411 33476
rect 5353 33467 5411 33473
rect 6270 33464 6276 33476
rect 6328 33464 6334 33516
rect 14458 33464 14464 33516
rect 14516 33464 14522 33516
rect 17310 33464 17316 33516
rect 17368 33464 17374 33516
rect 17402 33464 17408 33516
rect 17460 33464 17466 33516
rect 18874 33464 18880 33516
rect 18932 33504 18938 33516
rect 19409 33507 19467 33513
rect 19409 33504 19421 33507
rect 18932 33476 19421 33504
rect 18932 33464 18938 33476
rect 19409 33473 19421 33476
rect 19455 33473 19467 33507
rect 19409 33467 19467 33473
rect 21266 33464 21272 33516
rect 21324 33504 21330 33516
rect 21913 33507 21971 33513
rect 21913 33504 21925 33507
rect 21324 33476 21925 33504
rect 21324 33464 21330 33476
rect 21913 33473 21925 33476
rect 21959 33473 21971 33507
rect 21913 33467 21971 33473
rect 22180 33507 22238 33513
rect 22180 33473 22192 33507
rect 22226 33504 22238 33507
rect 22738 33504 22744 33516
rect 22226 33476 22744 33504
rect 22226 33473 22238 33476
rect 22180 33467 22238 33473
rect 22738 33464 22744 33476
rect 22796 33464 22802 33516
rect 24029 33507 24087 33513
rect 24029 33473 24041 33507
rect 24075 33504 24087 33507
rect 24394 33504 24400 33516
rect 24075 33476 24400 33504
rect 24075 33473 24087 33476
rect 24029 33467 24087 33473
rect 24394 33464 24400 33476
rect 24452 33464 24458 33516
rect 26694 33464 26700 33516
rect 26752 33464 26758 33516
rect 35986 33464 35992 33516
rect 36044 33504 36050 33516
rect 36173 33507 36231 33513
rect 36173 33504 36185 33507
rect 36044 33476 36185 33504
rect 36044 33464 36050 33476
rect 36173 33473 36185 33476
rect 36219 33473 36231 33507
rect 36173 33467 36231 33473
rect 19150 33396 19156 33448
rect 19208 33396 19214 33448
rect 24121 33439 24179 33445
rect 24121 33405 24133 33439
rect 24167 33405 24179 33439
rect 24121 33399 24179 33405
rect 24136 33368 24164 33399
rect 24302 33396 24308 33448
rect 24360 33396 24366 33448
rect 26326 33396 26332 33448
rect 26384 33436 26390 33448
rect 26973 33439 27031 33445
rect 26973 33436 26985 33439
rect 26384 33408 26985 33436
rect 26384 33396 26390 33408
rect 26973 33405 26985 33408
rect 27019 33405 27031 33439
rect 26973 33399 27031 33405
rect 26418 33368 26424 33380
rect 24136 33340 26424 33368
rect 26418 33328 26424 33340
rect 26476 33368 26482 33380
rect 26878 33368 26884 33380
rect 26476 33340 26884 33368
rect 26476 33328 26482 33340
rect 26878 33328 26884 33340
rect 26936 33328 26942 33380
rect 36354 33328 36360 33380
rect 36412 33328 36418 33380
rect 18782 33260 18788 33312
rect 18840 33260 18846 33312
rect 20254 33260 20260 33312
rect 20312 33300 20318 33312
rect 20533 33303 20591 33309
rect 20533 33300 20545 33303
rect 20312 33272 20545 33300
rect 20312 33260 20318 33272
rect 20533 33269 20545 33272
rect 20579 33269 20591 33303
rect 20533 33263 20591 33269
rect 22278 33260 22284 33312
rect 22336 33300 22342 33312
rect 23293 33303 23351 33309
rect 23293 33300 23305 33303
rect 22336 33272 23305 33300
rect 22336 33260 22342 33272
rect 23293 33269 23305 33272
rect 23339 33269 23351 33303
rect 23293 33263 23351 33269
rect 23661 33303 23719 33309
rect 23661 33269 23673 33303
rect 23707 33300 23719 33303
rect 24210 33300 24216 33312
rect 23707 33272 24216 33300
rect 23707 33269 23719 33272
rect 23661 33263 23719 33269
rect 24210 33260 24216 33272
rect 24268 33260 24274 33312
rect 28350 33260 28356 33312
rect 28408 33260 28414 33312
rect 1104 33210 36800 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 36800 33210
rect 1104 33136 36800 33158
rect 2682 33056 2688 33108
rect 2740 33096 2746 33108
rect 3053 33099 3111 33105
rect 3053 33096 3065 33099
rect 2740 33068 3065 33096
rect 2740 33056 2746 33068
rect 3053 33065 3065 33068
rect 3099 33096 3111 33099
rect 7374 33096 7380 33108
rect 3099 33068 4844 33096
rect 3099 33065 3111 33068
rect 3053 33059 3111 33065
rect 3786 32960 3792 32972
rect 3528 32932 3792 32960
rect 1673 32895 1731 32901
rect 1673 32861 1685 32895
rect 1719 32892 1731 32895
rect 3528 32892 3556 32932
rect 3786 32920 3792 32932
rect 3844 32920 3850 32972
rect 1719 32864 3556 32892
rect 1719 32861 1731 32864
rect 1673 32855 1731 32861
rect 3602 32852 3608 32904
rect 3660 32852 3666 32904
rect 4816 32892 4844 33068
rect 7116 33068 7380 33096
rect 6822 33028 6828 33040
rect 6656 33000 6828 33028
rect 6656 32969 6684 33000
rect 6822 32988 6828 33000
rect 6880 32988 6886 33040
rect 6641 32963 6699 32969
rect 6641 32929 6653 32963
rect 6687 32929 6699 32963
rect 7116 32960 7144 33068
rect 7374 33056 7380 33068
rect 7432 33096 7438 33108
rect 9490 33096 9496 33108
rect 7432 33068 9496 33096
rect 7432 33056 7438 33068
rect 9490 33056 9496 33068
rect 9548 33056 9554 33108
rect 9674 33056 9680 33108
rect 9732 33096 9738 33108
rect 9732 33068 11744 33096
rect 9732 33056 9738 33068
rect 7190 32988 7196 33040
rect 7248 33028 7254 33040
rect 7248 33000 7420 33028
rect 7248 32988 7254 33000
rect 7285 32963 7343 32969
rect 7285 32960 7297 32963
rect 7116 32932 7297 32960
rect 6641 32923 6699 32929
rect 7285 32929 7297 32932
rect 7331 32929 7343 32963
rect 7392 32960 7420 33000
rect 9858 32988 9864 33040
rect 9916 33028 9922 33040
rect 9916 33000 10824 33028
rect 9916 32988 9922 33000
rect 7561 32963 7619 32969
rect 7561 32960 7573 32963
rect 7392 32932 7573 32960
rect 7285 32923 7343 32929
rect 7561 32929 7573 32932
rect 7607 32929 7619 32963
rect 7561 32923 7619 32929
rect 7837 32963 7895 32969
rect 7837 32929 7849 32963
rect 7883 32960 7895 32963
rect 8018 32960 8024 32972
rect 7883 32932 8024 32960
rect 7883 32929 7895 32932
rect 7837 32923 7895 32929
rect 8018 32920 8024 32932
rect 8076 32920 8082 32972
rect 10686 32920 10692 32972
rect 10744 32920 10750 32972
rect 10796 32960 10824 33000
rect 11241 32963 11299 32969
rect 10796 32932 11008 32960
rect 10980 32904 11008 32932
rect 11241 32929 11253 32963
rect 11287 32960 11299 32963
rect 11422 32960 11428 32972
rect 11287 32932 11428 32960
rect 11287 32929 11299 32932
rect 11241 32923 11299 32929
rect 11422 32920 11428 32932
rect 11480 32920 11486 32972
rect 11716 32960 11744 33068
rect 11790 33056 11796 33108
rect 11848 33096 11854 33108
rect 14182 33096 14188 33108
rect 11848 33068 14188 33096
rect 11848 33056 11854 33068
rect 14182 33056 14188 33068
rect 14240 33056 14246 33108
rect 14277 33099 14335 33105
rect 14277 33065 14289 33099
rect 14323 33096 14335 33099
rect 14458 33096 14464 33108
rect 14323 33068 14464 33096
rect 14323 33065 14335 33068
rect 14277 33059 14335 33065
rect 14458 33056 14464 33068
rect 14516 33056 14522 33108
rect 15488 33068 16528 33096
rect 14829 32963 14887 32969
rect 14829 32960 14841 32963
rect 11716 32932 14841 32960
rect 14829 32929 14841 32932
rect 14875 32960 14887 32963
rect 15488 32960 15516 33068
rect 14875 32932 15516 32960
rect 16500 32960 16528 33068
rect 17310 33056 17316 33108
rect 17368 33096 17374 33108
rect 17497 33099 17555 33105
rect 17497 33096 17509 33099
rect 17368 33068 17509 33096
rect 17368 33056 17374 33068
rect 17497 33065 17509 33068
rect 17543 33065 17555 33099
rect 17497 33059 17555 33065
rect 18874 33056 18880 33108
rect 18932 33056 18938 33108
rect 22094 33096 22100 33108
rect 20180 33068 22100 33096
rect 17034 32988 17040 33040
rect 17092 33028 17098 33040
rect 18690 33028 18696 33040
rect 17092 33000 18696 33028
rect 17092 32988 17098 33000
rect 18690 32988 18696 33000
rect 18748 32988 18754 33040
rect 19337 33031 19395 33037
rect 19337 32997 19349 33031
rect 19383 32997 19395 33031
rect 19337 32991 19395 32997
rect 18046 32960 18052 32972
rect 16500 32932 18052 32960
rect 14875 32929 14887 32932
rect 14829 32923 14887 32929
rect 18046 32920 18052 32932
rect 18104 32920 18110 32972
rect 6822 32892 6828 32904
rect 4816 32864 6828 32892
rect 6822 32852 6828 32864
rect 6880 32852 6886 32904
rect 7650 32852 7656 32904
rect 7708 32901 7714 32904
rect 7708 32895 7736 32901
rect 7724 32861 7736 32895
rect 7708 32855 7736 32861
rect 7708 32852 7714 32855
rect 10042 32852 10048 32904
rect 10100 32852 10106 32904
rect 10226 32852 10232 32904
rect 10284 32852 10290 32904
rect 10962 32852 10968 32904
rect 11020 32852 11026 32904
rect 11054 32852 11060 32904
rect 11112 32901 11118 32904
rect 11112 32895 11140 32901
rect 11128 32861 11140 32895
rect 11112 32855 11140 32861
rect 11112 32852 11118 32855
rect 12434 32852 12440 32904
rect 12492 32852 12498 32904
rect 14645 32895 14703 32901
rect 14645 32861 14657 32895
rect 14691 32892 14703 32895
rect 15194 32892 15200 32904
rect 14691 32864 15200 32892
rect 14691 32861 14703 32864
rect 14645 32855 14703 32861
rect 15194 32852 15200 32864
rect 15252 32852 15258 32904
rect 15470 32852 15476 32904
rect 15528 32852 15534 32904
rect 17865 32895 17923 32901
rect 15580 32864 17080 32892
rect 1946 32833 1952 32836
rect 1940 32787 1952 32833
rect 1946 32784 1952 32787
rect 2004 32784 2010 32836
rect 4034 32827 4092 32833
rect 4034 32824 4046 32827
rect 3436 32796 4046 32824
rect 3436 32765 3464 32796
rect 4034 32793 4046 32796
rect 4080 32793 4092 32827
rect 4034 32787 4092 32793
rect 12894 32784 12900 32836
rect 12952 32824 12958 32836
rect 14737 32827 14795 32833
rect 14737 32824 14749 32827
rect 12952 32796 14749 32824
rect 12952 32784 12958 32796
rect 14737 32793 14749 32796
rect 14783 32793 14795 32827
rect 14737 32787 14795 32793
rect 3421 32759 3479 32765
rect 3421 32725 3433 32759
rect 3467 32725 3479 32759
rect 3421 32719 3479 32725
rect 4246 32716 4252 32768
rect 4304 32756 4310 32768
rect 5169 32759 5227 32765
rect 5169 32756 5181 32759
rect 4304 32728 5181 32756
rect 4304 32716 4310 32728
rect 5169 32725 5181 32728
rect 5215 32756 5227 32759
rect 7650 32756 7656 32768
rect 5215 32728 7656 32756
rect 5215 32725 5227 32728
rect 5169 32719 5227 32725
rect 7650 32716 7656 32728
rect 7708 32716 7714 32768
rect 8481 32759 8539 32765
rect 8481 32725 8493 32759
rect 8527 32756 8539 32759
rect 9582 32756 9588 32768
rect 8527 32728 9588 32756
rect 8527 32725 8539 32728
rect 8481 32719 8539 32725
rect 9582 32716 9588 32728
rect 9640 32716 9646 32768
rect 11514 32716 11520 32768
rect 11572 32756 11578 32768
rect 11885 32759 11943 32765
rect 11885 32756 11897 32759
rect 11572 32728 11897 32756
rect 11572 32716 11578 32728
rect 11885 32725 11897 32728
rect 11931 32725 11943 32759
rect 11885 32719 11943 32725
rect 12250 32716 12256 32768
rect 12308 32716 12314 32768
rect 13170 32716 13176 32768
rect 13228 32756 13234 32768
rect 15580 32756 15608 32864
rect 15740 32827 15798 32833
rect 15740 32793 15752 32827
rect 15786 32824 15798 32827
rect 16022 32824 16028 32836
rect 15786 32796 16028 32824
rect 15786 32793 15798 32796
rect 15740 32787 15798 32793
rect 16022 32784 16028 32796
rect 16080 32784 16086 32836
rect 16206 32784 16212 32836
rect 16264 32824 16270 32836
rect 17052 32824 17080 32864
rect 17865 32861 17877 32895
rect 17911 32892 17923 32895
rect 17954 32892 17960 32904
rect 17911 32864 17960 32892
rect 17911 32861 17923 32864
rect 17865 32855 17923 32861
rect 17954 32852 17960 32864
rect 18012 32892 18018 32904
rect 18782 32892 18788 32904
rect 18012 32864 18788 32892
rect 18012 32852 18018 32864
rect 18782 32852 18788 32864
rect 18840 32852 18846 32904
rect 19061 32895 19119 32901
rect 19061 32861 19073 32895
rect 19107 32892 19119 32895
rect 19352 32892 19380 32991
rect 19978 32920 19984 32972
rect 20036 32920 20042 32972
rect 20180 32969 20208 33068
rect 22094 33056 22100 33068
rect 22152 33056 22158 33108
rect 22186 33056 22192 33108
rect 22244 33096 22250 33108
rect 23937 33099 23995 33105
rect 23937 33096 23949 33099
rect 22244 33068 23949 33096
rect 22244 33056 22250 33068
rect 23937 33065 23949 33068
rect 23983 33065 23995 33099
rect 25682 33096 25688 33108
rect 23937 33059 23995 33065
rect 24596 33068 25688 33096
rect 20254 32988 20260 33040
rect 20312 33028 20318 33040
rect 20312 33000 20944 33028
rect 20312 32988 20318 33000
rect 20165 32963 20223 32969
rect 20165 32929 20177 32963
rect 20211 32929 20223 32963
rect 20165 32923 20223 32929
rect 20806 32920 20812 32972
rect 20864 32920 20870 32972
rect 20916 32960 20944 33000
rect 21744 33000 22876 33028
rect 21202 32963 21260 32969
rect 21202 32960 21214 32963
rect 20916 32932 21214 32960
rect 21202 32929 21214 32932
rect 21248 32960 21260 32963
rect 21744 32960 21772 33000
rect 21248 32932 21772 32960
rect 21248 32929 21260 32932
rect 21202 32923 21260 32929
rect 22094 32920 22100 32972
rect 22152 32920 22158 32972
rect 22278 32920 22284 32972
rect 22336 32920 22342 32972
rect 22646 32920 22652 32972
rect 22704 32960 22710 32972
rect 22741 32963 22799 32969
rect 22741 32960 22753 32963
rect 22704 32932 22753 32960
rect 22704 32920 22710 32932
rect 22741 32929 22753 32932
rect 22787 32929 22799 32963
rect 22848 32960 22876 33000
rect 23134 32963 23192 32969
rect 23134 32960 23146 32963
rect 22848 32932 23146 32960
rect 22741 32923 22799 32929
rect 23134 32929 23146 32932
rect 23180 32929 23192 32963
rect 23134 32923 23192 32929
rect 23293 32963 23351 32969
rect 23293 32929 23305 32963
rect 23339 32960 23351 32963
rect 23474 32960 23480 32972
rect 23339 32932 23480 32960
rect 23339 32929 23351 32932
rect 23293 32923 23351 32929
rect 23474 32920 23480 32932
rect 23532 32960 23538 32972
rect 24596 32960 24624 33068
rect 25682 33056 25688 33068
rect 25740 33096 25746 33108
rect 26142 33096 26148 33108
rect 25740 33068 26148 33096
rect 25740 33056 25746 33068
rect 26142 33056 26148 33068
rect 26200 33056 26206 33108
rect 26421 33099 26479 33105
rect 26421 33065 26433 33099
rect 26467 33096 26479 33099
rect 26694 33096 26700 33108
rect 26467 33068 26700 33096
rect 26467 33065 26479 33068
rect 26421 33059 26479 33065
rect 26694 33056 26700 33068
rect 26752 33056 26758 33108
rect 24688 33000 25268 33028
rect 24688 32969 24716 33000
rect 23532 32932 24624 32960
rect 24673 32963 24731 32969
rect 23532 32920 23538 32932
rect 24673 32929 24685 32963
rect 24719 32960 24731 32963
rect 24762 32960 24768 32972
rect 24719 32932 24768 32960
rect 24719 32929 24731 32932
rect 24673 32923 24731 32929
rect 24762 32920 24768 32932
rect 24820 32920 24826 32972
rect 25133 32963 25191 32969
rect 25133 32960 25145 32963
rect 24872 32932 25145 32960
rect 19107 32864 19380 32892
rect 19705 32895 19763 32901
rect 19107 32861 19119 32864
rect 19061 32855 19119 32861
rect 19705 32861 19717 32895
rect 19751 32892 19763 32895
rect 20254 32892 20260 32904
rect 19751 32864 20260 32892
rect 19751 32861 19763 32864
rect 19705 32855 19763 32861
rect 20254 32852 20260 32864
rect 20312 32852 20318 32904
rect 20349 32895 20407 32901
rect 20349 32861 20361 32895
rect 20395 32861 20407 32895
rect 20349 32855 20407 32861
rect 19150 32824 19156 32836
rect 16264 32796 16988 32824
rect 17052 32796 19156 32824
rect 16264 32784 16270 32796
rect 13228 32728 15608 32756
rect 13228 32716 13234 32728
rect 16850 32716 16856 32768
rect 16908 32716 16914 32768
rect 16960 32756 16988 32796
rect 19150 32784 19156 32796
rect 19208 32784 19214 32836
rect 17957 32759 18015 32765
rect 17957 32756 17969 32759
rect 16960 32728 17969 32756
rect 17957 32725 17969 32728
rect 18003 32725 18015 32759
rect 17957 32719 18015 32725
rect 18322 32716 18328 32768
rect 18380 32756 18386 32768
rect 18874 32756 18880 32768
rect 18380 32728 18880 32756
rect 18380 32716 18386 32728
rect 18874 32716 18880 32728
rect 18932 32716 18938 32768
rect 19797 32759 19855 32765
rect 19797 32725 19809 32759
rect 19843 32756 19855 32759
rect 19886 32756 19892 32768
rect 19843 32728 19892 32756
rect 19843 32725 19855 32728
rect 19797 32719 19855 32725
rect 19886 32716 19892 32728
rect 19944 32716 19950 32768
rect 20364 32756 20392 32855
rect 21082 32852 21088 32904
rect 21140 32852 21146 32904
rect 21358 32852 21364 32904
rect 21416 32852 21422 32904
rect 23014 32852 23020 32904
rect 23072 32852 23078 32904
rect 24210 32852 24216 32904
rect 24268 32852 24274 32904
rect 24486 32852 24492 32904
rect 24544 32852 24550 32904
rect 24872 32892 24900 32932
rect 25133 32929 25145 32932
rect 25179 32929 25191 32963
rect 25240 32960 25268 33000
rect 25240 32932 26832 32960
rect 25133 32923 25191 32929
rect 24688 32864 24900 32892
rect 22278 32824 22284 32836
rect 21836 32796 22284 32824
rect 21836 32756 21864 32796
rect 22278 32784 22284 32796
rect 22336 32784 22342 32836
rect 23934 32784 23940 32836
rect 23992 32824 23998 32836
rect 24688 32824 24716 32864
rect 25406 32852 25412 32904
rect 25464 32852 25470 32904
rect 25498 32852 25504 32904
rect 25556 32901 25562 32904
rect 25556 32895 25584 32901
rect 25572 32861 25584 32895
rect 25556 32855 25584 32861
rect 25556 32852 25562 32855
rect 25682 32852 25688 32904
rect 25740 32852 25746 32904
rect 26804 32901 26832 32932
rect 26878 32920 26884 32972
rect 26936 32920 26942 32972
rect 27065 32963 27123 32969
rect 27065 32929 27077 32963
rect 27111 32960 27123 32963
rect 27614 32960 27620 32972
rect 27111 32932 27620 32960
rect 27111 32929 27123 32932
rect 27065 32923 27123 32929
rect 27614 32920 27620 32932
rect 27672 32960 27678 32972
rect 28166 32960 28172 32972
rect 27672 32932 28172 32960
rect 27672 32920 27678 32932
rect 28166 32920 28172 32932
rect 28224 32920 28230 32972
rect 26789 32895 26847 32901
rect 26789 32861 26801 32895
rect 26835 32892 26847 32895
rect 28350 32892 28356 32904
rect 26835 32864 28356 32892
rect 26835 32861 26847 32864
rect 26789 32855 26847 32861
rect 28350 32852 28356 32864
rect 28408 32852 28414 32904
rect 23992 32796 24716 32824
rect 23992 32784 23998 32796
rect 20364 32728 21864 32756
rect 22002 32716 22008 32768
rect 22060 32716 22066 32768
rect 22094 32716 22100 32768
rect 22152 32756 22158 32768
rect 23014 32756 23020 32768
rect 22152 32728 23020 32756
rect 22152 32716 22158 32728
rect 23014 32716 23020 32728
rect 23072 32716 23078 32768
rect 24026 32716 24032 32768
rect 24084 32716 24090 32768
rect 24394 32716 24400 32768
rect 24452 32756 24458 32768
rect 25498 32756 25504 32768
rect 24452 32728 25504 32756
rect 24452 32716 24458 32728
rect 25498 32716 25504 32728
rect 25556 32716 25562 32768
rect 25682 32716 25688 32768
rect 25740 32756 25746 32768
rect 26329 32759 26387 32765
rect 26329 32756 26341 32759
rect 25740 32728 26341 32756
rect 25740 32716 25746 32728
rect 26329 32725 26341 32728
rect 26375 32725 26387 32759
rect 26329 32719 26387 32725
rect 1104 32666 36800 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 36800 32666
rect 1104 32592 36800 32614
rect 1946 32512 1952 32564
rect 2004 32512 2010 32564
rect 2682 32512 2688 32564
rect 2740 32512 2746 32564
rect 3602 32512 3608 32564
rect 3660 32552 3666 32564
rect 3881 32555 3939 32561
rect 3881 32552 3893 32555
rect 3660 32524 3893 32552
rect 3660 32512 3666 32524
rect 3881 32521 3893 32524
rect 3927 32521 3939 32555
rect 3881 32515 3939 32521
rect 4246 32512 4252 32564
rect 4304 32512 4310 32564
rect 6914 32552 6920 32564
rect 6472 32524 6920 32552
rect 2777 32487 2835 32493
rect 2777 32453 2789 32487
rect 2823 32484 2835 32487
rect 3326 32484 3332 32496
rect 2823 32456 3332 32484
rect 2823 32453 2835 32456
rect 2777 32447 2835 32453
rect 3326 32444 3332 32456
rect 3384 32484 3390 32496
rect 4341 32487 4399 32493
rect 4341 32484 4353 32487
rect 3384 32456 4353 32484
rect 3384 32444 3390 32456
rect 4341 32453 4353 32456
rect 4387 32453 4399 32487
rect 4341 32447 4399 32453
rect 1397 32419 1455 32425
rect 1397 32385 1409 32419
rect 1443 32416 1455 32419
rect 1486 32416 1492 32428
rect 1443 32388 1492 32416
rect 1443 32385 1455 32388
rect 1397 32379 1455 32385
rect 1486 32376 1492 32388
rect 1544 32376 1550 32428
rect 2133 32419 2191 32425
rect 2133 32385 2145 32419
rect 2179 32416 2191 32419
rect 2179 32388 2360 32416
rect 2179 32385 2191 32388
rect 2133 32379 2191 32385
rect 2332 32289 2360 32388
rect 2590 32376 2596 32428
rect 2648 32416 2654 32428
rect 6472 32425 6500 32524
rect 6914 32512 6920 32524
rect 6972 32512 6978 32564
rect 8202 32512 8208 32564
rect 8260 32552 8266 32564
rect 8938 32552 8944 32564
rect 8260 32524 8944 32552
rect 8260 32512 8266 32524
rect 8938 32512 8944 32524
rect 8996 32512 9002 32564
rect 9490 32512 9496 32564
rect 9548 32552 9554 32564
rect 13814 32552 13820 32564
rect 9548 32524 13820 32552
rect 9548 32512 9554 32524
rect 13814 32512 13820 32524
rect 13872 32512 13878 32564
rect 14274 32552 14280 32564
rect 13924 32524 14280 32552
rect 11238 32484 11244 32496
rect 8220 32456 11244 32484
rect 6457 32419 6515 32425
rect 2648 32388 4660 32416
rect 2648 32376 2654 32388
rect 2976 32357 3004 32388
rect 2961 32351 3019 32357
rect 2961 32317 2973 32351
rect 3007 32317 3019 32351
rect 2961 32311 3019 32317
rect 4525 32351 4583 32357
rect 4525 32317 4537 32351
rect 4571 32317 4583 32351
rect 4632 32348 4660 32388
rect 6457 32385 6469 32419
rect 6503 32385 6515 32419
rect 6457 32379 6515 32385
rect 6641 32419 6699 32425
rect 6641 32385 6653 32419
rect 6687 32416 6699 32419
rect 6822 32416 6828 32428
rect 6687 32388 6828 32416
rect 6687 32385 6699 32388
rect 6641 32379 6699 32385
rect 6822 32376 6828 32388
rect 6880 32376 6886 32428
rect 7558 32425 7564 32428
rect 7515 32419 7564 32425
rect 7515 32385 7527 32419
rect 7561 32385 7564 32419
rect 7515 32379 7564 32385
rect 7558 32376 7564 32379
rect 7616 32376 7622 32428
rect 4632 32320 6914 32348
rect 4525 32311 4583 32317
rect 2317 32283 2375 32289
rect 2317 32249 2329 32283
rect 2363 32249 2375 32283
rect 2317 32243 2375 32249
rect 934 32172 940 32224
rect 992 32212 998 32224
rect 1581 32215 1639 32221
rect 1581 32212 1593 32215
rect 992 32184 1593 32212
rect 992 32172 998 32184
rect 1581 32181 1593 32184
rect 1627 32181 1639 32215
rect 4540 32212 4568 32311
rect 6886 32292 6914 32320
rect 7190 32308 7196 32360
rect 7248 32348 7254 32360
rect 7377 32351 7435 32357
rect 7377 32348 7389 32351
rect 7248 32320 7389 32348
rect 7248 32308 7254 32320
rect 7377 32317 7389 32320
rect 7423 32317 7435 32351
rect 7377 32311 7435 32317
rect 7653 32351 7711 32357
rect 7653 32317 7665 32351
rect 7699 32348 7711 32351
rect 7834 32348 7840 32360
rect 7699 32320 7840 32348
rect 7699 32317 7711 32320
rect 7653 32311 7711 32317
rect 7834 32308 7840 32320
rect 7892 32348 7898 32360
rect 8220 32348 8248 32456
rect 11238 32444 11244 32456
rect 11296 32444 11302 32496
rect 12152 32487 12210 32493
rect 12152 32453 12164 32487
rect 12198 32484 12210 32487
rect 12250 32484 12256 32496
rect 12198 32456 12256 32484
rect 12198 32453 12210 32456
rect 12152 32447 12210 32453
rect 12250 32444 12256 32456
rect 12308 32444 12314 32496
rect 8478 32376 8484 32428
rect 8536 32416 8542 32428
rect 8645 32419 8703 32425
rect 8645 32416 8657 32419
rect 8536 32388 8657 32416
rect 8536 32376 8542 32388
rect 8645 32385 8657 32388
rect 8691 32385 8703 32419
rect 8645 32379 8703 32385
rect 8938 32376 8944 32428
rect 8996 32416 9002 32428
rect 8996 32388 9444 32416
rect 8996 32376 9002 32388
rect 7892 32320 8248 32348
rect 7892 32308 7898 32320
rect 8386 32308 8392 32360
rect 8444 32308 8450 32360
rect 6886 32252 6920 32292
rect 6914 32240 6920 32252
rect 6972 32240 6978 32292
rect 7098 32240 7104 32292
rect 7156 32240 7162 32292
rect 9416 32280 9444 32388
rect 9766 32376 9772 32428
rect 9824 32416 9830 32428
rect 9861 32419 9919 32425
rect 9861 32416 9873 32419
rect 9824 32388 9873 32416
rect 9824 32376 9830 32388
rect 9861 32385 9873 32388
rect 9907 32385 9919 32419
rect 9861 32379 9919 32385
rect 11885 32419 11943 32425
rect 11885 32385 11897 32419
rect 11931 32416 11943 32419
rect 11974 32416 11980 32428
rect 11931 32388 11980 32416
rect 11931 32385 11943 32388
rect 11885 32379 11943 32385
rect 11974 32376 11980 32388
rect 12032 32376 12038 32428
rect 13924 32425 13952 32524
rect 14274 32512 14280 32524
rect 14332 32552 14338 32564
rect 15194 32552 15200 32564
rect 14332 32524 15200 32552
rect 14332 32512 14338 32524
rect 15194 32512 15200 32524
rect 15252 32512 15258 32564
rect 16117 32555 16175 32561
rect 16117 32521 16129 32555
rect 16163 32552 16175 32555
rect 16850 32552 16856 32564
rect 16163 32524 16856 32552
rect 16163 32521 16175 32524
rect 16117 32515 16175 32521
rect 16850 32512 16856 32524
rect 16908 32512 16914 32564
rect 17954 32552 17960 32564
rect 17236 32524 17960 32552
rect 15470 32444 15476 32496
rect 15528 32444 15534 32496
rect 16206 32444 16212 32496
rect 16264 32444 16270 32496
rect 13909 32419 13967 32425
rect 13909 32385 13921 32419
rect 13955 32385 13967 32419
rect 13909 32379 13967 32385
rect 14734 32376 14740 32428
rect 14792 32425 14798 32428
rect 14792 32419 14820 32425
rect 14808 32385 14820 32419
rect 15488 32416 15516 32444
rect 15488 32388 16436 32416
rect 14792 32379 14820 32385
rect 14792 32376 14798 32379
rect 9490 32308 9496 32360
rect 9548 32348 9554 32360
rect 10137 32351 10195 32357
rect 10137 32348 10149 32351
rect 9548 32320 10149 32348
rect 9548 32308 9554 32320
rect 10137 32317 10149 32320
rect 10183 32317 10195 32351
rect 10137 32311 10195 32317
rect 12986 32308 12992 32360
rect 13044 32308 13050 32360
rect 13725 32351 13783 32357
rect 13725 32317 13737 32351
rect 13771 32348 13783 32351
rect 13998 32348 14004 32360
rect 13771 32320 14004 32348
rect 13771 32317 13783 32320
rect 13725 32311 13783 32317
rect 13998 32308 14004 32320
rect 14056 32308 14062 32360
rect 14642 32348 14648 32360
rect 14108 32320 14648 32348
rect 13004 32280 13032 32308
rect 14108 32280 14136 32320
rect 14642 32308 14648 32320
rect 14700 32308 14706 32360
rect 14921 32351 14979 32357
rect 14921 32317 14933 32351
rect 14967 32348 14979 32351
rect 16298 32348 16304 32360
rect 14967 32320 16304 32348
rect 14967 32317 14979 32320
rect 14921 32311 14979 32317
rect 16298 32308 16304 32320
rect 16356 32308 16362 32360
rect 16408 32357 16436 32388
rect 16393 32351 16451 32357
rect 16393 32317 16405 32351
rect 16439 32348 16451 32351
rect 16868 32348 16896 32512
rect 17236 32428 17264 32524
rect 17954 32512 17960 32524
rect 18012 32512 18018 32564
rect 18046 32512 18052 32564
rect 18104 32552 18110 32564
rect 19429 32555 19487 32561
rect 19429 32552 19441 32555
rect 18104 32524 19441 32552
rect 18104 32512 18110 32524
rect 19429 32521 19441 32524
rect 19475 32521 19487 32555
rect 19429 32515 19487 32521
rect 21082 32512 21088 32564
rect 21140 32552 21146 32564
rect 22094 32552 22100 32564
rect 21140 32524 22100 32552
rect 21140 32512 21146 32524
rect 22094 32512 22100 32524
rect 22152 32512 22158 32564
rect 22278 32512 22284 32564
rect 22336 32552 22342 32564
rect 22373 32555 22431 32561
rect 22373 32552 22385 32555
rect 22336 32524 22385 32552
rect 22336 32512 22342 32524
rect 22373 32521 22385 32524
rect 22419 32521 22431 32555
rect 22373 32515 22431 32521
rect 22738 32512 22744 32564
rect 22796 32552 22802 32564
rect 22833 32555 22891 32561
rect 22833 32552 22845 32555
rect 22796 32524 22845 32552
rect 22796 32512 22802 32524
rect 22833 32521 22845 32524
rect 22879 32521 22891 32555
rect 22833 32515 22891 32521
rect 24486 32512 24492 32564
rect 24544 32552 24550 32564
rect 26510 32552 26516 32564
rect 24544 32524 26516 32552
rect 24544 32512 24550 32524
rect 18874 32444 18880 32496
rect 18932 32444 18938 32496
rect 19886 32444 19892 32496
rect 19944 32484 19950 32496
rect 23376 32487 23434 32493
rect 19944 32456 22094 32484
rect 19944 32444 19950 32456
rect 17034 32376 17040 32428
rect 17092 32376 17098 32428
rect 17218 32376 17224 32428
rect 17276 32376 17282 32428
rect 17954 32376 17960 32428
rect 18012 32376 18018 32428
rect 19245 32419 19303 32425
rect 19245 32385 19257 32419
rect 19291 32385 19303 32419
rect 19245 32379 19303 32385
rect 19613 32419 19671 32425
rect 19613 32385 19625 32419
rect 19659 32416 19671 32419
rect 19978 32416 19984 32428
rect 19659 32388 19984 32416
rect 19659 32385 19671 32388
rect 19613 32379 19671 32385
rect 18046 32348 18052 32360
rect 18104 32357 18110 32360
rect 18104 32351 18132 32357
rect 16439 32320 16712 32348
rect 16868 32320 18052 32348
rect 16439 32317 16451 32320
rect 16393 32311 16451 32317
rect 9416 32252 11192 32280
rect 13004 32252 14136 32280
rect 14369 32283 14427 32289
rect 4614 32212 4620 32224
rect 4540 32184 4620 32212
rect 1581 32175 1639 32181
rect 4614 32172 4620 32184
rect 4672 32212 4678 32224
rect 8202 32212 8208 32224
rect 4672 32184 8208 32212
rect 4672 32172 4678 32184
rect 8202 32172 8208 32184
rect 8260 32172 8266 32224
rect 8297 32215 8355 32221
rect 8297 32181 8309 32215
rect 8343 32212 8355 32215
rect 8754 32212 8760 32224
rect 8343 32184 8760 32212
rect 8343 32181 8355 32184
rect 8297 32175 8355 32181
rect 8754 32172 8760 32184
rect 8812 32172 8818 32224
rect 9122 32172 9128 32224
rect 9180 32212 9186 32224
rect 9769 32215 9827 32221
rect 9769 32212 9781 32215
rect 9180 32184 9781 32212
rect 9180 32172 9186 32184
rect 9769 32181 9781 32184
rect 9815 32212 9827 32215
rect 11054 32212 11060 32224
rect 9815 32184 11060 32212
rect 9815 32181 9827 32184
rect 9769 32175 9827 32181
rect 11054 32172 11060 32184
rect 11112 32172 11118 32224
rect 11164 32212 11192 32252
rect 14369 32249 14381 32283
rect 14415 32249 14427 32283
rect 16684 32280 16712 32320
rect 18046 32308 18052 32320
rect 18120 32317 18132 32351
rect 18104 32311 18132 32317
rect 18233 32351 18291 32357
rect 18233 32317 18245 32351
rect 18279 32348 18291 32351
rect 18598 32348 18604 32360
rect 18279 32320 18604 32348
rect 18279 32317 18291 32320
rect 18233 32311 18291 32317
rect 18104 32308 18110 32311
rect 18598 32308 18604 32320
rect 18656 32308 18662 32360
rect 14369 32243 14427 32249
rect 15488 32252 16344 32280
rect 16684 32252 16804 32280
rect 12986 32212 12992 32224
rect 11164 32184 12992 32212
rect 12986 32172 12992 32184
rect 13044 32172 13050 32224
rect 13262 32172 13268 32224
rect 13320 32172 13326 32224
rect 14384 32212 14412 32243
rect 15488 32212 15516 32252
rect 14384 32184 15516 32212
rect 15562 32172 15568 32224
rect 15620 32172 15626 32224
rect 15749 32215 15807 32221
rect 15749 32181 15761 32215
rect 15795 32212 15807 32215
rect 16206 32212 16212 32224
rect 15795 32184 16212 32212
rect 15795 32181 15807 32184
rect 15749 32175 15807 32181
rect 16206 32172 16212 32184
rect 16264 32172 16270 32224
rect 16316 32212 16344 32252
rect 16666 32212 16672 32224
rect 16316 32184 16672 32212
rect 16666 32172 16672 32184
rect 16724 32172 16730 32224
rect 16776 32212 16804 32252
rect 16850 32240 16856 32292
rect 16908 32280 16914 32292
rect 17494 32280 17500 32292
rect 16908 32252 17500 32280
rect 16908 32240 16914 32252
rect 17494 32240 17500 32252
rect 17552 32280 17558 32292
rect 17681 32283 17739 32289
rect 17681 32280 17693 32283
rect 17552 32252 17693 32280
rect 17552 32240 17558 32252
rect 17681 32249 17693 32252
rect 17727 32249 17739 32283
rect 19260 32280 19288 32379
rect 19978 32376 19984 32388
rect 20036 32376 20042 32428
rect 22066 32416 22094 32456
rect 23376 32453 23388 32487
rect 23422 32484 23434 32487
rect 24026 32484 24032 32496
rect 23422 32456 24032 32484
rect 23422 32453 23434 32456
rect 23376 32447 23434 32453
rect 24026 32444 24032 32456
rect 24084 32444 24090 32496
rect 24596 32425 24624 32524
rect 26510 32512 26516 32524
rect 26568 32512 26574 32564
rect 27709 32555 27767 32561
rect 27709 32521 27721 32555
rect 27755 32521 27767 32555
rect 27709 32515 27767 32521
rect 27724 32484 27752 32515
rect 28230 32487 28288 32493
rect 28230 32484 28242 32487
rect 27724 32456 28242 32484
rect 28230 32453 28242 32456
rect 28276 32453 28288 32487
rect 28230 32447 28288 32453
rect 22465 32419 22523 32425
rect 22465 32416 22477 32419
rect 22066 32388 22477 32416
rect 22465 32385 22477 32388
rect 22511 32385 22523 32419
rect 23017 32419 23075 32425
rect 23017 32416 23029 32419
rect 22465 32379 22523 32385
rect 22572 32388 23029 32416
rect 22005 32283 22063 32289
rect 19260 32252 21312 32280
rect 17681 32243 17739 32249
rect 19797 32215 19855 32221
rect 19797 32212 19809 32215
rect 16776 32184 19809 32212
rect 19797 32181 19809 32184
rect 19843 32181 19855 32215
rect 21284 32212 21312 32252
rect 22005 32249 22017 32283
rect 22051 32280 22063 32283
rect 22572 32280 22600 32388
rect 23017 32385 23029 32388
rect 23063 32385 23075 32419
rect 23017 32379 23075 32385
rect 24581 32419 24639 32425
rect 24581 32385 24593 32419
rect 24627 32385 24639 32419
rect 24581 32379 24639 32385
rect 24762 32376 24768 32428
rect 24820 32376 24826 32428
rect 25590 32376 25596 32428
rect 25648 32425 25654 32428
rect 25648 32419 25676 32425
rect 25664 32385 25676 32419
rect 25648 32379 25676 32385
rect 27893 32419 27951 32425
rect 27893 32385 27905 32419
rect 27939 32416 27951 32419
rect 28534 32416 28540 32428
rect 27939 32388 28540 32416
rect 27939 32385 27951 32388
rect 27893 32379 27951 32385
rect 25648 32376 25654 32379
rect 28534 32376 28540 32388
rect 28592 32376 28598 32428
rect 22649 32351 22707 32357
rect 22649 32317 22661 32351
rect 22695 32348 22707 32351
rect 22695 32320 22784 32348
rect 22695 32317 22707 32320
rect 22649 32311 22707 32317
rect 22051 32252 22600 32280
rect 22051 32249 22063 32252
rect 22005 32243 22063 32249
rect 22756 32212 22784 32320
rect 22830 32308 22836 32360
rect 22888 32348 22894 32360
rect 23109 32351 23167 32357
rect 23109 32348 23121 32351
rect 22888 32320 23121 32348
rect 22888 32308 22894 32320
rect 23109 32317 23121 32320
rect 23155 32317 23167 32351
rect 23109 32311 23167 32317
rect 25498 32308 25504 32360
rect 25556 32308 25562 32360
rect 25774 32308 25780 32360
rect 25832 32308 25838 32360
rect 26878 32308 26884 32360
rect 26936 32348 26942 32360
rect 27985 32351 28043 32357
rect 27985 32348 27997 32351
rect 26936 32320 27997 32348
rect 26936 32308 26942 32320
rect 27985 32317 27997 32320
rect 28031 32317 28043 32351
rect 27985 32311 28043 32317
rect 24394 32240 24400 32292
rect 24452 32280 24458 32292
rect 24489 32283 24547 32289
rect 24489 32280 24501 32283
rect 24452 32252 24501 32280
rect 24452 32240 24458 32252
rect 24489 32249 24501 32252
rect 24535 32249 24547 32283
rect 24489 32243 24547 32249
rect 25222 32240 25228 32292
rect 25280 32240 25286 32292
rect 27614 32280 27620 32292
rect 26206 32252 27620 32280
rect 26206 32212 26234 32252
rect 27614 32240 27620 32252
rect 27672 32240 27678 32292
rect 21284 32184 26234 32212
rect 26421 32215 26479 32221
rect 19797 32175 19855 32181
rect 26421 32181 26433 32215
rect 26467 32212 26479 32215
rect 27246 32212 27252 32224
rect 26467 32184 27252 32212
rect 26467 32181 26479 32184
rect 26421 32175 26479 32181
rect 27246 32172 27252 32184
rect 27304 32172 27310 32224
rect 28000 32212 28028 32311
rect 29270 32212 29276 32224
rect 28000 32184 29276 32212
rect 29270 32172 29276 32184
rect 29328 32172 29334 32224
rect 29362 32172 29368 32224
rect 29420 32172 29426 32224
rect 1104 32122 36800 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 36800 32122
rect 1104 32048 36800 32070
rect 6638 31968 6644 32020
rect 6696 32008 6702 32020
rect 7834 32008 7840 32020
rect 6696 31980 7840 32008
rect 6696 31968 6702 31980
rect 7834 31968 7840 31980
rect 7892 31968 7898 32020
rect 8389 32011 8447 32017
rect 8389 31977 8401 32011
rect 8435 32008 8447 32011
rect 8478 32008 8484 32020
rect 8435 31980 8484 32008
rect 8435 31977 8447 31980
rect 8389 31971 8447 31977
rect 8478 31968 8484 31980
rect 8536 31968 8542 32020
rect 8588 31980 11652 32008
rect 7098 31940 7104 31952
rect 7024 31912 7104 31940
rect 4525 31875 4583 31881
rect 4525 31841 4537 31875
rect 4571 31872 4583 31875
rect 4614 31872 4620 31884
rect 4571 31844 4620 31872
rect 4571 31841 4583 31844
rect 4525 31835 4583 31841
rect 4614 31832 4620 31844
rect 4672 31832 4678 31884
rect 6089 31875 6147 31881
rect 6089 31841 6101 31875
rect 6135 31872 6147 31875
rect 7024 31872 7052 31912
rect 7098 31900 7104 31912
rect 7156 31940 7162 31952
rect 8588 31940 8616 31980
rect 7156 31912 8616 31940
rect 7156 31900 7162 31912
rect 9306 31900 9312 31952
rect 9364 31900 9370 31952
rect 10704 31949 10732 31980
rect 10689 31943 10747 31949
rect 10689 31909 10701 31943
rect 10735 31909 10747 31943
rect 11624 31940 11652 31980
rect 11790 31968 11796 32020
rect 11848 32008 11854 32020
rect 11885 32011 11943 32017
rect 11885 32008 11897 32011
rect 11848 31980 11897 32008
rect 11848 31968 11854 31980
rect 11885 31977 11897 31980
rect 11931 31977 11943 32011
rect 11885 31971 11943 31977
rect 12434 31968 12440 32020
rect 12492 31968 12498 32020
rect 13262 31968 13268 32020
rect 13320 32008 13326 32020
rect 14734 32008 14740 32020
rect 13320 31980 14740 32008
rect 13320 31968 13326 31980
rect 14734 31968 14740 31980
rect 14792 31968 14798 32020
rect 22646 32008 22652 32020
rect 14844 31980 22652 32008
rect 14844 31940 14872 31980
rect 22646 31968 22652 31980
rect 22704 32008 22710 32020
rect 23934 32008 23940 32020
rect 22704 31980 23940 32008
rect 22704 31968 22710 31980
rect 23934 31968 23940 31980
rect 23992 31968 23998 32020
rect 26206 31980 28028 32008
rect 11624 31912 14872 31940
rect 10689 31903 10747 31909
rect 15746 31900 15752 31952
rect 15804 31940 15810 31952
rect 15933 31943 15991 31949
rect 15933 31940 15945 31943
rect 15804 31912 15945 31940
rect 15804 31900 15810 31912
rect 15933 31909 15945 31912
rect 15979 31909 15991 31943
rect 15933 31903 15991 31909
rect 17681 31943 17739 31949
rect 17681 31909 17693 31943
rect 17727 31940 17739 31943
rect 17770 31940 17776 31952
rect 17727 31912 17776 31940
rect 17727 31909 17739 31912
rect 17681 31903 17739 31909
rect 17770 31900 17776 31912
rect 17828 31900 17834 31952
rect 18708 31912 19012 31940
rect 6135 31844 7052 31872
rect 6135 31841 6147 31844
rect 6089 31835 6147 31841
rect 7190 31832 7196 31884
rect 7248 31872 7254 31884
rect 7374 31872 7380 31884
rect 7248 31844 7380 31872
rect 7248 31832 7254 31844
rect 7374 31832 7380 31844
rect 7432 31832 7438 31884
rect 9033 31875 9091 31881
rect 9033 31872 9045 31875
rect 8404 31844 9045 31872
rect 5350 31764 5356 31816
rect 5408 31804 5414 31816
rect 5445 31807 5503 31813
rect 5445 31804 5457 31807
rect 5408 31776 5457 31804
rect 5408 31764 5414 31776
rect 5445 31773 5457 31776
rect 5491 31773 5503 31807
rect 5445 31767 5503 31773
rect 5629 31807 5687 31813
rect 5629 31773 5641 31807
rect 5675 31773 5687 31807
rect 5629 31767 5687 31773
rect 2774 31696 2780 31748
rect 2832 31736 2838 31748
rect 4341 31739 4399 31745
rect 4341 31736 4353 31739
rect 2832 31708 4353 31736
rect 2832 31696 2838 31708
rect 4341 31705 4353 31708
rect 4387 31705 4399 31739
rect 4341 31699 4399 31705
rect 5644 31680 5672 31767
rect 6362 31764 6368 31816
rect 6420 31764 6426 31816
rect 6454 31764 6460 31816
rect 6512 31813 6518 31816
rect 6512 31807 6540 31813
rect 6528 31773 6540 31807
rect 6512 31767 6540 31773
rect 6512 31764 6518 31767
rect 6638 31764 6644 31816
rect 6696 31764 6702 31816
rect 7285 31807 7343 31813
rect 7285 31773 7297 31807
rect 7331 31804 7343 31807
rect 7466 31804 7472 31816
rect 7331 31776 7472 31804
rect 7331 31773 7343 31776
rect 7285 31767 7343 31773
rect 7466 31764 7472 31776
rect 7524 31764 7530 31816
rect 8404 31813 8432 31844
rect 9033 31841 9045 31844
rect 9079 31841 9091 31875
rect 9861 31875 9919 31881
rect 9861 31872 9873 31875
rect 9033 31835 9091 31841
rect 9324 31844 9873 31872
rect 8389 31807 8447 31813
rect 8389 31773 8401 31807
rect 8435 31773 8447 31807
rect 8389 31767 8447 31773
rect 8665 31807 8723 31813
rect 8665 31773 8677 31807
rect 8711 31804 8723 31807
rect 8938 31804 8944 31816
rect 8711 31776 8944 31804
rect 8711 31773 8723 31776
rect 8665 31767 8723 31773
rect 8938 31764 8944 31776
rect 8996 31764 9002 31816
rect 9122 31764 9128 31816
rect 9180 31764 9186 31816
rect 9324 31813 9352 31844
rect 9861 31841 9873 31844
rect 9907 31841 9919 31875
rect 9861 31835 9919 31841
rect 10042 31832 10048 31884
rect 10100 31832 10106 31884
rect 10962 31832 10968 31884
rect 11020 31832 11026 31884
rect 11054 31832 11060 31884
rect 11112 31881 11118 31884
rect 11112 31875 11140 31881
rect 11128 31841 11140 31875
rect 11112 31835 11140 31841
rect 11112 31832 11118 31835
rect 11238 31832 11244 31884
rect 11296 31872 11302 31884
rect 11296 31844 11836 31872
rect 11296 31832 11302 31844
rect 9309 31807 9367 31813
rect 9309 31773 9321 31807
rect 9355 31773 9367 31807
rect 9309 31767 9367 31773
rect 9585 31807 9643 31813
rect 9585 31773 9597 31807
rect 9631 31804 9643 31807
rect 9674 31804 9680 31816
rect 9631 31776 9680 31804
rect 9631 31773 9643 31776
rect 9585 31767 9643 31773
rect 9674 31764 9680 31776
rect 9732 31804 9738 31816
rect 9769 31807 9827 31813
rect 9769 31804 9781 31807
rect 9732 31776 9781 31804
rect 9732 31764 9738 31776
rect 9769 31773 9781 31776
rect 9815 31773 9827 31807
rect 9769 31767 9827 31773
rect 9953 31807 10011 31813
rect 9953 31773 9965 31807
rect 9999 31773 10011 31807
rect 9953 31767 10011 31773
rect 9968 31736 9996 31767
rect 10226 31764 10232 31816
rect 10284 31764 10290 31816
rect 11808 31804 11836 31844
rect 12894 31832 12900 31884
rect 12952 31832 12958 31884
rect 12986 31832 12992 31884
rect 13044 31872 13050 31884
rect 13044 31844 13308 31872
rect 13044 31832 13050 31844
rect 13170 31804 13176 31816
rect 11808 31776 13176 31804
rect 13170 31764 13176 31776
rect 13228 31764 13234 31816
rect 10244 31736 10272 31764
rect 9968 31708 10272 31736
rect 3418 31628 3424 31680
rect 3476 31668 3482 31680
rect 3881 31671 3939 31677
rect 3881 31668 3893 31671
rect 3476 31640 3893 31668
rect 3476 31628 3482 31640
rect 3881 31637 3893 31640
rect 3927 31637 3939 31671
rect 3881 31631 3939 31637
rect 4249 31671 4307 31677
rect 4249 31637 4261 31671
rect 4295 31668 4307 31671
rect 5534 31668 5540 31680
rect 4295 31640 5540 31668
rect 4295 31637 4307 31640
rect 4249 31631 4307 31637
rect 5534 31628 5540 31640
rect 5592 31628 5598 31680
rect 5626 31628 5632 31680
rect 5684 31628 5690 31680
rect 8570 31628 8576 31680
rect 8628 31668 8634 31680
rect 9493 31671 9551 31677
rect 9493 31668 9505 31671
rect 8628 31640 9505 31668
rect 8628 31628 8634 31640
rect 9493 31637 9505 31640
rect 9539 31637 9551 31671
rect 9493 31631 9551 31637
rect 12805 31671 12863 31677
rect 12805 31637 12817 31671
rect 12851 31668 12863 31671
rect 13170 31668 13176 31680
rect 12851 31640 13176 31668
rect 12851 31637 12863 31640
rect 12805 31631 12863 31637
rect 13170 31628 13176 31640
rect 13228 31628 13234 31680
rect 13280 31668 13308 31844
rect 13998 31832 14004 31884
rect 14056 31872 14062 31884
rect 14093 31875 14151 31881
rect 14093 31872 14105 31875
rect 14056 31844 14105 31872
rect 14056 31832 14062 31844
rect 14093 31841 14105 31844
rect 14139 31841 14151 31875
rect 14093 31835 14151 31841
rect 14274 31832 14280 31884
rect 14332 31832 14338 31884
rect 14734 31832 14740 31884
rect 14792 31832 14798 31884
rect 14826 31832 14832 31884
rect 14884 31872 14890 31884
rect 15130 31875 15188 31881
rect 15130 31872 15142 31875
rect 14884 31844 15142 31872
rect 14884 31832 14890 31844
rect 15130 31841 15142 31844
rect 15176 31841 15188 31875
rect 15130 31835 15188 31841
rect 17034 31832 17040 31884
rect 17092 31832 17098 31884
rect 17218 31832 17224 31884
rect 17276 31832 17282 31884
rect 17954 31832 17960 31884
rect 18012 31832 18018 31884
rect 18046 31832 18052 31884
rect 18104 31881 18110 31884
rect 18104 31875 18132 31881
rect 18120 31841 18132 31875
rect 18708 31872 18736 31912
rect 18104 31835 18132 31841
rect 18248 31844 18736 31872
rect 18104 31832 18110 31835
rect 18248 31816 18276 31844
rect 18782 31832 18788 31884
rect 18840 31872 18846 31884
rect 18877 31875 18935 31881
rect 18877 31872 18889 31875
rect 18840 31844 18889 31872
rect 18840 31832 18846 31844
rect 18877 31841 18889 31844
rect 18923 31841 18935 31875
rect 18984 31872 19012 31912
rect 19150 31900 19156 31952
rect 19208 31940 19214 31952
rect 23474 31940 23480 31952
rect 19208 31912 23480 31940
rect 19208 31900 19214 31912
rect 23474 31900 23480 31912
rect 23532 31900 23538 31952
rect 24302 31900 24308 31952
rect 24360 31940 24366 31952
rect 26206 31940 26234 31980
rect 24360 31912 26234 31940
rect 28000 31940 28028 31980
rect 28534 31968 28540 32020
rect 28592 31968 28598 32020
rect 31846 32008 31852 32020
rect 29288 31980 31852 32008
rect 29288 31940 29316 31980
rect 31846 31968 31852 31980
rect 31904 31968 31910 32020
rect 28000 31912 29316 31940
rect 24360 31900 24366 31912
rect 25774 31872 25780 31884
rect 18984 31844 25780 31872
rect 18877 31835 18935 31841
rect 25774 31832 25780 31844
rect 25832 31832 25838 31884
rect 28626 31832 28632 31884
rect 28684 31872 28690 31884
rect 29181 31875 29239 31881
rect 28684 31844 29132 31872
rect 28684 31832 28690 31844
rect 15010 31764 15016 31816
rect 15068 31764 15074 31816
rect 15286 31764 15292 31816
rect 15344 31764 15350 31816
rect 16022 31764 16028 31816
rect 16080 31764 16086 31816
rect 16206 31764 16212 31816
rect 16264 31764 16270 31816
rect 16298 31764 16304 31816
rect 16356 31804 16362 31816
rect 16356 31776 16574 31804
rect 16356 31764 16362 31776
rect 15102 31668 15108 31680
rect 13280 31640 15108 31668
rect 15102 31628 15108 31640
rect 15160 31628 15166 31680
rect 16040 31677 16068 31764
rect 16025 31671 16083 31677
rect 16025 31637 16037 31671
rect 16071 31637 16083 31671
rect 16546 31668 16574 31776
rect 18230 31764 18236 31816
rect 18288 31764 18294 31816
rect 26878 31764 26884 31816
rect 26936 31804 26942 31816
rect 27065 31807 27123 31813
rect 27065 31804 27077 31807
rect 26936 31776 27077 31804
rect 26936 31764 26942 31776
rect 27065 31773 27077 31776
rect 27111 31773 27123 31807
rect 27065 31767 27123 31773
rect 28074 31764 28080 31816
rect 28132 31804 28138 31816
rect 28997 31807 29055 31813
rect 28997 31804 29009 31807
rect 28132 31776 29009 31804
rect 28132 31764 28138 31776
rect 28997 31773 29009 31776
rect 29043 31773 29055 31807
rect 29104 31804 29132 31844
rect 29181 31841 29193 31875
rect 29227 31872 29239 31875
rect 29288 31872 29316 31912
rect 30745 31943 30803 31949
rect 30745 31909 30757 31943
rect 30791 31940 30803 31943
rect 31938 31940 31944 31952
rect 30791 31912 31944 31940
rect 30791 31909 30803 31912
rect 30745 31903 30803 31909
rect 31938 31900 31944 31912
rect 31996 31900 32002 31952
rect 31389 31875 31447 31881
rect 31389 31872 31401 31875
rect 29227 31844 29316 31872
rect 29380 31844 31401 31872
rect 29227 31841 29239 31844
rect 29181 31835 29239 31841
rect 29380 31804 29408 31844
rect 31389 31841 31401 31844
rect 31435 31872 31447 31875
rect 32582 31872 32588 31884
rect 31435 31844 32588 31872
rect 31435 31841 31447 31844
rect 31389 31835 31447 31841
rect 32582 31832 32588 31844
rect 32640 31832 32646 31884
rect 29104 31776 29408 31804
rect 28997 31767 29055 31773
rect 29822 31764 29828 31816
rect 29880 31764 29886 31816
rect 31202 31764 31208 31816
rect 31260 31764 31266 31816
rect 27338 31745 27344 31748
rect 27332 31699 27344 31745
rect 27338 31696 27344 31699
rect 27396 31696 27402 31748
rect 28905 31739 28963 31745
rect 28905 31705 28917 31739
rect 28951 31736 28963 31739
rect 29362 31736 29368 31748
rect 28951 31708 29368 31736
rect 28951 31705 28963 31708
rect 28905 31699 28963 31705
rect 29362 31696 29368 31708
rect 29420 31696 29426 31748
rect 18506 31668 18512 31680
rect 16546 31640 18512 31668
rect 16025 31631 16083 31637
rect 18506 31628 18512 31640
rect 18564 31628 18570 31680
rect 27890 31628 27896 31680
rect 27948 31668 27954 31680
rect 28445 31671 28503 31677
rect 28445 31668 28457 31671
rect 27948 31640 28457 31668
rect 27948 31628 27954 31640
rect 28445 31637 28457 31640
rect 28491 31637 28503 31671
rect 28445 31631 28503 31637
rect 29638 31628 29644 31680
rect 29696 31628 29702 31680
rect 30006 31628 30012 31680
rect 30064 31668 30070 31680
rect 31113 31671 31171 31677
rect 31113 31668 31125 31671
rect 30064 31640 31125 31668
rect 30064 31628 30070 31640
rect 31113 31637 31125 31640
rect 31159 31637 31171 31671
rect 31113 31631 31171 31637
rect 1104 31578 36800 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 36800 31578
rect 1104 31504 36800 31526
rect 3237 31467 3295 31473
rect 3237 31433 3249 31467
rect 3283 31433 3295 31467
rect 3237 31427 3295 31433
rect 1762 31396 1768 31408
rect 1596 31368 1768 31396
rect 1596 31337 1624 31368
rect 1762 31356 1768 31368
rect 1820 31396 1826 31408
rect 3252 31396 3280 31427
rect 10226 31424 10232 31476
rect 10284 31464 10290 31476
rect 10689 31467 10747 31473
rect 10689 31464 10701 31467
rect 10284 31436 10701 31464
rect 10284 31424 10290 31436
rect 10689 31433 10701 31436
rect 10735 31433 10747 31467
rect 10689 31427 10747 31433
rect 23474 31424 23480 31476
rect 23532 31464 23538 31476
rect 24489 31467 24547 31473
rect 24489 31464 24501 31467
rect 23532 31436 24501 31464
rect 23532 31424 23538 31436
rect 24489 31433 24501 31436
rect 24535 31433 24547 31467
rect 27249 31467 27307 31473
rect 24489 31427 24547 31433
rect 25148 31436 26648 31464
rect 3758 31399 3816 31405
rect 3758 31396 3770 31399
rect 1820 31368 1992 31396
rect 3252 31368 3770 31396
rect 1820 31356 1826 31368
rect 1854 31337 1860 31340
rect 1581 31331 1639 31337
rect 1581 31297 1593 31331
rect 1627 31297 1639 31331
rect 1581 31291 1639 31297
rect 1848 31291 1860 31337
rect 1854 31288 1860 31291
rect 1912 31288 1918 31340
rect 1964 31328 1992 31368
rect 3758 31365 3770 31368
rect 3804 31365 3816 31399
rect 3758 31359 3816 31365
rect 7282 31356 7288 31408
rect 7340 31396 7346 31408
rect 7340 31368 7512 31396
rect 7340 31356 7346 31368
rect 1964 31300 2774 31328
rect 2746 31260 2774 31300
rect 3418 31288 3424 31340
rect 3476 31288 3482 31340
rect 7374 31288 7380 31340
rect 7432 31288 7438 31340
rect 7484 31337 7512 31368
rect 9306 31356 9312 31408
rect 9364 31396 9370 31408
rect 9554 31399 9612 31405
rect 9554 31396 9566 31399
rect 9364 31368 9566 31396
rect 9364 31356 9370 31368
rect 9554 31365 9566 31368
rect 9600 31365 9612 31399
rect 9554 31359 9612 31365
rect 7469 31331 7527 31337
rect 7469 31297 7481 31331
rect 7515 31328 7527 31331
rect 7650 31328 7656 31340
rect 7515 31300 7656 31328
rect 7515 31297 7527 31300
rect 7469 31291 7527 31297
rect 7650 31288 7656 31300
rect 7708 31288 7714 31340
rect 9398 31328 9404 31340
rect 9324 31300 9404 31328
rect 3510 31260 3516 31272
rect 2746 31232 3516 31260
rect 3510 31220 3516 31232
rect 3568 31220 3574 31272
rect 7558 31220 7564 31272
rect 7616 31220 7622 31272
rect 8386 31220 8392 31272
rect 8444 31260 8450 31272
rect 9324 31269 9352 31300
rect 9398 31288 9404 31300
rect 9456 31288 9462 31340
rect 19886 31288 19892 31340
rect 19944 31288 19950 31340
rect 23109 31331 23167 31337
rect 23109 31297 23121 31331
rect 23155 31328 23167 31331
rect 23842 31328 23848 31340
rect 23155 31300 23848 31328
rect 23155 31297 23167 31300
rect 23109 31291 23167 31297
rect 23842 31288 23848 31300
rect 23900 31288 23906 31340
rect 24305 31331 24363 31337
rect 24305 31297 24317 31331
rect 24351 31328 24363 31331
rect 24762 31328 24768 31340
rect 24351 31300 24768 31328
rect 24351 31297 24363 31300
rect 24305 31291 24363 31297
rect 24762 31288 24768 31300
rect 24820 31288 24826 31340
rect 25148 31337 25176 31436
rect 26620 31396 26648 31436
rect 27249 31433 27261 31467
rect 27295 31464 27307 31467
rect 27338 31464 27344 31476
rect 27295 31436 27344 31464
rect 27295 31433 27307 31436
rect 27249 31427 27307 31433
rect 27338 31424 27344 31436
rect 27396 31424 27402 31476
rect 27890 31424 27896 31476
rect 27948 31424 27954 31476
rect 27908 31396 27936 31424
rect 26620 31368 27936 31396
rect 27985 31399 28043 31405
rect 27985 31365 27997 31399
rect 28031 31396 28043 31399
rect 28074 31396 28080 31408
rect 28031 31368 28080 31396
rect 28031 31365 28043 31368
rect 27985 31359 28043 31365
rect 28074 31356 28080 31368
rect 28132 31356 28138 31408
rect 29638 31405 29644 31408
rect 29632 31359 29644 31405
rect 29638 31356 29644 31359
rect 29696 31356 29702 31408
rect 25133 31331 25191 31337
rect 25133 31297 25145 31331
rect 25179 31328 25191 31331
rect 25314 31328 25320 31340
rect 25179 31300 25320 31328
rect 25179 31297 25191 31300
rect 25133 31291 25191 31297
rect 25314 31288 25320 31300
rect 25372 31288 25378 31340
rect 26142 31288 26148 31340
rect 26200 31288 26206 31340
rect 27433 31331 27491 31337
rect 27433 31297 27445 31331
rect 27479 31328 27491 31331
rect 27479 31300 27568 31328
rect 27479 31297 27491 31300
rect 27433 31291 27491 31297
rect 9309 31263 9367 31269
rect 9309 31260 9321 31263
rect 8444 31232 9321 31260
rect 8444 31220 8450 31232
rect 9309 31229 9321 31232
rect 9355 31229 9367 31263
rect 9309 31223 9367 31229
rect 24946 31220 24952 31272
rect 25004 31220 25010 31272
rect 26050 31269 26056 31272
rect 25869 31263 25927 31269
rect 25869 31260 25881 31263
rect 25700 31232 25881 31260
rect 4893 31195 4951 31201
rect 4893 31161 4905 31195
rect 4939 31192 4951 31195
rect 5534 31192 5540 31204
rect 4939 31164 5540 31192
rect 4939 31161 4951 31164
rect 4893 31155 4951 31161
rect 5534 31152 5540 31164
rect 5592 31192 5598 31204
rect 6454 31192 6460 31204
rect 5592 31164 6460 31192
rect 5592 31152 5598 31164
rect 6454 31152 6460 31164
rect 6512 31152 6518 31204
rect 23290 31152 23296 31204
rect 23348 31152 23354 31204
rect 23934 31152 23940 31204
rect 23992 31192 23998 31204
rect 24121 31195 24179 31201
rect 24121 31192 24133 31195
rect 23992 31164 24133 31192
rect 23992 31152 23998 31164
rect 24121 31161 24133 31164
rect 24167 31192 24179 31195
rect 25593 31195 25651 31201
rect 25593 31192 25605 31195
rect 24167 31164 25605 31192
rect 24167 31161 24179 31164
rect 24121 31155 24179 31161
rect 25593 31161 25605 31164
rect 25639 31161 25651 31195
rect 25593 31155 25651 31161
rect 2682 31084 2688 31136
rect 2740 31124 2746 31136
rect 2961 31127 3019 31133
rect 2961 31124 2973 31127
rect 2740 31096 2973 31124
rect 2740 31084 2746 31096
rect 2961 31093 2973 31096
rect 3007 31124 3019 31127
rect 5626 31124 5632 31136
rect 3007 31096 5632 31124
rect 3007 31093 3019 31096
rect 2961 31087 3019 31093
rect 5626 31084 5632 31096
rect 5684 31084 5690 31136
rect 7009 31127 7067 31133
rect 7009 31093 7021 31127
rect 7055 31124 7067 31127
rect 8018 31124 8024 31136
rect 7055 31096 8024 31124
rect 7055 31093 7067 31096
rect 7009 31087 7067 31093
rect 8018 31084 8024 31096
rect 8076 31084 8082 31136
rect 19702 31084 19708 31136
rect 19760 31084 19766 31136
rect 25700 31124 25728 31232
rect 25869 31229 25881 31232
rect 25915 31229 25927 31263
rect 25869 31223 25927 31229
rect 26007 31263 26056 31269
rect 26007 31229 26019 31263
rect 26053 31229 26056 31263
rect 26007 31223 26056 31229
rect 26050 31220 26056 31223
rect 26108 31260 26114 31272
rect 26108 31232 27476 31260
rect 26108 31220 26114 31232
rect 26050 31124 26056 31136
rect 25700 31096 26056 31124
rect 26050 31084 26056 31096
rect 26108 31084 26114 31136
rect 26510 31084 26516 31136
rect 26568 31124 26574 31136
rect 26789 31127 26847 31133
rect 26789 31124 26801 31127
rect 26568 31096 26801 31124
rect 26568 31084 26574 31096
rect 26789 31093 26801 31096
rect 26835 31093 26847 31127
rect 27448 31124 27476 31232
rect 27540 31201 27568 31300
rect 29270 31288 29276 31340
rect 29328 31328 29334 31340
rect 29365 31331 29423 31337
rect 29365 31328 29377 31331
rect 29328 31300 29377 31328
rect 29328 31288 29334 31300
rect 29365 31297 29377 31300
rect 29411 31328 29423 31331
rect 30190 31328 30196 31340
rect 29411 31300 30196 31328
rect 29411 31297 29423 31300
rect 29365 31291 29423 31297
rect 30190 31288 30196 31300
rect 30248 31328 30254 31340
rect 31113 31331 31171 31337
rect 31113 31328 31125 31331
rect 30248 31300 31125 31328
rect 30248 31288 30254 31300
rect 31113 31297 31125 31300
rect 31159 31297 31171 31331
rect 31113 31291 31171 31297
rect 31938 31288 31944 31340
rect 31996 31288 32002 31340
rect 28166 31220 28172 31272
rect 28224 31260 28230 31272
rect 28534 31260 28540 31272
rect 28224 31232 28540 31260
rect 28224 31220 28230 31232
rect 28534 31220 28540 31232
rect 28592 31220 28598 31272
rect 30558 31220 30564 31272
rect 30616 31260 30622 31272
rect 30837 31263 30895 31269
rect 30837 31260 30849 31263
rect 30616 31232 30849 31260
rect 30616 31220 30622 31232
rect 30837 31229 30849 31232
rect 30883 31229 30895 31263
rect 30837 31223 30895 31229
rect 27525 31195 27583 31201
rect 27525 31161 27537 31195
rect 27571 31161 27583 31195
rect 27525 31155 27583 31161
rect 29362 31124 29368 31136
rect 27448 31096 29368 31124
rect 26789 31087 26847 31093
rect 29362 31084 29368 31096
rect 29420 31084 29426 31136
rect 30742 31084 30748 31136
rect 30800 31084 30806 31136
rect 31754 31084 31760 31136
rect 31812 31084 31818 31136
rect 1104 31034 36800 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 36800 31034
rect 1104 30960 36800 30982
rect 1854 30880 1860 30932
rect 1912 30920 1918 30932
rect 1949 30923 2007 30929
rect 1949 30920 1961 30923
rect 1912 30892 1961 30920
rect 1912 30880 1918 30892
rect 1949 30889 1961 30892
rect 1995 30889 2007 30923
rect 1949 30883 2007 30889
rect 7374 30880 7380 30932
rect 7432 30920 7438 30932
rect 8573 30923 8631 30929
rect 8573 30920 8585 30923
rect 7432 30892 8585 30920
rect 7432 30880 7438 30892
rect 8573 30889 8585 30892
rect 8619 30889 8631 30923
rect 8573 30883 8631 30889
rect 26050 30880 26056 30932
rect 26108 30920 26114 30932
rect 29733 30923 29791 30929
rect 26108 30892 26740 30920
rect 26108 30880 26114 30892
rect 2317 30855 2375 30861
rect 2317 30821 2329 30855
rect 2363 30821 2375 30855
rect 2317 30815 2375 30821
rect 2133 30719 2191 30725
rect 2133 30685 2145 30719
rect 2179 30716 2191 30719
rect 2332 30716 2360 30815
rect 25222 30812 25228 30864
rect 25280 30852 25286 30864
rect 26712 30852 26740 30892
rect 29733 30889 29745 30923
rect 29779 30920 29791 30923
rect 29822 30920 29828 30932
rect 29779 30892 29828 30920
rect 29779 30889 29791 30892
rect 29733 30883 29791 30889
rect 29822 30880 29828 30892
rect 29880 30880 29886 30932
rect 30742 30852 30748 30864
rect 25280 30824 25820 30852
rect 26712 30824 30748 30852
rect 25280 30812 25286 30824
rect 25792 30796 25820 30824
rect 2590 30744 2596 30796
rect 2648 30784 2654 30796
rect 2869 30787 2927 30793
rect 2869 30784 2881 30787
rect 2648 30756 2881 30784
rect 2648 30744 2654 30756
rect 2869 30753 2881 30756
rect 2915 30753 2927 30787
rect 2869 30747 2927 30753
rect 5261 30787 5319 30793
rect 5261 30753 5273 30787
rect 5307 30784 5319 30787
rect 5350 30784 5356 30796
rect 5307 30756 5356 30784
rect 5307 30753 5319 30756
rect 5261 30747 5319 30753
rect 5350 30744 5356 30756
rect 5408 30744 5414 30796
rect 5445 30787 5503 30793
rect 5445 30753 5457 30787
rect 5491 30784 5503 30787
rect 5626 30784 5632 30796
rect 5491 30756 5632 30784
rect 5491 30753 5503 30756
rect 5445 30747 5503 30753
rect 5626 30744 5632 30756
rect 5684 30744 5690 30796
rect 5810 30744 5816 30796
rect 5868 30784 5874 30796
rect 5905 30787 5963 30793
rect 5905 30784 5917 30787
rect 5868 30756 5917 30784
rect 5868 30744 5874 30756
rect 5905 30753 5917 30756
rect 5951 30753 5963 30787
rect 5905 30747 5963 30753
rect 6178 30744 6184 30796
rect 6236 30744 6242 30796
rect 6362 30793 6368 30796
rect 6319 30787 6368 30793
rect 6319 30753 6331 30787
rect 6365 30753 6368 30787
rect 6319 30747 6368 30753
rect 6362 30744 6368 30747
rect 6420 30744 6426 30796
rect 6457 30787 6515 30793
rect 6457 30753 6469 30787
rect 6503 30784 6515 30787
rect 6638 30784 6644 30796
rect 6503 30756 6644 30784
rect 6503 30753 6515 30756
rect 6457 30747 6515 30753
rect 6638 30744 6644 30756
rect 6696 30784 6702 30796
rect 21269 30787 21327 30793
rect 21269 30784 21281 30787
rect 6696 30756 7328 30784
rect 6696 30744 6702 30756
rect 2179 30688 2360 30716
rect 2179 30685 2191 30688
rect 2133 30679 2191 30685
rect 2682 30676 2688 30728
rect 2740 30676 2746 30728
rect 2774 30676 2780 30728
rect 2832 30676 2838 30728
rect 5169 30719 5227 30725
rect 5169 30685 5181 30719
rect 5215 30685 5227 30719
rect 5169 30679 5227 30685
rect 5184 30648 5212 30679
rect 7190 30676 7196 30728
rect 7248 30676 7254 30728
rect 7300 30716 7328 30756
rect 20456 30756 21281 30784
rect 11330 30716 11336 30728
rect 7300 30688 11336 30716
rect 11330 30676 11336 30688
rect 11388 30676 11394 30728
rect 11977 30719 12035 30725
rect 11977 30685 11989 30719
rect 12023 30716 12035 30719
rect 12066 30716 12072 30728
rect 12023 30688 12072 30716
rect 12023 30685 12035 30688
rect 11977 30679 12035 30685
rect 12066 30676 12072 30688
rect 12124 30676 12130 30728
rect 14274 30676 14280 30728
rect 14332 30676 14338 30728
rect 15470 30676 15476 30728
rect 15528 30716 15534 30728
rect 17313 30719 17371 30725
rect 17313 30716 17325 30719
rect 15528 30688 17325 30716
rect 15528 30676 15534 30688
rect 17313 30685 17325 30688
rect 17359 30685 17371 30719
rect 17313 30679 17371 30685
rect 19426 30676 19432 30728
rect 19484 30676 19490 30728
rect 19702 30725 19708 30728
rect 19696 30716 19708 30725
rect 19663 30688 19708 30716
rect 19696 30679 19708 30688
rect 19702 30676 19708 30679
rect 19760 30676 19766 30728
rect 20456 30716 20484 30756
rect 21269 30753 21281 30756
rect 21315 30753 21327 30787
rect 21269 30747 21327 30753
rect 20272 30688 20484 30716
rect 5258 30648 5264 30660
rect 5184 30620 5264 30648
rect 5258 30608 5264 30620
rect 5316 30608 5322 30660
rect 7460 30651 7518 30657
rect 7460 30617 7472 30651
rect 7506 30648 7518 30651
rect 7834 30648 7840 30660
rect 7506 30620 7840 30648
rect 7506 30617 7518 30620
rect 7460 30611 7518 30617
rect 7834 30608 7840 30620
rect 7892 30608 7898 30660
rect 12244 30651 12302 30657
rect 12244 30617 12256 30651
rect 12290 30648 12302 30651
rect 12342 30648 12348 30660
rect 12290 30620 12348 30648
rect 12290 30617 12302 30620
rect 12244 30611 12302 30617
rect 12342 30608 12348 30620
rect 12400 30608 12406 30660
rect 19444 30648 19472 30676
rect 20272 30648 20300 30688
rect 21174 30676 21180 30728
rect 21232 30676 21238 30728
rect 21284 30716 21312 30747
rect 25314 30744 25320 30796
rect 25372 30744 25378 30796
rect 25774 30744 25780 30796
rect 25832 30744 25838 30796
rect 25866 30744 25872 30796
rect 25924 30784 25930 30796
rect 30208 30793 30236 30824
rect 30742 30812 30748 30824
rect 30800 30812 30806 30864
rect 26329 30787 26387 30793
rect 26329 30784 26341 30787
rect 25924 30756 26341 30784
rect 25924 30744 25930 30756
rect 26329 30753 26341 30756
rect 26375 30753 26387 30787
rect 26329 30747 26387 30753
rect 30193 30787 30251 30793
rect 30193 30753 30205 30787
rect 30239 30753 30251 30787
rect 30193 30747 30251 30753
rect 30282 30744 30288 30796
rect 30340 30744 30346 30796
rect 22646 30716 22652 30728
rect 21284 30688 22652 30716
rect 22646 30676 22652 30688
rect 22704 30716 22710 30728
rect 22833 30719 22891 30725
rect 22833 30716 22845 30719
rect 22704 30688 22845 30716
rect 22704 30676 22710 30688
rect 22833 30685 22845 30688
rect 22879 30685 22891 30719
rect 22833 30679 22891 30685
rect 24578 30676 24584 30728
rect 24636 30676 24642 30728
rect 24946 30676 24952 30728
rect 25004 30716 25010 30728
rect 25130 30716 25136 30728
rect 25004 30688 25136 30716
rect 25004 30676 25010 30688
rect 25130 30676 25136 30688
rect 25188 30676 25194 30728
rect 26050 30676 26056 30728
rect 26108 30676 26114 30728
rect 26142 30676 26148 30728
rect 26200 30725 26206 30728
rect 26200 30719 26228 30725
rect 26216 30685 26228 30719
rect 26200 30679 26228 30685
rect 26200 30676 26206 30679
rect 21514 30651 21572 30657
rect 21514 30648 21526 30651
rect 19444 30620 20300 30648
rect 21008 30620 21526 30648
rect 4798 30540 4804 30592
rect 4856 30580 4862 30592
rect 4985 30583 5043 30589
rect 4985 30580 4997 30583
rect 4856 30552 4997 30580
rect 4856 30540 4862 30552
rect 4985 30549 4997 30552
rect 5031 30549 5043 30583
rect 4985 30543 5043 30549
rect 7098 30540 7104 30592
rect 7156 30540 7162 30592
rect 13354 30540 13360 30592
rect 13412 30540 13418 30592
rect 14090 30540 14096 30592
rect 14148 30540 14154 30592
rect 17218 30540 17224 30592
rect 17276 30580 17282 30592
rect 17405 30583 17463 30589
rect 17405 30580 17417 30583
rect 17276 30552 17417 30580
rect 17276 30540 17282 30552
rect 17405 30549 17417 30552
rect 17451 30549 17463 30583
rect 17405 30543 17463 30549
rect 20714 30540 20720 30592
rect 20772 30580 20778 30592
rect 21008 30589 21036 30620
rect 21514 30617 21526 30620
rect 21560 30617 21572 30651
rect 21514 30611 21572 30617
rect 23100 30651 23158 30657
rect 23100 30617 23112 30651
rect 23146 30648 23158 30651
rect 30300 30648 30328 30744
rect 30374 30676 30380 30728
rect 30432 30716 30438 30728
rect 30745 30719 30803 30725
rect 30745 30716 30757 30719
rect 30432 30688 30757 30716
rect 30432 30676 30438 30688
rect 30745 30685 30757 30688
rect 30791 30685 30803 30719
rect 30745 30679 30803 30685
rect 31012 30719 31070 30725
rect 31012 30685 31024 30719
rect 31058 30716 31070 30719
rect 31754 30716 31760 30728
rect 31058 30688 31760 30716
rect 31058 30685 31070 30688
rect 31012 30679 31070 30685
rect 31754 30676 31760 30688
rect 31812 30676 31818 30728
rect 32398 30648 32404 30660
rect 23146 30620 24440 30648
rect 30300 30620 32404 30648
rect 23146 30617 23158 30620
rect 23100 30611 23158 30617
rect 20809 30583 20867 30589
rect 20809 30580 20821 30583
rect 20772 30552 20821 30580
rect 20772 30540 20778 30552
rect 20809 30549 20821 30552
rect 20855 30549 20867 30583
rect 20809 30543 20867 30549
rect 20993 30583 21051 30589
rect 20993 30549 21005 30583
rect 21039 30549 21051 30583
rect 20993 30543 21051 30549
rect 22186 30540 22192 30592
rect 22244 30580 22250 30592
rect 22649 30583 22707 30589
rect 22649 30580 22661 30583
rect 22244 30552 22661 30580
rect 22244 30540 22250 30552
rect 22649 30549 22661 30552
rect 22695 30549 22707 30583
rect 22649 30543 22707 30549
rect 24210 30540 24216 30592
rect 24268 30540 24274 30592
rect 24412 30589 24440 30620
rect 32398 30608 32404 30620
rect 32456 30608 32462 30660
rect 24397 30583 24455 30589
rect 24397 30549 24409 30583
rect 24443 30549 24455 30583
rect 24397 30543 24455 30549
rect 25774 30540 25780 30592
rect 25832 30580 25838 30592
rect 26234 30580 26240 30592
rect 25832 30552 26240 30580
rect 25832 30540 25838 30552
rect 26234 30540 26240 30552
rect 26292 30540 26298 30592
rect 26602 30540 26608 30592
rect 26660 30580 26666 30592
rect 26973 30583 27031 30589
rect 26973 30580 26985 30583
rect 26660 30552 26985 30580
rect 26660 30540 26666 30552
rect 26973 30549 26985 30552
rect 27019 30549 27031 30583
rect 26973 30543 27031 30549
rect 29822 30540 29828 30592
rect 29880 30580 29886 30592
rect 30006 30580 30012 30592
rect 29880 30552 30012 30580
rect 29880 30540 29886 30552
rect 30006 30540 30012 30552
rect 30064 30580 30070 30592
rect 30101 30583 30159 30589
rect 30101 30580 30113 30583
rect 30064 30552 30113 30580
rect 30064 30540 30070 30552
rect 30101 30549 30113 30552
rect 30147 30549 30159 30583
rect 30101 30543 30159 30549
rect 31202 30540 31208 30592
rect 31260 30580 31266 30592
rect 32125 30583 32183 30589
rect 32125 30580 32137 30583
rect 31260 30552 32137 30580
rect 31260 30540 31266 30552
rect 32125 30549 32137 30552
rect 32171 30549 32183 30583
rect 32125 30543 32183 30549
rect 1104 30490 36800 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 36800 30490
rect 1104 30416 36800 30438
rect 4724 30348 5028 30376
rect 3510 30200 3516 30252
rect 3568 30240 3574 30252
rect 4617 30243 4675 30249
rect 4617 30240 4629 30243
rect 3568 30212 4629 30240
rect 3568 30200 3574 30212
rect 4617 30209 4629 30212
rect 4663 30240 4675 30243
rect 4724 30240 4752 30348
rect 4798 30268 4804 30320
rect 4856 30308 4862 30320
rect 5000 30308 5028 30348
rect 7834 30336 7840 30388
rect 7892 30336 7898 30388
rect 11330 30336 11336 30388
rect 11388 30376 11394 30388
rect 11882 30376 11888 30388
rect 11388 30348 11888 30376
rect 11388 30336 11394 30348
rect 11882 30336 11888 30348
rect 11940 30336 11946 30388
rect 12342 30336 12348 30388
rect 12400 30336 12406 30388
rect 13081 30379 13139 30385
rect 13081 30345 13093 30379
rect 13127 30376 13139 30379
rect 13354 30376 13360 30388
rect 13127 30348 13360 30376
rect 13127 30345 13139 30348
rect 13081 30339 13139 30345
rect 13354 30336 13360 30348
rect 13412 30336 13418 30388
rect 16945 30379 17003 30385
rect 16945 30345 16957 30379
rect 16991 30345 17003 30379
rect 16945 30339 17003 30345
rect 7190 30308 7196 30320
rect 4856 30280 4936 30308
rect 5000 30280 7196 30308
rect 4856 30268 4862 30280
rect 4908 30249 4936 30280
rect 7190 30268 7196 30280
rect 7248 30268 7254 30320
rect 12158 30308 12164 30320
rect 9968 30280 12164 30308
rect 4663 30212 4752 30240
rect 4884 30243 4942 30249
rect 4663 30209 4675 30212
rect 4617 30203 4675 30209
rect 4884 30209 4896 30243
rect 4930 30209 4942 30243
rect 4884 30203 4942 30209
rect 6917 30243 6975 30249
rect 6917 30209 6929 30243
rect 6963 30240 6975 30243
rect 7006 30240 7012 30252
rect 6963 30212 7012 30240
rect 6963 30209 6975 30212
rect 6917 30203 6975 30209
rect 7006 30200 7012 30212
rect 7064 30200 7070 30252
rect 7208 30181 7236 30268
rect 8018 30200 8024 30252
rect 8076 30200 8082 30252
rect 8748 30243 8806 30249
rect 8748 30209 8760 30243
rect 8794 30240 8806 30243
rect 9122 30240 9128 30252
rect 8794 30212 9128 30240
rect 8794 30209 8806 30212
rect 8748 30203 8806 30209
rect 9122 30200 9128 30212
rect 9180 30200 9186 30252
rect 9968 30249 9996 30280
rect 12158 30268 12164 30280
rect 12216 30308 12222 30320
rect 13900 30311 13958 30317
rect 12216 30280 13676 30308
rect 12216 30268 12222 30280
rect 10226 30249 10232 30252
rect 9953 30243 10011 30249
rect 9953 30209 9965 30243
rect 9999 30209 10011 30243
rect 10220 30240 10232 30249
rect 10187 30212 10232 30240
rect 9953 30203 10011 30209
rect 10220 30203 10232 30212
rect 10226 30200 10232 30203
rect 10284 30200 10290 30252
rect 10502 30200 10508 30252
rect 10560 30240 10566 30252
rect 11517 30243 11575 30249
rect 11517 30240 11529 30243
rect 10560 30212 11529 30240
rect 10560 30200 10566 30212
rect 11517 30209 11529 30212
rect 11563 30209 11575 30243
rect 11517 30203 11575 30209
rect 11701 30243 11759 30249
rect 11701 30209 11713 30243
rect 11747 30209 11759 30243
rect 11701 30203 11759 30209
rect 12529 30243 12587 30249
rect 12529 30209 12541 30243
rect 12575 30240 12587 30243
rect 12575 30212 12664 30240
rect 12575 30209 12587 30212
rect 12529 30203 12587 30209
rect 7193 30175 7251 30181
rect 7193 30141 7205 30175
rect 7239 30141 7251 30175
rect 7193 30135 7251 30141
rect 8386 30132 8392 30184
rect 8444 30172 8450 30184
rect 8481 30175 8539 30181
rect 8481 30172 8493 30175
rect 8444 30144 8493 30172
rect 8444 30132 8450 30144
rect 8481 30141 8493 30144
rect 8527 30141 8539 30175
rect 11716 30172 11744 30203
rect 8481 30135 8539 30141
rect 11348 30144 11744 30172
rect 5350 29996 5356 30048
rect 5408 30036 5414 30048
rect 5997 30039 6055 30045
rect 5997 30036 6009 30039
rect 5408 30008 6009 30036
rect 5408 29996 5414 30008
rect 5997 30005 6009 30008
rect 6043 30005 6055 30039
rect 5997 29999 6055 30005
rect 9858 29996 9864 30048
rect 9916 29996 9922 30048
rect 10134 29996 10140 30048
rect 10192 30036 10198 30048
rect 11348 30045 11376 30144
rect 12636 30113 12664 30212
rect 12986 30200 12992 30252
rect 13044 30200 13050 30252
rect 13648 30249 13676 30280
rect 13900 30277 13912 30311
rect 13946 30308 13958 30311
rect 14090 30308 14096 30320
rect 13946 30280 14096 30308
rect 13946 30277 13958 30280
rect 13900 30271 13958 30277
rect 14090 30268 14096 30280
rect 14148 30268 14154 30320
rect 16960 30308 16988 30339
rect 19886 30336 19892 30388
rect 19944 30336 19950 30388
rect 20349 30379 20407 30385
rect 20349 30345 20361 30379
rect 20395 30376 20407 30379
rect 20714 30376 20720 30388
rect 20395 30348 20720 30376
rect 20395 30345 20407 30348
rect 20349 30339 20407 30345
rect 20714 30336 20720 30348
rect 20772 30336 20778 30388
rect 21174 30336 21180 30388
rect 21232 30376 21238 30388
rect 21821 30379 21879 30385
rect 21821 30376 21833 30379
rect 21232 30348 21833 30376
rect 21232 30336 21238 30348
rect 21821 30345 21833 30348
rect 21867 30345 21879 30379
rect 22186 30376 22192 30388
rect 21821 30339 21879 30345
rect 22066 30348 22192 30376
rect 17466 30311 17524 30317
rect 17466 30308 17478 30311
rect 15304 30280 16804 30308
rect 16960 30280 17478 30308
rect 13633 30243 13691 30249
rect 13633 30209 13645 30243
rect 13679 30240 13691 30243
rect 15304 30240 15332 30280
rect 13679 30212 15332 30240
rect 15372 30243 15430 30249
rect 13679 30209 13691 30212
rect 13633 30203 13691 30209
rect 15372 30209 15384 30243
rect 15418 30240 15430 30243
rect 15418 30212 16712 30240
rect 15418 30209 15430 30212
rect 15372 30203 15430 30209
rect 13262 30132 13268 30184
rect 13320 30132 13326 30184
rect 15105 30175 15163 30181
rect 15105 30141 15117 30175
rect 15151 30141 15163 30175
rect 15105 30135 15163 30141
rect 12621 30107 12679 30113
rect 12621 30073 12633 30107
rect 12667 30073 12679 30107
rect 12621 30067 12679 30073
rect 11333 30039 11391 30045
rect 11333 30036 11345 30039
rect 10192 30008 11345 30036
rect 10192 29996 10198 30008
rect 11333 30005 11345 30008
rect 11379 30005 11391 30039
rect 11333 29999 11391 30005
rect 11514 29996 11520 30048
rect 11572 29996 11578 30048
rect 14550 29996 14556 30048
rect 14608 30036 14614 30048
rect 15013 30039 15071 30045
rect 15013 30036 15025 30039
rect 14608 30008 15025 30036
rect 14608 29996 14614 30008
rect 15013 30005 15025 30008
rect 15059 30005 15071 30039
rect 15120 30036 15148 30135
rect 16684 30113 16712 30212
rect 16776 30172 16804 30280
rect 17466 30277 17478 30280
rect 17512 30277 17524 30311
rect 17466 30271 17524 30277
rect 19536 30280 20576 30308
rect 16850 30200 16856 30252
rect 16908 30200 16914 30252
rect 17126 30200 17132 30252
rect 17184 30200 17190 30252
rect 19536 30249 19564 30280
rect 18785 30243 18843 30249
rect 18785 30209 18797 30243
rect 18831 30209 18843 30243
rect 18785 30203 18843 30209
rect 19521 30243 19579 30249
rect 19521 30209 19533 30243
rect 19567 30209 19579 30243
rect 19521 30203 19579 30209
rect 17218 30172 17224 30184
rect 16776 30144 17224 30172
rect 17218 30132 17224 30144
rect 17276 30132 17282 30184
rect 16669 30107 16727 30113
rect 16669 30073 16681 30107
rect 16715 30073 16727 30107
rect 18800 30104 18828 30203
rect 20254 30200 20260 30252
rect 20312 30200 20318 30252
rect 20548 30181 20576 30280
rect 20622 30268 20628 30320
rect 20680 30308 20686 30320
rect 22066 30308 22094 30348
rect 22186 30336 22192 30348
rect 22244 30336 22250 30388
rect 23753 30379 23811 30385
rect 23753 30345 23765 30379
rect 23799 30376 23811 30379
rect 24578 30376 24584 30388
rect 23799 30348 24584 30376
rect 23799 30345 23811 30348
rect 23753 30339 23811 30345
rect 24578 30336 24584 30348
rect 24636 30336 24642 30388
rect 25130 30336 25136 30388
rect 25188 30376 25194 30388
rect 31202 30376 31208 30388
rect 25188 30348 31208 30376
rect 25188 30336 25194 30348
rect 31202 30336 31208 30348
rect 31260 30336 31266 30388
rect 20680 30280 22094 30308
rect 20680 30268 20686 30280
rect 22278 30268 22284 30320
rect 22336 30268 22342 30320
rect 24762 30308 24768 30320
rect 23216 30280 24768 30308
rect 23216 30249 23244 30280
rect 24762 30268 24768 30280
rect 24820 30268 24826 30320
rect 26142 30308 26148 30320
rect 24872 30280 26148 30308
rect 23201 30243 23259 30249
rect 22066 30212 23152 30240
rect 20533 30175 20591 30181
rect 20533 30141 20545 30175
rect 20579 30172 20591 30175
rect 22066 30172 22094 30212
rect 20579 30144 22094 30172
rect 20579 30141 20591 30144
rect 20533 30135 20591 30141
rect 22462 30132 22468 30184
rect 22520 30132 22526 30184
rect 23124 30172 23152 30212
rect 23201 30209 23213 30243
rect 23247 30209 23259 30243
rect 23201 30203 23259 30209
rect 23750 30200 23756 30252
rect 23808 30240 23814 30252
rect 24026 30240 24032 30252
rect 23808 30212 24032 30240
rect 23808 30200 23814 30212
rect 24026 30200 24032 30212
rect 24084 30240 24090 30252
rect 24121 30243 24179 30249
rect 24121 30240 24133 30243
rect 24084 30212 24133 30240
rect 24084 30200 24090 30212
rect 24121 30209 24133 30212
rect 24167 30209 24179 30243
rect 24121 30203 24179 30209
rect 24210 30200 24216 30252
rect 24268 30240 24274 30252
rect 24394 30240 24400 30252
rect 24268 30212 24400 30240
rect 24268 30200 24274 30212
rect 24394 30200 24400 30212
rect 24452 30200 24458 30252
rect 24305 30175 24363 30181
rect 24305 30172 24317 30175
rect 23124 30144 24317 30172
rect 24305 30141 24317 30144
rect 24351 30172 24363 30175
rect 24872 30172 24900 30280
rect 26142 30268 26148 30280
rect 26200 30268 26206 30320
rect 25038 30200 25044 30252
rect 25096 30200 25102 30252
rect 27341 30243 27399 30249
rect 27341 30209 27353 30243
rect 27387 30240 27399 30243
rect 27387 30212 27476 30240
rect 27387 30209 27399 30212
rect 27341 30203 27399 30209
rect 24351 30144 24900 30172
rect 24351 30141 24363 30144
rect 24305 30135 24363 30141
rect 24946 30132 24952 30184
rect 25004 30172 25010 30184
rect 25317 30175 25375 30181
rect 25317 30172 25329 30175
rect 25004 30144 25329 30172
rect 25004 30132 25010 30144
rect 25317 30141 25329 30144
rect 25363 30141 25375 30175
rect 25317 30135 25375 30141
rect 22480 30104 22508 30132
rect 18800 30076 22508 30104
rect 16669 30067 16727 30073
rect 23382 30064 23388 30116
rect 23440 30104 23446 30116
rect 27448 30113 27476 30212
rect 27798 30200 27804 30252
rect 27856 30200 27862 30252
rect 27893 30243 27951 30249
rect 27893 30209 27905 30243
rect 27939 30240 27951 30243
rect 28074 30240 28080 30252
rect 27939 30212 28080 30240
rect 27939 30209 27951 30212
rect 27893 30203 27951 30209
rect 28074 30200 28080 30212
rect 28132 30200 28138 30252
rect 36173 30243 36231 30249
rect 36173 30209 36185 30243
rect 36219 30240 36231 30243
rect 36538 30240 36544 30252
rect 36219 30212 36544 30240
rect 36219 30209 36231 30212
rect 36173 30203 36231 30209
rect 36538 30200 36544 30212
rect 36596 30200 36602 30252
rect 27982 30132 27988 30184
rect 28040 30132 28046 30184
rect 27433 30107 27491 30113
rect 23440 30076 27292 30104
rect 23440 30064 23446 30076
rect 15470 30036 15476 30048
rect 15120 30008 15476 30036
rect 15013 29999 15071 30005
rect 15470 29996 15476 30008
rect 15528 29996 15534 30048
rect 16485 30039 16543 30045
rect 16485 30005 16497 30039
rect 16531 30036 16543 30039
rect 16574 30036 16580 30048
rect 16531 30008 16580 30036
rect 16531 30005 16543 30008
rect 16485 29999 16543 30005
rect 16574 29996 16580 30008
rect 16632 29996 16638 30048
rect 17862 29996 17868 30048
rect 17920 30036 17926 30048
rect 18601 30039 18659 30045
rect 18601 30036 18613 30039
rect 17920 30008 18613 30036
rect 17920 29996 17926 30008
rect 18601 30005 18613 30008
rect 18647 30005 18659 30039
rect 18601 29999 18659 30005
rect 18874 29996 18880 30048
rect 18932 29996 18938 30048
rect 19702 29996 19708 30048
rect 19760 29996 19766 30048
rect 20254 29996 20260 30048
rect 20312 30036 20318 30048
rect 20898 30036 20904 30048
rect 20312 30008 20904 30036
rect 20312 29996 20318 30008
rect 20898 29996 20904 30008
rect 20956 30036 20962 30048
rect 22278 30036 22284 30048
rect 20956 30008 22284 30036
rect 20956 29996 20962 30008
rect 22278 29996 22284 30008
rect 22336 29996 22342 30048
rect 27154 29996 27160 30048
rect 27212 29996 27218 30048
rect 27264 30036 27292 30076
rect 27433 30073 27445 30107
rect 27479 30073 27491 30107
rect 27433 30067 27491 30073
rect 28442 30036 28448 30048
rect 27264 30008 28448 30036
rect 28442 29996 28448 30008
rect 28500 29996 28506 30048
rect 36354 29996 36360 30048
rect 36412 29996 36418 30048
rect 1104 29946 36800 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 36800 29946
rect 1104 29872 36800 29894
rect 5258 29792 5264 29844
rect 5316 29792 5322 29844
rect 9122 29792 9128 29844
rect 9180 29792 9186 29844
rect 10226 29792 10232 29844
rect 10284 29832 10290 29844
rect 10321 29835 10379 29841
rect 10321 29832 10333 29835
rect 10284 29804 10333 29832
rect 10284 29792 10290 29804
rect 10321 29801 10333 29804
rect 10367 29801 10379 29835
rect 10321 29795 10379 29801
rect 14093 29835 14151 29841
rect 14093 29801 14105 29835
rect 14139 29832 14151 29835
rect 14274 29832 14280 29844
rect 14139 29804 14280 29832
rect 14139 29801 14151 29804
rect 14093 29795 14151 29801
rect 14274 29792 14280 29804
rect 14332 29792 14338 29844
rect 16117 29835 16175 29841
rect 16117 29801 16129 29835
rect 16163 29832 16175 29835
rect 16850 29832 16856 29844
rect 16163 29804 16856 29832
rect 16163 29801 16175 29804
rect 16117 29795 16175 29801
rect 16850 29792 16856 29804
rect 16908 29792 16914 29844
rect 17126 29792 17132 29844
rect 17184 29832 17190 29844
rect 17405 29835 17463 29841
rect 17405 29832 17417 29835
rect 17184 29804 17417 29832
rect 17184 29792 17190 29804
rect 17405 29801 17417 29804
rect 17451 29801 17463 29835
rect 17405 29795 17463 29801
rect 27798 29792 27804 29844
rect 27856 29832 27862 29844
rect 28258 29832 28264 29844
rect 27856 29804 28264 29832
rect 27856 29792 27862 29804
rect 28258 29792 28264 29804
rect 28316 29792 28322 29844
rect 5169 29767 5227 29773
rect 5169 29733 5181 29767
rect 5215 29764 5227 29767
rect 5902 29764 5908 29776
rect 5215 29736 5908 29764
rect 5215 29733 5227 29736
rect 5169 29727 5227 29733
rect 5902 29724 5908 29736
rect 5960 29724 5966 29776
rect 7558 29764 7564 29776
rect 6288 29736 7564 29764
rect 3510 29656 3516 29708
rect 3568 29696 3574 29708
rect 3789 29699 3847 29705
rect 3789 29696 3801 29699
rect 3568 29668 3801 29696
rect 3568 29656 3574 29668
rect 3789 29665 3801 29668
rect 3835 29665 3847 29699
rect 3789 29659 3847 29665
rect 5718 29656 5724 29708
rect 5776 29656 5782 29708
rect 5813 29699 5871 29705
rect 5813 29665 5825 29699
rect 5859 29696 5871 29699
rect 6288 29696 6316 29736
rect 7558 29724 7564 29736
rect 7616 29724 7622 29776
rect 13262 29764 13268 29776
rect 8956 29736 13268 29764
rect 5859 29668 6316 29696
rect 5859 29665 5871 29668
rect 5813 29659 5871 29665
rect 6362 29656 6368 29708
rect 6420 29696 6426 29708
rect 7285 29699 7343 29705
rect 7285 29696 7297 29699
rect 6420 29668 7297 29696
rect 6420 29656 6426 29668
rect 7285 29665 7297 29668
rect 7331 29696 7343 29699
rect 8956 29696 8984 29736
rect 7331 29668 8984 29696
rect 7331 29665 7343 29668
rect 7285 29659 7343 29665
rect 3602 29588 3608 29640
rect 3660 29588 3666 29640
rect 5350 29588 5356 29640
rect 5408 29628 5414 29640
rect 5629 29631 5687 29637
rect 5629 29628 5641 29631
rect 5408 29600 5641 29628
rect 5408 29588 5414 29600
rect 5629 29597 5641 29600
rect 5675 29597 5687 29631
rect 5629 29591 5687 29597
rect 7101 29631 7159 29637
rect 7101 29597 7113 29631
rect 7147 29628 7159 29631
rect 7650 29628 7656 29640
rect 7147 29600 7656 29628
rect 7147 29597 7159 29600
rect 7101 29591 7159 29597
rect 7650 29588 7656 29600
rect 7708 29628 7714 29640
rect 8202 29628 8208 29640
rect 7708 29600 8208 29628
rect 7708 29588 7714 29600
rect 8202 29588 8208 29600
rect 8260 29588 8266 29640
rect 8956 29637 8984 29668
rect 9217 29699 9275 29705
rect 9217 29665 9229 29699
rect 9263 29696 9275 29699
rect 9677 29699 9735 29705
rect 9677 29696 9689 29699
rect 9263 29668 9689 29696
rect 9263 29665 9275 29668
rect 9217 29659 9275 29665
rect 9677 29665 9689 29668
rect 9723 29665 9735 29699
rect 9677 29659 9735 29665
rect 8941 29631 8999 29637
rect 8941 29597 8953 29631
rect 8987 29597 8999 29631
rect 8941 29591 8999 29597
rect 9033 29631 9091 29637
rect 9033 29597 9045 29631
rect 9079 29628 9091 29631
rect 9490 29628 9496 29640
rect 9079 29600 9496 29628
rect 9079 29597 9091 29600
rect 9033 29591 9091 29597
rect 9490 29588 9496 29600
rect 9548 29588 9554 29640
rect 9784 29637 9812 29736
rect 13262 29724 13268 29736
rect 13320 29764 13326 29776
rect 19702 29764 19708 29776
rect 13320 29736 19708 29764
rect 13320 29724 13326 29736
rect 11514 29696 11520 29708
rect 10336 29668 11520 29696
rect 10336 29637 10364 29668
rect 11514 29656 11520 29668
rect 11572 29656 11578 29708
rect 14645 29699 14703 29705
rect 14645 29696 14657 29699
rect 12406 29668 14657 29696
rect 9585 29631 9643 29637
rect 9585 29597 9597 29631
rect 9631 29597 9643 29631
rect 9585 29591 9643 29597
rect 9769 29631 9827 29637
rect 9769 29597 9781 29631
rect 9815 29597 9827 29631
rect 9769 29591 9827 29597
rect 10321 29631 10379 29637
rect 10321 29597 10333 29631
rect 10367 29597 10379 29631
rect 10321 29591 10379 29597
rect 4034 29563 4092 29569
rect 4034 29560 4046 29563
rect 3436 29532 4046 29560
rect 3436 29501 3464 29532
rect 4034 29529 4046 29532
rect 4080 29529 4092 29563
rect 4034 29523 4092 29529
rect 7558 29520 7564 29572
rect 7616 29560 7622 29572
rect 9600 29560 9628 29591
rect 10594 29588 10600 29640
rect 10652 29588 10658 29640
rect 9858 29560 9864 29572
rect 7616 29532 9536 29560
rect 9600 29532 9864 29560
rect 7616 29520 7622 29532
rect 3421 29495 3479 29501
rect 3421 29461 3433 29495
rect 3467 29461 3479 29495
rect 3421 29455 3479 29461
rect 6178 29452 6184 29504
rect 6236 29492 6242 29504
rect 6733 29495 6791 29501
rect 6733 29492 6745 29495
rect 6236 29464 6745 29492
rect 6236 29452 6242 29464
rect 6733 29461 6745 29464
rect 6779 29461 6791 29495
rect 6733 29455 6791 29461
rect 7193 29495 7251 29501
rect 7193 29461 7205 29495
rect 7239 29492 7251 29495
rect 7834 29492 7840 29504
rect 7239 29464 7840 29492
rect 7239 29461 7251 29464
rect 7193 29455 7251 29461
rect 7834 29452 7840 29464
rect 7892 29452 7898 29504
rect 9508 29492 9536 29532
rect 9858 29520 9864 29532
rect 9916 29560 9922 29572
rect 10962 29560 10968 29572
rect 9916 29532 10968 29560
rect 9916 29520 9922 29532
rect 10962 29520 10968 29532
rect 11020 29520 11026 29572
rect 10502 29492 10508 29504
rect 9508 29464 10508 29492
rect 10502 29452 10508 29464
rect 10560 29492 10566 29504
rect 12406 29492 12434 29668
rect 14645 29665 14657 29668
rect 14691 29665 14703 29699
rect 14645 29659 14703 29665
rect 14461 29631 14519 29637
rect 14461 29597 14473 29631
rect 14507 29628 14519 29631
rect 14550 29628 14556 29640
rect 14507 29600 14556 29628
rect 14507 29597 14519 29600
rect 14461 29591 14519 29597
rect 14550 29588 14556 29600
rect 14608 29588 14614 29640
rect 14660 29628 14688 29659
rect 16574 29656 16580 29708
rect 16632 29656 16638 29708
rect 16776 29705 16804 29736
rect 19702 29724 19708 29736
rect 19760 29724 19766 29776
rect 16761 29699 16819 29705
rect 16761 29665 16773 29699
rect 16807 29665 16819 29699
rect 16761 29659 16819 29665
rect 17957 29699 18015 29705
rect 17957 29665 17969 29699
rect 18003 29696 18015 29699
rect 18874 29696 18880 29708
rect 18003 29668 18880 29696
rect 18003 29665 18015 29668
rect 17957 29659 18015 29665
rect 17972 29628 18000 29659
rect 18874 29656 18880 29668
rect 18932 29656 18938 29708
rect 22646 29656 22652 29708
rect 22704 29696 22710 29708
rect 24946 29696 24952 29708
rect 22704 29668 24952 29696
rect 22704 29656 22710 29668
rect 24946 29656 24952 29668
rect 25004 29656 25010 29708
rect 26878 29656 26884 29708
rect 26936 29656 26942 29708
rect 14660 29600 18000 29628
rect 21082 29588 21088 29640
rect 21140 29628 21146 29640
rect 23290 29628 23296 29640
rect 21140 29600 23296 29628
rect 21140 29588 21146 29600
rect 23290 29588 23296 29600
rect 23348 29588 23354 29640
rect 24854 29588 24860 29640
rect 24912 29588 24918 29640
rect 27154 29637 27160 29640
rect 27148 29628 27160 29637
rect 27115 29600 27160 29628
rect 27148 29591 27160 29600
rect 27154 29588 27160 29591
rect 27212 29588 27218 29640
rect 29362 29588 29368 29640
rect 29420 29588 29426 29640
rect 29549 29631 29607 29637
rect 29549 29597 29561 29631
rect 29595 29628 29607 29631
rect 30190 29628 30196 29640
rect 29595 29600 30196 29628
rect 29595 29597 29607 29600
rect 29549 29591 29607 29597
rect 30190 29588 30196 29600
rect 30248 29588 30254 29640
rect 31202 29588 31208 29640
rect 31260 29588 31266 29640
rect 16942 29520 16948 29572
rect 17000 29560 17006 29572
rect 17770 29560 17776 29572
rect 17000 29532 17776 29560
rect 17000 29520 17006 29532
rect 17770 29520 17776 29532
rect 17828 29520 17834 29572
rect 25194 29563 25252 29569
rect 25194 29560 25206 29563
rect 24688 29532 25206 29560
rect 10560 29464 12434 29492
rect 10560 29452 10566 29464
rect 12986 29452 12992 29504
rect 13044 29492 13050 29504
rect 14553 29495 14611 29501
rect 14553 29492 14565 29495
rect 13044 29464 14565 29492
rect 13044 29452 13050 29464
rect 14553 29461 14565 29464
rect 14599 29461 14611 29495
rect 14553 29455 14611 29461
rect 16485 29495 16543 29501
rect 16485 29461 16497 29495
rect 16531 29492 16543 29495
rect 17310 29492 17316 29504
rect 16531 29464 17316 29492
rect 16531 29461 16543 29464
rect 16485 29455 16543 29461
rect 17310 29452 17316 29464
rect 17368 29492 17374 29504
rect 17678 29492 17684 29504
rect 17368 29464 17684 29492
rect 17368 29452 17374 29464
rect 17678 29452 17684 29464
rect 17736 29492 17742 29504
rect 17865 29495 17923 29501
rect 17865 29492 17877 29495
rect 17736 29464 17877 29492
rect 17736 29452 17742 29464
rect 17865 29461 17877 29464
rect 17911 29461 17923 29495
rect 17865 29455 17923 29461
rect 20438 29452 20444 29504
rect 20496 29492 20502 29504
rect 20806 29492 20812 29504
rect 20496 29464 20812 29492
rect 20496 29452 20502 29464
rect 20806 29452 20812 29464
rect 20864 29452 20870 29504
rect 24688 29501 24716 29532
rect 25194 29529 25206 29532
rect 25240 29529 25252 29563
rect 29794 29563 29852 29569
rect 29794 29560 29806 29563
rect 25194 29523 25252 29529
rect 29196 29532 29806 29560
rect 24673 29495 24731 29501
rect 24673 29461 24685 29495
rect 24719 29461 24731 29495
rect 24673 29455 24731 29461
rect 25498 29452 25504 29504
rect 25556 29492 25562 29504
rect 29196 29501 29224 29532
rect 29794 29529 29806 29532
rect 29840 29529 29852 29563
rect 29794 29523 29852 29529
rect 26329 29495 26387 29501
rect 26329 29492 26341 29495
rect 25556 29464 26341 29492
rect 25556 29452 25562 29464
rect 26329 29461 26341 29464
rect 26375 29461 26387 29495
rect 26329 29455 26387 29461
rect 29181 29495 29239 29501
rect 29181 29461 29193 29495
rect 29227 29461 29239 29495
rect 29181 29455 29239 29461
rect 29914 29452 29920 29504
rect 29972 29492 29978 29504
rect 30929 29495 30987 29501
rect 30929 29492 30941 29495
rect 29972 29464 30941 29492
rect 29972 29452 29978 29464
rect 30929 29461 30941 29464
rect 30975 29461 30987 29495
rect 30929 29455 30987 29461
rect 31018 29452 31024 29504
rect 31076 29452 31082 29504
rect 1104 29402 36800 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 36800 29402
rect 1104 29328 36800 29350
rect 3602 29248 3608 29300
rect 3660 29288 3666 29300
rect 4249 29291 4307 29297
rect 4249 29288 4261 29291
rect 3660 29260 4261 29288
rect 3660 29248 3666 29260
rect 4249 29257 4261 29260
rect 4295 29257 4307 29291
rect 4249 29251 4307 29257
rect 4617 29291 4675 29297
rect 4617 29257 4629 29291
rect 4663 29288 4675 29291
rect 4706 29288 4712 29300
rect 4663 29260 4712 29288
rect 4663 29257 4675 29260
rect 4617 29251 4675 29257
rect 4706 29248 4712 29260
rect 4764 29288 4770 29300
rect 5718 29288 5724 29300
rect 4764 29260 5724 29288
rect 4764 29248 4770 29260
rect 5718 29248 5724 29260
rect 5776 29248 5782 29300
rect 5997 29291 6055 29297
rect 5997 29257 6009 29291
rect 6043 29257 6055 29291
rect 5997 29251 6055 29257
rect 6012 29220 6040 29251
rect 7834 29248 7840 29300
rect 7892 29248 7898 29300
rect 9490 29248 9496 29300
rect 9548 29288 9554 29300
rect 10318 29288 10324 29300
rect 9548 29260 10324 29288
rect 9548 29248 9554 29260
rect 10318 29248 10324 29260
rect 10376 29288 10382 29300
rect 10594 29288 10600 29300
rect 10376 29260 10600 29288
rect 10376 29248 10382 29260
rect 10594 29248 10600 29260
rect 10652 29248 10658 29300
rect 20622 29288 20628 29300
rect 19812 29260 20628 29288
rect 6702 29223 6760 29229
rect 6702 29220 6714 29223
rect 6012 29192 6714 29220
rect 6702 29189 6714 29192
rect 6748 29189 6760 29223
rect 19426 29220 19432 29232
rect 6702 29183 6760 29189
rect 18340 29192 19432 29220
rect 1578 29112 1584 29164
rect 1636 29112 1642 29164
rect 1762 29112 1768 29164
rect 1820 29112 1826 29164
rect 2038 29161 2044 29164
rect 2032 29115 2044 29161
rect 2038 29112 2044 29115
rect 2096 29112 2102 29164
rect 4709 29155 4767 29161
rect 4709 29121 4721 29155
rect 4755 29152 4767 29155
rect 5902 29152 5908 29164
rect 4755 29124 5908 29152
rect 4755 29121 4767 29124
rect 4709 29115 4767 29121
rect 5902 29112 5908 29124
rect 5960 29112 5966 29164
rect 6178 29112 6184 29164
rect 6236 29112 6242 29164
rect 6457 29155 6515 29161
rect 6457 29121 6469 29155
rect 6503 29152 6515 29155
rect 8386 29152 8392 29164
rect 6503 29124 8392 29152
rect 6503 29121 6515 29124
rect 6457 29115 6515 29121
rect 8386 29112 8392 29124
rect 8444 29112 8450 29164
rect 12526 29112 12532 29164
rect 12584 29112 12590 29164
rect 18340 29161 18368 29192
rect 19426 29180 19432 29192
rect 19484 29180 19490 29232
rect 18325 29155 18383 29161
rect 18325 29121 18337 29155
rect 18371 29121 18383 29155
rect 18325 29115 18383 29121
rect 18592 29155 18650 29161
rect 18592 29121 18604 29155
rect 18638 29152 18650 29155
rect 19150 29152 19156 29164
rect 18638 29124 19156 29152
rect 18638 29121 18650 29124
rect 18592 29115 18650 29121
rect 19150 29112 19156 29124
rect 19208 29112 19214 29164
rect 19812 29161 19840 29260
rect 20622 29248 20628 29260
rect 20680 29248 20686 29300
rect 24854 29248 24860 29300
rect 24912 29288 24918 29300
rect 25133 29291 25191 29297
rect 25133 29288 25145 29291
rect 24912 29260 25145 29288
rect 24912 29248 24918 29260
rect 25133 29257 25145 29260
rect 25179 29257 25191 29291
rect 25133 29251 25191 29257
rect 25498 29248 25504 29300
rect 25556 29248 25562 29300
rect 27430 29288 27436 29300
rect 27264 29260 27436 29288
rect 22462 29180 22468 29232
rect 22520 29220 22526 29232
rect 22520 29192 23796 29220
rect 22520 29180 22526 29192
rect 19797 29155 19855 29161
rect 19797 29121 19809 29155
rect 19843 29121 19855 29155
rect 19797 29115 19855 29121
rect 20990 29112 20996 29164
rect 21048 29112 21054 29164
rect 22646 29112 22652 29164
rect 22704 29112 22710 29164
rect 22922 29161 22928 29164
rect 22916 29115 22928 29161
rect 22922 29112 22928 29115
rect 22980 29112 22986 29164
rect 23290 29112 23296 29164
rect 23348 29152 23354 29164
rect 23768 29152 23796 29192
rect 24486 29180 24492 29232
rect 24544 29220 24550 29232
rect 25516 29220 25544 29248
rect 24544 29192 25544 29220
rect 24544 29180 24550 29192
rect 27264 29161 27292 29260
rect 27430 29248 27436 29260
rect 27488 29288 27494 29300
rect 27488 29260 28948 29288
rect 27488 29248 27494 29260
rect 28920 29220 28948 29260
rect 29362 29248 29368 29300
rect 29420 29288 29426 29300
rect 29549 29291 29607 29297
rect 29549 29288 29561 29291
rect 29420 29260 29561 29288
rect 29420 29248 29426 29260
rect 29549 29257 29561 29260
rect 29595 29257 29607 29291
rect 29549 29251 29607 29257
rect 29914 29248 29920 29300
rect 29972 29248 29978 29300
rect 29932 29220 29960 29248
rect 28920 29192 29960 29220
rect 30828 29223 30886 29229
rect 30828 29189 30840 29223
rect 30874 29220 30886 29223
rect 31018 29220 31024 29232
rect 30874 29192 31024 29220
rect 30874 29189 30886 29192
rect 30828 29183 30886 29189
rect 31018 29180 31024 29192
rect 31076 29180 31082 29232
rect 27249 29155 27307 29161
rect 23348 29124 23704 29152
rect 23768 29124 25820 29152
rect 23348 29112 23354 29124
rect 4893 29087 4951 29093
rect 4893 29053 4905 29087
rect 4939 29084 4951 29087
rect 6362 29084 6368 29096
rect 4939 29056 6368 29084
rect 4939 29053 4951 29056
rect 4893 29047 4951 29053
rect 6362 29044 6368 29056
rect 6420 29044 6426 29096
rect 19981 29087 20039 29093
rect 19981 29053 19993 29087
rect 20027 29084 20039 29087
rect 20530 29084 20536 29096
rect 20027 29056 20536 29084
rect 20027 29053 20039 29056
rect 19981 29047 20039 29053
rect 20530 29044 20536 29056
rect 20588 29044 20594 29096
rect 20714 29044 20720 29096
rect 20772 29044 20778 29096
rect 20806 29044 20812 29096
rect 20864 29093 20870 29096
rect 20864 29087 20892 29093
rect 20880 29053 20892 29087
rect 20864 29047 20892 29053
rect 20864 29044 20870 29047
rect 21174 29044 21180 29096
rect 21232 29084 21238 29096
rect 21637 29087 21695 29093
rect 21637 29084 21649 29087
rect 21232 29056 21649 29084
rect 21232 29044 21238 29056
rect 21637 29053 21649 29056
rect 21683 29053 21695 29087
rect 21637 29047 21695 29053
rect 1397 29019 1455 29025
rect 1397 28985 1409 29019
rect 1443 29016 1455 29019
rect 1670 29016 1676 29028
rect 1443 28988 1676 29016
rect 1443 28985 1455 28988
rect 1397 28979 1455 28985
rect 1670 28976 1676 28988
rect 1728 28976 1734 29028
rect 12345 29019 12403 29025
rect 12345 28985 12357 29019
rect 12391 29016 12403 29019
rect 12434 29016 12440 29028
rect 12391 28988 12440 29016
rect 12391 28985 12403 28988
rect 12345 28979 12403 28985
rect 12434 28976 12440 28988
rect 12492 28976 12498 29028
rect 20438 29016 20444 29028
rect 19352 28988 20444 29016
rect 3142 28908 3148 28960
rect 3200 28908 3206 28960
rect 5810 28908 5816 28960
rect 5868 28948 5874 28960
rect 10686 28948 10692 28960
rect 5868 28920 10692 28948
rect 5868 28908 5874 28920
rect 10686 28908 10692 28920
rect 10744 28948 10750 28960
rect 19352 28948 19380 28988
rect 20438 28976 20444 28988
rect 20496 28976 20502 29028
rect 23676 29016 23704 29124
rect 24026 29044 24032 29096
rect 24084 29084 24090 29096
rect 25038 29084 25044 29096
rect 24084 29056 25044 29084
rect 24084 29044 24090 29056
rect 25038 29044 25044 29056
rect 25096 29084 25102 29096
rect 25792 29093 25820 29124
rect 27249 29121 27261 29155
rect 27295 29121 27307 29155
rect 27249 29115 27307 29121
rect 27356 29124 27660 29152
rect 25593 29087 25651 29093
rect 25593 29084 25605 29087
rect 25096 29056 25605 29084
rect 25096 29044 25102 29056
rect 25593 29053 25605 29056
rect 25639 29053 25651 29087
rect 25593 29047 25651 29053
rect 25777 29087 25835 29093
rect 25777 29053 25789 29087
rect 25823 29084 25835 29087
rect 27356 29084 27384 29124
rect 25823 29056 27384 29084
rect 27433 29087 27491 29093
rect 25823 29053 25835 29056
rect 25777 29047 25835 29053
rect 27433 29053 27445 29087
rect 27479 29084 27491 29087
rect 27522 29084 27528 29096
rect 27479 29056 27528 29084
rect 27479 29053 27491 29056
rect 27433 29047 27491 29053
rect 27522 29044 27528 29056
rect 27580 29044 27586 29096
rect 27632 29084 27660 29124
rect 28166 29112 28172 29164
rect 28224 29112 28230 29164
rect 28258 29112 28264 29164
rect 28316 29161 28322 29164
rect 28316 29155 28344 29161
rect 28332 29121 28344 29155
rect 28316 29115 28344 29121
rect 28316 29112 28322 29115
rect 28442 29112 28448 29164
rect 28500 29112 28506 29164
rect 29012 29124 30236 29152
rect 29012 29084 29040 29124
rect 27632 29056 29040 29084
rect 29822 29044 29828 29096
rect 29880 29084 29886 29096
rect 30208 29093 30236 29124
rect 30558 29112 30564 29164
rect 30616 29112 30622 29164
rect 30009 29087 30067 29093
rect 30009 29084 30021 29087
rect 29880 29056 30021 29084
rect 29880 29044 29886 29056
rect 30009 29053 30021 29056
rect 30055 29053 30067 29087
rect 30009 29047 30067 29053
rect 30193 29087 30251 29093
rect 30193 29053 30205 29087
rect 30239 29084 30251 29087
rect 30466 29084 30472 29096
rect 30239 29056 30472 29084
rect 30239 29053 30251 29056
rect 30193 29047 30251 29053
rect 30466 29044 30472 29056
rect 30524 29044 30530 29096
rect 27893 29019 27951 29025
rect 27893 29016 27905 29019
rect 23676 28988 27905 29016
rect 27893 28985 27905 28988
rect 27939 28985 27951 29019
rect 27893 28979 27951 28985
rect 29086 28976 29092 29028
rect 29144 28976 29150 29028
rect 10744 28920 19380 28948
rect 19705 28951 19763 28957
rect 10744 28908 10750 28920
rect 19705 28917 19717 28951
rect 19751 28948 19763 28951
rect 19886 28948 19892 28960
rect 19751 28920 19892 28948
rect 19751 28917 19763 28920
rect 19705 28911 19763 28917
rect 19886 28908 19892 28920
rect 19944 28948 19950 28960
rect 20806 28948 20812 28960
rect 19944 28920 20812 28948
rect 19944 28908 19950 28920
rect 20806 28908 20812 28920
rect 20864 28948 20870 28960
rect 21542 28948 21548 28960
rect 20864 28920 21548 28948
rect 20864 28908 20870 28920
rect 21542 28908 21548 28920
rect 21600 28908 21606 28960
rect 23658 28908 23664 28960
rect 23716 28948 23722 28960
rect 24029 28951 24087 28957
rect 24029 28948 24041 28951
rect 23716 28920 24041 28948
rect 23716 28908 23722 28920
rect 24029 28917 24041 28920
rect 24075 28948 24087 28951
rect 24578 28948 24584 28960
rect 24075 28920 24584 28948
rect 24075 28917 24087 28920
rect 24029 28911 24087 28917
rect 24578 28908 24584 28920
rect 24636 28948 24642 28960
rect 25498 28948 25504 28960
rect 24636 28920 25504 28948
rect 24636 28908 24642 28920
rect 25498 28908 25504 28920
rect 25556 28908 25562 28960
rect 28166 28908 28172 28960
rect 28224 28948 28230 28960
rect 28810 28948 28816 28960
rect 28224 28920 28816 28948
rect 28224 28908 28230 28920
rect 28810 28908 28816 28920
rect 28868 28908 28874 28960
rect 31938 28908 31944 28960
rect 31996 28908 32002 28960
rect 1104 28858 36800 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 36800 28858
rect 1104 28784 36800 28806
rect 2038 28704 2044 28756
rect 2096 28704 2102 28756
rect 17494 28744 17500 28756
rect 5092 28716 9260 28744
rect 2409 28679 2467 28685
rect 2409 28645 2421 28679
rect 2455 28645 2467 28679
rect 2409 28639 2467 28645
rect 2225 28543 2283 28549
rect 2225 28509 2237 28543
rect 2271 28540 2283 28543
rect 2424 28540 2452 28639
rect 3053 28611 3111 28617
rect 3053 28577 3065 28611
rect 3099 28608 3111 28611
rect 3510 28608 3516 28620
rect 3099 28580 3516 28608
rect 3099 28577 3111 28580
rect 3053 28571 3111 28577
rect 3510 28568 3516 28580
rect 3568 28608 3574 28620
rect 5092 28608 5120 28716
rect 5350 28676 5356 28688
rect 5184 28648 5356 28676
rect 5184 28617 5212 28648
rect 5350 28636 5356 28648
rect 5408 28636 5414 28688
rect 5810 28636 5816 28688
rect 5868 28636 5874 28688
rect 8938 28636 8944 28688
rect 8996 28636 9002 28688
rect 3568 28580 5120 28608
rect 5169 28611 5227 28617
rect 3568 28568 3574 28580
rect 5169 28577 5181 28611
rect 5215 28577 5227 28611
rect 5169 28571 5227 28577
rect 5902 28568 5908 28620
rect 5960 28608 5966 28620
rect 6089 28611 6147 28617
rect 6089 28608 6101 28611
rect 5960 28580 6101 28608
rect 5960 28568 5966 28580
rect 6089 28577 6101 28580
rect 6135 28577 6147 28611
rect 6089 28571 6147 28577
rect 6365 28611 6423 28617
rect 6365 28577 6377 28611
rect 6411 28608 6423 28611
rect 6546 28608 6552 28620
rect 6411 28580 6552 28608
rect 6411 28577 6423 28580
rect 6365 28571 6423 28577
rect 6546 28568 6552 28580
rect 6604 28568 6610 28620
rect 2271 28512 2452 28540
rect 2271 28509 2283 28512
rect 2225 28503 2283 28509
rect 5350 28500 5356 28552
rect 5408 28500 5414 28552
rect 6178 28500 6184 28552
rect 6236 28549 6242 28552
rect 9232 28549 9260 28716
rect 14752 28716 17500 28744
rect 13541 28679 13599 28685
rect 9784 28648 11008 28676
rect 9784 28552 9812 28648
rect 10870 28568 10876 28620
rect 10928 28568 10934 28620
rect 10980 28608 11008 28648
rect 13541 28645 13553 28679
rect 13587 28676 13599 28679
rect 14366 28676 14372 28688
rect 13587 28648 14372 28676
rect 13587 28645 13599 28648
rect 13541 28639 13599 28645
rect 14366 28636 14372 28648
rect 14424 28676 14430 28688
rect 14752 28685 14780 28716
rect 17494 28704 17500 28716
rect 17552 28744 17558 28756
rect 17552 28716 18644 28744
rect 17552 28704 17558 28716
rect 14737 28679 14795 28685
rect 14424 28648 14596 28676
rect 14424 28636 14430 28648
rect 11238 28608 11244 28620
rect 11296 28617 11302 28620
rect 11296 28611 11324 28617
rect 10980 28580 11244 28608
rect 11238 28568 11244 28580
rect 11312 28577 11324 28611
rect 11296 28571 11324 28577
rect 11425 28611 11483 28617
rect 11425 28577 11437 28611
rect 11471 28608 11483 28611
rect 11606 28608 11612 28620
rect 11471 28580 11612 28608
rect 11471 28577 11483 28580
rect 11425 28571 11483 28577
rect 11296 28568 11302 28571
rect 11606 28568 11612 28580
rect 11664 28568 11670 28620
rect 12158 28568 12164 28620
rect 12216 28568 12222 28620
rect 14090 28568 14096 28620
rect 14148 28608 14154 28620
rect 14458 28608 14464 28620
rect 14148 28580 14464 28608
rect 14148 28568 14154 28580
rect 14458 28568 14464 28580
rect 14516 28568 14522 28620
rect 14568 28608 14596 28648
rect 14737 28645 14749 28679
rect 14783 28645 14795 28679
rect 14737 28639 14795 28645
rect 16574 28636 16580 28688
rect 16632 28676 16638 28688
rect 18616 28676 18644 28716
rect 19150 28704 19156 28756
rect 19208 28744 19214 28756
rect 19245 28747 19303 28753
rect 19245 28744 19257 28747
rect 19208 28716 19257 28744
rect 19208 28704 19214 28716
rect 19245 28713 19257 28716
rect 19291 28713 19303 28747
rect 19245 28707 19303 28713
rect 20272 28716 22876 28744
rect 20272 28676 20300 28716
rect 16632 28648 17724 28676
rect 18616 28648 20116 28676
rect 16632 28636 16638 28648
rect 17696 28620 17724 28648
rect 15130 28611 15188 28617
rect 15130 28608 15142 28611
rect 14568 28580 15142 28608
rect 15130 28577 15142 28580
rect 15176 28577 15188 28611
rect 15130 28571 15188 28577
rect 15289 28611 15347 28617
rect 15289 28577 15301 28611
rect 15335 28608 15347 28611
rect 15335 28580 16896 28608
rect 15335 28577 15347 28580
rect 15289 28571 15347 28577
rect 6236 28543 6264 28549
rect 6252 28509 6264 28543
rect 6236 28503 6264 28509
rect 9217 28543 9275 28549
rect 9217 28509 9229 28543
rect 9263 28540 9275 28543
rect 9306 28540 9312 28552
rect 9263 28512 9312 28540
rect 9263 28509 9275 28512
rect 9217 28503 9275 28509
rect 6236 28500 6242 28503
rect 9306 28500 9312 28512
rect 9364 28500 9370 28552
rect 9493 28543 9551 28549
rect 9493 28509 9505 28543
rect 9539 28540 9551 28543
rect 9766 28540 9772 28552
rect 9539 28512 9772 28540
rect 9539 28509 9551 28512
rect 9493 28503 9551 28509
rect 9766 28500 9772 28512
rect 9824 28500 9830 28552
rect 10042 28500 10048 28552
rect 10100 28540 10106 28552
rect 10229 28543 10287 28549
rect 10229 28540 10241 28543
rect 10100 28512 10241 28540
rect 10100 28500 10106 28512
rect 10229 28509 10241 28512
rect 10275 28509 10287 28543
rect 10229 28503 10287 28509
rect 10410 28500 10416 28552
rect 10468 28500 10474 28552
rect 11146 28500 11152 28552
rect 11204 28500 11210 28552
rect 12434 28549 12440 28552
rect 12428 28503 12440 28549
rect 12434 28500 12440 28503
rect 12492 28500 12498 28552
rect 13906 28500 13912 28552
rect 13964 28540 13970 28552
rect 14277 28543 14335 28549
rect 14277 28540 14289 28543
rect 13964 28512 14289 28540
rect 13964 28500 13970 28512
rect 14277 28509 14289 28512
rect 14323 28509 14335 28543
rect 14277 28503 14335 28509
rect 15010 28500 15016 28552
rect 15068 28500 15074 28552
rect 2777 28475 2835 28481
rect 2777 28441 2789 28475
rect 2823 28472 2835 28475
rect 3142 28472 3148 28484
rect 2823 28444 3148 28472
rect 2823 28441 2835 28444
rect 2777 28435 2835 28441
rect 3142 28432 3148 28444
rect 3200 28472 3206 28484
rect 8941 28475 8999 28481
rect 3200 28444 4568 28472
rect 3200 28432 3206 28444
rect 2866 28364 2872 28416
rect 2924 28364 2930 28416
rect 4540 28404 4568 28444
rect 8941 28441 8953 28475
rect 8987 28472 8999 28475
rect 9401 28475 9459 28481
rect 9401 28472 9413 28475
rect 8987 28444 9413 28472
rect 8987 28441 8999 28444
rect 8941 28435 8999 28441
rect 9401 28441 9413 28444
rect 9447 28441 9459 28475
rect 9401 28435 9459 28441
rect 6086 28404 6092 28416
rect 4540 28376 6092 28404
rect 6086 28364 6092 28376
rect 6144 28364 6150 28416
rect 7009 28407 7067 28413
rect 7009 28373 7021 28407
rect 7055 28404 7067 28407
rect 7098 28404 7104 28416
rect 7055 28376 7104 28404
rect 7055 28373 7067 28376
rect 7009 28367 7067 28373
rect 7098 28364 7104 28376
rect 7156 28364 7162 28416
rect 8570 28364 8576 28416
rect 8628 28404 8634 28416
rect 9125 28407 9183 28413
rect 9125 28404 9137 28407
rect 8628 28376 9137 28404
rect 8628 28364 8634 28376
rect 9125 28373 9137 28376
rect 9171 28373 9183 28407
rect 9125 28367 9183 28373
rect 12066 28364 12072 28416
rect 12124 28364 12130 28416
rect 13354 28364 13360 28416
rect 13412 28404 13418 28416
rect 14274 28404 14280 28416
rect 13412 28376 14280 28404
rect 13412 28364 13418 28376
rect 14274 28364 14280 28376
rect 14332 28404 14338 28416
rect 15010 28404 15016 28416
rect 14332 28376 15016 28404
rect 14332 28364 14338 28376
rect 15010 28364 15016 28376
rect 15068 28364 15074 28416
rect 15286 28364 15292 28416
rect 15344 28404 15350 28416
rect 15933 28407 15991 28413
rect 15933 28404 15945 28407
rect 15344 28376 15945 28404
rect 15344 28364 15350 28376
rect 15933 28373 15945 28376
rect 15979 28373 15991 28407
rect 16868 28404 16896 28580
rect 16942 28568 16948 28620
rect 17000 28568 17006 28620
rect 17586 28568 17592 28620
rect 17644 28568 17650 28620
rect 17678 28568 17684 28620
rect 17736 28608 17742 28620
rect 17865 28611 17923 28617
rect 17865 28608 17877 28611
rect 17736 28580 17877 28608
rect 17736 28568 17742 28580
rect 17865 28577 17877 28580
rect 17911 28577 17923 28611
rect 17865 28571 17923 28577
rect 18690 28568 18696 28620
rect 18748 28608 18754 28620
rect 18748 28580 19840 28608
rect 18748 28568 18754 28580
rect 17126 28500 17132 28552
rect 17184 28500 17190 28552
rect 17954 28500 17960 28552
rect 18012 28549 18018 28552
rect 18012 28543 18040 28549
rect 18028 28509 18040 28543
rect 18012 28503 18040 28509
rect 18012 28500 18018 28503
rect 18138 28500 18144 28552
rect 18196 28500 18202 28552
rect 19429 28543 19487 28549
rect 19429 28509 19441 28543
rect 19475 28540 19487 28543
rect 19475 28512 19564 28540
rect 19475 28509 19487 28512
rect 19429 28503 19487 28509
rect 18046 28404 18052 28416
rect 16868 28376 18052 28404
rect 15933 28367 15991 28373
rect 18046 28364 18052 28376
rect 18104 28404 18110 28416
rect 18598 28404 18604 28416
rect 18104 28376 18604 28404
rect 18104 28364 18110 28376
rect 18598 28364 18604 28376
rect 18656 28364 18662 28416
rect 18785 28407 18843 28413
rect 18785 28373 18797 28407
rect 18831 28404 18843 28407
rect 18874 28404 18880 28416
rect 18831 28376 18880 28404
rect 18831 28373 18843 28376
rect 18785 28367 18843 28373
rect 18874 28364 18880 28376
rect 18932 28364 18938 28416
rect 19536 28413 19564 28512
rect 19521 28407 19579 28413
rect 19521 28373 19533 28407
rect 19567 28373 19579 28407
rect 19812 28404 19840 28580
rect 19978 28568 19984 28620
rect 20036 28568 20042 28620
rect 19886 28500 19892 28552
rect 19944 28500 19950 28552
rect 20088 28540 20116 28648
rect 20180 28648 20300 28676
rect 20180 28620 20208 28648
rect 20714 28636 20720 28688
rect 20772 28676 20778 28688
rect 22848 28676 22876 28716
rect 22922 28704 22928 28756
rect 22980 28744 22986 28756
rect 23017 28747 23075 28753
rect 23017 28744 23029 28747
rect 22980 28716 23029 28744
rect 22980 28704 22986 28716
rect 23017 28713 23029 28716
rect 23063 28713 23075 28747
rect 23017 28707 23075 28713
rect 25409 28747 25467 28753
rect 25409 28713 25421 28747
rect 25455 28744 25467 28747
rect 25866 28744 25872 28756
rect 25455 28716 25872 28744
rect 25455 28713 25467 28716
rect 25409 28707 25467 28713
rect 25866 28704 25872 28716
rect 25924 28704 25930 28756
rect 26142 28704 26148 28756
rect 26200 28744 26206 28756
rect 30745 28747 30803 28753
rect 26200 28716 30696 28744
rect 26200 28704 26206 28716
rect 27982 28676 27988 28688
rect 20772 28648 21312 28676
rect 22848 28648 27988 28676
rect 20772 28636 20778 28648
rect 20162 28568 20168 28620
rect 20220 28568 20226 28620
rect 21082 28608 21088 28620
rect 20272 28580 21088 28608
rect 20272 28540 20300 28580
rect 21082 28568 21088 28580
rect 21140 28608 21146 28620
rect 21177 28611 21235 28617
rect 21177 28608 21189 28611
rect 21140 28580 21189 28608
rect 21140 28568 21146 28580
rect 21177 28577 21189 28580
rect 21223 28577 21235 28611
rect 21284 28608 21312 28648
rect 21453 28611 21511 28617
rect 21453 28608 21465 28611
rect 21284 28580 21465 28608
rect 21177 28571 21235 28577
rect 21453 28577 21465 28580
rect 21499 28577 21511 28611
rect 21453 28571 21511 28577
rect 21542 28568 21548 28620
rect 21600 28617 21606 28620
rect 21600 28611 21628 28617
rect 21616 28577 21628 28611
rect 23382 28608 23388 28620
rect 21600 28571 21628 28577
rect 21744 28580 23388 28608
rect 21600 28568 21606 28571
rect 21744 28552 21772 28580
rect 23382 28568 23388 28580
rect 23440 28568 23446 28620
rect 23952 28617 23980 28648
rect 27982 28636 27988 28648
rect 28040 28636 28046 28688
rect 30668 28676 30696 28716
rect 30745 28713 30757 28747
rect 30791 28744 30803 28747
rect 31202 28744 31208 28756
rect 30791 28716 31208 28744
rect 30791 28713 30803 28716
rect 30745 28707 30803 28713
rect 31202 28704 31208 28716
rect 31260 28704 31266 28756
rect 30668 28648 31340 28676
rect 23937 28611 23995 28617
rect 23937 28577 23949 28611
rect 23983 28577 23995 28611
rect 26418 28608 26424 28620
rect 23937 28571 23995 28577
rect 25148 28580 26424 28608
rect 20088 28512 20300 28540
rect 20533 28543 20591 28549
rect 20533 28509 20545 28543
rect 20579 28540 20591 28543
rect 20622 28540 20628 28552
rect 20579 28512 20628 28540
rect 20579 28509 20591 28512
rect 20533 28503 20591 28509
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 20714 28500 20720 28552
rect 20772 28500 20778 28552
rect 21726 28500 21732 28552
rect 21784 28500 21790 28552
rect 23201 28543 23259 28549
rect 23201 28509 23213 28543
rect 23247 28540 23259 28543
rect 23753 28543 23811 28549
rect 23247 28512 23336 28540
rect 23247 28509 23259 28512
rect 23201 28503 23259 28509
rect 21726 28404 21732 28416
rect 19812 28376 21732 28404
rect 19521 28367 19579 28373
rect 21726 28364 21732 28376
rect 21784 28364 21790 28416
rect 22370 28364 22376 28416
rect 22428 28364 22434 28416
rect 23308 28413 23336 28512
rect 23753 28509 23765 28543
rect 23799 28540 23811 28543
rect 25148 28540 25176 28580
rect 26418 28568 26424 28580
rect 26476 28568 26482 28620
rect 27430 28568 27436 28620
rect 27488 28568 27494 28620
rect 27522 28568 27528 28620
rect 27580 28608 27586 28620
rect 28077 28611 28135 28617
rect 28077 28608 28089 28611
rect 27580 28580 28089 28608
rect 27580 28568 27586 28580
rect 28077 28577 28089 28580
rect 28123 28577 28135 28611
rect 28077 28571 28135 28577
rect 28166 28568 28172 28620
rect 28224 28608 28230 28620
rect 28353 28611 28411 28617
rect 28353 28608 28365 28611
rect 28224 28580 28365 28608
rect 28224 28568 28230 28580
rect 28353 28577 28365 28580
rect 28399 28577 28411 28611
rect 28353 28571 28411 28577
rect 28442 28568 28448 28620
rect 28500 28617 28506 28620
rect 28500 28611 28528 28617
rect 28516 28577 28528 28611
rect 28500 28571 28528 28577
rect 28500 28568 28506 28571
rect 28810 28568 28816 28620
rect 28868 28608 28874 28620
rect 31312 28617 31340 28648
rect 31205 28611 31263 28617
rect 31205 28608 31217 28611
rect 28868 28580 31217 28608
rect 28868 28568 28874 28580
rect 31205 28577 31217 28580
rect 31251 28577 31263 28611
rect 31205 28571 31263 28577
rect 31297 28611 31355 28617
rect 31297 28577 31309 28611
rect 31343 28608 31355 28611
rect 32030 28608 32036 28620
rect 31343 28580 32036 28608
rect 31343 28577 31355 28580
rect 31297 28571 31355 28577
rect 23799 28512 25176 28540
rect 25225 28543 25283 28549
rect 23799 28509 23811 28512
rect 23753 28503 23811 28509
rect 25225 28509 25237 28543
rect 25271 28540 25283 28543
rect 25774 28540 25780 28552
rect 25271 28512 25780 28540
rect 25271 28509 25283 28512
rect 25225 28503 25283 28509
rect 23658 28432 23664 28484
rect 23716 28432 23722 28484
rect 23293 28407 23351 28413
rect 23293 28373 23305 28407
rect 23339 28373 23351 28407
rect 23293 28367 23351 28373
rect 23382 28364 23388 28416
rect 23440 28404 23446 28416
rect 25240 28404 25268 28503
rect 25774 28500 25780 28512
rect 25832 28540 25838 28552
rect 25832 28512 27568 28540
rect 25832 28500 25838 28512
rect 25869 28475 25927 28481
rect 25869 28441 25881 28475
rect 25915 28472 25927 28475
rect 26050 28472 26056 28484
rect 25915 28444 26056 28472
rect 25915 28441 25927 28444
rect 25869 28435 25927 28441
rect 26050 28432 26056 28444
rect 26108 28432 26114 28484
rect 23440 28376 25268 28404
rect 23440 28364 23446 28376
rect 25406 28364 25412 28416
rect 25464 28404 25470 28416
rect 25961 28407 26019 28413
rect 25961 28404 25973 28407
rect 25464 28376 25973 28404
rect 25464 28364 25470 28376
rect 25961 28373 25973 28376
rect 26007 28373 26019 28407
rect 27540 28404 27568 28512
rect 27614 28500 27620 28552
rect 27672 28500 27678 28552
rect 28626 28500 28632 28552
rect 28684 28500 28690 28552
rect 31220 28540 31248 28571
rect 32030 28568 32036 28580
rect 32088 28568 32094 28620
rect 31938 28540 31944 28552
rect 31220 28512 31944 28540
rect 31938 28500 31944 28512
rect 31996 28500 32002 28552
rect 28626 28404 28632 28416
rect 27540 28376 28632 28404
rect 25961 28367 26019 28373
rect 28626 28364 28632 28376
rect 28684 28364 28690 28416
rect 29270 28364 29276 28416
rect 29328 28364 29334 28416
rect 29822 28364 29828 28416
rect 29880 28404 29886 28416
rect 31113 28407 31171 28413
rect 31113 28404 31125 28407
rect 29880 28376 31125 28404
rect 29880 28364 29886 28376
rect 31113 28373 31125 28376
rect 31159 28373 31171 28407
rect 31113 28367 31171 28373
rect 1104 28314 36800 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 36800 28314
rect 1104 28240 36800 28262
rect 4985 28203 5043 28209
rect 4985 28169 4997 28203
rect 5031 28200 5043 28203
rect 5350 28200 5356 28212
rect 5031 28172 5356 28200
rect 5031 28169 5043 28172
rect 4985 28163 5043 28169
rect 5350 28160 5356 28172
rect 5408 28160 5414 28212
rect 9766 28160 9772 28212
rect 9824 28160 9830 28212
rect 12526 28160 12532 28212
rect 12584 28160 12590 28212
rect 12897 28203 12955 28209
rect 12897 28169 12909 28203
rect 12943 28200 12955 28203
rect 14366 28200 14372 28212
rect 12943 28172 14372 28200
rect 12943 28169 12955 28172
rect 12897 28163 12955 28169
rect 14366 28160 14372 28172
rect 14424 28160 14430 28212
rect 16114 28160 16120 28212
rect 16172 28200 16178 28212
rect 16209 28203 16267 28209
rect 16209 28200 16221 28203
rect 16172 28172 16221 28200
rect 16172 28160 16178 28172
rect 16209 28169 16221 28172
rect 16255 28169 16267 28203
rect 19705 28203 19763 28209
rect 19705 28200 19717 28203
rect 16209 28163 16267 28169
rect 16684 28172 19717 28200
rect 8656 28135 8714 28141
rect 8656 28101 8668 28135
rect 8702 28132 8714 28135
rect 8938 28132 8944 28144
rect 8702 28104 8944 28132
rect 8702 28101 8714 28104
rect 8656 28095 8714 28101
rect 8938 28092 8944 28104
rect 8996 28092 9002 28144
rect 9306 28092 9312 28144
rect 9364 28132 9370 28144
rect 16482 28132 16488 28144
rect 9364 28104 13216 28132
rect 9364 28092 9370 28104
rect 3878 28073 3884 28076
rect 3872 28027 3884 28073
rect 3878 28024 3884 28027
rect 3936 28024 3942 28076
rect 8386 28024 8392 28076
rect 8444 28024 8450 28076
rect 12894 28024 12900 28076
rect 12952 28064 12958 28076
rect 12989 28067 13047 28073
rect 12989 28064 13001 28067
rect 12952 28036 13001 28064
rect 12952 28024 12958 28036
rect 12989 28033 13001 28036
rect 13035 28033 13047 28067
rect 12989 28027 13047 28033
rect 3050 27956 3056 28008
rect 3108 27996 3114 28008
rect 13188 28005 13216 28104
rect 15580 28104 16488 28132
rect 13357 28067 13415 28073
rect 13357 28033 13369 28067
rect 13403 28064 13415 28067
rect 13403 28036 13768 28064
rect 13403 28033 13415 28036
rect 13357 28027 13415 28033
rect 3605 27999 3663 28005
rect 3605 27996 3617 27999
rect 3108 27968 3617 27996
rect 3108 27956 3114 27968
rect 3605 27965 3617 27968
rect 3651 27965 3663 27999
rect 3605 27959 3663 27965
rect 13173 27999 13231 28005
rect 13173 27965 13185 27999
rect 13219 27996 13231 27999
rect 13541 27999 13599 28005
rect 13219 27968 13492 27996
rect 13219 27965 13231 27968
rect 13173 27959 13231 27965
rect 13464 27860 13492 27968
rect 13541 27965 13553 27999
rect 13587 27965 13599 27999
rect 13740 27996 13768 28036
rect 14274 28024 14280 28076
rect 14332 28024 14338 28076
rect 14366 28024 14372 28076
rect 14424 28073 14430 28076
rect 14424 28067 14452 28073
rect 14440 28033 14452 28067
rect 14424 28027 14452 28033
rect 14424 28024 14430 28027
rect 14090 27996 14096 28008
rect 13740 27968 14096 27996
rect 13541 27959 13599 27965
rect 13556 27928 13584 27959
rect 14090 27956 14096 27968
rect 14148 27956 14154 28008
rect 14550 27956 14556 28008
rect 14608 27996 14614 28008
rect 15580 27996 15608 28104
rect 16482 28092 16488 28104
rect 16540 28092 16546 28144
rect 15657 28067 15715 28073
rect 15657 28033 15669 28067
rect 15703 28064 15715 28067
rect 16117 28067 16175 28073
rect 15703 28036 15792 28064
rect 15703 28033 15715 28036
rect 15657 28027 15715 28033
rect 14608 27968 15608 27996
rect 14608 27956 14614 27968
rect 13906 27928 13912 27940
rect 13556 27900 13912 27928
rect 13906 27888 13912 27900
rect 13964 27888 13970 27940
rect 13998 27888 14004 27940
rect 14056 27888 14062 27940
rect 15764 27937 15792 28036
rect 16117 28033 16129 28067
rect 16163 28064 16175 28067
rect 16574 28064 16580 28076
rect 16163 28036 16580 28064
rect 16163 28033 16175 28036
rect 16117 28027 16175 28033
rect 16574 28024 16580 28036
rect 16632 28024 16638 28076
rect 16393 27999 16451 28005
rect 16393 27965 16405 27999
rect 16439 27996 16451 27999
rect 16684 27996 16712 28172
rect 19705 28169 19717 28172
rect 19751 28169 19763 28203
rect 19705 28163 19763 28169
rect 20438 28160 20444 28212
rect 20496 28160 20502 28212
rect 20990 28160 20996 28212
rect 21048 28160 21054 28212
rect 23382 28200 23388 28212
rect 21468 28172 23388 28200
rect 16853 28067 16911 28073
rect 16853 28033 16865 28067
rect 16899 28064 16911 28067
rect 16942 28064 16948 28076
rect 16899 28036 16948 28064
rect 16899 28033 16911 28036
rect 16853 28027 16911 28033
rect 16942 28024 16948 28036
rect 17000 28024 17006 28076
rect 17770 28024 17776 28076
rect 17828 28024 17834 28076
rect 17862 28024 17868 28076
rect 17920 28073 17926 28076
rect 17920 28067 17948 28073
rect 17936 28033 17948 28067
rect 17920 28027 17948 28033
rect 17920 28024 17926 28027
rect 18046 28024 18052 28076
rect 18104 28024 18110 28076
rect 18877 28067 18935 28073
rect 18877 28033 18889 28067
rect 18923 28033 18935 28067
rect 18877 28027 18935 28033
rect 16439 27968 16712 27996
rect 17037 27999 17095 28005
rect 16439 27965 16451 27968
rect 16393 27959 16451 27965
rect 17037 27965 17049 27999
rect 17083 27996 17095 27999
rect 17126 27996 17132 28008
rect 17083 27968 17132 27996
rect 17083 27965 17095 27968
rect 17037 27959 17095 27965
rect 15749 27931 15807 27937
rect 14936 27900 15608 27928
rect 14936 27860 14964 27900
rect 13464 27832 14964 27860
rect 15194 27820 15200 27872
rect 15252 27820 15258 27872
rect 15470 27820 15476 27872
rect 15528 27820 15534 27872
rect 15580 27860 15608 27900
rect 15749 27897 15761 27931
rect 15795 27897 15807 27931
rect 15749 27891 15807 27897
rect 16408 27860 16436 27959
rect 17126 27956 17132 27968
rect 17184 27956 17190 28008
rect 17494 27956 17500 28008
rect 17552 27956 17558 28008
rect 18230 27956 18236 28008
rect 18288 27996 18294 28008
rect 18892 27996 18920 28027
rect 19334 28024 19340 28076
rect 19392 28024 19398 28076
rect 19521 28067 19579 28073
rect 19521 28033 19533 28067
rect 19567 28064 19579 28067
rect 20162 28064 20168 28076
rect 19567 28036 20168 28064
rect 19567 28033 19579 28036
rect 19521 28027 19579 28033
rect 20162 28024 20168 28036
rect 20220 28024 20226 28076
rect 20346 28024 20352 28076
rect 20404 28024 20410 28076
rect 20809 28067 20867 28073
rect 20809 28033 20821 28067
rect 20855 28064 20867 28067
rect 21468 28064 21496 28172
rect 23382 28160 23388 28172
rect 23440 28160 23446 28212
rect 24486 28200 24492 28212
rect 23492 28172 24492 28200
rect 21726 28092 21732 28144
rect 21784 28132 21790 28144
rect 22066 28135 22124 28141
rect 22066 28132 22078 28135
rect 21784 28104 22078 28132
rect 21784 28092 21790 28104
rect 22066 28101 22078 28104
rect 22112 28101 22124 28135
rect 22066 28095 22124 28101
rect 20855 28036 21496 28064
rect 20855 28033 20867 28036
rect 20809 28027 20867 28033
rect 21542 28024 21548 28076
rect 21600 28024 21606 28076
rect 23492 28073 23520 28172
rect 24486 28160 24492 28172
rect 24544 28160 24550 28212
rect 24946 28160 24952 28212
rect 25004 28200 25010 28212
rect 25004 28172 25176 28200
rect 25004 28160 25010 28172
rect 25148 28132 25176 28172
rect 26234 28160 26240 28212
rect 26292 28200 26298 28212
rect 27157 28203 27215 28209
rect 27157 28200 27169 28203
rect 26292 28172 27169 28200
rect 26292 28160 26298 28172
rect 27157 28169 27169 28172
rect 27203 28169 27215 28203
rect 27157 28163 27215 28169
rect 27065 28135 27123 28141
rect 27065 28132 27077 28135
rect 25148 28104 27077 28132
rect 27065 28101 27077 28104
rect 27111 28132 27123 28135
rect 27522 28132 27528 28144
rect 27111 28104 27528 28132
rect 27111 28101 27123 28104
rect 27065 28095 27123 28101
rect 27522 28092 27528 28104
rect 27580 28092 27586 28144
rect 27614 28092 27620 28144
rect 27672 28132 27678 28144
rect 28721 28135 28779 28141
rect 28721 28132 28733 28135
rect 27672 28104 28733 28132
rect 27672 28092 27678 28104
rect 28721 28101 28733 28104
rect 28767 28132 28779 28135
rect 28902 28132 28908 28144
rect 28767 28104 28908 28132
rect 28767 28101 28779 28104
rect 28721 28095 28779 28101
rect 28902 28092 28908 28104
rect 28960 28092 28966 28144
rect 23477 28067 23535 28073
rect 23477 28033 23489 28067
rect 23523 28033 23535 28067
rect 23477 28027 23535 28033
rect 24394 28024 24400 28076
rect 24452 28024 24458 28076
rect 24578 28073 24584 28076
rect 24535 28067 24584 28073
rect 24535 28033 24547 28067
rect 24581 28033 24584 28067
rect 24535 28027 24584 28033
rect 24578 28024 24584 28027
rect 24636 28024 24642 28076
rect 25676 28067 25734 28073
rect 25676 28033 25688 28067
rect 25722 28064 25734 28067
rect 25958 28064 25964 28076
rect 25722 28036 25964 28064
rect 25722 28033 25734 28036
rect 25676 28027 25734 28033
rect 25958 28024 25964 28036
rect 26016 28024 26022 28076
rect 21821 27999 21879 28005
rect 18288 27968 19196 27996
rect 18288 27956 18294 27968
rect 16482 27888 16488 27940
rect 16540 27928 16546 27940
rect 19168 27937 19196 27968
rect 21821 27965 21833 27999
rect 21867 27965 21879 27999
rect 21821 27959 21879 27965
rect 19153 27931 19211 27937
rect 16540 27900 17632 27928
rect 16540 27888 16546 27900
rect 15580 27832 16436 27860
rect 16666 27820 16672 27872
rect 16724 27860 16730 27872
rect 17494 27860 17500 27872
rect 16724 27832 17500 27860
rect 16724 27820 16730 27832
rect 17494 27820 17500 27832
rect 17552 27820 17558 27872
rect 17604 27860 17632 27900
rect 19153 27897 19165 27931
rect 19199 27897 19211 27931
rect 19153 27891 19211 27897
rect 19978 27888 19984 27940
rect 20036 27928 20042 27940
rect 20806 27928 20812 27940
rect 20036 27900 20812 27928
rect 20036 27888 20042 27900
rect 20806 27888 20812 27900
rect 20864 27888 20870 27940
rect 21361 27931 21419 27937
rect 21361 27897 21373 27931
rect 21407 27928 21419 27931
rect 21634 27928 21640 27940
rect 21407 27900 21640 27928
rect 21407 27897 21419 27900
rect 21361 27891 21419 27897
rect 21634 27888 21640 27900
rect 21692 27888 21698 27940
rect 21726 27888 21732 27940
rect 21784 27928 21790 27940
rect 21836 27928 21864 27959
rect 23658 27956 23664 28008
rect 23716 27956 23722 28008
rect 24673 27999 24731 28005
rect 24673 27965 24685 27999
rect 24719 27996 24731 27999
rect 24854 27996 24860 28008
rect 24719 27968 24860 27996
rect 24719 27965 24731 27968
rect 24673 27959 24731 27965
rect 24854 27956 24860 27968
rect 24912 27956 24918 28008
rect 25406 27996 25412 28008
rect 25056 27968 25412 27996
rect 21784 27900 21864 27928
rect 21784 27888 21790 27900
rect 23842 27888 23848 27940
rect 23900 27928 23906 27940
rect 24121 27931 24179 27937
rect 24121 27928 24133 27931
rect 23900 27900 24133 27928
rect 23900 27888 23906 27900
rect 24121 27897 24133 27900
rect 24167 27928 24179 27931
rect 24210 27928 24216 27940
rect 24167 27900 24216 27928
rect 24167 27897 24179 27900
rect 24121 27891 24179 27897
rect 24210 27888 24216 27900
rect 24268 27888 24274 27940
rect 18138 27860 18144 27872
rect 17604 27832 18144 27860
rect 18138 27820 18144 27832
rect 18196 27820 18202 27872
rect 18690 27820 18696 27872
rect 18748 27820 18754 27872
rect 18966 27820 18972 27872
rect 19024 27820 19030 27872
rect 20714 27820 20720 27872
rect 20772 27860 20778 27872
rect 23201 27863 23259 27869
rect 23201 27860 23213 27863
rect 20772 27832 23213 27860
rect 20772 27820 20778 27832
rect 23201 27829 23213 27832
rect 23247 27829 23259 27863
rect 23201 27823 23259 27829
rect 24026 27820 24032 27872
rect 24084 27860 24090 27872
rect 24854 27860 24860 27872
rect 24084 27832 24860 27860
rect 24084 27820 24090 27832
rect 24854 27820 24860 27832
rect 24912 27860 24918 27872
rect 25056 27860 25084 27968
rect 25406 27956 25412 27968
rect 25464 27956 25470 28008
rect 28810 27956 28816 28008
rect 28868 27956 28874 28008
rect 28905 27999 28963 28005
rect 28905 27965 28917 27999
rect 28951 27965 28963 27999
rect 28905 27959 28963 27965
rect 28626 27888 28632 27940
rect 28684 27928 28690 27940
rect 28920 27928 28948 27959
rect 28684 27900 28948 27928
rect 28684 27888 28690 27900
rect 24912 27832 25084 27860
rect 24912 27820 24918 27832
rect 25130 27820 25136 27872
rect 25188 27860 25194 27872
rect 25317 27863 25375 27869
rect 25317 27860 25329 27863
rect 25188 27832 25329 27860
rect 25188 27820 25194 27832
rect 25317 27829 25329 27832
rect 25363 27829 25375 27863
rect 25317 27823 25375 27829
rect 26786 27820 26792 27872
rect 26844 27820 26850 27872
rect 27890 27820 27896 27872
rect 27948 27860 27954 27872
rect 28353 27863 28411 27869
rect 28353 27860 28365 27863
rect 27948 27832 28365 27860
rect 27948 27820 27954 27832
rect 28353 27829 28365 27832
rect 28399 27829 28411 27863
rect 28353 27823 28411 27829
rect 1104 27770 36800 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 36800 27770
rect 1104 27696 36800 27718
rect 3878 27616 3884 27668
rect 3936 27616 3942 27668
rect 5736 27628 6592 27656
rect 4157 27591 4215 27597
rect 4157 27557 4169 27591
rect 4203 27557 4215 27591
rect 4157 27551 4215 27557
rect 5629 27591 5687 27597
rect 5629 27557 5641 27591
rect 5675 27588 5687 27591
rect 5736 27588 5764 27628
rect 5675 27560 5764 27588
rect 6564 27588 6592 27628
rect 10796 27628 11652 27656
rect 7282 27588 7288 27600
rect 6564 27560 7288 27588
rect 5675 27557 5687 27560
rect 5629 27551 5687 27557
rect 3510 27480 3516 27532
rect 3568 27480 3574 27532
rect 1397 27455 1455 27461
rect 1397 27421 1409 27455
rect 1443 27452 1455 27455
rect 3050 27452 3056 27464
rect 1443 27424 3056 27452
rect 1443 27421 1455 27424
rect 1397 27415 1455 27421
rect 3050 27412 3056 27424
rect 3108 27412 3114 27464
rect 3234 27412 3240 27464
rect 3292 27452 3298 27464
rect 3329 27455 3387 27461
rect 3329 27452 3341 27455
rect 3292 27424 3341 27452
rect 3292 27412 3298 27424
rect 3329 27421 3341 27424
rect 3375 27421 3387 27455
rect 3329 27415 3387 27421
rect 4065 27455 4123 27461
rect 4065 27421 4077 27455
rect 4111 27452 4123 27455
rect 4172 27452 4200 27551
rect 7282 27548 7288 27560
rect 7340 27548 7346 27600
rect 7374 27548 7380 27600
rect 7432 27548 7438 27600
rect 10796 27588 10824 27628
rect 9968 27560 10824 27588
rect 11624 27588 11652 27628
rect 13998 27616 14004 27668
rect 14056 27656 14062 27668
rect 16666 27656 16672 27668
rect 14056 27628 16672 27656
rect 14056 27616 14062 27628
rect 16666 27616 16672 27628
rect 16724 27616 16730 27668
rect 17126 27616 17132 27668
rect 17184 27656 17190 27668
rect 18598 27656 18604 27668
rect 17184 27628 18604 27656
rect 17184 27616 17190 27628
rect 18598 27616 18604 27628
rect 18656 27656 18662 27668
rect 18656 27628 18736 27656
rect 18656 27616 18662 27628
rect 14016 27588 14044 27616
rect 18708 27597 18736 27628
rect 19334 27616 19340 27668
rect 19392 27656 19398 27668
rect 21177 27659 21235 27665
rect 19392 27628 21128 27656
rect 19392 27616 19398 27628
rect 11624 27560 14044 27588
rect 18693 27591 18751 27597
rect 4798 27480 4804 27532
rect 4856 27480 4862 27532
rect 5169 27523 5227 27529
rect 5169 27520 5181 27523
rect 4908 27492 5181 27520
rect 4111 27424 4200 27452
rect 4525 27455 4583 27461
rect 4111 27421 4123 27424
rect 4065 27415 4123 27421
rect 4525 27421 4537 27455
rect 4571 27452 4583 27455
rect 4908 27452 4936 27492
rect 5169 27489 5181 27492
rect 5215 27520 5227 27523
rect 5350 27520 5356 27532
rect 5215 27492 5356 27520
rect 5215 27489 5227 27492
rect 5169 27483 5227 27489
rect 5350 27480 5356 27492
rect 5408 27480 5414 27532
rect 5902 27480 5908 27532
rect 5960 27480 5966 27532
rect 6086 27529 6092 27532
rect 6043 27523 6092 27529
rect 6043 27489 6055 27523
rect 6089 27489 6092 27523
rect 6043 27483 6092 27489
rect 6086 27480 6092 27483
rect 6144 27480 6150 27532
rect 6914 27480 6920 27532
rect 6972 27520 6978 27532
rect 7392 27520 7420 27548
rect 6972 27492 7420 27520
rect 7561 27523 7619 27529
rect 6972 27480 6978 27492
rect 7561 27489 7573 27523
rect 7607 27520 7619 27523
rect 9968 27520 9996 27560
rect 18693 27557 18705 27591
rect 18739 27557 18751 27591
rect 21100 27588 21128 27628
rect 21177 27625 21189 27659
rect 21223 27656 21235 27659
rect 21542 27656 21548 27668
rect 21223 27628 21548 27656
rect 21223 27625 21235 27628
rect 21177 27619 21235 27625
rect 21542 27616 21548 27628
rect 21600 27616 21606 27668
rect 21726 27656 21732 27668
rect 21652 27628 21732 27656
rect 21652 27588 21680 27628
rect 21726 27616 21732 27628
rect 21784 27656 21790 27668
rect 24026 27656 24032 27668
rect 21784 27628 24032 27656
rect 21784 27616 21790 27628
rect 24026 27616 24032 27628
rect 24084 27616 24090 27668
rect 24320 27628 26188 27656
rect 21100 27560 21680 27588
rect 18693 27551 18751 27557
rect 7607 27492 9996 27520
rect 7607 27489 7619 27492
rect 7561 27483 7619 27489
rect 10042 27480 10048 27532
rect 10100 27480 10106 27532
rect 10229 27523 10287 27529
rect 10229 27489 10241 27523
rect 10275 27520 10287 27523
rect 10410 27520 10416 27532
rect 10275 27492 10416 27520
rect 10275 27489 10287 27492
rect 10229 27483 10287 27489
rect 10410 27480 10416 27492
rect 10468 27480 10474 27532
rect 10686 27480 10692 27532
rect 10744 27480 10750 27532
rect 11054 27480 11060 27532
rect 11112 27529 11118 27532
rect 11112 27523 11140 27529
rect 11128 27489 11140 27523
rect 14550 27520 14556 27532
rect 11112 27483 11140 27489
rect 11808 27492 14556 27520
rect 11112 27480 11118 27483
rect 4571 27424 4936 27452
rect 4985 27455 5043 27461
rect 4571 27421 4583 27424
rect 4525 27415 4583 27421
rect 4985 27421 4997 27455
rect 5031 27452 5043 27455
rect 5074 27452 5080 27464
rect 5031 27424 5080 27452
rect 5031 27421 5043 27424
rect 4985 27415 5043 27421
rect 5074 27412 5080 27424
rect 5132 27412 5138 27464
rect 6178 27412 6184 27464
rect 6236 27412 6242 27464
rect 7006 27412 7012 27464
rect 7064 27452 7070 27464
rect 7101 27455 7159 27461
rect 7101 27452 7113 27455
rect 7064 27424 7113 27452
rect 7064 27412 7070 27424
rect 7101 27421 7113 27424
rect 7147 27421 7159 27455
rect 7101 27415 7159 27421
rect 7834 27412 7840 27464
rect 7892 27412 7898 27464
rect 7926 27412 7932 27464
rect 7984 27461 7990 27464
rect 7984 27455 8012 27461
rect 8000 27421 8012 27455
rect 7984 27415 8012 27421
rect 7984 27412 7990 27415
rect 8110 27412 8116 27464
rect 8168 27412 8174 27464
rect 10962 27412 10968 27464
rect 11020 27412 11026 27464
rect 11238 27412 11244 27464
rect 11296 27412 11302 27464
rect 1664 27387 1722 27393
rect 1664 27353 1676 27387
rect 1710 27384 1722 27387
rect 1762 27384 1768 27396
rect 1710 27356 1768 27384
rect 1710 27353 1722 27356
rect 1664 27347 1722 27353
rect 1762 27344 1768 27356
rect 1820 27344 1826 27396
rect 2792 27356 5212 27384
rect 2792 27325 2820 27356
rect 2777 27319 2835 27325
rect 2777 27285 2789 27319
rect 2823 27285 2835 27319
rect 2777 27279 2835 27285
rect 2866 27276 2872 27328
rect 2924 27276 2930 27328
rect 3252 27325 3280 27356
rect 3237 27319 3295 27325
rect 3237 27285 3249 27319
rect 3283 27285 3295 27319
rect 3237 27279 3295 27285
rect 4246 27276 4252 27328
rect 4304 27316 4310 27328
rect 4617 27319 4675 27325
rect 4617 27316 4629 27319
rect 4304 27288 4629 27316
rect 4304 27276 4310 27288
rect 4617 27285 4629 27288
rect 4663 27285 4675 27319
rect 5184 27316 5212 27356
rect 6748 27356 7144 27384
rect 6748 27316 6776 27356
rect 5184 27288 6776 27316
rect 4617 27279 4675 27285
rect 6822 27276 6828 27328
rect 6880 27276 6886 27328
rect 7116 27316 7144 27356
rect 8680 27356 10272 27384
rect 7650 27316 7656 27328
rect 7116 27288 7656 27316
rect 7650 27276 7656 27288
rect 7708 27316 7714 27328
rect 7926 27316 7932 27328
rect 7708 27288 7932 27316
rect 7708 27276 7714 27288
rect 7926 27276 7932 27288
rect 7984 27276 7990 27328
rect 8110 27276 8116 27328
rect 8168 27316 8174 27328
rect 8680 27316 8708 27356
rect 8168 27288 8708 27316
rect 8168 27276 8174 27288
rect 8754 27276 8760 27328
rect 8812 27276 8818 27328
rect 10244 27316 10272 27356
rect 11808 27316 11836 27492
rect 14550 27480 14556 27492
rect 14608 27480 14614 27532
rect 21821 27523 21879 27529
rect 21821 27489 21833 27523
rect 21867 27520 21879 27523
rect 23566 27520 23572 27532
rect 21867 27492 23572 27520
rect 21867 27489 21879 27492
rect 21821 27483 21879 27489
rect 14274 27412 14280 27464
rect 14332 27412 14338 27464
rect 15470 27461 15476 27464
rect 15197 27455 15255 27461
rect 15197 27421 15209 27455
rect 15243 27421 15255 27455
rect 15464 27452 15476 27461
rect 15431 27424 15476 27452
rect 15197 27415 15255 27421
rect 15464 27415 15476 27424
rect 13630 27344 13636 27396
rect 13688 27384 13694 27396
rect 15212 27384 15240 27415
rect 15470 27412 15476 27415
rect 15528 27412 15534 27464
rect 17313 27455 17371 27461
rect 17313 27421 17325 27455
rect 17359 27421 17371 27455
rect 17313 27415 17371 27421
rect 19245 27455 19303 27461
rect 19245 27421 19257 27455
rect 19291 27452 19303 27455
rect 21836 27452 21864 27483
rect 23566 27480 23572 27492
rect 23624 27480 23630 27532
rect 23658 27480 23664 27532
rect 23716 27520 23722 27532
rect 24320 27520 24348 27628
rect 24581 27523 24639 27529
rect 24581 27520 24593 27523
rect 23716 27492 24593 27520
rect 23716 27480 23722 27492
rect 24581 27489 24593 27492
rect 24627 27489 24639 27523
rect 24581 27483 24639 27489
rect 24946 27480 24952 27532
rect 25004 27520 25010 27532
rect 25498 27529 25504 27532
rect 25041 27523 25099 27529
rect 25041 27520 25053 27523
rect 25004 27492 25053 27520
rect 25004 27480 25010 27492
rect 25041 27489 25053 27492
rect 25087 27489 25099 27523
rect 25041 27483 25099 27489
rect 25455 27523 25504 27529
rect 25455 27489 25467 27523
rect 25501 27489 25504 27523
rect 25455 27483 25504 27489
rect 25498 27480 25504 27483
rect 25556 27480 25562 27532
rect 25593 27523 25651 27529
rect 25593 27489 25605 27523
rect 25639 27520 25651 27523
rect 25774 27520 25780 27532
rect 25639 27492 25780 27520
rect 25639 27489 25651 27492
rect 25593 27483 25651 27489
rect 25774 27480 25780 27492
rect 25832 27480 25838 27532
rect 19291 27424 21864 27452
rect 24397 27455 24455 27461
rect 19291 27421 19303 27424
rect 19245 27415 19303 27421
rect 24397 27421 24409 27455
rect 24443 27452 24455 27455
rect 24486 27452 24492 27464
rect 24443 27424 24492 27452
rect 24443 27421 24455 27424
rect 24397 27415 24455 27421
rect 17328 27384 17356 27415
rect 24486 27412 24492 27424
rect 24544 27412 24550 27464
rect 25314 27412 25320 27464
rect 25372 27412 25378 27464
rect 26160 27452 26188 27628
rect 28902 27616 28908 27668
rect 28960 27616 28966 27668
rect 27982 27548 27988 27600
rect 28040 27548 28046 27600
rect 28920 27588 28948 27616
rect 29365 27591 29423 27597
rect 29365 27588 29377 27591
rect 28920 27560 29377 27588
rect 29365 27557 29377 27560
rect 29411 27557 29423 27591
rect 31021 27591 31079 27597
rect 31021 27588 31033 27591
rect 29365 27551 29423 27557
rect 29472 27560 31033 27588
rect 26878 27480 26884 27532
rect 26936 27480 26942 27532
rect 28000 27520 28028 27548
rect 28000 27492 28120 27520
rect 26697 27455 26755 27461
rect 26697 27452 26709 27455
rect 26160 27424 26709 27452
rect 26697 27421 26709 27424
rect 26743 27452 26755 27455
rect 26786 27452 26792 27464
rect 26743 27424 26792 27452
rect 26743 27421 26755 27424
rect 26697 27415 26755 27421
rect 26786 27412 26792 27424
rect 26844 27412 26850 27464
rect 27890 27412 27896 27464
rect 27948 27412 27954 27464
rect 27982 27412 27988 27464
rect 28040 27412 28046 27464
rect 28092 27452 28120 27492
rect 29472 27452 29500 27560
rect 31021 27557 31033 27560
rect 31067 27557 31079 27591
rect 31021 27551 31079 27557
rect 31846 27548 31852 27600
rect 31904 27548 31910 27600
rect 30377 27523 30435 27529
rect 30377 27489 30389 27523
rect 30423 27520 30435 27523
rect 30926 27520 30932 27532
rect 30423 27492 30932 27520
rect 30423 27489 30435 27492
rect 30377 27483 30435 27489
rect 30926 27480 30932 27492
rect 30984 27520 30990 27532
rect 31205 27523 31263 27529
rect 31205 27520 31217 27523
rect 30984 27492 31217 27520
rect 30984 27480 30990 27492
rect 31205 27489 31217 27492
rect 31251 27489 31263 27523
rect 31205 27483 31263 27489
rect 31573 27455 31631 27461
rect 31573 27452 31585 27455
rect 28092 27424 29500 27452
rect 30760 27424 31585 27452
rect 17402 27384 17408 27396
rect 13688 27356 17408 27384
rect 13688 27344 13694 27356
rect 17402 27344 17408 27356
rect 17460 27344 17466 27396
rect 17586 27393 17592 27396
rect 17580 27347 17592 27393
rect 17586 27344 17592 27347
rect 17644 27344 17650 27396
rect 20714 27344 20720 27396
rect 20772 27384 20778 27396
rect 21545 27387 21603 27393
rect 21545 27384 21557 27387
rect 20772 27356 21557 27384
rect 20772 27344 20778 27356
rect 21545 27353 21557 27356
rect 21591 27353 21603 27387
rect 28230 27387 28288 27393
rect 28230 27384 28242 27387
rect 21545 27347 21603 27353
rect 27724 27356 28242 27384
rect 10244 27288 11836 27316
rect 11885 27319 11943 27325
rect 11885 27285 11897 27319
rect 11931 27316 11943 27319
rect 11974 27316 11980 27328
rect 11931 27288 11980 27316
rect 11931 27285 11943 27288
rect 11885 27279 11943 27285
rect 11974 27276 11980 27288
rect 12032 27276 12038 27328
rect 14090 27276 14096 27328
rect 14148 27276 14154 27328
rect 14734 27276 14740 27328
rect 14792 27316 14798 27328
rect 15562 27316 15568 27328
rect 14792 27288 15568 27316
rect 14792 27276 14798 27288
rect 15562 27276 15568 27288
rect 15620 27276 15626 27328
rect 16574 27276 16580 27328
rect 16632 27316 16638 27328
rect 17862 27316 17868 27328
rect 16632 27288 17868 27316
rect 16632 27276 16638 27288
rect 17862 27276 17868 27288
rect 17920 27276 17926 27328
rect 19426 27276 19432 27328
rect 19484 27276 19490 27328
rect 20622 27276 20628 27328
rect 20680 27316 20686 27328
rect 21637 27319 21695 27325
rect 21637 27316 21649 27319
rect 20680 27288 21649 27316
rect 20680 27276 20686 27288
rect 21637 27285 21649 27288
rect 21683 27285 21695 27319
rect 21637 27279 21695 27285
rect 24394 27276 24400 27328
rect 24452 27316 24458 27328
rect 25222 27316 25228 27328
rect 24452 27288 25228 27316
rect 24452 27276 24458 27288
rect 25222 27276 25228 27288
rect 25280 27276 25286 27328
rect 25866 27276 25872 27328
rect 25924 27316 25930 27328
rect 26237 27319 26295 27325
rect 26237 27316 26249 27319
rect 25924 27288 26249 27316
rect 25924 27276 25930 27288
rect 26237 27285 26249 27288
rect 26283 27285 26295 27319
rect 26237 27279 26295 27285
rect 26326 27276 26332 27328
rect 26384 27276 26390 27328
rect 26786 27276 26792 27328
rect 26844 27276 26850 27328
rect 27724 27325 27752 27356
rect 28230 27353 28242 27356
rect 28276 27353 28288 27387
rect 28230 27347 28288 27353
rect 30760 27328 30788 27424
rect 31573 27421 31585 27424
rect 31619 27421 31631 27455
rect 31573 27415 31631 27421
rect 35434 27412 35440 27464
rect 35492 27452 35498 27464
rect 36173 27455 36231 27461
rect 36173 27452 36185 27455
rect 35492 27424 36185 27452
rect 35492 27412 35498 27424
rect 36173 27421 36185 27424
rect 36219 27421 36231 27455
rect 36173 27415 36231 27421
rect 30837 27387 30895 27393
rect 30837 27353 30849 27387
rect 30883 27384 30895 27387
rect 31110 27384 31116 27396
rect 30883 27356 31116 27384
rect 30883 27353 30895 27356
rect 30837 27347 30895 27353
rect 31110 27344 31116 27356
rect 31168 27344 31174 27396
rect 31665 27387 31723 27393
rect 31665 27353 31677 27387
rect 31711 27384 31723 27387
rect 33318 27384 33324 27396
rect 31711 27356 33324 27384
rect 31711 27353 31723 27356
rect 31665 27347 31723 27353
rect 33318 27344 33324 27356
rect 33376 27344 33382 27396
rect 27709 27319 27767 27325
rect 27709 27285 27721 27319
rect 27755 27285 27767 27319
rect 27709 27279 27767 27285
rect 30650 27276 30656 27328
rect 30708 27276 30714 27328
rect 30742 27276 30748 27328
rect 30800 27276 30806 27328
rect 31481 27319 31539 27325
rect 31481 27285 31493 27319
rect 31527 27316 31539 27319
rect 31570 27316 31576 27328
rect 31527 27288 31576 27316
rect 31527 27285 31539 27288
rect 31481 27279 31539 27285
rect 31570 27276 31576 27288
rect 31628 27276 31634 27328
rect 36354 27276 36360 27328
rect 36412 27276 36418 27328
rect 1104 27226 36800 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 36800 27226
rect 1104 27152 36800 27174
rect 1762 27072 1768 27124
rect 1820 27072 1826 27124
rect 2777 27115 2835 27121
rect 2777 27081 2789 27115
rect 2823 27081 2835 27115
rect 2777 27075 2835 27081
rect 2792 27044 2820 27075
rect 10410 27072 10416 27124
rect 10468 27112 10474 27124
rect 11333 27115 11391 27121
rect 11333 27112 11345 27115
rect 10468 27084 11345 27112
rect 10468 27072 10474 27084
rect 11333 27081 11345 27084
rect 11379 27081 11391 27115
rect 11333 27075 11391 27081
rect 3298 27047 3356 27053
rect 3298 27044 3310 27047
rect 2792 27016 3310 27044
rect 3298 27013 3310 27016
rect 3344 27013 3356 27047
rect 11348 27044 11376 27075
rect 13998 27072 14004 27124
rect 14056 27112 14062 27124
rect 14458 27112 14464 27124
rect 14056 27084 14464 27112
rect 14056 27072 14062 27084
rect 14458 27072 14464 27084
rect 14516 27112 14522 27124
rect 15013 27115 15071 27121
rect 15013 27112 15025 27115
rect 14516 27084 15025 27112
rect 14516 27072 14522 27084
rect 15013 27081 15025 27084
rect 15059 27081 15071 27115
rect 15013 27075 15071 27081
rect 15102 27072 15108 27124
rect 15160 27112 15166 27124
rect 18230 27112 18236 27124
rect 15160 27084 18236 27112
rect 15160 27072 15166 27084
rect 18230 27072 18236 27084
rect 18288 27072 18294 27124
rect 18598 27072 18604 27124
rect 18656 27072 18662 27124
rect 23658 27072 23664 27124
rect 23716 27112 23722 27124
rect 24762 27112 24768 27124
rect 23716 27084 24768 27112
rect 23716 27072 23722 27084
rect 24762 27072 24768 27084
rect 24820 27072 24826 27124
rect 25958 27072 25964 27124
rect 26016 27072 26022 27124
rect 26326 27072 26332 27124
rect 26384 27072 26390 27124
rect 26418 27072 26424 27124
rect 26476 27072 26482 27124
rect 26878 27072 26884 27124
rect 26936 27112 26942 27124
rect 28626 27112 28632 27124
rect 26936 27084 28632 27112
rect 26936 27072 26942 27084
rect 28626 27072 28632 27084
rect 28684 27112 28690 27124
rect 30653 27115 30711 27121
rect 30653 27112 30665 27115
rect 28684 27084 30665 27112
rect 28684 27072 28690 27084
rect 30653 27081 30665 27084
rect 30699 27081 30711 27115
rect 30653 27075 30711 27081
rect 31110 27072 31116 27124
rect 31168 27072 31174 27124
rect 13900 27047 13958 27053
rect 11348 27016 11744 27044
rect 3298 27007 3356 27013
rect 1949 26979 2007 26985
rect 1949 26945 1961 26979
rect 1995 26976 2007 26979
rect 2866 26976 2872 26988
rect 1995 26948 2872 26976
rect 1995 26945 2007 26948
rect 1949 26939 2007 26945
rect 2866 26936 2872 26948
rect 2924 26936 2930 26988
rect 2958 26936 2964 26988
rect 3016 26936 3022 26988
rect 6825 26979 6883 26985
rect 6825 26976 6837 26979
rect 4448 26948 6837 26976
rect 3050 26868 3056 26920
rect 3108 26868 3114 26920
rect 4448 26849 4476 26948
rect 6825 26945 6837 26948
rect 6871 26976 6883 26979
rect 7006 26976 7012 26988
rect 6871 26948 7012 26976
rect 6871 26945 6883 26948
rect 6825 26939 6883 26945
rect 7006 26936 7012 26948
rect 7064 26936 7070 26988
rect 7558 26936 7564 26988
rect 7616 26936 7622 26988
rect 7650 26936 7656 26988
rect 7708 26985 7714 26988
rect 7708 26979 7736 26985
rect 7724 26945 7736 26979
rect 7708 26939 7736 26945
rect 7708 26936 7714 26939
rect 8478 26936 8484 26988
rect 8536 26976 8542 26988
rect 10226 26985 10232 26988
rect 9401 26979 9459 26985
rect 9401 26976 9413 26979
rect 8536 26948 9413 26976
rect 8536 26936 8542 26948
rect 9401 26945 9413 26948
rect 9447 26945 9459 26979
rect 10220 26976 10232 26985
rect 10187 26948 10232 26976
rect 9401 26939 9459 26945
rect 10220 26939 10232 26948
rect 10226 26936 10232 26939
rect 10284 26936 10290 26988
rect 11238 26936 11244 26988
rect 11296 26976 11302 26988
rect 11716 26985 11744 27016
rect 13900 27013 13912 27047
rect 13946 27044 13958 27047
rect 14090 27044 14096 27056
rect 13946 27016 14096 27044
rect 13946 27013 13958 27016
rect 13900 27007 13958 27013
rect 14090 27004 14096 27016
rect 14148 27004 14154 27056
rect 18966 27044 18972 27056
rect 17328 27016 18972 27044
rect 11517 26979 11575 26985
rect 11517 26976 11529 26979
rect 11296 26948 11529 26976
rect 11296 26936 11302 26948
rect 11517 26945 11529 26948
rect 11563 26945 11575 26979
rect 11517 26939 11575 26945
rect 11701 26979 11759 26985
rect 11701 26945 11713 26979
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 12434 26936 12440 26988
rect 12492 26936 12498 26988
rect 15010 26936 15016 26988
rect 15068 26976 15074 26988
rect 17328 26985 17356 27016
rect 18966 27004 18972 27016
rect 19024 27004 19030 27056
rect 19702 27004 19708 27056
rect 19760 27044 19766 27056
rect 20533 27047 20591 27053
rect 20533 27044 20545 27047
rect 19760 27016 20545 27044
rect 19760 27004 19766 27016
rect 20533 27013 20545 27016
rect 20579 27044 20591 27047
rect 20622 27044 20628 27056
rect 20579 27016 20628 27044
rect 20579 27013 20591 27016
rect 20533 27007 20591 27013
rect 20622 27004 20628 27016
rect 20680 27044 20686 27056
rect 20993 27047 21051 27053
rect 20993 27044 21005 27047
rect 20680 27016 21005 27044
rect 20680 27004 20686 27016
rect 20993 27013 21005 27016
rect 21039 27013 21051 27047
rect 20993 27007 21051 27013
rect 22830 27004 22836 27056
rect 22888 27044 22894 27056
rect 26344 27044 26372 27072
rect 22888 27016 23241 27044
rect 22888 27004 22894 27016
rect 17313 26979 17371 26985
rect 17313 26976 17325 26979
rect 15068 26948 17325 26976
rect 15068 26936 15074 26948
rect 17313 26945 17325 26948
rect 17359 26945 17371 26979
rect 17313 26939 17371 26945
rect 17402 26936 17408 26988
rect 17460 26976 17466 26988
rect 17589 26979 17647 26985
rect 17589 26976 17601 26979
rect 17460 26948 17601 26976
rect 17460 26936 17466 26948
rect 17589 26945 17601 26948
rect 17635 26945 17647 26979
rect 17589 26939 17647 26945
rect 19886 26936 19892 26988
rect 19944 26936 19950 26988
rect 20717 26979 20775 26985
rect 20717 26945 20729 26979
rect 20763 26976 20775 26979
rect 20806 26976 20812 26988
rect 20763 26948 20812 26976
rect 20763 26945 20775 26948
rect 20717 26939 20775 26945
rect 20806 26936 20812 26948
rect 20864 26936 20870 26988
rect 22738 26936 22744 26988
rect 22796 26976 22802 26988
rect 23213 26985 23241 27016
rect 26160 27016 26372 27044
rect 22925 26979 22983 26985
rect 22925 26976 22937 26979
rect 22796 26948 22937 26976
rect 22796 26936 22802 26948
rect 22925 26945 22937 26948
rect 22971 26945 22983 26979
rect 22925 26939 22983 26945
rect 23109 26979 23167 26985
rect 23109 26945 23121 26979
rect 23155 26945 23167 26979
rect 23109 26939 23167 26945
rect 23201 26979 23259 26985
rect 23201 26945 23213 26979
rect 23247 26945 23259 26979
rect 23201 26939 23259 26945
rect 6641 26911 6699 26917
rect 6641 26877 6653 26911
rect 6687 26908 6699 26911
rect 6914 26908 6920 26920
rect 6687 26880 6920 26908
rect 6687 26877 6699 26880
rect 6641 26871 6699 26877
rect 6914 26868 6920 26880
rect 6972 26868 6978 26920
rect 7837 26911 7895 26917
rect 7837 26908 7849 26911
rect 7024 26880 7849 26908
rect 4433 26843 4491 26849
rect 4433 26809 4445 26843
rect 4479 26840 4491 26843
rect 4614 26840 4620 26852
rect 4479 26812 4620 26840
rect 4479 26809 4491 26812
rect 4433 26803 4491 26809
rect 4614 26800 4620 26812
rect 4672 26800 4678 26852
rect 6178 26800 6184 26852
rect 6236 26840 6242 26852
rect 7024 26840 7052 26880
rect 7837 26877 7849 26880
rect 7883 26877 7895 26911
rect 7837 26871 7895 26877
rect 9953 26911 10011 26917
rect 9953 26877 9965 26911
rect 9999 26877 10011 26911
rect 9953 26871 10011 26877
rect 6236 26812 7052 26840
rect 6236 26800 6242 26812
rect 7282 26800 7288 26852
rect 7340 26800 7346 26852
rect 7650 26732 7656 26784
rect 7708 26772 7714 26784
rect 8481 26775 8539 26781
rect 8481 26772 8493 26775
rect 7708 26744 8493 26772
rect 7708 26732 7714 26744
rect 8481 26741 8493 26744
rect 8527 26741 8539 26775
rect 8481 26735 8539 26741
rect 9490 26732 9496 26784
rect 9548 26732 9554 26784
rect 9968 26772 9996 26871
rect 11330 26868 11336 26920
rect 11388 26908 11394 26920
rect 13630 26908 13636 26920
rect 11388 26880 13636 26908
rect 11388 26868 11394 26880
rect 13630 26868 13636 26880
rect 13688 26868 13694 26920
rect 17678 26868 17684 26920
rect 17736 26908 17742 26920
rect 18693 26911 18751 26917
rect 18693 26908 18705 26911
rect 17736 26880 18705 26908
rect 17736 26868 17742 26880
rect 18693 26877 18705 26880
rect 18739 26877 18751 26911
rect 18693 26871 18751 26877
rect 18785 26911 18843 26917
rect 18785 26877 18797 26911
rect 18831 26908 18843 26911
rect 19426 26908 19432 26920
rect 18831 26880 19432 26908
rect 18831 26877 18843 26880
rect 18785 26871 18843 26877
rect 10962 26800 10968 26852
rect 11020 26840 11026 26852
rect 11020 26812 12434 26840
rect 11020 26800 11026 26812
rect 11330 26772 11336 26784
rect 9968 26744 11336 26772
rect 11330 26732 11336 26744
rect 11388 26732 11394 26784
rect 11514 26732 11520 26784
rect 11572 26732 11578 26784
rect 12158 26732 12164 26784
rect 12216 26772 12222 26784
rect 12253 26775 12311 26781
rect 12253 26772 12265 26775
rect 12216 26744 12265 26772
rect 12216 26732 12222 26744
rect 12253 26741 12265 26744
rect 12299 26741 12311 26775
rect 12406 26772 12434 26812
rect 14642 26800 14648 26852
rect 14700 26840 14706 26852
rect 18800 26840 18828 26871
rect 19426 26868 19432 26880
rect 19484 26868 19490 26920
rect 14700 26812 18828 26840
rect 23124 26840 23152 26939
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 26160 26985 26188 27016
rect 32582 27004 32588 27056
rect 32640 27004 32646 27056
rect 25041 26979 25099 26985
rect 25041 26976 25053 26979
rect 24820 26948 25053 26976
rect 24820 26936 24826 26948
rect 25041 26945 25053 26948
rect 25087 26945 25099 26979
rect 25041 26939 25099 26945
rect 26145 26979 26203 26985
rect 26145 26945 26157 26979
rect 26191 26945 26203 26979
rect 26145 26939 26203 26945
rect 26329 26979 26387 26985
rect 26329 26945 26341 26979
rect 26375 26976 26387 26979
rect 26786 26976 26792 26988
rect 26375 26948 26792 26976
rect 26375 26945 26387 26948
rect 26329 26939 26387 26945
rect 25056 26908 25084 26939
rect 26344 26908 26372 26939
rect 26786 26936 26792 26948
rect 26844 26936 26850 26988
rect 28353 26979 28411 26985
rect 28353 26945 28365 26979
rect 28399 26976 28411 26979
rect 28810 26976 28816 26988
rect 28399 26948 28816 26976
rect 28399 26945 28411 26948
rect 28353 26939 28411 26945
rect 28810 26936 28816 26948
rect 28868 26976 28874 26988
rect 29641 26979 29699 26985
rect 29641 26976 29653 26979
rect 28868 26948 29653 26976
rect 28868 26936 28874 26948
rect 29641 26945 29653 26948
rect 29687 26976 29699 26979
rect 30190 26976 30196 26988
rect 29687 26948 30196 26976
rect 29687 26945 29699 26948
rect 29641 26939 29699 26945
rect 30190 26936 30196 26948
rect 30248 26936 30254 26988
rect 30834 26936 30840 26988
rect 30892 26976 30898 26988
rect 31021 26979 31079 26985
rect 31021 26976 31033 26979
rect 30892 26948 31033 26976
rect 30892 26936 30898 26948
rect 31021 26945 31033 26948
rect 31067 26945 31079 26979
rect 31021 26939 31079 26945
rect 31205 26979 31263 26985
rect 31205 26945 31217 26979
rect 31251 26976 31263 26979
rect 31294 26976 31300 26988
rect 31251 26948 31300 26976
rect 31251 26945 31263 26948
rect 31205 26939 31263 26945
rect 31294 26936 31300 26948
rect 31352 26936 31358 26988
rect 31662 26936 31668 26988
rect 31720 26976 31726 26988
rect 32125 26979 32183 26985
rect 32125 26976 32137 26979
rect 31720 26948 32137 26976
rect 31720 26936 31726 26948
rect 32125 26945 32137 26948
rect 32171 26945 32183 26979
rect 32125 26939 32183 26945
rect 32677 26979 32735 26985
rect 32677 26945 32689 26979
rect 32723 26945 32735 26979
rect 32677 26939 32735 26945
rect 25056 26880 26372 26908
rect 30469 26911 30527 26917
rect 30469 26877 30481 26911
rect 30515 26908 30527 26911
rect 30742 26908 30748 26920
rect 30515 26880 30748 26908
rect 30515 26877 30527 26880
rect 30469 26871 30527 26877
rect 30742 26868 30748 26880
rect 30800 26908 30806 26920
rect 30926 26908 30932 26920
rect 30800 26880 30932 26908
rect 30800 26868 30806 26880
rect 30926 26868 30932 26880
rect 30984 26868 30990 26920
rect 31846 26868 31852 26920
rect 31904 26908 31910 26920
rect 32692 26908 32720 26939
rect 33318 26936 33324 26988
rect 33376 26936 33382 26988
rect 33505 26979 33563 26985
rect 33505 26945 33517 26979
rect 33551 26945 33563 26979
rect 33505 26939 33563 26945
rect 31904 26880 32720 26908
rect 31904 26868 31910 26880
rect 32858 26868 32864 26920
rect 32916 26908 32922 26920
rect 33520 26908 33548 26939
rect 32916 26880 33548 26908
rect 32916 26868 32922 26880
rect 29086 26840 29092 26852
rect 23124 26812 29092 26840
rect 14700 26800 14706 26812
rect 29086 26800 29092 26812
rect 29144 26800 29150 26852
rect 29822 26800 29828 26852
rect 29880 26800 29886 26852
rect 15102 26772 15108 26784
rect 12406 26744 15108 26772
rect 12253 26735 12311 26741
rect 15102 26732 15108 26744
rect 15160 26732 15166 26784
rect 17770 26732 17776 26784
rect 17828 26772 17834 26784
rect 18233 26775 18291 26781
rect 18233 26772 18245 26775
rect 17828 26744 18245 26772
rect 17828 26732 17834 26744
rect 18233 26741 18245 26744
rect 18279 26741 18291 26775
rect 18233 26735 18291 26741
rect 19610 26732 19616 26784
rect 19668 26772 19674 26784
rect 19705 26775 19763 26781
rect 19705 26772 19717 26775
rect 19668 26744 19717 26772
rect 19668 26732 19674 26744
rect 19705 26741 19717 26744
rect 19751 26741 19763 26775
rect 19705 26735 19763 26741
rect 20990 26732 20996 26784
rect 21048 26772 21054 26784
rect 21085 26775 21143 26781
rect 21085 26772 21097 26775
rect 21048 26744 21097 26772
rect 21048 26732 21054 26744
rect 21085 26741 21097 26744
rect 21131 26741 21143 26775
rect 21085 26735 21143 26741
rect 22741 26775 22799 26781
rect 22741 26741 22753 26775
rect 22787 26772 22799 26775
rect 23474 26772 23480 26784
rect 22787 26744 23480 26772
rect 22787 26741 22799 26744
rect 22741 26735 22799 26741
rect 23474 26732 23480 26744
rect 23532 26732 23538 26784
rect 25038 26732 25044 26784
rect 25096 26772 25102 26784
rect 25133 26775 25191 26781
rect 25133 26772 25145 26775
rect 25096 26744 25145 26772
rect 25096 26732 25102 26744
rect 25133 26741 25145 26744
rect 25179 26741 25191 26775
rect 25133 26735 25191 26741
rect 28074 26732 28080 26784
rect 28132 26772 28138 26784
rect 28442 26772 28448 26784
rect 28132 26744 28448 26772
rect 28132 26732 28138 26744
rect 28442 26732 28448 26744
rect 28500 26732 28506 26784
rect 1104 26682 36800 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 36800 26682
rect 1104 26608 36800 26630
rect 2958 26528 2964 26580
rect 3016 26568 3022 26580
rect 4157 26571 4215 26577
rect 4157 26568 4169 26571
rect 3016 26540 4169 26568
rect 3016 26528 3022 26540
rect 4157 26537 4169 26540
rect 4203 26537 4215 26571
rect 4157 26531 4215 26537
rect 10137 26571 10195 26577
rect 10137 26537 10149 26571
rect 10183 26568 10195 26571
rect 10226 26568 10232 26580
rect 10183 26540 10232 26568
rect 10183 26537 10195 26540
rect 10137 26531 10195 26537
rect 10226 26528 10232 26540
rect 10284 26528 10290 26580
rect 12894 26528 12900 26580
rect 12952 26568 12958 26580
rect 13633 26571 13691 26577
rect 13633 26568 13645 26571
rect 12952 26540 13645 26568
rect 12952 26528 12958 26540
rect 13633 26537 13645 26540
rect 13679 26537 13691 26571
rect 13633 26531 13691 26537
rect 14093 26571 14151 26577
rect 14093 26537 14105 26571
rect 14139 26568 14151 26571
rect 14274 26568 14280 26580
rect 14139 26540 14280 26568
rect 14139 26537 14151 26540
rect 14093 26531 14151 26537
rect 14274 26528 14280 26540
rect 14332 26528 14338 26580
rect 16114 26528 16120 26580
rect 16172 26568 16178 26580
rect 17405 26571 17463 26577
rect 17405 26568 17417 26571
rect 16172 26540 17417 26568
rect 16172 26528 16178 26540
rect 17405 26537 17417 26540
rect 17451 26537 17463 26571
rect 17405 26531 17463 26537
rect 17586 26528 17592 26580
rect 17644 26528 17650 26580
rect 21266 26528 21272 26580
rect 21324 26568 21330 26580
rect 22370 26568 22376 26580
rect 21324 26540 22376 26568
rect 21324 26528 21330 26540
rect 22370 26528 22376 26540
rect 22428 26528 22434 26580
rect 32398 26528 32404 26580
rect 32456 26528 32462 26580
rect 7282 26460 7288 26512
rect 7340 26500 7346 26512
rect 7926 26500 7932 26512
rect 7340 26472 7932 26500
rect 7340 26460 7346 26472
rect 7926 26460 7932 26472
rect 7984 26460 7990 26512
rect 10962 26500 10968 26512
rect 8956 26472 10968 26500
rect 4614 26432 4620 26444
rect 4540 26404 4620 26432
rect 4540 26373 4568 26404
rect 4614 26392 4620 26404
rect 4672 26392 4678 26444
rect 4798 26392 4804 26444
rect 4856 26392 4862 26444
rect 8570 26392 8576 26444
rect 8628 26432 8634 26444
rect 8956 26441 8984 26472
rect 10962 26460 10968 26472
rect 11020 26460 11026 26512
rect 22738 26500 22744 26512
rect 21468 26472 22744 26500
rect 8757 26435 8815 26441
rect 8757 26432 8769 26435
rect 8628 26404 8769 26432
rect 8628 26392 8634 26404
rect 8757 26401 8769 26404
rect 8803 26401 8815 26435
rect 8757 26395 8815 26401
rect 8941 26435 8999 26441
rect 8941 26401 8953 26435
rect 8987 26401 8999 26435
rect 11514 26432 11520 26444
rect 8941 26395 8999 26401
rect 10336 26404 11520 26432
rect 4525 26367 4583 26373
rect 4525 26333 4537 26367
rect 4571 26333 4583 26367
rect 4816 26364 4844 26392
rect 4816 26336 9168 26364
rect 4525 26327 4583 26333
rect 4614 26256 4620 26308
rect 4672 26256 4678 26308
rect 8478 26256 8484 26308
rect 8536 26296 8542 26308
rect 8573 26299 8631 26305
rect 8573 26296 8585 26299
rect 8536 26268 8585 26296
rect 8536 26256 8542 26268
rect 8573 26265 8585 26268
rect 8619 26296 8631 26299
rect 9140 26296 9168 26336
rect 9214 26324 9220 26376
rect 9272 26324 9278 26376
rect 10137 26367 10195 26373
rect 10137 26333 10149 26367
rect 10183 26358 10195 26367
rect 10336 26364 10364 26404
rect 11514 26392 11520 26404
rect 11572 26392 11578 26444
rect 14642 26432 14648 26444
rect 14384 26404 14648 26432
rect 10244 26358 10364 26364
rect 10183 26336 10364 26358
rect 10413 26367 10471 26373
rect 10183 26333 10272 26336
rect 10137 26330 10272 26333
rect 10413 26333 10425 26367
rect 10459 26364 10471 26367
rect 11238 26364 11244 26376
rect 10459 26336 11244 26364
rect 10459 26333 10471 26336
rect 10137 26327 10195 26330
rect 10413 26327 10471 26333
rect 10428 26296 10456 26327
rect 11238 26324 11244 26336
rect 11296 26324 11302 26376
rect 11330 26324 11336 26376
rect 11388 26364 11394 26376
rect 11882 26364 11888 26376
rect 11388 26336 11888 26364
rect 11388 26324 11394 26336
rect 11882 26324 11888 26336
rect 11940 26324 11946 26376
rect 12158 26373 12164 26376
rect 12152 26364 12164 26373
rect 12119 26336 12164 26364
rect 12152 26327 12164 26336
rect 12158 26324 12164 26327
rect 12216 26324 12222 26376
rect 14384 26364 14412 26404
rect 14642 26392 14648 26404
rect 14700 26392 14706 26444
rect 17129 26435 17187 26441
rect 17129 26401 17141 26435
rect 17175 26432 17187 26435
rect 17310 26432 17316 26444
rect 17175 26404 17316 26432
rect 17175 26401 17187 26404
rect 17129 26395 17187 26401
rect 17310 26392 17316 26404
rect 17368 26392 17374 26444
rect 21468 26441 21496 26472
rect 22738 26460 22744 26472
rect 22796 26460 22802 26512
rect 31938 26500 31944 26512
rect 30300 26472 31944 26500
rect 21453 26435 21511 26441
rect 21453 26432 21465 26435
rect 21100 26404 21465 26432
rect 12406 26336 14412 26364
rect 8619 26268 9076 26296
rect 9140 26268 10456 26296
rect 11256 26296 11284 26324
rect 12406 26296 12434 26336
rect 14458 26324 14464 26376
rect 14516 26324 14522 26376
rect 17770 26324 17776 26376
rect 17828 26324 17834 26376
rect 19334 26324 19340 26376
rect 19392 26324 19398 26376
rect 19610 26373 19616 26376
rect 19604 26364 19616 26373
rect 19571 26336 19616 26364
rect 19604 26327 19616 26336
rect 19610 26324 19616 26327
rect 19668 26324 19674 26376
rect 21100 26373 21128 26404
rect 21453 26401 21465 26404
rect 21499 26401 21511 26435
rect 21453 26395 21511 26401
rect 21818 26392 21824 26444
rect 21876 26392 21882 26444
rect 23198 26392 23204 26444
rect 23256 26432 23262 26444
rect 23845 26435 23903 26441
rect 23845 26432 23857 26435
rect 23256 26404 23857 26432
rect 23256 26392 23262 26404
rect 23845 26401 23857 26404
rect 23891 26401 23903 26435
rect 25590 26432 25596 26444
rect 23845 26395 23903 26401
rect 24504 26404 25596 26432
rect 21085 26367 21143 26373
rect 21085 26364 21097 26367
rect 19720 26336 21097 26364
rect 11256 26268 12434 26296
rect 8619 26265 8631 26268
rect 8573 26259 8631 26265
rect 9048 26228 9076 26268
rect 13354 26256 13360 26308
rect 13412 26296 13418 26308
rect 13541 26299 13599 26305
rect 13541 26296 13553 26299
rect 13412 26268 13553 26296
rect 13412 26256 13418 26268
rect 13541 26265 13553 26268
rect 13587 26296 13599 26299
rect 14553 26299 14611 26305
rect 14553 26296 14565 26299
rect 13587 26268 14565 26296
rect 13587 26265 13599 26268
rect 13541 26259 13599 26265
rect 14553 26265 14565 26268
rect 14599 26265 14611 26299
rect 14553 26259 14611 26265
rect 16850 26256 16856 26308
rect 16908 26296 16914 26308
rect 16945 26299 17003 26305
rect 16945 26296 16957 26299
rect 16908 26268 16957 26296
rect 16908 26256 16914 26268
rect 16945 26265 16957 26268
rect 16991 26296 17003 26299
rect 17313 26299 17371 26305
rect 17313 26296 17325 26299
rect 16991 26268 17325 26296
rect 16991 26265 17003 26268
rect 16945 26259 17003 26265
rect 17313 26265 17325 26268
rect 17359 26296 17371 26299
rect 17678 26296 17684 26308
rect 17359 26268 17684 26296
rect 17359 26265 17371 26268
rect 17313 26259 17371 26265
rect 17678 26256 17684 26268
rect 17736 26256 17742 26308
rect 17862 26256 17868 26308
rect 17920 26296 17926 26308
rect 19720 26296 19748 26336
rect 21085 26333 21097 26336
rect 21131 26333 21143 26367
rect 21085 26327 21143 26333
rect 21358 26324 21364 26376
rect 21416 26324 21422 26376
rect 21910 26324 21916 26376
rect 21968 26324 21974 26376
rect 23385 26367 23443 26373
rect 23385 26364 23397 26367
rect 22572 26336 23397 26364
rect 17920 26268 19748 26296
rect 20901 26299 20959 26305
rect 17920 26256 17926 26268
rect 20901 26265 20913 26299
rect 20947 26296 20959 26299
rect 21174 26296 21180 26308
rect 20947 26268 21180 26296
rect 20947 26265 20959 26268
rect 20901 26259 20959 26265
rect 21174 26256 21180 26268
rect 21232 26256 21238 26308
rect 21542 26256 21548 26308
rect 21600 26296 21606 26308
rect 22097 26299 22155 26305
rect 22097 26296 22109 26299
rect 21600 26268 22109 26296
rect 21600 26256 21606 26268
rect 22097 26265 22109 26268
rect 22143 26265 22155 26299
rect 22097 26259 22155 26265
rect 22462 26256 22468 26308
rect 22520 26296 22526 26308
rect 22572 26305 22600 26336
rect 23385 26333 23397 26336
rect 23431 26333 23443 26367
rect 23385 26327 23443 26333
rect 23753 26367 23811 26373
rect 23753 26333 23765 26367
rect 23799 26364 23811 26367
rect 24504 26364 24532 26404
rect 25590 26392 25596 26404
rect 25648 26392 25654 26444
rect 30300 26441 30328 26472
rect 31938 26460 31944 26472
rect 31996 26500 32002 26512
rect 32858 26500 32864 26512
rect 31996 26472 32864 26500
rect 31996 26460 32002 26472
rect 32858 26460 32864 26472
rect 32916 26460 32922 26512
rect 30285 26435 30343 26441
rect 30285 26401 30297 26435
rect 30331 26401 30343 26435
rect 30285 26395 30343 26401
rect 30650 26392 30656 26444
rect 30708 26432 30714 26444
rect 31202 26432 31208 26444
rect 30708 26404 31208 26432
rect 30708 26392 30714 26404
rect 31202 26392 31208 26404
rect 31260 26432 31266 26444
rect 31662 26432 31668 26444
rect 31260 26404 31668 26432
rect 31260 26392 31266 26404
rect 31662 26392 31668 26404
rect 31720 26432 31726 26444
rect 33318 26432 33324 26444
rect 31720 26404 31984 26432
rect 31720 26392 31726 26404
rect 23799 26336 24532 26364
rect 23799 26333 23811 26336
rect 23753 26327 23811 26333
rect 24578 26324 24584 26376
rect 24636 26324 24642 26376
rect 28534 26324 28540 26376
rect 28592 26364 28598 26376
rect 30469 26367 30527 26373
rect 30469 26364 30481 26367
rect 28592 26336 30481 26364
rect 28592 26324 28598 26336
rect 30469 26333 30481 26336
rect 30515 26333 30527 26367
rect 30469 26327 30527 26333
rect 30929 26367 30987 26373
rect 30929 26333 30941 26367
rect 30975 26364 30987 26367
rect 31481 26367 31539 26373
rect 31481 26364 31493 26367
rect 30975 26336 31493 26364
rect 30975 26333 30987 26336
rect 30929 26327 30987 26333
rect 31481 26333 31493 26336
rect 31527 26333 31539 26367
rect 31481 26327 31539 26333
rect 22557 26299 22615 26305
rect 22557 26296 22569 26299
rect 22520 26268 22569 26296
rect 22520 26256 22526 26268
rect 22557 26265 22569 26268
rect 22603 26265 22615 26299
rect 22557 26259 22615 26265
rect 22922 26256 22928 26308
rect 22980 26296 22986 26308
rect 24029 26299 24087 26305
rect 24029 26296 24041 26299
rect 22980 26268 24041 26296
rect 22980 26256 22986 26268
rect 24029 26265 24041 26268
rect 24075 26265 24087 26299
rect 24029 26259 24087 26265
rect 30834 26256 30840 26308
rect 30892 26256 30898 26308
rect 31021 26299 31079 26305
rect 31021 26265 31033 26299
rect 31067 26296 31079 26299
rect 31294 26296 31300 26308
rect 31067 26268 31300 26296
rect 31067 26265 31079 26268
rect 31021 26259 31079 26265
rect 31294 26256 31300 26268
rect 31352 26256 31358 26308
rect 31496 26296 31524 26327
rect 31570 26324 31576 26376
rect 31628 26364 31634 26376
rect 31846 26364 31852 26376
rect 31628 26336 31852 26364
rect 31628 26324 31634 26336
rect 31846 26324 31852 26336
rect 31904 26324 31910 26376
rect 31956 26373 31984 26404
rect 32048 26404 33324 26432
rect 31941 26367 31999 26373
rect 31941 26333 31953 26367
rect 31987 26333 31999 26367
rect 31941 26327 31999 26333
rect 32048 26296 32076 26404
rect 33318 26392 33324 26404
rect 33376 26392 33382 26444
rect 32677 26367 32735 26373
rect 32677 26333 32689 26367
rect 32723 26364 32735 26367
rect 32858 26364 32864 26376
rect 32723 26336 32864 26364
rect 32723 26333 32735 26336
rect 32677 26327 32735 26333
rect 32858 26324 32864 26336
rect 32916 26324 32922 26376
rect 31496 26268 32076 26296
rect 10321 26231 10379 26237
rect 10321 26228 10333 26231
rect 9048 26200 10333 26228
rect 10321 26197 10333 26200
rect 10367 26197 10379 26231
rect 10321 26191 10379 26197
rect 13170 26188 13176 26240
rect 13228 26228 13234 26240
rect 13265 26231 13323 26237
rect 13265 26228 13277 26231
rect 13228 26200 13277 26228
rect 13228 26188 13234 26200
rect 13265 26197 13277 26200
rect 13311 26197 13323 26231
rect 13265 26191 13323 26197
rect 20714 26188 20720 26240
rect 20772 26188 20778 26240
rect 21266 26188 21272 26240
rect 21324 26188 21330 26240
rect 24394 26188 24400 26240
rect 24452 26188 24458 26240
rect 1104 26138 36800 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 36800 26138
rect 1104 26064 36800 26086
rect 2225 26027 2283 26033
rect 2225 25993 2237 26027
rect 2271 25993 2283 26027
rect 2225 25987 2283 25993
rect 2041 25891 2099 25897
rect 2041 25857 2053 25891
rect 2087 25888 2099 25891
rect 2240 25888 2268 25987
rect 6822 25984 6828 26036
rect 6880 25984 6886 26036
rect 9398 26024 9404 26036
rect 6932 25996 9404 26024
rect 2685 25959 2743 25965
rect 2685 25925 2697 25959
rect 2731 25956 2743 25959
rect 2774 25956 2780 25968
rect 2731 25928 2780 25956
rect 2731 25925 2743 25928
rect 2685 25919 2743 25925
rect 2774 25916 2780 25928
rect 2832 25916 2838 25968
rect 4982 25916 4988 25968
rect 5040 25956 5046 25968
rect 6932 25956 6960 25996
rect 9398 25984 9404 25996
rect 9456 25984 9462 26036
rect 12434 25984 12440 26036
rect 12492 25984 12498 26036
rect 12805 26027 12863 26033
rect 12805 25993 12817 26027
rect 12851 26024 12863 26027
rect 12986 26024 12992 26036
rect 12851 25996 12992 26024
rect 12851 25993 12863 25996
rect 12805 25987 12863 25993
rect 12986 25984 12992 25996
rect 13044 26024 13050 26036
rect 13538 26024 13544 26036
rect 13044 25996 13544 26024
rect 13044 25984 13050 25996
rect 13538 25984 13544 25996
rect 13596 25984 13602 26036
rect 17037 26027 17095 26033
rect 17037 25993 17049 26027
rect 17083 26024 17095 26027
rect 17310 26024 17316 26036
rect 17083 25996 17316 26024
rect 17083 25993 17095 25996
rect 17037 25987 17095 25993
rect 17310 25984 17316 25996
rect 17368 25984 17374 26036
rect 18690 25984 18696 26036
rect 18748 26024 18754 26036
rect 18969 26027 19027 26033
rect 18969 26024 18981 26027
rect 18748 25996 18981 26024
rect 18748 25984 18754 25996
rect 18969 25993 18981 25996
rect 19015 25993 19027 26027
rect 18969 25987 19027 25993
rect 19886 25984 19892 26036
rect 19944 25984 19950 26036
rect 20349 26027 20407 26033
rect 20349 25993 20361 26027
rect 20395 26024 20407 26027
rect 20714 26024 20720 26036
rect 20395 25996 20720 26024
rect 20395 25993 20407 25996
rect 20349 25987 20407 25993
rect 20714 25984 20720 25996
rect 20772 25984 20778 26036
rect 22738 25984 22744 26036
rect 22796 26024 22802 26036
rect 22925 26027 22983 26033
rect 22925 26024 22937 26027
rect 22796 25996 22937 26024
rect 22796 25984 22802 25996
rect 22925 25993 22937 25996
rect 22971 25993 22983 26027
rect 26510 26024 26516 26036
rect 22925 25987 22983 25993
rect 24044 25996 26516 26024
rect 8481 25959 8539 25965
rect 8481 25956 8493 25959
rect 5040 25928 6960 25956
rect 7944 25928 8493 25956
rect 5040 25916 5046 25928
rect 2087 25860 2268 25888
rect 2593 25891 2651 25897
rect 2087 25857 2099 25860
rect 2041 25851 2099 25857
rect 2593 25857 2605 25891
rect 2639 25888 2651 25891
rect 2866 25888 2872 25900
rect 2639 25860 2872 25888
rect 2639 25857 2651 25860
rect 2593 25851 2651 25857
rect 2866 25848 2872 25860
rect 2924 25848 2930 25900
rect 6362 25848 6368 25900
rect 6420 25888 6426 25900
rect 6733 25891 6791 25897
rect 6733 25888 6745 25891
rect 6420 25860 6745 25888
rect 6420 25848 6426 25860
rect 6733 25857 6745 25860
rect 6779 25857 6791 25891
rect 6733 25851 6791 25857
rect 7558 25848 7564 25900
rect 7616 25888 7622 25900
rect 7944 25897 7972 25928
rect 8481 25925 8493 25928
rect 8527 25956 8539 25959
rect 8527 25928 12020 25956
rect 8527 25925 8539 25928
rect 8481 25919 8539 25925
rect 7929 25891 7987 25897
rect 7929 25888 7941 25891
rect 7616 25860 7941 25888
rect 7616 25848 7622 25860
rect 7929 25857 7941 25860
rect 7975 25857 7987 25891
rect 7929 25851 7987 25857
rect 8202 25848 8208 25900
rect 8260 25888 8266 25900
rect 9122 25897 9128 25900
rect 8297 25891 8355 25897
rect 8297 25888 8309 25891
rect 8260 25860 8309 25888
rect 8260 25848 8266 25860
rect 8297 25857 8309 25860
rect 8343 25857 8355 25891
rect 8297 25851 8355 25857
rect 9116 25851 9128 25897
rect 9122 25848 9128 25851
rect 9180 25848 9186 25900
rect 9398 25848 9404 25900
rect 9456 25888 9462 25900
rect 9456 25860 10263 25888
rect 9456 25848 9462 25860
rect 2777 25823 2835 25829
rect 2777 25789 2789 25823
rect 2823 25820 2835 25823
rect 3142 25820 3148 25832
rect 2823 25792 3148 25820
rect 2823 25789 2835 25792
rect 2777 25783 2835 25789
rect 3142 25780 3148 25792
rect 3200 25780 3206 25832
rect 7009 25823 7067 25829
rect 7009 25789 7021 25823
rect 7055 25789 7067 25823
rect 7009 25783 7067 25789
rect 7024 25752 7052 25783
rect 7282 25780 7288 25832
rect 7340 25820 7346 25832
rect 7469 25823 7527 25829
rect 7469 25820 7481 25823
rect 7340 25792 7481 25820
rect 7340 25780 7346 25792
rect 7469 25789 7481 25792
rect 7515 25789 7527 25823
rect 7469 25783 7527 25789
rect 7837 25823 7895 25829
rect 7837 25789 7849 25823
rect 7883 25820 7895 25823
rect 8662 25820 8668 25832
rect 7883 25792 8668 25820
rect 7883 25789 7895 25792
rect 7837 25783 7895 25789
rect 8662 25780 8668 25792
rect 8720 25780 8726 25832
rect 8849 25823 8907 25829
rect 8849 25789 8861 25823
rect 8895 25789 8907 25823
rect 10235 25820 10263 25860
rect 10318 25848 10324 25900
rect 10376 25848 10382 25900
rect 10505 25891 10563 25897
rect 10505 25857 10517 25891
rect 10551 25857 10563 25891
rect 10505 25851 10563 25857
rect 10520 25820 10548 25851
rect 11790 25848 11796 25900
rect 11848 25888 11854 25900
rect 11885 25891 11943 25897
rect 11885 25888 11897 25891
rect 11848 25860 11897 25888
rect 11848 25848 11854 25860
rect 11885 25857 11897 25860
rect 11931 25857 11943 25891
rect 11885 25851 11943 25857
rect 10235 25792 10548 25820
rect 8849 25783 8907 25789
rect 8202 25752 8208 25764
rect 7024 25724 8208 25752
rect 8202 25712 8208 25724
rect 8260 25712 8266 25764
rect 8864 25752 8892 25783
rect 8680 25724 8892 25752
rect 10520 25752 10548 25792
rect 11514 25780 11520 25832
rect 11572 25780 11578 25832
rect 11992 25829 12020 25928
rect 14844 25928 17356 25956
rect 12406 25860 13124 25888
rect 11977 25823 12035 25829
rect 11977 25789 11989 25823
rect 12023 25820 12035 25823
rect 12158 25820 12164 25832
rect 12023 25792 12164 25820
rect 12023 25789 12035 25792
rect 11977 25783 12035 25789
rect 12158 25780 12164 25792
rect 12216 25780 12222 25832
rect 12406 25752 12434 25860
rect 13096 25829 13124 25860
rect 13354 25848 13360 25900
rect 13412 25888 13418 25900
rect 13449 25891 13507 25897
rect 13449 25888 13461 25891
rect 13412 25860 13461 25888
rect 13412 25848 13418 25860
rect 13449 25857 13461 25860
rect 13495 25857 13507 25891
rect 14844 25888 14872 25928
rect 13449 25851 13507 25857
rect 13602 25860 14872 25888
rect 12897 25823 12955 25829
rect 12897 25789 12909 25823
rect 12943 25789 12955 25823
rect 12897 25783 12955 25789
rect 13081 25823 13139 25829
rect 13081 25789 13093 25823
rect 13127 25820 13139 25823
rect 13602 25820 13630 25860
rect 15102 25848 15108 25900
rect 15160 25848 15166 25900
rect 15372 25891 15430 25897
rect 15372 25857 15384 25891
rect 15418 25888 15430 25891
rect 15838 25888 15844 25900
rect 15418 25860 15844 25888
rect 15418 25857 15430 25860
rect 15372 25851 15430 25857
rect 15838 25848 15844 25860
rect 15896 25848 15902 25900
rect 13127 25792 13630 25820
rect 14369 25823 14427 25829
rect 13127 25789 13139 25792
rect 13081 25783 13139 25789
rect 14369 25789 14381 25823
rect 14415 25789 14427 25823
rect 14369 25783 14427 25789
rect 10520 25724 12434 25752
rect 12912 25752 12940 25783
rect 13170 25752 13176 25764
rect 12912 25724 13176 25752
rect 8680 25696 8708 25724
rect 13170 25712 13176 25724
rect 13228 25712 13234 25764
rect 14384 25752 14412 25783
rect 14734 25780 14740 25832
rect 14792 25780 14798 25832
rect 14829 25823 14887 25829
rect 14829 25789 14841 25823
rect 14875 25820 14887 25823
rect 14918 25820 14924 25832
rect 14875 25792 14924 25820
rect 14875 25789 14887 25792
rect 14829 25783 14887 25789
rect 14918 25780 14924 25792
rect 14976 25780 14982 25832
rect 17126 25820 17132 25832
rect 16500 25792 17132 25820
rect 16500 25761 16528 25792
rect 17126 25780 17132 25792
rect 17184 25780 17190 25832
rect 17328 25829 17356 25928
rect 18322 25916 18328 25968
rect 18380 25916 18386 25968
rect 21358 25956 21364 25968
rect 18708 25928 21364 25956
rect 17497 25891 17555 25897
rect 17497 25857 17509 25891
rect 17543 25888 17555 25891
rect 18233 25891 18291 25897
rect 17543 25860 18184 25888
rect 17543 25857 17555 25860
rect 17497 25851 17555 25857
rect 17313 25823 17371 25829
rect 17313 25789 17325 25823
rect 17359 25820 17371 25823
rect 17862 25820 17868 25832
rect 17359 25792 17724 25820
rect 17359 25789 17371 25792
rect 17313 25783 17371 25789
rect 17696 25761 17724 25792
rect 17788 25792 17868 25820
rect 16485 25755 16543 25761
rect 14384 25724 15173 25752
rect 1762 25644 1768 25696
rect 1820 25684 1826 25696
rect 1857 25687 1915 25693
rect 1857 25684 1869 25687
rect 1820 25656 1869 25684
rect 1820 25644 1826 25656
rect 1857 25653 1869 25656
rect 1903 25653 1915 25687
rect 1857 25647 1915 25653
rect 6365 25687 6423 25693
rect 6365 25653 6377 25687
rect 6411 25684 6423 25687
rect 6638 25684 6644 25696
rect 6411 25656 6644 25684
rect 6411 25653 6423 25656
rect 6365 25647 6423 25653
rect 6638 25644 6644 25656
rect 6696 25644 6702 25696
rect 7374 25644 7380 25696
rect 7432 25684 7438 25696
rect 8113 25687 8171 25693
rect 8113 25684 8125 25687
rect 7432 25656 8125 25684
rect 7432 25644 7438 25656
rect 8113 25653 8125 25656
rect 8159 25653 8171 25687
rect 8113 25647 8171 25653
rect 8662 25644 8668 25696
rect 8720 25684 8726 25696
rect 9214 25684 9220 25696
rect 8720 25656 9220 25684
rect 8720 25644 8726 25656
rect 9214 25644 9220 25656
rect 9272 25644 9278 25696
rect 10229 25687 10287 25693
rect 10229 25653 10241 25687
rect 10275 25684 10287 25687
rect 10318 25684 10324 25696
rect 10275 25656 10324 25684
rect 10275 25653 10287 25656
rect 10229 25647 10287 25653
rect 10318 25644 10324 25656
rect 10376 25644 10382 25696
rect 10410 25644 10416 25696
rect 10468 25644 10474 25696
rect 10686 25644 10692 25696
rect 10744 25684 10750 25696
rect 12161 25687 12219 25693
rect 12161 25684 12173 25687
rect 10744 25656 12173 25684
rect 10744 25644 10750 25656
rect 12161 25653 12173 25656
rect 12207 25653 12219 25687
rect 12161 25647 12219 25653
rect 13538 25644 13544 25696
rect 13596 25644 13602 25696
rect 14642 25644 14648 25696
rect 14700 25684 14706 25696
rect 15013 25687 15071 25693
rect 15013 25684 15025 25687
rect 14700 25656 15025 25684
rect 14700 25644 14706 25656
rect 15013 25653 15025 25656
rect 15059 25653 15071 25687
rect 15145 25684 15173 25724
rect 16485 25721 16497 25755
rect 16531 25721 16543 25755
rect 17681 25755 17739 25761
rect 16485 25715 16543 25721
rect 16592 25724 17632 25752
rect 16592 25684 16620 25724
rect 15145 25656 16620 25684
rect 15013 25647 15071 25653
rect 16666 25644 16672 25696
rect 16724 25644 16730 25696
rect 17604 25684 17632 25724
rect 17681 25721 17693 25755
rect 17727 25721 17739 25755
rect 17681 25715 17739 25721
rect 17788 25684 17816 25792
rect 17862 25780 17868 25792
rect 17920 25780 17926 25832
rect 18156 25752 18184 25860
rect 18233 25857 18245 25891
rect 18279 25888 18291 25891
rect 18340 25888 18368 25916
rect 18279 25860 18368 25888
rect 18279 25857 18291 25860
rect 18233 25851 18291 25857
rect 18322 25780 18328 25832
rect 18380 25820 18386 25832
rect 18708 25820 18736 25928
rect 18785 25891 18843 25897
rect 18785 25857 18797 25891
rect 18831 25888 18843 25891
rect 18966 25888 18972 25900
rect 18831 25860 18972 25888
rect 18831 25857 18843 25860
rect 18785 25851 18843 25857
rect 18966 25848 18972 25860
rect 19024 25848 19030 25900
rect 19076 25897 19104 25928
rect 21358 25916 21364 25928
rect 21416 25956 21422 25968
rect 22830 25956 22836 25968
rect 21416 25928 22836 25956
rect 21416 25916 21422 25928
rect 22830 25916 22836 25928
rect 22888 25916 22894 25968
rect 19061 25891 19119 25897
rect 19061 25857 19073 25891
rect 19107 25857 19119 25891
rect 19061 25851 19119 25857
rect 20257 25891 20315 25897
rect 20257 25857 20269 25891
rect 20303 25888 20315 25891
rect 20990 25888 20996 25900
rect 20303 25860 20996 25888
rect 20303 25857 20315 25860
rect 20257 25851 20315 25857
rect 20990 25848 20996 25860
rect 21048 25888 21054 25900
rect 21726 25888 21732 25900
rect 21048 25860 21732 25888
rect 21048 25848 21054 25860
rect 21726 25848 21732 25860
rect 21784 25848 21790 25900
rect 22094 25848 22100 25900
rect 22152 25888 22158 25900
rect 22649 25891 22707 25897
rect 22649 25888 22661 25891
rect 22152 25860 22661 25888
rect 22152 25848 22158 25860
rect 22649 25857 22661 25860
rect 22695 25857 22707 25891
rect 22649 25851 22707 25857
rect 23293 25891 23351 25897
rect 23293 25857 23305 25891
rect 23339 25888 23351 25891
rect 24044 25888 24072 25996
rect 26510 25984 26516 25996
rect 26568 25984 26574 26036
rect 26973 26027 27031 26033
rect 26973 25993 26985 26027
rect 27019 25993 27031 26027
rect 26973 25987 27031 25993
rect 24394 25965 24400 25968
rect 24388 25956 24400 25965
rect 24355 25928 24400 25956
rect 24388 25919 24400 25928
rect 24394 25916 24400 25919
rect 24452 25916 24458 25968
rect 23339 25860 24072 25888
rect 24121 25891 24179 25897
rect 23339 25857 23351 25860
rect 23293 25851 23351 25857
rect 24121 25857 24133 25891
rect 24167 25888 24179 25891
rect 24854 25888 24860 25900
rect 24167 25860 24860 25888
rect 24167 25857 24179 25860
rect 24121 25851 24179 25857
rect 24854 25848 24860 25860
rect 24912 25888 24918 25900
rect 25958 25888 25964 25900
rect 24912 25860 25964 25888
rect 24912 25848 24918 25860
rect 25958 25848 25964 25860
rect 26016 25848 26022 25900
rect 26329 25891 26387 25897
rect 26329 25857 26341 25891
rect 26375 25888 26387 25891
rect 26988 25888 27016 25987
rect 33318 25984 33324 26036
rect 33376 25984 33382 26036
rect 26375 25860 27016 25888
rect 26375 25857 26387 25860
rect 26329 25851 26387 25857
rect 27338 25848 27344 25900
rect 27396 25848 27402 25900
rect 28074 25848 28080 25900
rect 28132 25848 28138 25900
rect 31294 25848 31300 25900
rect 31352 25888 31358 25900
rect 31389 25891 31447 25897
rect 31389 25888 31401 25891
rect 31352 25860 31401 25888
rect 31352 25848 31358 25860
rect 31389 25857 31401 25860
rect 31435 25857 31447 25891
rect 31389 25851 31447 25857
rect 32125 25891 32183 25897
rect 32125 25857 32137 25891
rect 32171 25888 32183 25891
rect 33134 25888 33140 25900
rect 32171 25860 33140 25888
rect 32171 25857 32183 25860
rect 32125 25851 32183 25857
rect 33134 25848 33140 25860
rect 33192 25888 33198 25900
rect 33505 25891 33563 25897
rect 33505 25888 33517 25891
rect 33192 25860 33517 25888
rect 33192 25848 33198 25860
rect 33505 25857 33517 25860
rect 33551 25857 33563 25891
rect 33505 25851 33563 25857
rect 18380 25792 18736 25820
rect 18984 25820 19012 25848
rect 20162 25820 20168 25832
rect 18984 25792 20168 25820
rect 18380 25780 18386 25792
rect 20162 25780 20168 25792
rect 20220 25780 20226 25832
rect 20530 25780 20536 25832
rect 20588 25780 20594 25832
rect 23385 25823 23443 25829
rect 23385 25789 23397 25823
rect 23431 25789 23443 25823
rect 23385 25783 23443 25789
rect 20548 25752 20576 25780
rect 23198 25752 23204 25764
rect 18156 25724 20576 25752
rect 22066 25724 23204 25752
rect 17604 25656 17816 25684
rect 18506 25644 18512 25696
rect 18564 25644 18570 25696
rect 18598 25644 18604 25696
rect 18656 25644 18662 25696
rect 20806 25644 20812 25696
rect 20864 25684 20870 25696
rect 21910 25684 21916 25696
rect 20864 25656 21916 25684
rect 20864 25644 20870 25656
rect 21910 25644 21916 25656
rect 21968 25684 21974 25696
rect 22066 25684 22094 25724
rect 23198 25712 23204 25724
rect 23256 25752 23262 25764
rect 23400 25752 23428 25783
rect 26418 25780 26424 25832
rect 26476 25820 26482 25832
rect 27433 25823 27491 25829
rect 27433 25820 27445 25823
rect 26476 25792 27445 25820
rect 26476 25780 26482 25792
rect 27433 25789 27445 25792
rect 27479 25789 27491 25823
rect 27433 25783 27491 25789
rect 27522 25780 27528 25832
rect 27580 25780 27586 25832
rect 30006 25780 30012 25832
rect 30064 25820 30070 25832
rect 32309 25823 32367 25829
rect 30064 25792 31754 25820
rect 30064 25780 30070 25792
rect 23256 25724 23428 25752
rect 23256 25712 23262 25724
rect 31110 25712 31116 25764
rect 31168 25752 31174 25764
rect 31726 25752 31754 25792
rect 32309 25789 32321 25823
rect 32355 25789 32367 25823
rect 32309 25783 32367 25789
rect 32324 25752 32352 25783
rect 32398 25780 32404 25832
rect 32456 25820 32462 25832
rect 32585 25823 32643 25829
rect 32585 25820 32597 25823
rect 32456 25792 32597 25820
rect 32456 25780 32462 25792
rect 32585 25789 32597 25792
rect 32631 25789 32643 25823
rect 32585 25783 32643 25789
rect 32677 25823 32735 25829
rect 32677 25789 32689 25823
rect 32723 25820 32735 25823
rect 32950 25820 32956 25832
rect 32723 25792 32956 25820
rect 32723 25789 32735 25792
rect 32677 25783 32735 25789
rect 32950 25780 32956 25792
rect 33008 25780 33014 25832
rect 31168 25724 31616 25752
rect 31726 25724 32352 25752
rect 31168 25712 31174 25724
rect 21968 25656 22094 25684
rect 21968 25644 21974 25656
rect 23566 25644 23572 25696
rect 23624 25644 23630 25696
rect 25498 25644 25504 25696
rect 25556 25644 25562 25696
rect 26145 25687 26203 25693
rect 26145 25653 26157 25687
rect 26191 25684 26203 25687
rect 26234 25684 26240 25696
rect 26191 25656 26240 25684
rect 26191 25653 26203 25656
rect 26145 25647 26203 25653
rect 26234 25644 26240 25656
rect 26292 25644 26298 25696
rect 27890 25644 27896 25696
rect 27948 25644 27954 25696
rect 31202 25644 31208 25696
rect 31260 25684 31266 25696
rect 31481 25687 31539 25693
rect 31481 25684 31493 25687
rect 31260 25656 31493 25684
rect 31260 25644 31266 25656
rect 31481 25653 31493 25656
rect 31527 25653 31539 25687
rect 31588 25684 31616 25724
rect 33870 25712 33876 25764
rect 33928 25712 33934 25764
rect 33965 25687 34023 25693
rect 33965 25684 33977 25687
rect 31588 25656 33977 25684
rect 31481 25647 31539 25653
rect 33965 25653 33977 25656
rect 34011 25653 34023 25687
rect 33965 25647 34023 25653
rect 1104 25594 36800 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 36800 25594
rect 1104 25520 36800 25542
rect 2866 25440 2872 25492
rect 2924 25440 2930 25492
rect 7190 25480 7196 25492
rect 5552 25452 7196 25480
rect 2884 25344 2912 25440
rect 4709 25347 4767 25353
rect 2884 25316 4200 25344
rect 1762 25285 1768 25288
rect 1489 25279 1547 25285
rect 1489 25245 1501 25279
rect 1535 25245 1547 25279
rect 1756 25276 1768 25285
rect 1723 25248 1768 25276
rect 1489 25239 1547 25245
rect 1756 25239 1768 25248
rect 1504 25208 1532 25239
rect 1762 25236 1768 25239
rect 1820 25236 1826 25288
rect 3973 25279 4031 25285
rect 3973 25245 3985 25279
rect 4019 25276 4031 25279
rect 4172 25276 4200 25316
rect 4709 25313 4721 25347
rect 4755 25344 4767 25347
rect 4982 25344 4988 25356
rect 4755 25316 4988 25344
rect 4755 25313 4767 25316
rect 4709 25307 4767 25313
rect 4982 25304 4988 25316
rect 5040 25344 5046 25356
rect 5442 25344 5448 25356
rect 5040 25316 5448 25344
rect 5040 25304 5046 25316
rect 5442 25304 5448 25316
rect 5500 25304 5506 25356
rect 5552 25353 5580 25452
rect 7190 25440 7196 25452
rect 7248 25440 7254 25492
rect 8018 25480 8024 25492
rect 7392 25452 8024 25480
rect 5537 25347 5595 25353
rect 5537 25313 5549 25347
rect 5583 25313 5595 25347
rect 5537 25307 5595 25313
rect 5810 25304 5816 25356
rect 5868 25304 5874 25356
rect 6089 25347 6147 25353
rect 6089 25313 6101 25347
rect 6135 25344 6147 25347
rect 7392 25344 7420 25452
rect 8018 25440 8024 25452
rect 8076 25440 8082 25492
rect 9122 25440 9128 25492
rect 9180 25480 9186 25492
rect 9309 25483 9367 25489
rect 9309 25480 9321 25483
rect 9180 25452 9321 25480
rect 9180 25440 9186 25452
rect 9309 25449 9321 25452
rect 9355 25449 9367 25483
rect 11514 25480 11520 25492
rect 9309 25443 9367 25449
rect 9416 25452 11520 25480
rect 9416 25412 9444 25452
rect 11514 25440 11520 25452
rect 11572 25480 11578 25492
rect 17678 25480 17684 25492
rect 11572 25452 17684 25480
rect 11572 25440 11578 25452
rect 17678 25440 17684 25452
rect 17736 25440 17742 25492
rect 20806 25480 20812 25492
rect 19260 25452 20812 25480
rect 7944 25384 9444 25412
rect 6135 25316 7420 25344
rect 6135 25313 6147 25316
rect 6089 25307 6147 25313
rect 7466 25304 7472 25356
rect 7524 25304 7530 25356
rect 7558 25304 7564 25356
rect 7616 25304 7622 25356
rect 4798 25276 4804 25288
rect 4019 25248 4108 25276
rect 4172 25248 4804 25276
rect 4019 25245 4031 25248
rect 3973 25239 4031 25245
rect 2866 25208 2872 25220
rect 1504 25180 2872 25208
rect 2866 25168 2872 25180
rect 2924 25168 2930 25220
rect 3786 25100 3792 25152
rect 3844 25100 3850 25152
rect 4080 25149 4108 25248
rect 4798 25236 4804 25248
rect 4856 25276 4862 25288
rect 4893 25279 4951 25285
rect 4893 25276 4905 25279
rect 4856 25248 4905 25276
rect 4856 25236 4862 25248
rect 4893 25245 4905 25248
rect 4939 25245 4951 25279
rect 4893 25239 4951 25245
rect 5077 25279 5135 25285
rect 5077 25245 5089 25279
rect 5123 25276 5135 25279
rect 5258 25276 5264 25288
rect 5123 25248 5264 25276
rect 5123 25245 5135 25248
rect 5077 25239 5135 25245
rect 5258 25236 5264 25248
rect 5316 25236 5322 25288
rect 5902 25236 5908 25288
rect 5960 25285 5966 25288
rect 5960 25279 5988 25285
rect 5976 25245 5988 25279
rect 5960 25239 5988 25245
rect 7101 25279 7159 25285
rect 7101 25245 7113 25279
rect 7147 25276 7159 25279
rect 7282 25276 7288 25288
rect 7147 25248 7288 25276
rect 7147 25245 7159 25248
rect 7101 25239 7159 25245
rect 5960 25236 5966 25239
rect 7282 25236 7288 25248
rect 7340 25276 7346 25288
rect 7944 25285 7972 25384
rect 10410 25372 10416 25424
rect 10468 25372 10474 25424
rect 10781 25415 10839 25421
rect 10781 25412 10793 25415
rect 10520 25384 10793 25412
rect 9306 25344 9312 25356
rect 9140 25316 9312 25344
rect 9140 25285 9168 25316
rect 9306 25304 9312 25316
rect 9364 25304 9370 25356
rect 9401 25347 9459 25353
rect 9401 25313 9413 25347
rect 9447 25344 9459 25347
rect 10428 25344 10456 25372
rect 9447 25316 10456 25344
rect 9447 25313 9459 25316
rect 9401 25307 9459 25313
rect 7929 25279 7987 25285
rect 7929 25276 7941 25279
rect 7340 25248 7941 25276
rect 7340 25236 7346 25248
rect 7929 25245 7941 25248
rect 7975 25245 7987 25279
rect 7929 25239 7987 25245
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25245 9183 25279
rect 9125 25239 9183 25245
rect 9217 25279 9275 25285
rect 9217 25245 9229 25279
rect 9263 25276 9275 25279
rect 9490 25276 9496 25288
rect 9263 25248 9496 25276
rect 9263 25245 9275 25248
rect 9217 25239 9275 25245
rect 9490 25236 9496 25248
rect 9548 25236 9554 25288
rect 10321 25279 10379 25285
rect 10321 25245 10333 25279
rect 10367 25245 10379 25279
rect 10321 25239 10379 25245
rect 10413 25279 10471 25285
rect 10413 25245 10425 25279
rect 10459 25276 10471 25279
rect 10520 25276 10548 25384
rect 10781 25381 10793 25384
rect 10827 25381 10839 25415
rect 10781 25375 10839 25381
rect 12158 25372 12164 25424
rect 12216 25412 12222 25424
rect 19260 25412 19288 25452
rect 20806 25440 20812 25452
rect 20864 25440 20870 25492
rect 24489 25483 24547 25489
rect 24489 25449 24501 25483
rect 24535 25480 24547 25483
rect 24578 25480 24584 25492
rect 24535 25452 24584 25480
rect 24535 25449 24547 25452
rect 24489 25443 24547 25449
rect 24578 25440 24584 25452
rect 24636 25440 24642 25492
rect 24670 25440 24676 25492
rect 24728 25480 24734 25492
rect 27338 25480 27344 25492
rect 24728 25452 27344 25480
rect 24728 25440 24734 25452
rect 27338 25440 27344 25452
rect 27396 25440 27402 25492
rect 27982 25480 27988 25492
rect 27632 25452 27988 25480
rect 12216 25384 19288 25412
rect 12216 25372 12222 25384
rect 10597 25347 10655 25353
rect 10597 25313 10609 25347
rect 10643 25344 10655 25347
rect 11238 25344 11244 25356
rect 10643 25316 11244 25344
rect 10643 25313 10655 25316
rect 10597 25307 10655 25313
rect 11238 25304 11244 25316
rect 11296 25304 11302 25356
rect 11425 25347 11483 25353
rect 11425 25313 11437 25347
rect 11471 25344 11483 25347
rect 11514 25344 11520 25356
rect 11471 25316 11520 25344
rect 11471 25313 11483 25316
rect 11425 25307 11483 25313
rect 11514 25304 11520 25316
rect 11572 25304 11578 25356
rect 18966 25344 18972 25356
rect 15764 25316 18972 25344
rect 10459 25248 10548 25276
rect 10459 25245 10471 25248
rect 10413 25239 10471 25245
rect 4433 25211 4491 25217
rect 4433 25177 4445 25211
rect 4479 25208 4491 25211
rect 4706 25208 4712 25220
rect 4479 25180 4712 25208
rect 4479 25177 4491 25180
rect 4433 25171 4491 25177
rect 4706 25168 4712 25180
rect 4764 25168 4770 25220
rect 7006 25168 7012 25220
rect 7064 25208 7070 25220
rect 8113 25211 8171 25217
rect 8113 25208 8125 25211
rect 7064 25180 8125 25208
rect 7064 25168 7070 25180
rect 8113 25177 8125 25180
rect 8159 25208 8171 25211
rect 10336 25208 10364 25239
rect 10686 25236 10692 25288
rect 10744 25236 10750 25288
rect 14829 25279 14887 25285
rect 14829 25276 14841 25279
rect 11164 25248 14841 25276
rect 11164 25208 11192 25248
rect 14829 25245 14841 25248
rect 14875 25245 14887 25279
rect 14829 25239 14887 25245
rect 8159 25180 11192 25208
rect 11241 25211 11299 25217
rect 8159 25177 8171 25180
rect 8113 25171 8171 25177
rect 11241 25177 11253 25211
rect 11287 25208 11299 25211
rect 12066 25208 12072 25220
rect 11287 25180 12072 25208
rect 11287 25177 11299 25180
rect 11241 25171 11299 25177
rect 12066 25168 12072 25180
rect 12124 25168 12130 25220
rect 4065 25143 4123 25149
rect 4065 25109 4077 25143
rect 4111 25109 4123 25143
rect 4065 25103 4123 25109
rect 4522 25100 4528 25152
rect 4580 25140 4586 25152
rect 5810 25140 5816 25152
rect 4580 25112 5816 25140
rect 4580 25100 4586 25112
rect 5810 25100 5816 25112
rect 5868 25100 5874 25152
rect 6733 25143 6791 25149
rect 6733 25109 6745 25143
rect 6779 25140 6791 25143
rect 6914 25140 6920 25152
rect 6779 25112 6920 25140
rect 6779 25109 6791 25112
rect 6733 25103 6791 25109
rect 6914 25100 6920 25112
rect 6972 25100 6978 25152
rect 7190 25100 7196 25152
rect 7248 25140 7254 25152
rect 7745 25143 7803 25149
rect 7745 25140 7757 25143
rect 7248 25112 7757 25140
rect 7248 25100 7254 25112
rect 7745 25109 7757 25112
rect 7791 25109 7803 25143
rect 7745 25103 7803 25109
rect 9950 25100 9956 25152
rect 10008 25140 10014 25152
rect 10137 25143 10195 25149
rect 10137 25140 10149 25143
rect 10008 25112 10149 25140
rect 10008 25100 10014 25112
rect 10137 25109 10149 25112
rect 10183 25109 10195 25143
rect 10137 25103 10195 25109
rect 11146 25100 11152 25152
rect 11204 25100 11210 25152
rect 14458 25100 14464 25152
rect 14516 25140 14522 25152
rect 14645 25143 14703 25149
rect 14645 25140 14657 25143
rect 14516 25112 14657 25140
rect 14516 25100 14522 25112
rect 14645 25109 14657 25112
rect 14691 25109 14703 25143
rect 14844 25140 14872 25239
rect 14918 25236 14924 25288
rect 14976 25276 14982 25288
rect 15105 25279 15163 25285
rect 15105 25276 15117 25279
rect 14976 25248 15117 25276
rect 14976 25236 14982 25248
rect 15105 25245 15117 25248
rect 15151 25245 15163 25279
rect 15105 25239 15163 25245
rect 15013 25211 15071 25217
rect 15013 25177 15025 25211
rect 15059 25208 15071 25211
rect 15286 25208 15292 25220
rect 15059 25180 15292 25208
rect 15059 25177 15071 25180
rect 15013 25171 15071 25177
rect 15286 25168 15292 25180
rect 15344 25168 15350 25220
rect 15764 25140 15792 25316
rect 18966 25304 18972 25316
rect 19024 25304 19030 25356
rect 19076 25316 19380 25344
rect 16117 25279 16175 25285
rect 16117 25245 16129 25279
rect 16163 25276 16175 25279
rect 16666 25276 16672 25288
rect 16163 25248 16672 25276
rect 16163 25245 16175 25248
rect 16117 25239 16175 25245
rect 16666 25236 16672 25248
rect 16724 25236 16730 25288
rect 19076 25285 19104 25316
rect 19352 25288 19380 25316
rect 20530 25304 20536 25356
rect 20588 25344 20594 25356
rect 27632 25353 27660 25452
rect 27982 25440 27988 25452
rect 28040 25480 28046 25492
rect 28040 25452 29592 25480
rect 28040 25440 28046 25452
rect 25133 25347 25191 25353
rect 25133 25344 25145 25347
rect 20588 25316 25145 25344
rect 20588 25304 20594 25316
rect 25133 25313 25145 25316
rect 25179 25344 25191 25347
rect 27617 25347 27675 25353
rect 25179 25316 25636 25344
rect 25179 25313 25191 25316
rect 25133 25307 25191 25313
rect 19061 25279 19119 25285
rect 19061 25245 19073 25279
rect 19107 25245 19119 25279
rect 19061 25239 19119 25245
rect 19242 25236 19248 25288
rect 19300 25236 19306 25288
rect 19334 25236 19340 25288
rect 19392 25236 19398 25288
rect 24949 25279 25007 25285
rect 24949 25245 24961 25279
rect 24995 25276 25007 25279
rect 25498 25276 25504 25288
rect 24995 25248 25504 25276
rect 24995 25245 25007 25248
rect 24949 25239 25007 25245
rect 25498 25236 25504 25248
rect 25556 25236 25562 25288
rect 15838 25168 15844 25220
rect 15896 25208 15902 25220
rect 19490 25211 19548 25217
rect 19490 25208 19502 25211
rect 15896 25180 15976 25208
rect 15896 25168 15902 25180
rect 15948 25149 15976 25180
rect 18892 25180 19502 25208
rect 18892 25149 18920 25180
rect 19490 25177 19502 25180
rect 19536 25177 19548 25211
rect 22094 25208 22100 25220
rect 19490 25171 19548 25177
rect 19628 25180 22100 25208
rect 14844 25112 15792 25140
rect 15933 25143 15991 25149
rect 14645 25103 14703 25109
rect 15933 25109 15945 25143
rect 15979 25109 15991 25143
rect 15933 25103 15991 25109
rect 18877 25143 18935 25149
rect 18877 25109 18889 25143
rect 18923 25109 18935 25143
rect 18877 25103 18935 25109
rect 18966 25100 18972 25152
rect 19024 25140 19030 25152
rect 19628 25140 19656 25180
rect 22094 25168 22100 25180
rect 22152 25168 22158 25220
rect 25608 25208 25636 25316
rect 27617 25313 27629 25347
rect 27663 25313 27675 25347
rect 27617 25307 27675 25313
rect 25958 25236 25964 25288
rect 26016 25236 26022 25288
rect 26234 25285 26240 25288
rect 26228 25276 26240 25285
rect 26195 25248 26240 25276
rect 26228 25239 26240 25248
rect 26234 25236 26240 25239
rect 26292 25236 26298 25288
rect 27890 25285 27896 25288
rect 27884 25276 27896 25285
rect 27851 25248 27896 25276
rect 27884 25239 27896 25248
rect 27890 25236 27896 25239
rect 27948 25236 27954 25288
rect 29362 25236 29368 25288
rect 29420 25236 29426 25288
rect 29564 25285 29592 25452
rect 30466 25440 30472 25492
rect 30524 25480 30530 25492
rect 31665 25483 31723 25489
rect 31665 25480 31677 25483
rect 30524 25452 31677 25480
rect 30524 25440 30530 25452
rect 31665 25449 31677 25452
rect 31711 25449 31723 25483
rect 31665 25443 31723 25449
rect 32306 25440 32312 25492
rect 32364 25440 32370 25492
rect 32398 25412 32404 25424
rect 31864 25384 32404 25412
rect 31110 25304 31116 25356
rect 31168 25344 31174 25356
rect 31864 25353 31892 25384
rect 32398 25372 32404 25384
rect 32456 25412 32462 25424
rect 32456 25384 32996 25412
rect 32456 25372 32462 25384
rect 32968 25356 32996 25384
rect 31389 25347 31447 25353
rect 31389 25344 31401 25347
rect 31168 25316 31401 25344
rect 31168 25304 31174 25316
rect 31389 25313 31401 25316
rect 31435 25313 31447 25347
rect 31389 25307 31447 25313
rect 31849 25347 31907 25353
rect 31849 25313 31861 25347
rect 31895 25313 31907 25347
rect 31849 25307 31907 25313
rect 32766 25304 32772 25356
rect 32824 25304 32830 25356
rect 32950 25304 32956 25356
rect 33008 25344 33014 25356
rect 33965 25347 34023 25353
rect 33965 25344 33977 25347
rect 33008 25316 33977 25344
rect 33008 25304 33014 25316
rect 33965 25313 33977 25316
rect 34011 25313 34023 25347
rect 33965 25307 34023 25313
rect 29549 25279 29607 25285
rect 29549 25245 29561 25279
rect 29595 25276 29607 25279
rect 30374 25276 30380 25288
rect 29595 25248 30380 25276
rect 29595 25245 29607 25248
rect 29549 25239 29607 25245
rect 30374 25236 30380 25248
rect 30432 25236 30438 25288
rect 30742 25236 30748 25288
rect 30800 25276 30806 25288
rect 31481 25279 31539 25285
rect 31481 25276 31493 25279
rect 30800 25248 31493 25276
rect 30800 25236 30806 25248
rect 31481 25245 31493 25248
rect 31527 25245 31539 25279
rect 31481 25239 31539 25245
rect 32217 25279 32275 25285
rect 32217 25245 32229 25279
rect 32263 25245 32275 25279
rect 32217 25239 32275 25245
rect 29086 25208 29092 25220
rect 25608 25180 29092 25208
rect 29086 25168 29092 25180
rect 29144 25168 29150 25220
rect 29794 25211 29852 25217
rect 29794 25208 29806 25211
rect 29196 25180 29806 25208
rect 19024 25112 19656 25140
rect 19024 25100 19030 25112
rect 19978 25100 19984 25152
rect 20036 25140 20042 25152
rect 20625 25143 20683 25149
rect 20625 25140 20637 25143
rect 20036 25112 20637 25140
rect 20036 25100 20042 25112
rect 20625 25109 20637 25112
rect 20671 25109 20683 25143
rect 20625 25103 20683 25109
rect 24857 25143 24915 25149
rect 24857 25109 24869 25143
rect 24903 25140 24915 25143
rect 25038 25140 25044 25152
rect 24903 25112 25044 25140
rect 24903 25109 24915 25112
rect 24857 25103 24915 25109
rect 25038 25100 25044 25112
rect 25096 25100 25102 25152
rect 28258 25100 28264 25152
rect 28316 25140 28322 25152
rect 29196 25149 29224 25180
rect 29794 25177 29806 25180
rect 29840 25177 29852 25211
rect 29794 25171 29852 25177
rect 31021 25211 31079 25217
rect 31021 25177 31033 25211
rect 31067 25208 31079 25211
rect 31386 25208 31392 25220
rect 31067 25180 31392 25208
rect 31067 25177 31079 25180
rect 31021 25171 31079 25177
rect 31386 25168 31392 25180
rect 31444 25168 31450 25220
rect 32232 25208 32260 25239
rect 33042 25236 33048 25288
rect 33100 25236 33106 25288
rect 33689 25279 33747 25285
rect 33689 25245 33701 25279
rect 33735 25276 33747 25279
rect 33870 25276 33876 25288
rect 33735 25248 33876 25276
rect 33735 25245 33747 25248
rect 33689 25239 33747 25245
rect 33870 25236 33876 25248
rect 33928 25236 33934 25288
rect 33134 25208 33140 25220
rect 32232 25180 33140 25208
rect 33134 25168 33140 25180
rect 33192 25168 33198 25220
rect 28997 25143 29055 25149
rect 28997 25140 29009 25143
rect 28316 25112 29009 25140
rect 28316 25100 28322 25112
rect 28997 25109 29009 25112
rect 29043 25109 29055 25143
rect 28997 25103 29055 25109
rect 29181 25143 29239 25149
rect 29181 25109 29193 25143
rect 29227 25109 29239 25143
rect 29181 25103 29239 25109
rect 30926 25100 30932 25152
rect 30984 25100 30990 25152
rect 31297 25143 31355 25149
rect 31297 25109 31309 25143
rect 31343 25140 31355 25143
rect 31570 25140 31576 25152
rect 31343 25112 31576 25140
rect 31343 25109 31355 25112
rect 31297 25103 31355 25109
rect 31570 25100 31576 25112
rect 31628 25100 31634 25152
rect 32030 25100 32036 25152
rect 32088 25100 32094 25152
rect 1104 25050 36800 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 36800 25050
rect 1104 24976 36800 24998
rect 4522 24896 4528 24948
rect 4580 24936 4586 24948
rect 4709 24939 4767 24945
rect 4709 24936 4721 24939
rect 4580 24908 4721 24936
rect 4580 24896 4586 24908
rect 4709 24905 4721 24908
rect 4755 24905 4767 24939
rect 4709 24899 4767 24905
rect 8202 24896 8208 24948
rect 8260 24936 8266 24948
rect 11514 24936 11520 24948
rect 8260 24908 11520 24936
rect 8260 24896 8266 24908
rect 11514 24896 11520 24908
rect 11572 24936 11578 24948
rect 18966 24936 18972 24948
rect 11572 24908 18972 24936
rect 11572 24896 11578 24908
rect 18966 24896 18972 24908
rect 19024 24896 19030 24948
rect 19334 24896 19340 24948
rect 19392 24936 19398 24948
rect 19613 24939 19671 24945
rect 19613 24936 19625 24939
rect 19392 24908 19625 24936
rect 19392 24896 19398 24908
rect 19613 24905 19625 24908
rect 19659 24905 19671 24939
rect 19613 24899 19671 24905
rect 19978 24896 19984 24948
rect 20036 24896 20042 24948
rect 20073 24939 20131 24945
rect 20073 24905 20085 24939
rect 20119 24936 20131 24939
rect 20898 24936 20904 24948
rect 20119 24908 20904 24936
rect 20119 24905 20131 24908
rect 20073 24899 20131 24905
rect 20898 24896 20904 24908
rect 20956 24896 20962 24948
rect 23661 24939 23719 24945
rect 23661 24936 23673 24939
rect 22664 24908 23673 24936
rect 3596 24871 3654 24877
rect 3596 24837 3608 24871
rect 3642 24868 3654 24871
rect 3786 24868 3792 24880
rect 3642 24840 3792 24868
rect 3642 24837 3654 24840
rect 3596 24831 3654 24837
rect 3786 24828 3792 24840
rect 3844 24828 3850 24880
rect 7561 24871 7619 24877
rect 7561 24837 7573 24871
rect 7607 24868 7619 24871
rect 7742 24868 7748 24880
rect 7607 24840 7748 24868
rect 7607 24837 7619 24840
rect 7561 24831 7619 24837
rect 7742 24828 7748 24840
rect 7800 24828 7806 24880
rect 18598 24868 18604 24880
rect 17880 24840 18604 24868
rect 1394 24760 1400 24812
rect 1452 24760 1458 24812
rect 6549 24803 6607 24809
rect 6549 24769 6561 24803
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 1673 24735 1731 24741
rect 1673 24701 1685 24735
rect 1719 24732 1731 24735
rect 1854 24732 1860 24744
rect 1719 24704 1860 24732
rect 1719 24701 1731 24704
rect 1673 24695 1731 24701
rect 1854 24692 1860 24704
rect 1912 24692 1918 24744
rect 2866 24692 2872 24744
rect 2924 24732 2930 24744
rect 3326 24732 3332 24744
rect 2924 24704 3332 24732
rect 2924 24692 2930 24704
rect 3326 24692 3332 24704
rect 3384 24692 3390 24744
rect 6564 24732 6592 24763
rect 6638 24760 6644 24812
rect 6696 24760 6702 24812
rect 6917 24803 6975 24809
rect 6917 24769 6929 24803
rect 6963 24800 6975 24803
rect 7190 24800 7196 24812
rect 6963 24772 7196 24800
rect 6963 24769 6975 24772
rect 6917 24763 6975 24769
rect 7190 24760 7196 24772
rect 7248 24760 7254 24812
rect 7650 24760 7656 24812
rect 7708 24760 7714 24812
rect 11882 24760 11888 24812
rect 11940 24800 11946 24812
rect 12342 24809 12348 24812
rect 12069 24803 12127 24809
rect 12069 24800 12081 24803
rect 11940 24772 12081 24800
rect 11940 24760 11946 24772
rect 12069 24769 12081 24772
rect 12115 24769 12127 24803
rect 12069 24763 12127 24769
rect 12336 24763 12348 24809
rect 12342 24760 12348 24763
rect 12400 24760 12406 24812
rect 12618 24760 12624 24812
rect 12676 24800 12682 24812
rect 13633 24803 13691 24809
rect 13633 24800 13645 24803
rect 12676 24772 13645 24800
rect 12676 24760 12682 24772
rect 13633 24769 13645 24772
rect 13679 24769 13691 24803
rect 13633 24763 13691 24769
rect 14369 24803 14427 24809
rect 14369 24769 14381 24803
rect 14415 24769 14427 24803
rect 14369 24763 14427 24769
rect 7006 24732 7012 24744
rect 6564 24704 7012 24732
rect 7006 24692 7012 24704
rect 7064 24692 7070 24744
rect 7837 24735 7895 24741
rect 7837 24701 7849 24735
rect 7883 24732 7895 24735
rect 8202 24732 8208 24744
rect 7883 24704 8208 24732
rect 7883 24701 7895 24704
rect 7837 24695 7895 24701
rect 8202 24692 8208 24704
rect 8260 24692 8266 24744
rect 14093 24735 14151 24741
rect 14093 24701 14105 24735
rect 14139 24732 14151 24735
rect 14384 24732 14412 24763
rect 14458 24760 14464 24812
rect 14516 24760 14522 24812
rect 14737 24803 14795 24809
rect 14737 24769 14749 24803
rect 14783 24800 14795 24803
rect 17589 24803 17647 24809
rect 14783 24772 15332 24800
rect 14783 24769 14795 24772
rect 14737 24763 14795 24769
rect 14139 24704 14412 24732
rect 14139 24701 14151 24704
rect 14093 24695 14151 24701
rect 14642 24692 14648 24744
rect 14700 24692 14706 24744
rect 14826 24692 14832 24744
rect 14884 24692 14890 24744
rect 15304 24741 15332 24772
rect 17589 24769 17601 24803
rect 17635 24769 17647 24803
rect 17589 24763 17647 24769
rect 17681 24803 17739 24809
rect 17681 24769 17693 24803
rect 17727 24800 17739 24803
rect 17880 24800 17908 24840
rect 18598 24828 18604 24840
rect 18656 24828 18662 24880
rect 21008 24840 21956 24868
rect 17727 24772 17908 24800
rect 17727 24769 17739 24772
rect 17681 24763 17739 24769
rect 15289 24735 15347 24741
rect 15289 24701 15301 24735
rect 15335 24701 15347 24735
rect 15289 24695 15347 24701
rect 6825 24667 6883 24673
rect 6825 24633 6837 24667
rect 6871 24664 6883 24667
rect 7558 24664 7564 24676
rect 6871 24636 7564 24664
rect 6871 24633 6883 24636
rect 6825 24627 6883 24633
rect 7558 24624 7564 24636
rect 7616 24624 7622 24676
rect 10870 24624 10876 24676
rect 10928 24664 10934 24676
rect 11882 24664 11888 24676
rect 10928 24636 11888 24664
rect 10928 24624 10934 24636
rect 11882 24624 11888 24636
rect 11940 24624 11946 24676
rect 13998 24624 14004 24676
rect 14056 24624 14062 24676
rect 14458 24624 14464 24676
rect 14516 24664 14522 24676
rect 15105 24667 15163 24673
rect 15105 24664 15117 24667
rect 14516 24636 15117 24664
rect 14516 24624 14522 24636
rect 15105 24633 15117 24636
rect 15151 24633 15163 24667
rect 15105 24627 15163 24633
rect 16482 24624 16488 24676
rect 16540 24664 16546 24676
rect 17604 24664 17632 24763
rect 17954 24760 17960 24812
rect 18012 24760 18018 24812
rect 18049 24803 18107 24809
rect 18049 24769 18061 24803
rect 18095 24800 18107 24803
rect 18095 24772 20116 24800
rect 18095 24769 18107 24772
rect 18049 24763 18107 24769
rect 17865 24735 17923 24741
rect 17865 24701 17877 24735
rect 17911 24732 17923 24735
rect 18506 24732 18512 24744
rect 17911 24704 18512 24732
rect 17911 24701 17923 24704
rect 17865 24695 17923 24701
rect 18506 24692 18512 24704
rect 18564 24692 18570 24744
rect 18598 24664 18604 24676
rect 16540 24636 17540 24664
rect 17604 24636 18604 24664
rect 16540 24624 16546 24636
rect 6270 24556 6276 24608
rect 6328 24596 6334 24608
rect 6365 24599 6423 24605
rect 6365 24596 6377 24599
rect 6328 24568 6377 24596
rect 6328 24556 6334 24568
rect 6365 24565 6377 24568
rect 6411 24565 6423 24599
rect 6365 24559 6423 24565
rect 7098 24556 7104 24608
rect 7156 24596 7162 24608
rect 7193 24599 7251 24605
rect 7193 24596 7205 24599
rect 7156 24568 7205 24596
rect 7156 24556 7162 24568
rect 7193 24565 7205 24568
rect 7239 24565 7251 24599
rect 7193 24559 7251 24565
rect 12986 24556 12992 24608
rect 13044 24596 13050 24608
rect 13449 24599 13507 24605
rect 13449 24596 13461 24599
rect 13044 24568 13461 24596
rect 13044 24556 13050 24568
rect 13449 24565 13461 24568
rect 13495 24565 13507 24599
rect 13449 24559 13507 24565
rect 14090 24556 14096 24608
rect 14148 24596 14154 24608
rect 14185 24599 14243 24605
rect 14185 24596 14197 24599
rect 14148 24568 14197 24596
rect 14148 24556 14154 24568
rect 14185 24565 14197 24568
rect 14231 24565 14243 24599
rect 14185 24559 14243 24565
rect 16666 24556 16672 24608
rect 16724 24596 16730 24608
rect 17405 24599 17463 24605
rect 17405 24596 17417 24599
rect 16724 24568 17417 24596
rect 16724 24556 16730 24568
rect 17405 24565 17417 24568
rect 17451 24565 17463 24599
rect 17512 24596 17540 24636
rect 18598 24624 18604 24636
rect 18656 24624 18662 24676
rect 20088 24664 20116 24772
rect 20162 24760 20168 24812
rect 20220 24800 20226 24812
rect 21008 24800 21036 24840
rect 20220 24772 21036 24800
rect 21085 24803 21143 24809
rect 20220 24760 20226 24772
rect 21085 24769 21097 24803
rect 21131 24769 21143 24803
rect 21085 24763 21143 24769
rect 20257 24735 20315 24741
rect 20257 24701 20269 24735
rect 20303 24701 20315 24735
rect 21100 24732 21128 24763
rect 21174 24760 21180 24812
rect 21232 24760 21238 24812
rect 21453 24803 21511 24809
rect 21453 24769 21465 24803
rect 21499 24800 21511 24803
rect 21818 24800 21824 24812
rect 21499 24772 21824 24800
rect 21499 24769 21511 24772
rect 21453 24763 21511 24769
rect 21818 24760 21824 24772
rect 21876 24760 21882 24812
rect 21928 24800 21956 24840
rect 22664 24809 22692 24908
rect 23661 24905 23673 24908
rect 23707 24905 23719 24939
rect 23661 24899 23719 24905
rect 24121 24939 24179 24945
rect 24121 24905 24133 24939
rect 24167 24936 24179 24939
rect 25130 24936 25136 24948
rect 24167 24908 25136 24936
rect 24167 24905 24179 24908
rect 24121 24899 24179 24905
rect 25130 24896 25136 24908
rect 25188 24896 25194 24948
rect 27893 24939 27951 24945
rect 27893 24905 27905 24939
rect 27939 24936 27951 24939
rect 28074 24936 28080 24948
rect 27939 24908 28080 24936
rect 27939 24905 27951 24908
rect 27893 24899 27951 24905
rect 28074 24896 28080 24908
rect 28132 24896 28138 24948
rect 28258 24896 28264 24948
rect 28316 24896 28322 24948
rect 29362 24896 29368 24948
rect 29420 24936 29426 24948
rect 29457 24939 29515 24945
rect 29457 24936 29469 24939
rect 29420 24908 29469 24936
rect 29420 24896 29426 24908
rect 29457 24905 29469 24908
rect 29503 24905 29515 24939
rect 29457 24899 29515 24905
rect 29822 24896 29828 24948
rect 29880 24896 29886 24948
rect 30561 24939 30619 24945
rect 30561 24905 30573 24939
rect 30607 24936 30619 24939
rect 31570 24936 31576 24948
rect 30607 24908 31576 24936
rect 30607 24905 30619 24908
rect 30561 24899 30619 24905
rect 31570 24896 31576 24908
rect 31628 24936 31634 24948
rect 32030 24936 32036 24948
rect 31628 24908 32036 24936
rect 31628 24896 31634 24908
rect 32030 24896 32036 24908
rect 32088 24896 32094 24948
rect 33870 24896 33876 24948
rect 33928 24896 33934 24948
rect 24029 24871 24087 24877
rect 24029 24837 24041 24871
rect 24075 24868 24087 24871
rect 25222 24868 25228 24880
rect 24075 24840 25228 24868
rect 24075 24837 24087 24840
rect 24029 24831 24087 24837
rect 25222 24828 25228 24840
rect 25280 24828 25286 24880
rect 33042 24868 33048 24880
rect 29840 24840 31064 24868
rect 22557 24803 22615 24809
rect 22557 24800 22569 24803
rect 21928 24772 22569 24800
rect 22557 24769 22569 24772
rect 22603 24769 22615 24803
rect 22557 24763 22615 24769
rect 22649 24803 22707 24809
rect 22649 24769 22661 24803
rect 22695 24769 22707 24803
rect 22649 24763 22707 24769
rect 22922 24760 22928 24812
rect 22980 24760 22986 24812
rect 23106 24760 23112 24812
rect 23164 24800 23170 24812
rect 27522 24800 27528 24812
rect 23164 24772 24072 24800
rect 23164 24760 23170 24772
rect 21266 24732 21272 24744
rect 21100 24704 21272 24732
rect 20257 24695 20315 24701
rect 20272 24664 20300 24695
rect 21266 24692 21272 24704
rect 21324 24692 21330 24744
rect 21361 24735 21419 24741
rect 21361 24701 21373 24735
rect 21407 24732 21419 24735
rect 21542 24732 21548 24744
rect 21407 24704 21548 24732
rect 21407 24701 21419 24704
rect 21361 24695 21419 24701
rect 21542 24692 21548 24704
rect 21600 24692 21606 24744
rect 23017 24735 23075 24741
rect 23017 24701 23029 24735
rect 23063 24732 23075 24735
rect 23198 24732 23204 24744
rect 23063 24704 23204 24732
rect 23063 24701 23075 24704
rect 23017 24695 23075 24701
rect 23198 24692 23204 24704
rect 23256 24692 23262 24744
rect 23934 24732 23940 24744
rect 23400 24704 23940 24732
rect 23400 24673 23428 24704
rect 23934 24692 23940 24704
rect 23992 24692 23998 24744
rect 24044 24732 24072 24772
rect 25976 24772 27528 24800
rect 24213 24735 24271 24741
rect 24213 24732 24225 24735
rect 24044 24704 24225 24732
rect 24213 24701 24225 24704
rect 24259 24701 24271 24735
rect 25976 24732 26004 24772
rect 27522 24760 27528 24772
rect 27580 24800 27586 24812
rect 29840 24800 29868 24840
rect 27580 24772 29868 24800
rect 29917 24803 29975 24809
rect 27580 24760 27586 24772
rect 24213 24695 24271 24701
rect 25332 24704 26004 24732
rect 23385 24667 23443 24673
rect 20088 24636 23336 24664
rect 18233 24599 18291 24605
rect 18233 24596 18245 24599
rect 17512 24568 18245 24596
rect 17405 24559 17463 24565
rect 18233 24565 18245 24568
rect 18279 24565 18291 24599
rect 18233 24559 18291 24565
rect 20898 24556 20904 24608
rect 20956 24556 20962 24608
rect 20990 24556 20996 24608
rect 21048 24596 21054 24608
rect 21542 24596 21548 24608
rect 21048 24568 21548 24596
rect 21048 24556 21054 24568
rect 21542 24556 21548 24568
rect 21600 24556 21606 24608
rect 22370 24556 22376 24608
rect 22428 24556 22434 24608
rect 22830 24556 22836 24608
rect 22888 24556 22894 24608
rect 23308 24596 23336 24636
rect 23385 24633 23397 24667
rect 23431 24633 23443 24667
rect 23385 24627 23443 24633
rect 23477 24667 23535 24673
rect 23477 24633 23489 24667
rect 23523 24664 23535 24667
rect 23750 24664 23756 24676
rect 23523 24636 23756 24664
rect 23523 24633 23535 24636
rect 23477 24627 23535 24633
rect 23750 24624 23756 24636
rect 23808 24624 23814 24676
rect 25332 24596 25360 24704
rect 26050 24692 26056 24744
rect 26108 24732 26114 24744
rect 28166 24732 28172 24744
rect 26108 24704 28172 24732
rect 26108 24692 26114 24704
rect 28166 24692 28172 24704
rect 28224 24692 28230 24744
rect 28350 24692 28356 24744
rect 28408 24692 28414 24744
rect 28460 24741 28488 24772
rect 29917 24769 29929 24803
rect 29963 24800 29975 24803
rect 30926 24800 30932 24812
rect 29963 24772 30932 24800
rect 29963 24769 29975 24772
rect 29917 24763 29975 24769
rect 28445 24735 28503 24741
rect 28445 24701 28457 24735
rect 28491 24701 28503 24735
rect 28445 24695 28503 24701
rect 27522 24624 27528 24676
rect 27580 24664 27586 24676
rect 29932 24664 29960 24763
rect 30926 24760 30932 24772
rect 30984 24760 30990 24812
rect 31036 24809 31064 24840
rect 32416 24840 33048 24868
rect 31021 24803 31079 24809
rect 31021 24769 31033 24803
rect 31067 24769 31079 24803
rect 31021 24763 31079 24769
rect 32214 24760 32220 24812
rect 32272 24800 32278 24812
rect 32416 24809 32444 24840
rect 33042 24828 33048 24840
rect 33100 24828 33106 24880
rect 32401 24803 32459 24809
rect 32401 24800 32413 24803
rect 32272 24772 32413 24800
rect 32272 24760 32278 24772
rect 32401 24769 32413 24772
rect 32447 24769 32459 24803
rect 32401 24763 32459 24769
rect 32582 24760 32588 24812
rect 32640 24800 32646 24812
rect 32749 24803 32807 24809
rect 32749 24800 32761 24803
rect 32640 24772 32761 24800
rect 32640 24760 32646 24772
rect 32749 24769 32761 24772
rect 32795 24769 32807 24803
rect 32749 24763 32807 24769
rect 30006 24692 30012 24744
rect 30064 24692 30070 24744
rect 30285 24735 30343 24741
rect 30285 24701 30297 24735
rect 30331 24701 30343 24735
rect 30285 24695 30343 24701
rect 27580 24636 29960 24664
rect 27580 24624 27586 24636
rect 23308 24568 25360 24596
rect 25406 24556 25412 24608
rect 25464 24596 25470 24608
rect 27798 24596 27804 24608
rect 25464 24568 27804 24596
rect 25464 24556 25470 24568
rect 27798 24556 27804 24568
rect 27856 24556 27862 24608
rect 29086 24556 29092 24608
rect 29144 24596 29150 24608
rect 30024 24596 30052 24692
rect 30300 24664 30328 24695
rect 30650 24692 30656 24744
rect 30708 24692 30714 24744
rect 30742 24692 30748 24744
rect 30800 24692 30806 24744
rect 31113 24735 31171 24741
rect 31113 24701 31125 24735
rect 31159 24732 31171 24735
rect 31294 24732 31300 24744
rect 31159 24704 31300 24732
rect 31159 24701 31171 24704
rect 31113 24695 31171 24701
rect 31294 24692 31300 24704
rect 31352 24692 31358 24744
rect 31386 24692 31392 24744
rect 31444 24692 31450 24744
rect 32493 24735 32551 24741
rect 32493 24732 32505 24735
rect 32232 24704 32505 24732
rect 31404 24664 31432 24692
rect 30300 24636 31432 24664
rect 29144 24568 30052 24596
rect 29144 24556 29150 24568
rect 30374 24556 30380 24608
rect 30432 24596 30438 24608
rect 32232 24605 32260 24704
rect 32493 24701 32505 24704
rect 32539 24701 32551 24735
rect 32493 24695 32551 24701
rect 32217 24599 32275 24605
rect 32217 24596 32229 24599
rect 30432 24568 32229 24596
rect 30432 24556 30438 24568
rect 32217 24565 32229 24568
rect 32263 24565 32275 24599
rect 32217 24559 32275 24565
rect 1104 24506 36800 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 36800 24506
rect 1104 24432 36800 24454
rect 3326 24352 3332 24404
rect 3384 24392 3390 24404
rect 3384 24364 8800 24392
rect 3384 24352 3390 24364
rect 2498 24284 2504 24336
rect 2556 24324 2562 24336
rect 2777 24327 2835 24333
rect 2777 24324 2789 24327
rect 2556 24296 2789 24324
rect 2556 24284 2562 24296
rect 2777 24293 2789 24296
rect 2823 24293 2835 24327
rect 2777 24287 2835 24293
rect 2792 24256 2820 24287
rect 5258 24284 5264 24336
rect 5316 24324 5322 24336
rect 5445 24327 5503 24333
rect 5445 24324 5457 24327
rect 5316 24296 5457 24324
rect 5316 24284 5322 24296
rect 5445 24293 5457 24296
rect 5491 24293 5503 24327
rect 5445 24287 5503 24293
rect 4985 24259 5043 24265
rect 4985 24256 4997 24259
rect 2792 24228 4997 24256
rect 4985 24225 4997 24228
rect 5031 24256 5043 24259
rect 5166 24256 5172 24268
rect 5031 24228 5172 24256
rect 5031 24225 5043 24228
rect 4985 24219 5043 24225
rect 5166 24216 5172 24228
rect 5224 24216 5230 24268
rect 5718 24216 5724 24268
rect 5776 24216 5782 24268
rect 7282 24216 7288 24268
rect 7340 24216 7346 24268
rect 8772 24265 8800 24364
rect 11238 24352 11244 24404
rect 11296 24392 11302 24404
rect 11517 24395 11575 24401
rect 11517 24392 11529 24395
rect 11296 24364 11529 24392
rect 11296 24352 11302 24364
rect 11517 24361 11529 24364
rect 11563 24361 11575 24395
rect 11517 24355 11575 24361
rect 12342 24352 12348 24404
rect 12400 24352 12406 24404
rect 14826 24392 14832 24404
rect 12544 24364 14832 24392
rect 11425 24327 11483 24333
rect 11425 24293 11437 24327
rect 11471 24324 11483 24327
rect 11698 24324 11704 24336
rect 11471 24296 11704 24324
rect 11471 24293 11483 24296
rect 11425 24287 11483 24293
rect 11698 24284 11704 24296
rect 11756 24284 11762 24336
rect 12544 24324 12572 24364
rect 14826 24352 14832 24364
rect 14884 24352 14890 24404
rect 17954 24352 17960 24404
rect 18012 24392 18018 24404
rect 18049 24395 18107 24401
rect 18049 24392 18061 24395
rect 18012 24364 18061 24392
rect 18012 24352 18018 24364
rect 18049 24361 18061 24364
rect 18095 24361 18107 24395
rect 18049 24355 18107 24361
rect 18598 24352 18604 24404
rect 18656 24352 18662 24404
rect 21266 24352 21272 24404
rect 21324 24352 21330 24404
rect 21818 24352 21824 24404
rect 21876 24352 21882 24404
rect 22094 24352 22100 24404
rect 22152 24392 22158 24404
rect 23106 24392 23112 24404
rect 22152 24364 23112 24392
rect 22152 24352 22158 24364
rect 23106 24352 23112 24364
rect 23164 24352 23170 24404
rect 23566 24352 23572 24404
rect 23624 24392 23630 24404
rect 23661 24395 23719 24401
rect 23661 24392 23673 24395
rect 23624 24364 23673 24392
rect 23624 24352 23630 24364
rect 23661 24361 23673 24364
rect 23707 24361 23719 24395
rect 23661 24355 23719 24361
rect 23934 24352 23940 24404
rect 23992 24392 23998 24404
rect 28445 24395 28503 24401
rect 28445 24392 28457 24395
rect 23992 24364 28457 24392
rect 23992 24352 23998 24364
rect 28445 24361 28457 24364
rect 28491 24361 28503 24395
rect 28445 24355 28503 24361
rect 32401 24395 32459 24401
rect 32401 24361 32413 24395
rect 32447 24392 32459 24395
rect 32582 24392 32588 24404
rect 32447 24364 32588 24392
rect 32447 24361 32459 24364
rect 32401 24355 32459 24361
rect 32582 24352 32588 24364
rect 32640 24352 32646 24404
rect 12406 24296 12572 24324
rect 12621 24327 12679 24333
rect 8757 24259 8815 24265
rect 8757 24225 8769 24259
rect 8803 24256 8815 24259
rect 8941 24259 8999 24265
rect 8941 24256 8953 24259
rect 8803 24228 8953 24256
rect 8803 24225 8815 24228
rect 8757 24219 8815 24225
rect 8941 24225 8953 24228
rect 8987 24225 8999 24259
rect 8941 24219 8999 24225
rect 11057 24259 11115 24265
rect 11057 24225 11069 24259
rect 11103 24256 11115 24259
rect 12406 24256 12434 24296
rect 12621 24293 12633 24327
rect 12667 24293 12679 24327
rect 12621 24287 12679 24293
rect 11103 24228 12434 24256
rect 11103 24225 11115 24228
rect 11057 24219 11115 24225
rect 1397 24191 1455 24197
rect 1397 24157 1409 24191
rect 1443 24188 1455 24191
rect 2958 24188 2964 24200
rect 1443 24160 2964 24188
rect 1443 24157 1455 24160
rect 1397 24151 1455 24157
rect 2958 24148 2964 24160
rect 3016 24148 3022 24200
rect 4798 24148 4804 24200
rect 4856 24148 4862 24200
rect 5810 24148 5816 24200
rect 5868 24197 5874 24200
rect 5868 24191 5896 24197
rect 5884 24157 5896 24191
rect 5868 24151 5896 24157
rect 5868 24148 5874 24151
rect 5994 24148 6000 24200
rect 6052 24148 6058 24200
rect 7006 24148 7012 24200
rect 7064 24148 7070 24200
rect 7098 24148 7104 24200
rect 7156 24148 7162 24200
rect 7374 24148 7380 24200
rect 7432 24148 7438 24200
rect 8573 24191 8631 24197
rect 8573 24157 8585 24191
rect 8619 24188 8631 24191
rect 8662 24188 8668 24200
rect 8619 24160 8668 24188
rect 8619 24157 8631 24160
rect 8573 24151 8631 24157
rect 8662 24148 8668 24160
rect 8720 24148 8726 24200
rect 12529 24191 12587 24197
rect 12529 24157 12541 24191
rect 12575 24188 12587 24191
rect 12636 24188 12664 24287
rect 12894 24216 12900 24268
rect 12952 24256 12958 24268
rect 13078 24256 13084 24268
rect 12952 24228 13084 24256
rect 12952 24216 12958 24228
rect 13078 24216 13084 24228
rect 13136 24216 13142 24268
rect 13265 24259 13323 24265
rect 13265 24225 13277 24259
rect 13311 24225 13323 24259
rect 14844 24256 14872 24352
rect 17862 24284 17868 24336
rect 17920 24284 17926 24336
rect 18506 24284 18512 24336
rect 18564 24284 18570 24336
rect 21177 24327 21235 24333
rect 21177 24293 21189 24327
rect 21223 24324 21235 24327
rect 21358 24324 21364 24336
rect 21223 24296 21364 24324
rect 21223 24293 21235 24296
rect 21177 24287 21235 24293
rect 21358 24284 21364 24296
rect 21416 24284 21422 24336
rect 21634 24284 21640 24336
rect 21692 24284 21698 24336
rect 25314 24324 25320 24336
rect 21744 24296 25320 24324
rect 17589 24259 17647 24265
rect 17589 24256 17601 24259
rect 14844 24228 17601 24256
rect 13265 24219 13323 24225
rect 17589 24225 17601 24228
rect 17635 24256 17647 24259
rect 17635 24228 21404 24256
rect 17635 24225 17647 24228
rect 17589 24219 17647 24225
rect 12575 24160 12664 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 12986 24148 12992 24200
rect 13044 24148 13050 24200
rect 13280 24188 13308 24219
rect 16482 24188 16488 24200
rect 13280 24160 16488 24188
rect 1664 24123 1722 24129
rect 1664 24089 1676 24123
rect 1710 24120 1722 24123
rect 1762 24120 1768 24132
rect 1710 24092 1768 24120
rect 1710 24089 1722 24092
rect 1664 24083 1722 24089
rect 1762 24080 1768 24092
rect 1820 24080 1826 24132
rect 8846 24080 8852 24132
rect 8904 24120 8910 24132
rect 9186 24123 9244 24129
rect 9186 24120 9198 24123
rect 8904 24092 9198 24120
rect 8904 24080 8910 24092
rect 9186 24089 9198 24092
rect 9232 24089 9244 24123
rect 9186 24083 9244 24089
rect 9306 24080 9312 24132
rect 9364 24120 9370 24132
rect 12618 24120 12624 24132
rect 9364 24092 12624 24120
rect 9364 24080 9370 24092
rect 12618 24080 12624 24092
rect 12676 24080 12682 24132
rect 12710 24080 12716 24132
rect 12768 24120 12774 24132
rect 13280 24120 13308 24160
rect 16482 24148 16488 24160
rect 16540 24148 16546 24200
rect 16942 24148 16948 24200
rect 17000 24188 17006 24200
rect 20438 24188 20444 24200
rect 17000 24160 20444 24188
rect 17000 24148 17006 24160
rect 20438 24148 20444 24160
rect 20496 24148 20502 24200
rect 21376 24197 21404 24228
rect 21450 24216 21456 24268
rect 21508 24256 21514 24268
rect 21744 24256 21772 24296
rect 25314 24284 25320 24296
rect 25372 24284 25378 24336
rect 25406 24284 25412 24336
rect 25464 24284 25470 24336
rect 32214 24324 32220 24336
rect 31726 24296 32220 24324
rect 21508 24228 21772 24256
rect 21508 24216 21514 24228
rect 24670 24216 24676 24268
rect 24728 24216 24734 24268
rect 25424 24256 25452 24284
rect 24780 24228 25881 24256
rect 21361 24191 21419 24197
rect 21361 24157 21373 24191
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 21913 24191 21971 24197
rect 21913 24157 21925 24191
rect 21959 24188 21971 24191
rect 22281 24191 22339 24197
rect 22281 24188 22293 24191
rect 21959 24160 22293 24188
rect 21959 24157 21971 24160
rect 21913 24151 21971 24157
rect 22281 24157 22293 24160
rect 22327 24188 22339 24191
rect 22462 24188 22468 24200
rect 22327 24160 22468 24188
rect 22327 24157 22339 24160
rect 22281 24151 22339 24157
rect 12768 24092 13308 24120
rect 12768 24080 12774 24092
rect 17126 24080 17132 24132
rect 17184 24120 17190 24132
rect 17586 24120 17592 24132
rect 17184 24092 17592 24120
rect 17184 24080 17190 24092
rect 17586 24080 17592 24092
rect 17644 24080 17650 24132
rect 18141 24123 18199 24129
rect 18141 24089 18153 24123
rect 18187 24120 18199 24123
rect 20809 24123 20867 24129
rect 20809 24120 20821 24123
rect 18187 24092 20821 24120
rect 18187 24089 18199 24092
rect 18141 24083 18199 24089
rect 20809 24089 20821 24092
rect 20855 24089 20867 24123
rect 21376 24120 21404 24151
rect 22462 24148 22468 24160
rect 22520 24148 22526 24200
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24188 22615 24191
rect 23198 24188 23204 24200
rect 22603 24160 23204 24188
rect 22603 24157 22615 24160
rect 22557 24151 22615 24157
rect 22572 24120 22600 24151
rect 23198 24148 23204 24160
rect 23256 24148 23262 24200
rect 23382 24148 23388 24200
rect 23440 24148 23446 24200
rect 23474 24148 23480 24200
rect 23532 24148 23538 24200
rect 23750 24148 23756 24200
rect 23808 24148 23814 24200
rect 23934 24148 23940 24200
rect 23992 24188 23998 24200
rect 24780 24188 24808 24228
rect 23992 24160 24808 24188
rect 23992 24148 23998 24160
rect 24854 24148 24860 24200
rect 24912 24148 24918 24200
rect 25590 24148 25596 24200
rect 25648 24148 25654 24200
rect 25682 24148 25688 24200
rect 25740 24197 25746 24200
rect 25853 24197 25881 24228
rect 26234 24216 26240 24268
rect 26292 24256 26298 24268
rect 27249 24259 27307 24265
rect 27249 24256 27261 24259
rect 26292 24228 27261 24256
rect 26292 24216 26298 24228
rect 27249 24225 27261 24228
rect 27295 24225 27307 24259
rect 27249 24219 27307 24225
rect 27522 24216 27528 24268
rect 27580 24216 27586 24268
rect 27663 24259 27721 24265
rect 27663 24225 27675 24259
rect 27709 24256 27721 24259
rect 27982 24256 27988 24268
rect 27709 24228 27988 24256
rect 27709 24225 27721 24228
rect 27663 24219 27721 24225
rect 27982 24216 27988 24228
rect 28040 24216 28046 24268
rect 28166 24216 28172 24268
rect 28224 24256 28230 24268
rect 31726 24256 31754 24296
rect 32214 24284 32220 24296
rect 32272 24284 32278 24336
rect 28224 24228 31754 24256
rect 28224 24216 28230 24228
rect 25740 24191 25768 24197
rect 25756 24157 25768 24191
rect 25853 24191 25927 24197
rect 25853 24160 25881 24191
rect 25740 24151 25768 24157
rect 25869 24157 25881 24160
rect 25915 24157 25927 24191
rect 25869 24151 25927 24157
rect 26605 24191 26663 24197
rect 26605 24157 26617 24191
rect 26651 24157 26663 24191
rect 26605 24151 26663 24157
rect 25740 24148 25746 24151
rect 21376 24092 22600 24120
rect 20809 24083 20867 24089
rect 6638 24012 6644 24064
rect 6696 24012 6702 24064
rect 6730 24012 6736 24064
rect 6788 24052 6794 24064
rect 6825 24055 6883 24061
rect 6825 24052 6837 24055
rect 6788 24024 6837 24052
rect 6788 24012 6794 24024
rect 6825 24021 6837 24024
rect 6871 24021 6883 24055
rect 6825 24015 6883 24021
rect 9858 24012 9864 24064
rect 9916 24052 9922 24064
rect 10321 24055 10379 24061
rect 10321 24052 10333 24055
rect 9916 24024 10333 24052
rect 9916 24012 9922 24024
rect 10321 24021 10333 24024
rect 10367 24021 10379 24055
rect 12636 24052 12664 24080
rect 18156 24052 18184 24083
rect 12636 24024 18184 24052
rect 20824 24052 20852 24083
rect 21726 24052 21732 24064
rect 20824 24024 21732 24052
rect 10321 24015 10379 24021
rect 21726 24012 21732 24024
rect 21784 24012 21790 24064
rect 23014 24012 23020 24064
rect 23072 24052 23078 24064
rect 23201 24055 23259 24061
rect 23201 24052 23213 24055
rect 23072 24024 23213 24052
rect 23072 24012 23078 24024
rect 23201 24021 23213 24024
rect 23247 24021 23259 24055
rect 23201 24015 23259 24021
rect 24026 24012 24032 24064
rect 24084 24052 24090 24064
rect 26513 24055 26571 24061
rect 26513 24052 26525 24055
rect 24084 24024 26525 24052
rect 24084 24012 24090 24024
rect 26513 24021 26525 24024
rect 26559 24021 26571 24055
rect 26620 24052 26648 24151
rect 26786 24148 26792 24200
rect 26844 24148 26850 24200
rect 27798 24148 27804 24200
rect 27856 24148 27862 24200
rect 32122 24148 32128 24200
rect 32180 24188 32186 24200
rect 32585 24191 32643 24197
rect 32585 24188 32597 24191
rect 32180 24160 32597 24188
rect 32180 24148 32186 24160
rect 32585 24157 32597 24160
rect 32631 24157 32643 24191
rect 32585 24151 32643 24157
rect 36078 24148 36084 24200
rect 36136 24188 36142 24200
rect 36173 24191 36231 24197
rect 36173 24188 36185 24191
rect 36136 24160 36185 24188
rect 36136 24148 36142 24160
rect 36173 24157 36185 24160
rect 36219 24157 36231 24191
rect 36173 24151 36231 24157
rect 26970 24052 26976 24064
rect 26620 24024 26976 24052
rect 26513 24015 26571 24021
rect 26970 24012 26976 24024
rect 27028 24052 27034 24064
rect 28258 24052 28264 24064
rect 27028 24024 28264 24052
rect 27028 24012 27034 24024
rect 28258 24012 28264 24024
rect 28316 24012 28322 24064
rect 36354 24012 36360 24064
rect 36412 24012 36418 24064
rect 1104 23962 36800 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 36800 23962
rect 1104 23888 36800 23910
rect 1762 23808 1768 23860
rect 1820 23808 1826 23860
rect 2133 23851 2191 23857
rect 2133 23817 2145 23851
rect 2179 23817 2191 23851
rect 2133 23811 2191 23817
rect 1949 23715 2007 23721
rect 1949 23681 1961 23715
rect 1995 23712 2007 23715
rect 2148 23712 2176 23811
rect 2498 23808 2504 23860
rect 2556 23808 2562 23860
rect 7009 23851 7067 23857
rect 7009 23817 7021 23851
rect 7055 23848 7067 23851
rect 7282 23848 7288 23860
rect 7055 23820 7288 23848
rect 7055 23817 7067 23820
rect 7009 23811 7067 23817
rect 7282 23808 7288 23820
rect 7340 23808 7346 23860
rect 7558 23808 7564 23860
rect 7616 23808 7622 23860
rect 8487 23851 8545 23857
rect 8487 23817 8499 23851
rect 8533 23848 8545 23851
rect 8846 23848 8852 23860
rect 8533 23820 8852 23848
rect 8533 23817 8545 23820
rect 8487 23811 8545 23817
rect 8846 23808 8852 23820
rect 8904 23808 8910 23860
rect 9646 23820 11192 23848
rect 3142 23740 3148 23792
rect 3200 23780 3206 23792
rect 3200 23752 7236 23780
rect 3200 23740 3206 23752
rect 1995 23684 2176 23712
rect 2593 23715 2651 23721
rect 1995 23681 2007 23684
rect 1949 23675 2007 23681
rect 2593 23681 2605 23715
rect 2639 23712 2651 23715
rect 2866 23712 2872 23724
rect 2639 23684 2872 23712
rect 2639 23681 2651 23684
rect 2593 23675 2651 23681
rect 2866 23672 2872 23684
rect 2924 23672 2930 23724
rect 2958 23672 2964 23724
rect 3016 23672 3022 23724
rect 3228 23715 3286 23721
rect 3228 23681 3240 23715
rect 3274 23712 3286 23715
rect 3786 23712 3792 23724
rect 3274 23684 3792 23712
rect 3274 23681 3286 23684
rect 3228 23675 3286 23681
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23712 6607 23715
rect 7208 23712 7236 23752
rect 8386 23740 8392 23792
rect 8444 23740 8450 23792
rect 9646 23780 9674 23820
rect 8680 23752 9674 23780
rect 11164 23780 11192 23820
rect 11514 23808 11520 23860
rect 11572 23848 11578 23860
rect 11701 23851 11759 23857
rect 11701 23848 11713 23851
rect 11572 23820 11713 23848
rect 11572 23808 11578 23820
rect 11701 23817 11713 23820
rect 11747 23848 11759 23851
rect 13814 23848 13820 23860
rect 11747 23820 13820 23848
rect 11747 23817 11759 23820
rect 11701 23811 11759 23817
rect 13814 23808 13820 23820
rect 13872 23848 13878 23860
rect 13872 23820 14412 23848
rect 13872 23808 13878 23820
rect 12710 23780 12716 23792
rect 11164 23752 12716 23780
rect 6595 23684 7144 23712
rect 7208 23684 8530 23712
rect 6595 23681 6607 23684
rect 6549 23675 6607 23681
rect 2682 23604 2688 23656
rect 2740 23604 2746 23656
rect 6638 23604 6644 23656
rect 6696 23644 6702 23656
rect 7116 23653 7144 23684
rect 7101 23647 7159 23653
rect 6696 23616 7052 23644
rect 6696 23604 6702 23616
rect 6178 23536 6184 23588
rect 6236 23576 6242 23588
rect 6825 23579 6883 23585
rect 6825 23576 6837 23579
rect 6236 23548 6837 23576
rect 6236 23536 6242 23548
rect 6825 23545 6837 23548
rect 6871 23545 6883 23579
rect 7024 23576 7052 23616
rect 7101 23613 7113 23647
rect 7147 23644 7159 23647
rect 8502 23644 8530 23684
rect 8570 23672 8576 23724
rect 8628 23672 8634 23724
rect 8680 23721 8708 23752
rect 9048 23721 9076 23752
rect 12710 23740 12716 23752
rect 12768 23740 12774 23792
rect 14384 23780 14412 23820
rect 14458 23808 14464 23860
rect 14516 23808 14522 23860
rect 17770 23848 17776 23860
rect 16868 23820 17776 23848
rect 16868 23780 16896 23820
rect 17770 23808 17776 23820
rect 17828 23808 17834 23860
rect 17862 23808 17868 23860
rect 17920 23848 17926 23860
rect 18509 23851 18567 23857
rect 18509 23848 18521 23851
rect 17920 23820 18521 23848
rect 17920 23808 17926 23820
rect 18509 23817 18521 23820
rect 18555 23817 18567 23851
rect 18509 23811 18567 23817
rect 20438 23808 20444 23860
rect 20496 23848 20502 23860
rect 21450 23848 21456 23860
rect 20496 23820 21456 23848
rect 20496 23808 20502 23820
rect 21450 23808 21456 23820
rect 21508 23808 21514 23860
rect 21634 23808 21640 23860
rect 21692 23808 21698 23860
rect 21726 23808 21732 23860
rect 21784 23848 21790 23860
rect 22373 23851 22431 23857
rect 22373 23848 22385 23851
rect 21784 23820 22385 23848
rect 21784 23808 21790 23820
rect 22373 23817 22385 23820
rect 22419 23848 22431 23851
rect 22419 23820 23152 23848
rect 22419 23817 22431 23820
rect 22373 23811 22431 23817
rect 14384 23752 16896 23780
rect 19978 23740 19984 23792
rect 20036 23740 20042 23792
rect 23124 23789 23152 23820
rect 23382 23808 23388 23860
rect 23440 23848 23446 23860
rect 23569 23851 23627 23857
rect 23569 23848 23581 23851
rect 23440 23820 23581 23848
rect 23440 23808 23446 23820
rect 23569 23817 23581 23820
rect 23615 23817 23627 23851
rect 23569 23811 23627 23817
rect 24854 23808 24860 23860
rect 24912 23848 24918 23860
rect 26142 23848 26148 23860
rect 24912 23820 26148 23848
rect 24912 23808 24918 23820
rect 26142 23808 26148 23820
rect 26200 23808 26206 23860
rect 27982 23808 27988 23860
rect 28040 23848 28046 23860
rect 29914 23848 29920 23860
rect 28040 23820 29920 23848
rect 28040 23808 28046 23820
rect 29914 23808 29920 23820
rect 29972 23848 29978 23860
rect 30285 23851 30343 23857
rect 30285 23848 30297 23851
rect 29972 23820 30297 23848
rect 29972 23808 29978 23820
rect 30285 23817 30297 23820
rect 30331 23817 30343 23851
rect 33226 23848 33232 23860
rect 30285 23811 30343 23817
rect 31726 23820 33232 23848
rect 23109 23783 23167 23789
rect 23109 23749 23121 23783
rect 23155 23749 23167 23783
rect 23109 23743 23167 23749
rect 23198 23740 23204 23792
rect 23256 23780 23262 23792
rect 23661 23783 23719 23789
rect 23661 23780 23673 23783
rect 23256 23752 23673 23780
rect 23256 23740 23262 23752
rect 23661 23749 23673 23752
rect 23707 23749 23719 23783
rect 23661 23743 23719 23749
rect 8665 23715 8723 23721
rect 8665 23681 8677 23715
rect 8711 23681 8723 23715
rect 8665 23675 8723 23681
rect 9033 23715 9091 23721
rect 9033 23681 9045 23715
rect 9079 23681 9091 23715
rect 9033 23675 9091 23681
rect 8680 23644 8708 23675
rect 9122 23672 9128 23724
rect 9180 23672 9186 23724
rect 9217 23715 9275 23721
rect 9217 23681 9229 23715
rect 9263 23712 9275 23715
rect 9493 23715 9551 23721
rect 9493 23712 9505 23715
rect 9263 23684 9505 23712
rect 9263 23681 9275 23684
rect 9217 23675 9275 23681
rect 9493 23681 9505 23684
rect 9539 23712 9551 23715
rect 9858 23712 9864 23724
rect 9539 23684 9864 23712
rect 9539 23681 9551 23684
rect 9493 23675 9551 23681
rect 9858 23672 9864 23684
rect 9916 23672 9922 23724
rect 11606 23672 11612 23724
rect 11664 23672 11670 23724
rect 11882 23672 11888 23724
rect 11940 23672 11946 23724
rect 12526 23672 12532 23724
rect 12584 23712 12590 23724
rect 12621 23715 12679 23721
rect 12621 23712 12633 23715
rect 12584 23684 12633 23712
rect 12584 23672 12590 23684
rect 12621 23681 12633 23684
rect 12667 23712 12679 23715
rect 12986 23712 12992 23724
rect 12667 23684 12992 23712
rect 12667 23681 12679 23684
rect 12621 23675 12679 23681
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 13814 23672 13820 23724
rect 13872 23672 13878 23724
rect 15010 23672 15016 23724
rect 15068 23712 15074 23724
rect 15105 23715 15163 23721
rect 15105 23712 15117 23715
rect 15068 23684 15117 23712
rect 15068 23672 15074 23684
rect 15105 23681 15117 23684
rect 15151 23681 15163 23715
rect 15105 23675 15163 23681
rect 15372 23715 15430 23721
rect 15372 23681 15384 23715
rect 15418 23712 15430 23715
rect 15654 23712 15660 23724
rect 15418 23684 15660 23712
rect 15418 23681 15430 23684
rect 15372 23675 15430 23681
rect 15654 23672 15660 23684
rect 15712 23672 15718 23724
rect 17586 23672 17592 23724
rect 17644 23672 17650 23724
rect 17862 23672 17868 23724
rect 17920 23672 17926 23724
rect 19337 23715 19395 23721
rect 19337 23681 19349 23715
rect 19383 23681 19395 23715
rect 19337 23675 19395 23681
rect 19429 23715 19487 23721
rect 19429 23681 19441 23715
rect 19475 23712 19487 23715
rect 19702 23712 19708 23724
rect 19475 23684 19708 23712
rect 19475 23681 19487 23684
rect 19429 23675 19487 23681
rect 7147 23616 8156 23644
rect 8502 23616 8708 23644
rect 9677 23647 9735 23653
rect 7147 23613 7159 23616
rect 7101 23607 7159 23613
rect 7377 23579 7435 23585
rect 7377 23576 7389 23579
rect 7024 23548 7389 23576
rect 6825 23539 6883 23545
rect 7377 23545 7389 23548
rect 7423 23545 7435 23579
rect 8128 23576 8156 23616
rect 9677 23613 9689 23647
rect 9723 23644 9735 23647
rect 10042 23644 10048 23656
rect 9723 23616 10048 23644
rect 9723 23613 9735 23616
rect 9677 23607 9735 23613
rect 10042 23604 10048 23616
rect 10100 23604 10106 23656
rect 10410 23604 10416 23656
rect 10468 23604 10474 23656
rect 10594 23653 10600 23656
rect 10551 23647 10600 23653
rect 10551 23613 10563 23647
rect 10597 23613 10600 23647
rect 10551 23607 10600 23613
rect 10594 23604 10600 23607
rect 10652 23604 10658 23656
rect 10686 23604 10692 23656
rect 10744 23604 10750 23656
rect 11054 23604 11060 23656
rect 11112 23604 11118 23656
rect 12805 23647 12863 23653
rect 12805 23613 12817 23647
rect 12851 23644 12863 23647
rect 12894 23644 12900 23656
rect 12851 23616 12900 23644
rect 12851 23613 12863 23616
rect 12805 23607 12863 23613
rect 12894 23604 12900 23616
rect 12952 23604 12958 23656
rect 13170 23604 13176 23656
rect 13228 23644 13234 23656
rect 13541 23647 13599 23653
rect 13541 23644 13553 23647
rect 13228 23616 13553 23644
rect 13228 23604 13234 23616
rect 13541 23613 13553 23616
rect 13587 23613 13599 23647
rect 13541 23607 13599 23613
rect 13630 23604 13636 23656
rect 13688 23653 13694 23656
rect 13688 23647 13716 23653
rect 13704 23613 13716 23647
rect 13688 23607 13716 23613
rect 13688 23604 13694 23607
rect 16206 23604 16212 23656
rect 16264 23644 16270 23656
rect 16669 23647 16727 23653
rect 16669 23644 16681 23647
rect 16264 23616 16681 23644
rect 16264 23604 16270 23616
rect 16669 23613 16681 23616
rect 16715 23613 16727 23647
rect 16669 23607 16727 23613
rect 16758 23604 16764 23656
rect 16816 23644 16822 23656
rect 16853 23647 16911 23653
rect 16853 23644 16865 23647
rect 16816 23616 16865 23644
rect 16816 23604 16822 23616
rect 16853 23613 16865 23616
rect 16899 23613 16911 23647
rect 17706 23647 17764 23653
rect 17706 23644 17718 23647
rect 16853 23607 16911 23613
rect 17420 23616 17718 23644
rect 9306 23576 9312 23588
rect 8128 23548 9312 23576
rect 7377 23539 7435 23545
rect 9306 23536 9312 23548
rect 9364 23536 9370 23588
rect 10137 23579 10195 23585
rect 10137 23545 10149 23579
rect 10183 23576 10195 23579
rect 10226 23576 10232 23588
rect 10183 23548 10232 23576
rect 10183 23545 10195 23548
rect 10137 23539 10195 23545
rect 10226 23536 10232 23548
rect 10284 23536 10290 23588
rect 11072 23576 11100 23604
rect 13265 23579 13323 23585
rect 11072 23548 12112 23576
rect 4341 23511 4399 23517
rect 4341 23477 4353 23511
rect 4387 23508 4399 23511
rect 4706 23508 4712 23520
rect 4387 23480 4712 23508
rect 4387 23477 4399 23480
rect 4341 23471 4399 23477
rect 4706 23468 4712 23480
rect 4764 23508 4770 23520
rect 5810 23508 5816 23520
rect 4764 23480 5816 23508
rect 4764 23468 4770 23480
rect 5810 23468 5816 23480
rect 5868 23468 5874 23520
rect 8570 23468 8576 23520
rect 8628 23508 8634 23520
rect 8938 23508 8944 23520
rect 8628 23480 8944 23508
rect 8628 23468 8634 23480
rect 8938 23468 8944 23480
rect 8996 23468 9002 23520
rect 10410 23468 10416 23520
rect 10468 23508 10474 23520
rect 10778 23508 10784 23520
rect 10468 23480 10784 23508
rect 10468 23468 10474 23480
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 10870 23468 10876 23520
rect 10928 23508 10934 23520
rect 12084 23517 12112 23548
rect 13265 23545 13277 23579
rect 13311 23545 13323 23579
rect 16942 23576 16948 23588
rect 13265 23539 13323 23545
rect 16040 23548 16948 23576
rect 11333 23511 11391 23517
rect 11333 23508 11345 23511
rect 10928 23480 11345 23508
rect 10928 23468 10934 23480
rect 11333 23477 11345 23480
rect 11379 23477 11391 23511
rect 11333 23471 11391 23477
rect 12069 23511 12127 23517
rect 12069 23477 12081 23511
rect 12115 23508 12127 23511
rect 13280 23508 13308 23539
rect 16040 23508 16068 23548
rect 16942 23536 16948 23548
rect 17000 23576 17006 23588
rect 17313 23579 17371 23585
rect 17313 23576 17325 23579
rect 17000 23548 17325 23576
rect 17000 23536 17006 23548
rect 17313 23545 17325 23548
rect 17359 23545 17371 23579
rect 17313 23539 17371 23545
rect 12115 23480 16068 23508
rect 12115 23477 12127 23480
rect 12069 23471 12127 23477
rect 16206 23468 16212 23520
rect 16264 23508 16270 23520
rect 16485 23511 16543 23517
rect 16485 23508 16497 23511
rect 16264 23480 16497 23508
rect 16264 23468 16270 23480
rect 16485 23477 16497 23480
rect 16531 23477 16543 23511
rect 16485 23471 16543 23477
rect 17218 23468 17224 23520
rect 17276 23508 17282 23520
rect 17420 23508 17448 23616
rect 17706 23613 17718 23616
rect 17752 23613 17764 23647
rect 17880 23644 17908 23672
rect 17880 23616 19288 23644
rect 17706 23607 17764 23613
rect 17276 23480 17448 23508
rect 17276 23468 17282 23480
rect 18966 23468 18972 23520
rect 19024 23468 19030 23520
rect 19260 23508 19288 23616
rect 19352 23576 19380 23675
rect 19702 23672 19708 23684
rect 19760 23672 19766 23724
rect 19794 23672 19800 23724
rect 19852 23712 19858 23724
rect 19996 23712 20024 23740
rect 19852 23684 20024 23712
rect 19852 23672 19858 23684
rect 20714 23672 20720 23724
rect 20772 23672 20778 23724
rect 22281 23715 22339 23721
rect 22281 23681 22293 23715
rect 22327 23712 22339 23715
rect 22462 23712 22468 23724
rect 22327 23684 22468 23712
rect 22327 23681 22339 23684
rect 22281 23675 22339 23681
rect 22462 23672 22468 23684
rect 22520 23672 22526 23724
rect 22830 23672 22836 23724
rect 22888 23712 22894 23724
rect 22888 23684 24164 23712
rect 22888 23672 22894 23684
rect 19610 23604 19616 23656
rect 19668 23604 19674 23656
rect 19981 23647 20039 23653
rect 19981 23613 19993 23647
rect 20027 23644 20039 23647
rect 20070 23644 20076 23656
rect 20027 23616 20076 23644
rect 20027 23613 20039 23616
rect 19981 23607 20039 23613
rect 20070 23604 20076 23616
rect 20128 23604 20134 23656
rect 20806 23644 20812 23656
rect 20864 23653 20870 23656
rect 20864 23647 20892 23653
rect 20272 23616 20812 23644
rect 19886 23576 19892 23588
rect 19352 23548 19892 23576
rect 19886 23536 19892 23548
rect 19944 23576 19950 23588
rect 20272 23576 20300 23616
rect 20806 23604 20812 23616
rect 20880 23613 20892 23647
rect 20864 23607 20892 23613
rect 20993 23647 21051 23653
rect 20993 23613 21005 23647
rect 21039 23644 21051 23647
rect 23934 23644 23940 23656
rect 21039 23616 23940 23644
rect 21039 23613 21051 23616
rect 20993 23607 21051 23613
rect 20864 23604 20870 23607
rect 19944 23548 20300 23576
rect 19944 23536 19950 23548
rect 20438 23536 20444 23588
rect 20496 23536 20502 23588
rect 21376 23508 21404 23616
rect 23934 23604 23940 23616
rect 23992 23604 23998 23656
rect 24136 23653 24164 23684
rect 24670 23672 24676 23724
rect 24728 23672 24734 23724
rect 24872 23721 24900 23808
rect 26786 23740 26792 23792
rect 26844 23780 26850 23792
rect 31726 23780 31754 23820
rect 33226 23808 33232 23820
rect 33284 23848 33290 23860
rect 33413 23851 33471 23857
rect 33413 23848 33425 23851
rect 33284 23820 33425 23848
rect 33284 23808 33290 23820
rect 33413 23817 33425 23820
rect 33459 23817 33471 23851
rect 33413 23811 33471 23817
rect 26844 23752 27200 23780
rect 26844 23740 26850 23752
rect 24857 23715 24915 23721
rect 24857 23681 24869 23715
rect 24903 23681 24915 23715
rect 24857 23675 24915 23681
rect 25590 23672 25596 23724
rect 25648 23672 25654 23724
rect 25682 23672 25688 23724
rect 25740 23721 25746 23724
rect 25740 23715 25768 23721
rect 25756 23681 25768 23715
rect 25740 23675 25768 23681
rect 25740 23672 25746 23675
rect 26970 23672 26976 23724
rect 27028 23672 27034 23724
rect 27172 23721 27200 23752
rect 28920 23752 31754 23780
rect 28920 23724 28948 23752
rect 33042 23740 33048 23792
rect 33100 23780 33106 23792
rect 33321 23783 33379 23789
rect 33321 23780 33333 23783
rect 33100 23752 33333 23780
rect 33100 23740 33106 23752
rect 33321 23749 33333 23752
rect 33367 23749 33379 23783
rect 33321 23743 33379 23749
rect 27157 23715 27215 23721
rect 27157 23681 27169 23715
rect 27203 23681 27215 23715
rect 27157 23675 27215 23681
rect 24121 23647 24179 23653
rect 24121 23613 24133 23647
rect 24167 23613 24179 23647
rect 24121 23607 24179 23613
rect 25869 23647 25927 23653
rect 25869 23613 25881 23647
rect 25915 23644 25927 23647
rect 26050 23644 26056 23656
rect 25915 23616 26056 23644
rect 25915 23613 25927 23616
rect 25869 23607 25927 23613
rect 26050 23604 26056 23616
rect 26108 23644 26114 23656
rect 27172 23644 27200 23675
rect 27890 23672 27896 23724
rect 27948 23672 27954 23724
rect 27982 23672 27988 23724
rect 28040 23721 28046 23724
rect 28040 23715 28068 23721
rect 28056 23681 28068 23715
rect 28040 23675 28068 23681
rect 28040 23672 28046 23675
rect 28902 23672 28908 23724
rect 28960 23672 28966 23724
rect 29178 23721 29184 23724
rect 29172 23675 29184 23721
rect 29178 23672 29184 23675
rect 29236 23672 29242 23724
rect 27522 23644 27528 23656
rect 26108 23616 26740 23644
rect 27172 23616 27528 23644
rect 26108 23604 26114 23616
rect 23382 23536 23388 23588
rect 23440 23536 23446 23588
rect 24026 23536 24032 23588
rect 24084 23536 24090 23588
rect 25314 23536 25320 23588
rect 25372 23536 25378 23588
rect 19260 23480 21404 23508
rect 21542 23468 21548 23520
rect 21600 23508 21606 23520
rect 22278 23508 22284 23520
rect 21600 23480 22284 23508
rect 21600 23468 21606 23480
rect 22278 23468 22284 23480
rect 22336 23468 22342 23520
rect 25130 23468 25136 23520
rect 25188 23508 25194 23520
rect 26513 23511 26571 23517
rect 26513 23508 26525 23511
rect 25188 23480 26525 23508
rect 25188 23468 25194 23480
rect 26513 23477 26525 23480
rect 26559 23477 26571 23511
rect 26712 23508 26740 23616
rect 27522 23604 27528 23616
rect 27580 23604 27586 23656
rect 28169 23647 28227 23653
rect 28169 23644 28181 23647
rect 27724 23616 28181 23644
rect 27614 23536 27620 23588
rect 27672 23536 27678 23588
rect 27724 23508 27752 23616
rect 28169 23613 28181 23616
rect 28215 23613 28227 23647
rect 28169 23607 28227 23613
rect 26712 23480 27752 23508
rect 26513 23471 26571 23477
rect 27982 23468 27988 23520
rect 28040 23508 28046 23520
rect 28813 23511 28871 23517
rect 28813 23508 28825 23511
rect 28040 23480 28825 23508
rect 28040 23468 28046 23480
rect 28813 23477 28825 23480
rect 28859 23477 28871 23511
rect 28813 23471 28871 23477
rect 1104 23418 36800 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 36800 23418
rect 1104 23344 36800 23366
rect 3786 23264 3792 23316
rect 3844 23264 3850 23316
rect 10962 23304 10968 23316
rect 10520 23276 10968 23304
rect 2869 23239 2927 23245
rect 2869 23205 2881 23239
rect 2915 23205 2927 23239
rect 3602 23236 3608 23248
rect 2869 23199 2927 23205
rect 3344 23208 3608 23236
rect 2884 23100 2912 23199
rect 3344 23177 3372 23208
rect 3602 23196 3608 23208
rect 3660 23236 3666 23248
rect 4062 23236 4068 23248
rect 3660 23208 4068 23236
rect 3660 23196 3666 23208
rect 4062 23196 4068 23208
rect 4120 23196 4126 23248
rect 4338 23196 4344 23248
rect 4396 23236 4402 23248
rect 5077 23239 5135 23245
rect 5077 23236 5089 23239
rect 4396 23208 5089 23236
rect 4396 23196 4402 23208
rect 5077 23205 5089 23208
rect 5123 23205 5135 23239
rect 5077 23199 5135 23205
rect 5442 23196 5448 23248
rect 5500 23196 5506 23248
rect 3329 23171 3387 23177
rect 3329 23137 3341 23171
rect 3375 23137 3387 23171
rect 3329 23131 3387 23137
rect 3513 23171 3571 23177
rect 3513 23137 3525 23171
rect 3559 23168 3571 23171
rect 4154 23168 4160 23180
rect 3559 23140 4160 23168
rect 3559 23137 3571 23140
rect 3513 23131 3571 23137
rect 4154 23128 4160 23140
rect 4212 23128 4218 23180
rect 5460 23168 5488 23196
rect 5629 23171 5687 23177
rect 5629 23168 5641 23171
rect 5460 23140 5641 23168
rect 5629 23137 5641 23140
rect 5675 23137 5687 23171
rect 5629 23131 5687 23137
rect 9858 23128 9864 23180
rect 9916 23128 9922 23180
rect 10042 23128 10048 23180
rect 10100 23128 10106 23180
rect 10520 23177 10548 23276
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 11054 23264 11060 23316
rect 11112 23304 11118 23316
rect 11514 23304 11520 23316
rect 11112 23276 11520 23304
rect 11112 23264 11118 23276
rect 11514 23264 11520 23276
rect 11572 23264 11578 23316
rect 11698 23264 11704 23316
rect 11756 23264 11762 23316
rect 13170 23264 13176 23316
rect 13228 23304 13234 23316
rect 13446 23304 13452 23316
rect 13228 23276 13452 23304
rect 13228 23264 13234 23276
rect 13446 23264 13452 23276
rect 13504 23264 13510 23316
rect 15654 23264 15660 23316
rect 15712 23264 15718 23316
rect 20456 23276 21404 23304
rect 11882 23196 11888 23248
rect 11940 23236 11946 23248
rect 18598 23236 18604 23248
rect 11940 23208 18604 23236
rect 11940 23196 11946 23208
rect 18598 23196 18604 23208
rect 18656 23196 18662 23248
rect 20254 23196 20260 23248
rect 20312 23236 20318 23248
rect 20456 23245 20484 23276
rect 20441 23239 20499 23245
rect 20441 23236 20453 23239
rect 20312 23208 20453 23236
rect 20312 23196 20318 23208
rect 20441 23205 20453 23208
rect 20487 23205 20499 23239
rect 20441 23199 20499 23205
rect 10505 23171 10563 23177
rect 10505 23137 10517 23171
rect 10551 23137 10563 23171
rect 10505 23131 10563 23137
rect 10594 23128 10600 23180
rect 10652 23168 10658 23180
rect 10898 23171 10956 23177
rect 10898 23168 10910 23171
rect 10652 23140 10910 23168
rect 10652 23128 10658 23140
rect 10898 23137 10910 23140
rect 10944 23137 10956 23171
rect 10898 23131 10956 23137
rect 16114 23128 16120 23180
rect 16172 23168 16178 23180
rect 16393 23171 16451 23177
rect 16393 23168 16405 23171
rect 16172 23140 16405 23168
rect 16172 23128 16178 23140
rect 16393 23137 16405 23140
rect 16439 23137 16451 23171
rect 16393 23131 16451 23137
rect 16482 23128 16488 23180
rect 16540 23128 16546 23180
rect 19794 23128 19800 23180
rect 19852 23128 19858 23180
rect 19981 23171 20039 23177
rect 19981 23137 19993 23171
rect 20027 23168 20039 23171
rect 20070 23168 20076 23180
rect 20027 23140 20076 23168
rect 20027 23137 20039 23140
rect 19981 23131 20039 23137
rect 20070 23128 20076 23140
rect 20128 23128 20134 23180
rect 20714 23128 20720 23180
rect 20772 23128 20778 23180
rect 20806 23128 20812 23180
rect 20864 23177 20870 23180
rect 20864 23171 20892 23177
rect 20880 23137 20892 23171
rect 21376 23168 21404 23276
rect 21450 23264 21456 23316
rect 21508 23304 21514 23316
rect 21508 23276 22094 23304
rect 21508 23264 21514 23276
rect 22066 23236 22094 23276
rect 24964 23276 28764 23304
rect 24964 23236 24992 23276
rect 22066 23208 24992 23236
rect 24964 23177 24992 23208
rect 24949 23171 25007 23177
rect 21376 23140 24716 23168
rect 20864 23131 20892 23137
rect 20864 23128 20870 23131
rect 3973 23103 4031 23109
rect 3973 23100 3985 23103
rect 2884 23072 3985 23100
rect 3973 23069 3985 23072
rect 4019 23069 4031 23103
rect 3973 23063 4031 23069
rect 5442 23060 5448 23112
rect 5500 23100 5506 23112
rect 5537 23103 5595 23109
rect 5537 23100 5549 23103
rect 5500 23072 5549 23100
rect 5500 23060 5506 23072
rect 5537 23069 5549 23072
rect 5583 23069 5595 23103
rect 5537 23063 5595 23069
rect 10778 23060 10784 23112
rect 10836 23060 10842 23112
rect 11054 23060 11060 23112
rect 11112 23060 11118 23112
rect 14458 23060 14464 23112
rect 14516 23060 14522 23112
rect 15841 23103 15899 23109
rect 15841 23069 15853 23103
rect 15887 23100 15899 23103
rect 15887 23072 15976 23100
rect 15887 23069 15899 23072
rect 15841 23063 15899 23069
rect 3237 23035 3295 23041
rect 3237 23001 3249 23035
rect 3283 23032 3295 23035
rect 4706 23032 4712 23044
rect 3283 23004 4712 23032
rect 3283 23001 3295 23004
rect 3237 22995 3295 23001
rect 4706 22992 4712 23004
rect 4764 22992 4770 23044
rect 4801 23035 4859 23041
rect 4801 23001 4813 23035
rect 4847 23032 4859 23035
rect 7558 23032 7564 23044
rect 4847 23004 7564 23032
rect 4847 23001 4859 23004
rect 4801 22995 4859 23001
rect 7558 22992 7564 23004
rect 7616 22992 7622 23044
rect 4062 22924 4068 22976
rect 4120 22964 4126 22976
rect 4893 22967 4951 22973
rect 4893 22964 4905 22967
rect 4120 22936 4905 22964
rect 4120 22924 4126 22936
rect 4893 22933 4905 22936
rect 4939 22933 4951 22967
rect 4893 22927 4951 22933
rect 5445 22967 5503 22973
rect 5445 22933 5457 22967
rect 5491 22964 5503 22967
rect 7098 22964 7104 22976
rect 5491 22936 7104 22964
rect 5491 22933 5503 22936
rect 5445 22927 5503 22933
rect 7098 22924 7104 22936
rect 7156 22964 7162 22976
rect 8110 22964 8116 22976
rect 7156 22936 8116 22964
rect 7156 22924 7162 22936
rect 8110 22924 8116 22936
rect 8168 22924 8174 22976
rect 14274 22924 14280 22976
rect 14332 22924 14338 22976
rect 15948 22973 15976 23072
rect 18966 23060 18972 23112
rect 19024 23060 19030 23112
rect 19245 23103 19303 23109
rect 19245 23069 19257 23103
rect 19291 23100 19303 23103
rect 19610 23100 19616 23112
rect 19291 23072 19616 23100
rect 19291 23069 19303 23072
rect 19245 23063 19303 23069
rect 19610 23060 19616 23072
rect 19668 23060 19674 23112
rect 20990 23060 20996 23112
rect 21048 23060 21054 23112
rect 23937 23103 23995 23109
rect 23937 23069 23949 23103
rect 23983 23100 23995 23103
rect 23983 23072 24440 23100
rect 23983 23069 23995 23072
rect 23937 23063 23995 23069
rect 16482 22992 16488 23044
rect 16540 23032 16546 23044
rect 16540 23004 19472 23032
rect 16540 22992 16546 23004
rect 15933 22967 15991 22973
rect 15933 22933 15945 22967
rect 15979 22933 15991 22967
rect 15933 22927 15991 22933
rect 16206 22924 16212 22976
rect 16264 22964 16270 22976
rect 16301 22967 16359 22973
rect 16301 22964 16313 22967
rect 16264 22936 16313 22964
rect 16264 22924 16270 22936
rect 16301 22933 16313 22936
rect 16347 22933 16359 22967
rect 16301 22927 16359 22933
rect 18782 22924 18788 22976
rect 18840 22924 18846 22976
rect 19444 22973 19472 23004
rect 19429 22967 19487 22973
rect 19429 22933 19441 22967
rect 19475 22933 19487 22967
rect 19429 22927 19487 22933
rect 19610 22924 19616 22976
rect 19668 22964 19674 22976
rect 21450 22964 21456 22976
rect 19668 22936 21456 22964
rect 19668 22924 19674 22936
rect 21450 22924 21456 22936
rect 21508 22924 21514 22976
rect 21634 22924 21640 22976
rect 21692 22924 21698 22976
rect 23750 22924 23756 22976
rect 23808 22924 23814 22976
rect 24412 22973 24440 23072
rect 24688 23032 24716 23140
rect 24949 23137 24961 23171
rect 24995 23137 25007 23171
rect 24949 23131 25007 23137
rect 26329 23171 26387 23177
rect 26329 23137 26341 23171
rect 26375 23168 26387 23171
rect 26418 23168 26424 23180
rect 26375 23140 26424 23168
rect 26375 23137 26387 23140
rect 26329 23131 26387 23137
rect 26418 23128 26424 23140
rect 26476 23128 26482 23180
rect 26510 23128 26516 23180
rect 26568 23128 26574 23180
rect 28736 23168 28764 23276
rect 29178 23264 29184 23316
rect 29236 23264 29242 23316
rect 34517 23307 34575 23313
rect 34517 23304 34529 23307
rect 32784 23276 34529 23304
rect 31662 23236 31668 23248
rect 30392 23208 31668 23236
rect 30392 23177 30420 23208
rect 31662 23196 31668 23208
rect 31720 23196 31726 23248
rect 32784 23245 32812 23276
rect 34517 23273 34529 23276
rect 34563 23273 34575 23307
rect 34517 23267 34575 23273
rect 32769 23239 32827 23245
rect 32769 23205 32781 23239
rect 32815 23236 32827 23239
rect 32858 23236 32864 23248
rect 32815 23208 32864 23236
rect 32815 23205 32827 23208
rect 32769 23199 32827 23205
rect 32858 23196 32864 23208
rect 32916 23196 32922 23248
rect 30101 23171 30159 23177
rect 30101 23168 30113 23171
rect 28736 23140 30113 23168
rect 30101 23137 30113 23140
rect 30147 23137 30159 23171
rect 30101 23131 30159 23137
rect 30377 23171 30435 23177
rect 30377 23137 30389 23171
rect 30423 23137 30435 23171
rect 32033 23171 32091 23177
rect 32033 23168 32045 23171
rect 30377 23131 30435 23137
rect 30484 23140 32045 23168
rect 24765 23103 24823 23109
rect 24765 23069 24777 23103
rect 24811 23100 24823 23103
rect 24854 23100 24860 23112
rect 24811 23072 24860 23100
rect 24811 23069 24823 23072
rect 24765 23063 24823 23069
rect 24854 23060 24860 23072
rect 24912 23100 24918 23112
rect 25682 23100 25688 23112
rect 24912 23072 25688 23100
rect 24912 23060 24918 23072
rect 25682 23060 25688 23072
rect 25740 23060 25746 23112
rect 27614 23060 27620 23112
rect 27672 23060 27678 23112
rect 27709 23103 27767 23109
rect 27709 23069 27721 23103
rect 27755 23100 27767 23103
rect 27798 23100 27804 23112
rect 27755 23072 27804 23100
rect 27755 23069 27767 23072
rect 27709 23063 27767 23069
rect 27798 23060 27804 23072
rect 27856 23100 27862 23112
rect 28902 23100 28908 23112
rect 27856 23072 28908 23100
rect 27856 23060 27862 23072
rect 28902 23060 28908 23072
rect 28960 23060 28966 23112
rect 29365 23103 29423 23109
rect 29365 23069 29377 23103
rect 29411 23100 29423 23103
rect 29411 23072 29592 23100
rect 29411 23069 29423 23072
rect 29365 23063 29423 23069
rect 25314 23032 25320 23044
rect 24688 23004 25320 23032
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 27954 23035 28012 23041
rect 27954 23032 27966 23035
rect 27448 23004 27966 23032
rect 24397 22967 24455 22973
rect 24397 22933 24409 22967
rect 24443 22933 24455 22967
rect 24397 22927 24455 22933
rect 24670 22924 24676 22976
rect 24728 22964 24734 22976
rect 24857 22967 24915 22973
rect 24857 22964 24869 22967
rect 24728 22936 24869 22964
rect 24728 22924 24734 22936
rect 24857 22933 24869 22936
rect 24903 22933 24915 22967
rect 24857 22927 24915 22933
rect 25498 22924 25504 22976
rect 25556 22964 25562 22976
rect 25869 22967 25927 22973
rect 25869 22964 25881 22967
rect 25556 22936 25881 22964
rect 25556 22924 25562 22936
rect 25869 22933 25881 22936
rect 25915 22933 25927 22967
rect 25869 22927 25927 22933
rect 26234 22924 26240 22976
rect 26292 22924 26298 22976
rect 27448 22973 27476 23004
rect 27954 23001 27966 23004
rect 28000 23001 28012 23035
rect 27954 22995 28012 23001
rect 27433 22967 27491 22973
rect 27433 22933 27445 22967
rect 27479 22933 27491 22967
rect 27433 22927 27491 22933
rect 28350 22924 28356 22976
rect 28408 22964 28414 22976
rect 29564 22973 29592 23072
rect 29914 23060 29920 23112
rect 29972 23060 29978 23112
rect 30116 23100 30144 23131
rect 30484 23100 30512 23140
rect 32033 23137 32045 23140
rect 32079 23137 32091 23171
rect 32033 23131 32091 23137
rect 32398 23128 32404 23180
rect 32456 23128 32462 23180
rect 30116 23072 30512 23100
rect 30650 23060 30656 23112
rect 30708 23100 30714 23112
rect 31021 23103 31079 23109
rect 31021 23100 31033 23103
rect 30708 23072 31033 23100
rect 30708 23060 30714 23072
rect 31021 23069 31033 23072
rect 31067 23100 31079 23103
rect 31757 23103 31815 23109
rect 31757 23100 31769 23103
rect 31067 23072 31769 23100
rect 31067 23069 31079 23072
rect 31021 23063 31079 23069
rect 31757 23069 31769 23072
rect 31803 23100 31815 23103
rect 33137 23103 33195 23109
rect 31803 23072 32352 23100
rect 31803 23069 31815 23072
rect 31757 23063 31815 23069
rect 31113 23035 31171 23041
rect 31113 23032 31125 23035
rect 30668 23004 31125 23032
rect 30668 22976 30696 23004
rect 31113 23001 31125 23004
rect 31159 23001 31171 23035
rect 31113 22995 31171 23001
rect 31297 23035 31355 23041
rect 31297 23001 31309 23035
rect 31343 23032 31355 23035
rect 31846 23032 31852 23044
rect 31343 23004 31852 23032
rect 31343 23001 31355 23004
rect 31297 22995 31355 23001
rect 29089 22967 29147 22973
rect 29089 22964 29101 22967
rect 28408 22936 29101 22964
rect 28408 22924 28414 22936
rect 29089 22933 29101 22936
rect 29135 22933 29147 22967
rect 29089 22927 29147 22933
rect 29549 22967 29607 22973
rect 29549 22933 29561 22967
rect 29595 22933 29607 22967
rect 29549 22927 29607 22933
rect 30009 22967 30067 22973
rect 30009 22933 30021 22967
rect 30055 22964 30067 22967
rect 30190 22964 30196 22976
rect 30055 22936 30196 22964
rect 30055 22933 30067 22936
rect 30009 22927 30067 22933
rect 30190 22924 30196 22936
rect 30248 22924 30254 22976
rect 30558 22924 30564 22976
rect 30616 22924 30622 22976
rect 30650 22924 30656 22976
rect 30708 22924 30714 22976
rect 30926 22924 30932 22976
rect 30984 22924 30990 22976
rect 31128 22964 31156 22995
rect 31846 22992 31852 23004
rect 31904 22992 31910 23044
rect 31386 22964 31392 22976
rect 31128 22936 31392 22964
rect 31386 22924 31392 22936
rect 31444 22964 31450 22976
rect 31573 22967 31631 22973
rect 31573 22964 31585 22967
rect 31444 22936 31585 22964
rect 31444 22924 31450 22936
rect 31573 22933 31585 22936
rect 31619 22933 31631 22967
rect 31573 22927 31631 22933
rect 31665 22967 31723 22973
rect 31665 22933 31677 22967
rect 31711 22964 31723 22967
rect 32214 22964 32220 22976
rect 31711 22936 32220 22964
rect 31711 22933 31723 22936
rect 31665 22927 31723 22933
rect 32214 22924 32220 22936
rect 32272 22924 32278 22976
rect 32324 22964 32352 23072
rect 33137 23069 33149 23103
rect 33183 23100 33195 23103
rect 33226 23100 33232 23112
rect 33183 23072 33232 23100
rect 33183 23069 33195 23072
rect 33137 23063 33195 23069
rect 33226 23060 33232 23072
rect 33284 23060 33290 23112
rect 33404 23035 33462 23041
rect 33404 23001 33416 23035
rect 33450 23032 33462 23035
rect 33778 23032 33784 23044
rect 33450 23004 33784 23032
rect 33450 23001 33462 23004
rect 33404 22995 33462 23001
rect 33778 22992 33784 23004
rect 33836 22992 33842 23044
rect 32861 22967 32919 22973
rect 32861 22964 32873 22967
rect 32324 22936 32873 22964
rect 32861 22933 32873 22936
rect 32907 22933 32919 22967
rect 32861 22927 32919 22933
rect 1104 22874 36800 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 36800 22874
rect 1104 22800 36800 22822
rect 4338 22720 4344 22772
rect 4396 22760 4402 22772
rect 4798 22760 4804 22772
rect 4396 22732 4804 22760
rect 4396 22720 4402 22732
rect 4798 22720 4804 22732
rect 4856 22720 4862 22772
rect 5442 22720 5448 22772
rect 5500 22720 5506 22772
rect 19886 22720 19892 22772
rect 19944 22720 19950 22772
rect 20806 22720 20812 22772
rect 20864 22760 20870 22772
rect 21082 22760 21088 22772
rect 20864 22732 21088 22760
rect 20864 22720 20870 22732
rect 21082 22720 21088 22732
rect 21140 22720 21146 22772
rect 24765 22763 24823 22769
rect 24765 22729 24777 22763
rect 24811 22760 24823 22763
rect 24854 22760 24860 22772
rect 24811 22732 24860 22760
rect 24811 22729 24823 22732
rect 24765 22723 24823 22729
rect 24854 22720 24860 22732
rect 24912 22720 24918 22772
rect 27614 22720 27620 22772
rect 27672 22760 27678 22772
rect 27985 22763 28043 22769
rect 27985 22760 27997 22763
rect 27672 22732 27997 22760
rect 27672 22720 27678 22732
rect 27985 22729 27997 22732
rect 28031 22729 28043 22763
rect 27985 22723 28043 22729
rect 30466 22720 30472 22772
rect 30524 22760 30530 22772
rect 30926 22760 30932 22772
rect 30524 22732 30932 22760
rect 30524 22720 30530 22732
rect 30926 22720 30932 22732
rect 30984 22720 30990 22772
rect 32306 22720 32312 22772
rect 32364 22720 32370 22772
rect 32398 22720 32404 22772
rect 32456 22720 32462 22772
rect 33778 22720 33784 22772
rect 33836 22720 33842 22772
rect 7650 22692 7656 22704
rect 1412 22664 7656 22692
rect 1412 22633 1440 22664
rect 7650 22652 7656 22664
rect 7708 22652 7714 22704
rect 8570 22692 8576 22704
rect 7760 22664 8576 22692
rect 1397 22627 1455 22633
rect 1397 22593 1409 22627
rect 1443 22593 1455 22627
rect 1397 22587 1455 22593
rect 2958 22584 2964 22636
rect 3016 22624 3022 22636
rect 4062 22624 4068 22636
rect 3016 22596 4068 22624
rect 3016 22584 3022 22596
rect 4062 22584 4068 22596
rect 4120 22584 4126 22636
rect 4332 22627 4390 22633
rect 4332 22593 4344 22627
rect 4378 22624 4390 22627
rect 4614 22624 4620 22636
rect 4378 22596 4620 22624
rect 4378 22593 4390 22596
rect 4332 22587 4390 22593
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 7558 22584 7564 22636
rect 7616 22624 7622 22636
rect 7760 22624 7788 22664
rect 8570 22652 8576 22664
rect 8628 22652 8634 22704
rect 9048 22664 12434 22692
rect 7834 22633 7840 22636
rect 7616 22596 7788 22624
rect 7616 22584 7622 22596
rect 7828 22587 7840 22633
rect 7834 22584 7840 22587
rect 7892 22584 7898 22636
rect 8386 22584 8392 22636
rect 8444 22624 8450 22636
rect 9048 22633 9076 22664
rect 9033 22627 9091 22633
rect 9033 22624 9045 22627
rect 8444 22596 9045 22624
rect 8444 22584 8450 22596
rect 9033 22593 9045 22596
rect 9079 22593 9091 22627
rect 9033 22587 9091 22593
rect 9217 22627 9275 22633
rect 9217 22593 9229 22627
rect 9263 22624 9275 22627
rect 10594 22624 10600 22636
rect 9263 22596 10600 22624
rect 9263 22593 9275 22596
rect 9217 22587 9275 22593
rect 9232 22556 9260 22587
rect 10594 22584 10600 22596
rect 10652 22584 10658 22636
rect 8956 22528 9260 22556
rect 12406 22556 12434 22664
rect 14274 22652 14280 22704
rect 14332 22692 14338 22704
rect 18782 22701 18788 22704
rect 14706 22695 14764 22701
rect 14706 22692 14718 22695
rect 14332 22664 14718 22692
rect 14332 22652 14338 22664
rect 14706 22661 14718 22664
rect 14752 22661 14764 22695
rect 18776 22692 18788 22701
rect 18743 22664 18788 22692
rect 14706 22655 14764 22661
rect 18776 22655 18788 22664
rect 18782 22652 18788 22655
rect 18840 22652 18846 22704
rect 23652 22695 23710 22701
rect 23652 22661 23664 22695
rect 23698 22692 23710 22695
rect 23750 22692 23756 22704
rect 23698 22664 23756 22692
rect 23698 22661 23710 22664
rect 23652 22655 23710 22661
rect 23750 22652 23756 22664
rect 23808 22652 23814 22704
rect 23860 22664 26556 22692
rect 12526 22584 12532 22636
rect 12584 22584 12590 22636
rect 13446 22584 13452 22636
rect 13504 22584 13510 22636
rect 13630 22633 13636 22636
rect 13587 22627 13636 22633
rect 13587 22593 13599 22627
rect 13633 22593 13636 22627
rect 13587 22587 13636 22593
rect 13630 22584 13636 22587
rect 13688 22584 13694 22636
rect 14461 22627 14519 22633
rect 14461 22593 14473 22627
rect 14507 22624 14519 22627
rect 15010 22624 15016 22636
rect 14507 22596 15016 22624
rect 14507 22593 14519 22596
rect 14461 22587 14519 22593
rect 15010 22584 15016 22596
rect 15068 22584 15074 22636
rect 18141 22627 18199 22633
rect 18141 22593 18153 22627
rect 18187 22624 18199 22627
rect 22830 22624 22836 22636
rect 18187 22596 22836 22624
rect 18187 22593 18199 22596
rect 18141 22587 18199 22593
rect 22830 22584 22836 22596
rect 22888 22624 22894 22636
rect 23860 22624 23888 22664
rect 26528 22636 26556 22664
rect 27706 22652 27712 22704
rect 27764 22692 27770 22704
rect 28350 22692 28356 22704
rect 27764 22664 28356 22692
rect 27764 22652 27770 22664
rect 28350 22652 28356 22664
rect 28408 22652 28414 22704
rect 32416 22692 32444 22720
rect 31864 22664 32444 22692
rect 22888 22596 23888 22624
rect 25685 22627 25743 22633
rect 22888 22584 22894 22596
rect 25685 22593 25697 22627
rect 25731 22624 25743 22627
rect 25958 22624 25964 22636
rect 25731 22596 25964 22624
rect 25731 22593 25743 22596
rect 25685 22587 25743 22593
rect 25958 22584 25964 22596
rect 26016 22584 26022 22636
rect 26510 22584 26516 22636
rect 26568 22624 26574 22636
rect 26568 22596 28672 22624
rect 26568 22584 26574 22596
rect 12618 22556 12624 22568
rect 12406 22528 12624 22556
rect 934 22448 940 22500
rect 992 22488 998 22500
rect 8956 22497 8984 22528
rect 12618 22516 12624 22528
rect 12676 22516 12682 22568
rect 12713 22559 12771 22565
rect 12713 22525 12725 22559
rect 12759 22556 12771 22559
rect 12894 22556 12900 22568
rect 12759 22528 12900 22556
rect 12759 22525 12771 22528
rect 12713 22519 12771 22525
rect 12894 22516 12900 22528
rect 12952 22556 12958 22568
rect 12952 22528 13308 22556
rect 12952 22516 12958 22528
rect 1581 22491 1639 22497
rect 1581 22488 1593 22491
rect 992 22460 1593 22488
rect 992 22448 998 22460
rect 1581 22457 1593 22460
rect 1627 22457 1639 22491
rect 1581 22451 1639 22457
rect 8941 22491 8999 22497
rect 8941 22457 8953 22491
rect 8987 22457 8999 22491
rect 8941 22451 8999 22457
rect 13170 22448 13176 22500
rect 13228 22448 13234 22500
rect 3878 22380 3884 22432
rect 3936 22420 3942 22432
rect 4430 22420 4436 22432
rect 3936 22392 4436 22420
rect 3936 22380 3942 22392
rect 4430 22380 4436 22392
rect 4488 22380 4494 22432
rect 9030 22380 9036 22432
rect 9088 22380 9094 22432
rect 13280 22420 13308 22528
rect 13722 22516 13728 22568
rect 13780 22516 13786 22568
rect 18509 22559 18567 22565
rect 18509 22525 18521 22559
rect 18555 22525 18567 22559
rect 23106 22556 23112 22568
rect 18509 22519 18567 22525
rect 21192 22528 23112 22556
rect 14274 22448 14280 22500
rect 14332 22488 14338 22500
rect 14332 22460 14504 22488
rect 14332 22448 14338 22460
rect 14292 22420 14320 22448
rect 13280 22392 14320 22420
rect 14366 22380 14372 22432
rect 14424 22380 14430 22432
rect 14476 22420 14504 22460
rect 15841 22423 15899 22429
rect 15841 22420 15853 22423
rect 14476 22392 15853 22420
rect 15841 22389 15853 22392
rect 15887 22389 15899 22423
rect 15841 22383 15899 22389
rect 16758 22380 16764 22432
rect 16816 22420 16822 22432
rect 17402 22420 17408 22432
rect 16816 22392 17408 22420
rect 16816 22380 16822 22392
rect 17402 22380 17408 22392
rect 17460 22380 17466 22432
rect 17862 22380 17868 22432
rect 17920 22420 17926 22432
rect 18325 22423 18383 22429
rect 18325 22420 18337 22423
rect 17920 22392 18337 22420
rect 17920 22380 17926 22392
rect 18325 22389 18337 22392
rect 18371 22389 18383 22423
rect 18524 22420 18552 22519
rect 21192 22432 21220 22528
rect 23106 22516 23112 22528
rect 23164 22556 23170 22568
rect 23385 22559 23443 22565
rect 23385 22556 23397 22559
rect 23164 22528 23397 22556
rect 23164 22516 23170 22528
rect 23385 22525 23397 22528
rect 23431 22525 23443 22559
rect 23385 22519 23443 22525
rect 28442 22516 28448 22568
rect 28500 22516 28506 22568
rect 28644 22565 28672 22596
rect 30834 22584 30840 22636
rect 30892 22624 30898 22636
rect 31864 22633 31892 22664
rect 31021 22627 31079 22633
rect 31021 22624 31033 22627
rect 30892 22596 31033 22624
rect 30892 22584 30898 22596
rect 31021 22593 31033 22596
rect 31067 22593 31079 22627
rect 31021 22587 31079 22593
rect 31665 22627 31723 22633
rect 31665 22593 31677 22627
rect 31711 22593 31723 22627
rect 31665 22587 31723 22593
rect 31849 22627 31907 22633
rect 31849 22593 31861 22627
rect 31895 22593 31907 22627
rect 31849 22587 31907 22593
rect 32125 22627 32183 22633
rect 32125 22593 32137 22627
rect 32171 22624 32183 22627
rect 32214 22624 32220 22636
rect 32171 22596 32220 22624
rect 32171 22593 32183 22596
rect 32125 22587 32183 22593
rect 28629 22559 28687 22565
rect 28629 22525 28641 22559
rect 28675 22556 28687 22559
rect 30558 22556 30564 22568
rect 28675 22528 30564 22556
rect 28675 22525 28687 22528
rect 28629 22519 28687 22525
rect 30558 22516 30564 22528
rect 30616 22516 30622 22568
rect 30745 22559 30803 22565
rect 30745 22525 30757 22559
rect 30791 22556 30803 22559
rect 30926 22556 30932 22568
rect 30791 22528 30932 22556
rect 30791 22525 30803 22528
rect 30745 22519 30803 22525
rect 30926 22516 30932 22528
rect 30984 22516 30990 22568
rect 31680 22556 31708 22587
rect 32214 22584 32220 22596
rect 32272 22584 32278 22636
rect 32306 22584 32312 22636
rect 32364 22584 32370 22636
rect 32401 22627 32459 22633
rect 32401 22593 32413 22627
rect 32447 22624 32459 22627
rect 32490 22624 32496 22636
rect 32447 22596 32496 22624
rect 32447 22593 32459 22596
rect 32401 22587 32459 22593
rect 32490 22584 32496 22596
rect 32548 22584 32554 22636
rect 32858 22584 32864 22636
rect 32916 22584 32922 22636
rect 33226 22584 33232 22636
rect 33284 22624 33290 22636
rect 33965 22627 34023 22633
rect 33965 22624 33977 22627
rect 33284 22596 33977 22624
rect 33284 22584 33290 22596
rect 33965 22593 33977 22596
rect 34011 22593 34023 22627
rect 33965 22587 34023 22593
rect 33134 22556 33140 22568
rect 31680 22528 33140 22556
rect 33134 22516 33140 22528
rect 33192 22516 33198 22568
rect 30944 22488 30972 22516
rect 31846 22488 31852 22500
rect 30944 22460 31852 22488
rect 31846 22448 31852 22460
rect 31904 22488 31910 22500
rect 32490 22488 32496 22500
rect 31904 22460 32496 22488
rect 31904 22448 31910 22460
rect 32490 22448 32496 22460
rect 32548 22448 32554 22500
rect 21174 22420 21180 22432
rect 18524 22392 21180 22420
rect 18325 22383 18383 22389
rect 21174 22380 21180 22392
rect 21232 22380 21238 22432
rect 25590 22380 25596 22432
rect 25648 22420 25654 22432
rect 25777 22423 25835 22429
rect 25777 22420 25789 22423
rect 25648 22392 25789 22420
rect 25648 22380 25654 22392
rect 25777 22389 25789 22392
rect 25823 22389 25835 22423
rect 25777 22383 25835 22389
rect 31662 22380 31668 22432
rect 31720 22380 31726 22432
rect 1104 22330 36800 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 36800 22330
rect 1104 22256 36800 22278
rect 4614 22176 4620 22228
rect 4672 22176 4678 22228
rect 7834 22176 7840 22228
rect 7892 22216 7898 22228
rect 7929 22219 7987 22225
rect 7929 22216 7941 22219
rect 7892 22188 7941 22216
rect 7892 22176 7898 22188
rect 7929 22185 7941 22188
rect 7975 22185 7987 22219
rect 7929 22179 7987 22185
rect 10134 22176 10140 22228
rect 10192 22216 10198 22228
rect 10597 22219 10655 22225
rect 10597 22216 10609 22219
rect 10192 22188 10609 22216
rect 10192 22176 10198 22188
rect 10597 22185 10609 22188
rect 10643 22185 10655 22219
rect 10597 22179 10655 22185
rect 2958 22148 2964 22160
rect 2792 22120 2964 22148
rect 2792 22080 2820 22120
rect 2958 22108 2964 22120
rect 3016 22108 3022 22160
rect 6914 22108 6920 22160
rect 6972 22108 6978 22160
rect 2700 22052 2820 22080
rect 1486 21972 1492 22024
rect 1544 22012 1550 22024
rect 1581 22015 1639 22021
rect 1581 22012 1593 22015
rect 1544 21984 1593 22012
rect 1544 21972 1550 21984
rect 1581 21981 1593 21984
rect 1627 22012 1639 22015
rect 2700 22012 2728 22052
rect 4154 22040 4160 22092
rect 4212 22080 4218 22092
rect 8294 22080 8300 22092
rect 4212 22052 8300 22080
rect 4212 22040 4218 22052
rect 1627 21984 2728 22012
rect 1627 21981 1639 21984
rect 1581 21975 1639 21981
rect 4798 21972 4804 22024
rect 4856 21972 4862 22024
rect 8220 22021 8248 22052
rect 8294 22040 8300 22052
rect 8352 22040 8358 22092
rect 8570 22040 8576 22092
rect 8628 22080 8634 22092
rect 9217 22083 9275 22089
rect 9217 22080 9229 22083
rect 8628 22052 9229 22080
rect 8628 22040 8634 22052
rect 9217 22049 9229 22052
rect 9263 22049 9275 22083
rect 10612 22080 10640 22179
rect 12618 22176 12624 22228
rect 12676 22216 12682 22228
rect 14185 22219 14243 22225
rect 12676 22188 13584 22216
rect 12676 22176 12682 22188
rect 12805 22151 12863 22157
rect 12805 22117 12817 22151
rect 12851 22117 12863 22151
rect 12805 22111 12863 22117
rect 13556 22148 13584 22188
rect 14185 22185 14197 22219
rect 14231 22216 14243 22219
rect 14458 22216 14464 22228
rect 14231 22188 14464 22216
rect 14231 22185 14243 22188
rect 14185 22179 14243 22185
rect 14458 22176 14464 22188
rect 14516 22176 14522 22228
rect 14734 22176 14740 22228
rect 14792 22216 14798 22228
rect 17862 22216 17868 22228
rect 14792 22188 17868 22216
rect 14792 22176 14798 22188
rect 17862 22176 17868 22188
rect 17920 22176 17926 22228
rect 26234 22176 26240 22228
rect 26292 22216 26298 22228
rect 26973 22219 27031 22225
rect 26973 22216 26985 22219
rect 26292 22188 26985 22216
rect 26292 22176 26298 22188
rect 26973 22185 26985 22188
rect 27019 22185 27031 22219
rect 26973 22179 27031 22185
rect 31386 22176 31392 22228
rect 31444 22216 31450 22228
rect 32306 22216 32312 22228
rect 31444 22188 32312 22216
rect 31444 22176 31450 22188
rect 32306 22176 32312 22188
rect 32364 22176 32370 22228
rect 16482 22148 16488 22160
rect 13556 22120 16488 22148
rect 10612 22052 10916 22080
rect 9217 22043 9275 22049
rect 10888 22021 10916 22052
rect 8205 22015 8263 22021
rect 8205 21981 8217 22015
rect 8251 21981 8263 22015
rect 10689 22015 10747 22021
rect 10689 22012 10701 22015
rect 8205 21975 8263 21981
rect 9692 21984 10701 22012
rect 9692 21956 9720 21984
rect 10689 21981 10701 21984
rect 10735 21981 10747 22015
rect 10689 21975 10747 21981
rect 10873 22015 10931 22021
rect 10873 21981 10885 22015
rect 10919 21981 10931 22015
rect 10873 21975 10931 21981
rect 11425 22015 11483 22021
rect 11425 21981 11437 22015
rect 11471 22012 11483 22015
rect 11974 22012 11980 22024
rect 11471 21984 11980 22012
rect 11471 21981 11483 21984
rect 11425 21975 11483 21981
rect 11974 21972 11980 21984
rect 12032 21972 12038 22024
rect 12820 22012 12848 22111
rect 13556 22089 13584 22120
rect 16482 22108 16488 22120
rect 16540 22108 16546 22160
rect 32674 22108 32680 22160
rect 32732 22148 32738 22160
rect 32732 22120 33548 22148
rect 32732 22108 32738 22120
rect 13541 22083 13599 22089
rect 13541 22049 13553 22083
rect 13587 22080 13599 22083
rect 13587 22052 13621 22080
rect 13587 22049 13599 22052
rect 13541 22043 13599 22049
rect 14734 22040 14740 22092
rect 14792 22040 14798 22092
rect 16206 22040 16212 22092
rect 16264 22040 16270 22092
rect 16393 22083 16451 22089
rect 16393 22049 16405 22083
rect 16439 22080 16451 22083
rect 16758 22080 16764 22092
rect 16439 22052 16764 22080
rect 16439 22049 16451 22052
rect 16393 22043 16451 22049
rect 16758 22040 16764 22052
rect 16816 22040 16822 22092
rect 16853 22083 16911 22089
rect 16853 22049 16865 22083
rect 16899 22080 16911 22083
rect 16942 22080 16948 22092
rect 16899 22052 16948 22080
rect 16899 22049 16911 22052
rect 16853 22043 16911 22049
rect 16942 22040 16948 22052
rect 17000 22040 17006 22092
rect 17126 22040 17132 22092
rect 17184 22040 17190 22092
rect 17218 22040 17224 22092
rect 17276 22089 17282 22092
rect 17276 22083 17304 22089
rect 17292 22049 17304 22083
rect 17276 22043 17304 22049
rect 17405 22083 17463 22089
rect 17405 22049 17417 22083
rect 17451 22080 17463 22083
rect 17586 22080 17592 22092
rect 17451 22052 17592 22080
rect 17451 22049 17463 22052
rect 17405 22043 17463 22049
rect 17276 22040 17282 22043
rect 17586 22040 17592 22052
rect 17644 22080 17650 22092
rect 20162 22080 20168 22092
rect 17644 22052 20168 22080
rect 17644 22040 17650 22052
rect 20162 22040 20168 22052
rect 20220 22040 20226 22092
rect 21174 22040 21180 22092
rect 21232 22080 21238 22092
rect 21361 22083 21419 22089
rect 21361 22080 21373 22083
rect 21232 22052 21373 22080
rect 21232 22040 21238 22052
rect 21361 22049 21373 22052
rect 21407 22049 21419 22083
rect 21361 22043 21419 22049
rect 23106 22040 23112 22092
rect 23164 22080 23170 22092
rect 25590 22080 25596 22092
rect 23164 22052 25596 22080
rect 23164 22040 23170 22052
rect 25590 22040 25596 22052
rect 25648 22040 25654 22092
rect 30653 22083 30711 22089
rect 30653 22049 30665 22083
rect 30699 22080 30711 22083
rect 30742 22080 30748 22092
rect 30699 22052 30748 22080
rect 30699 22049 30711 22052
rect 30653 22043 30711 22049
rect 30742 22040 30748 22052
rect 30800 22040 30806 22092
rect 32784 22089 32812 22120
rect 33520 22089 33548 22120
rect 31297 22083 31355 22089
rect 31297 22080 31309 22083
rect 30852 22052 31309 22080
rect 13265 22015 13323 22021
rect 13265 22012 13277 22015
rect 12820 21984 13277 22012
rect 13265 21981 13277 21984
rect 13311 22012 13323 22015
rect 13630 22012 13636 22024
rect 13311 21984 13636 22012
rect 13311 21981 13323 21984
rect 13265 21975 13323 21981
rect 13630 21972 13636 21984
rect 13688 21972 13694 22024
rect 14274 21972 14280 22024
rect 14332 22012 14338 22024
rect 14553 22015 14611 22021
rect 14553 22012 14565 22015
rect 14332 21984 14565 22012
rect 14332 21972 14338 21984
rect 14553 21981 14565 21984
rect 14599 21981 14611 22015
rect 14553 21975 14611 21981
rect 21266 21972 21272 22024
rect 21324 21972 21330 22024
rect 25498 21972 25504 22024
rect 25556 21972 25562 22024
rect 30466 21972 30472 22024
rect 30524 22012 30530 22024
rect 30852 22012 30880 22052
rect 31297 22049 31309 22052
rect 31343 22049 31355 22083
rect 31297 22043 31355 22049
rect 32769 22083 32827 22089
rect 32769 22049 32781 22083
rect 32815 22080 32827 22083
rect 33505 22083 33563 22089
rect 32815 22052 32849 22080
rect 32815 22049 32827 22052
rect 32769 22043 32827 22049
rect 33505 22049 33517 22083
rect 33551 22080 33563 22083
rect 33551 22052 33585 22080
rect 33551 22049 33563 22052
rect 33505 22043 33563 22049
rect 30524 21984 30880 22012
rect 31021 22015 31079 22021
rect 30524 21972 30530 21984
rect 31021 21981 31033 22015
rect 31067 21981 31079 22015
rect 31021 21975 31079 21981
rect 1848 21947 1906 21953
rect 1848 21913 1860 21947
rect 1894 21944 1906 21947
rect 1946 21944 1952 21956
rect 1894 21916 1952 21944
rect 1894 21913 1906 21916
rect 1848 21907 1906 21913
rect 1946 21904 1952 21916
rect 2004 21904 2010 21956
rect 6641 21947 6699 21953
rect 6641 21913 6653 21947
rect 6687 21944 6699 21947
rect 7374 21944 7380 21956
rect 6687 21916 7380 21944
rect 6687 21913 6699 21916
rect 6641 21907 6699 21913
rect 7374 21904 7380 21916
rect 7432 21904 7438 21956
rect 7929 21947 7987 21953
rect 7929 21913 7941 21947
rect 7975 21944 7987 21947
rect 9030 21944 9036 21956
rect 7975 21916 9036 21944
rect 7975 21913 7987 21916
rect 7929 21907 7987 21913
rect 9030 21904 9036 21916
rect 9088 21904 9094 21956
rect 9306 21904 9312 21956
rect 9364 21944 9370 21956
rect 9462 21947 9520 21953
rect 9462 21944 9474 21947
rect 9364 21916 9474 21944
rect 9364 21904 9370 21916
rect 9462 21913 9474 21916
rect 9508 21913 9520 21947
rect 9462 21907 9520 21913
rect 9674 21904 9680 21956
rect 9732 21904 9738 21956
rect 11692 21947 11750 21953
rect 11692 21913 11704 21947
rect 11738 21944 11750 21947
rect 11790 21944 11796 21956
rect 11738 21916 11796 21944
rect 11738 21913 11750 21916
rect 11692 21907 11750 21913
rect 11790 21904 11796 21916
rect 11848 21904 11854 21956
rect 13078 21904 13084 21956
rect 13136 21944 13142 21956
rect 14645 21947 14703 21953
rect 14645 21944 14657 21947
rect 13136 21916 14657 21944
rect 13136 21904 13142 21916
rect 14645 21913 14657 21916
rect 14691 21913 14703 21947
rect 21606 21947 21664 21953
rect 21606 21944 21618 21947
rect 14645 21907 14703 21913
rect 21100 21916 21618 21944
rect 2958 21836 2964 21888
rect 3016 21836 3022 21888
rect 4798 21836 4804 21888
rect 4856 21876 4862 21888
rect 5258 21876 5264 21888
rect 4856 21848 5264 21876
rect 4856 21836 4862 21848
rect 5258 21836 5264 21848
rect 5316 21836 5322 21888
rect 7006 21836 7012 21888
rect 7064 21876 7070 21888
rect 7101 21879 7159 21885
rect 7101 21876 7113 21879
rect 7064 21848 7113 21876
rect 7064 21836 7070 21848
rect 7101 21845 7113 21848
rect 7147 21845 7159 21879
rect 7101 21839 7159 21845
rect 7834 21836 7840 21888
rect 7892 21876 7898 21888
rect 8113 21879 8171 21885
rect 8113 21876 8125 21879
rect 7892 21848 8125 21876
rect 7892 21836 7898 21848
rect 8113 21845 8125 21848
rect 8159 21876 8171 21879
rect 8478 21876 8484 21888
rect 8159 21848 8484 21876
rect 8159 21845 8171 21848
rect 8113 21839 8171 21845
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 10778 21836 10784 21888
rect 10836 21836 10842 21888
rect 12894 21836 12900 21888
rect 12952 21836 12958 21888
rect 13262 21836 13268 21888
rect 13320 21876 13326 21888
rect 13357 21879 13415 21885
rect 13357 21876 13369 21879
rect 13320 21848 13369 21876
rect 13320 21836 13326 21848
rect 13357 21845 13369 21848
rect 13403 21876 13415 21879
rect 13446 21876 13452 21888
rect 13403 21848 13452 21876
rect 13403 21845 13415 21848
rect 13357 21839 13415 21845
rect 13446 21836 13452 21848
rect 13504 21836 13510 21888
rect 15010 21836 15016 21888
rect 15068 21876 15074 21888
rect 17034 21876 17040 21888
rect 15068 21848 17040 21876
rect 15068 21836 15074 21848
rect 17034 21836 17040 21848
rect 17092 21836 17098 21888
rect 17126 21836 17132 21888
rect 17184 21876 17190 21888
rect 21100 21885 21128 21916
rect 21606 21913 21618 21916
rect 21652 21913 21664 21947
rect 25838 21947 25896 21953
rect 25838 21944 25850 21947
rect 21606 21907 21664 21913
rect 25332 21916 25850 21944
rect 18049 21879 18107 21885
rect 18049 21876 18061 21879
rect 17184 21848 18061 21876
rect 17184 21836 17190 21848
rect 18049 21845 18061 21848
rect 18095 21845 18107 21879
rect 18049 21839 18107 21845
rect 21085 21879 21143 21885
rect 21085 21845 21097 21879
rect 21131 21845 21143 21879
rect 21085 21839 21143 21845
rect 22186 21836 22192 21888
rect 22244 21876 22250 21888
rect 25332 21885 25360 21916
rect 25838 21913 25850 21916
rect 25884 21913 25896 21947
rect 25838 21907 25896 21913
rect 30193 21947 30251 21953
rect 30193 21913 30205 21947
rect 30239 21944 30251 21947
rect 30650 21944 30656 21956
rect 30239 21916 30656 21944
rect 30239 21913 30251 21916
rect 30193 21907 30251 21913
rect 30650 21904 30656 21916
rect 30708 21904 30714 21956
rect 30742 21904 30748 21956
rect 30800 21944 30806 21956
rect 31036 21944 31064 21975
rect 32398 21972 32404 22024
rect 32456 22012 32462 22024
rect 32493 22015 32551 22021
rect 32493 22012 32505 22015
rect 32456 21984 32505 22012
rect 32456 21972 32462 21984
rect 32493 21981 32505 21984
rect 32539 21981 32551 22015
rect 32493 21975 32551 21981
rect 33134 21972 33140 22024
rect 33192 22012 33198 22024
rect 33321 22015 33379 22021
rect 33321 22012 33333 22015
rect 33192 21984 33333 22012
rect 33192 21972 33198 21984
rect 33321 21981 33333 21984
rect 33367 21981 33379 22015
rect 33321 21975 33379 21981
rect 30800 21916 31064 21944
rect 30800 21904 30806 21916
rect 22741 21879 22799 21885
rect 22741 21876 22753 21879
rect 22244 21848 22753 21876
rect 22244 21836 22250 21848
rect 22741 21845 22753 21848
rect 22787 21845 22799 21879
rect 22741 21839 22799 21845
rect 25317 21879 25375 21885
rect 25317 21845 25329 21879
rect 25363 21845 25375 21879
rect 25317 21839 25375 21845
rect 30558 21836 30564 21888
rect 30616 21836 30622 21888
rect 30834 21836 30840 21888
rect 30892 21836 30898 21888
rect 32122 21836 32128 21888
rect 32180 21836 32186 21888
rect 32582 21836 32588 21888
rect 32640 21836 32646 21888
rect 32953 21879 33011 21885
rect 32953 21845 32965 21879
rect 32999 21876 33011 21879
rect 33226 21876 33232 21888
rect 32999 21848 33232 21876
rect 32999 21845 33011 21848
rect 32953 21839 33011 21845
rect 33226 21836 33232 21848
rect 33284 21836 33290 21888
rect 33410 21836 33416 21888
rect 33468 21836 33474 21888
rect 1104 21786 36800 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 36800 21786
rect 1104 21712 36800 21734
rect 1946 21632 1952 21684
rect 2004 21632 2010 21684
rect 2225 21675 2283 21681
rect 2225 21641 2237 21675
rect 2271 21641 2283 21675
rect 2225 21635 2283 21641
rect 2685 21675 2743 21681
rect 2685 21641 2697 21675
rect 2731 21672 2743 21675
rect 2774 21672 2780 21684
rect 2731 21644 2780 21672
rect 2731 21641 2743 21644
rect 2685 21635 2743 21641
rect 2133 21539 2191 21545
rect 2133 21505 2145 21539
rect 2179 21536 2191 21539
rect 2240 21536 2268 21635
rect 2774 21632 2780 21644
rect 2832 21672 2838 21684
rect 3234 21672 3240 21684
rect 2832 21644 3240 21672
rect 2832 21632 2838 21644
rect 3234 21632 3240 21644
rect 3292 21632 3298 21684
rect 6178 21632 6184 21684
rect 6236 21632 6242 21684
rect 7282 21632 7288 21684
rect 7340 21672 7346 21684
rect 7929 21675 7987 21681
rect 7929 21672 7941 21675
rect 7340 21644 7941 21672
rect 7340 21632 7346 21644
rect 7929 21641 7941 21644
rect 7975 21641 7987 21675
rect 7929 21635 7987 21641
rect 11790 21632 11796 21684
rect 11848 21632 11854 21684
rect 11974 21632 11980 21684
rect 12032 21672 12038 21684
rect 15010 21672 15016 21684
rect 12032 21644 15016 21672
rect 12032 21632 12038 21644
rect 15010 21632 15016 21644
rect 15068 21632 15074 21684
rect 16761 21675 16819 21681
rect 16761 21641 16773 21675
rect 16807 21672 16819 21675
rect 16807 21644 17172 21672
rect 16807 21641 16819 21644
rect 16761 21635 16819 21641
rect 4062 21564 4068 21616
rect 4120 21604 4126 21616
rect 9309 21607 9367 21613
rect 4120 21576 4568 21604
rect 4120 21564 4126 21576
rect 2179 21508 2268 21536
rect 2593 21539 2651 21545
rect 2179 21505 2191 21508
rect 2133 21499 2191 21505
rect 2593 21505 2605 21539
rect 2639 21536 2651 21539
rect 2958 21536 2964 21548
rect 2639 21508 2964 21536
rect 2639 21505 2651 21508
rect 2593 21499 2651 21505
rect 2958 21496 2964 21508
rect 3016 21536 3022 21548
rect 4540 21545 4568 21576
rect 7392 21576 8892 21604
rect 7392 21548 7420 21576
rect 4525 21539 4583 21545
rect 3016 21508 4384 21536
rect 3016 21496 3022 21508
rect 2869 21471 2927 21477
rect 2869 21437 2881 21471
rect 2915 21468 2927 21471
rect 3142 21468 3148 21480
rect 2915 21440 3148 21468
rect 2915 21437 2927 21440
rect 2869 21431 2927 21437
rect 3142 21428 3148 21440
rect 3200 21428 3206 21480
rect 4356 21477 4384 21508
rect 4525 21505 4537 21539
rect 4571 21505 4583 21539
rect 4525 21499 4583 21505
rect 5258 21496 5264 21548
rect 5316 21496 5322 21548
rect 7190 21496 7196 21548
rect 7248 21496 7254 21548
rect 7285 21540 7343 21545
rect 7374 21540 7380 21548
rect 7285 21539 7380 21540
rect 7285 21505 7297 21539
rect 7331 21512 7380 21539
rect 7331 21505 7343 21512
rect 7285 21499 7343 21505
rect 7374 21496 7380 21512
rect 7432 21496 7438 21548
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21505 7803 21539
rect 7745 21499 7803 21505
rect 5442 21477 5448 21480
rect 4341 21471 4399 21477
rect 4341 21437 4353 21471
rect 4387 21437 4399 21471
rect 4341 21431 4399 21437
rect 5399 21471 5448 21477
rect 5399 21437 5411 21471
rect 5445 21437 5448 21471
rect 5399 21431 5448 21437
rect 4356 21400 4384 21431
rect 5442 21428 5448 21431
rect 5500 21428 5506 21480
rect 5537 21471 5595 21477
rect 5537 21437 5549 21471
rect 5583 21468 5595 21471
rect 6178 21468 6184 21480
rect 5583 21440 6184 21468
rect 5583 21437 5595 21440
rect 5537 21431 5595 21437
rect 6012 21412 6040 21440
rect 6178 21428 6184 21440
rect 6236 21428 6242 21480
rect 6825 21471 6883 21477
rect 6825 21437 6837 21471
rect 6871 21468 6883 21471
rect 7760 21468 7788 21499
rect 8018 21496 8024 21548
rect 8076 21496 8082 21548
rect 8662 21468 8668 21480
rect 6871 21440 8668 21468
rect 6871 21437 6883 21440
rect 6825 21431 6883 21437
rect 8662 21428 8668 21440
rect 8720 21428 8726 21480
rect 8864 21468 8892 21576
rect 9309 21573 9321 21607
rect 9355 21604 9367 21607
rect 10778 21604 10784 21616
rect 9355 21576 10784 21604
rect 9355 21573 9367 21576
rect 9309 21567 9367 21573
rect 10778 21564 10784 21576
rect 10836 21564 10842 21616
rect 14734 21604 14740 21616
rect 10888 21576 14740 21604
rect 8938 21496 8944 21548
rect 8996 21536 9002 21548
rect 9122 21536 9128 21548
rect 8996 21508 9128 21536
rect 8996 21496 9002 21508
rect 9122 21496 9128 21508
rect 9180 21536 9186 21548
rect 9493 21539 9551 21545
rect 9493 21536 9505 21539
rect 9180 21508 9505 21536
rect 9180 21496 9186 21508
rect 9493 21505 9505 21508
rect 9539 21505 9551 21539
rect 9493 21499 9551 21505
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 9674 21536 9680 21548
rect 9631 21508 9680 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 9674 21496 9680 21508
rect 9732 21536 9738 21548
rect 10888 21536 10916 21576
rect 14734 21564 14740 21576
rect 14792 21564 14798 21616
rect 17144 21604 17172 21644
rect 17770 21632 17776 21684
rect 17828 21672 17834 21684
rect 18417 21675 18475 21681
rect 18417 21672 18429 21675
rect 17828 21644 18429 21672
rect 17828 21632 17834 21644
rect 18417 21641 18429 21644
rect 18463 21641 18475 21675
rect 18417 21635 18475 21641
rect 21266 21632 21272 21684
rect 21324 21672 21330 21684
rect 21821 21675 21879 21681
rect 21821 21672 21833 21675
rect 21324 21644 21833 21672
rect 21324 21632 21330 21644
rect 21821 21641 21833 21644
rect 21867 21641 21879 21675
rect 22186 21672 22192 21684
rect 21821 21635 21879 21641
rect 22066 21644 22192 21672
rect 17282 21607 17340 21613
rect 17282 21604 17294 21607
rect 17144 21576 17294 21604
rect 17282 21573 17294 21576
rect 17328 21573 17340 21607
rect 17282 21567 17340 21573
rect 20070 21564 20076 21616
rect 20128 21604 20134 21616
rect 22066 21604 22094 21644
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 22278 21632 22284 21684
rect 22336 21632 22342 21684
rect 25041 21675 25099 21681
rect 25041 21641 25053 21675
rect 25087 21672 25099 21675
rect 26326 21672 26332 21684
rect 25087 21644 26332 21672
rect 25087 21641 25099 21644
rect 25041 21635 25099 21641
rect 26326 21632 26332 21644
rect 26384 21632 26390 21684
rect 28442 21632 28448 21684
rect 28500 21672 28506 21684
rect 28721 21675 28779 21681
rect 28721 21672 28733 21675
rect 28500 21644 28733 21672
rect 28500 21632 28506 21644
rect 28721 21641 28733 21644
rect 28767 21641 28779 21675
rect 28721 21635 28779 21641
rect 25314 21604 25320 21616
rect 20128 21576 22094 21604
rect 22388 21576 25320 21604
rect 20128 21564 20134 21576
rect 9732 21508 10916 21536
rect 11977 21539 12035 21545
rect 9732 21496 9738 21508
rect 11977 21505 11989 21539
rect 12023 21536 12035 21539
rect 12894 21536 12900 21548
rect 12023 21508 12900 21536
rect 12023 21505 12035 21508
rect 11977 21499 12035 21505
rect 12894 21496 12900 21508
rect 12952 21496 12958 21548
rect 15933 21539 15991 21545
rect 15933 21505 15945 21539
rect 15979 21536 15991 21539
rect 16850 21536 16856 21548
rect 15979 21508 16856 21536
rect 15979 21505 15991 21508
rect 15933 21499 15991 21505
rect 16850 21496 16856 21508
rect 16908 21496 16914 21548
rect 16942 21496 16948 21548
rect 17000 21496 17006 21548
rect 17034 21496 17040 21548
rect 17092 21496 17098 21548
rect 19702 21536 19708 21548
rect 17144 21508 19708 21536
rect 11514 21468 11520 21480
rect 8864 21440 11520 21468
rect 11514 21428 11520 21440
rect 11572 21428 11578 21480
rect 14274 21428 14280 21480
rect 14332 21468 14338 21480
rect 14332 21440 15976 21468
rect 14332 21428 14338 21440
rect 4614 21400 4620 21412
rect 4356 21372 4620 21400
rect 4614 21360 4620 21372
rect 4672 21360 4678 21412
rect 4798 21360 4804 21412
rect 4856 21400 4862 21412
rect 4985 21403 5043 21409
rect 4985 21400 4997 21403
rect 4856 21372 4997 21400
rect 4856 21360 4862 21372
rect 4985 21369 4997 21372
rect 5031 21369 5043 21403
rect 4985 21363 5043 21369
rect 5994 21360 6000 21412
rect 6052 21360 6058 21412
rect 9306 21360 9312 21412
rect 9364 21360 9370 21412
rect 14182 21360 14188 21412
rect 14240 21400 14246 21412
rect 15948 21400 15976 21440
rect 16022 21428 16028 21480
rect 16080 21428 16086 21480
rect 16209 21471 16267 21477
rect 16209 21437 16221 21471
rect 16255 21468 16267 21471
rect 16482 21468 16488 21480
rect 16255 21440 16488 21468
rect 16255 21437 16267 21440
rect 16209 21431 16267 21437
rect 16482 21428 16488 21440
rect 16540 21428 16546 21480
rect 17144 21468 17172 21508
rect 19702 21496 19708 21508
rect 19760 21536 19766 21548
rect 20625 21539 20683 21545
rect 19760 21508 20392 21536
rect 19760 21496 19766 21508
rect 20257 21471 20315 21477
rect 20257 21468 20269 21471
rect 17052 21440 17172 21468
rect 18064 21440 20269 21468
rect 17052 21400 17080 21440
rect 14240 21372 15700 21400
rect 15948 21372 17080 21400
rect 14240 21360 14246 21372
rect 5442 21292 5448 21344
rect 5500 21332 5506 21344
rect 5626 21332 5632 21344
rect 5500 21304 5632 21332
rect 5500 21292 5506 21304
rect 5626 21292 5632 21304
rect 5684 21292 5690 21344
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 7469 21335 7527 21341
rect 7469 21332 7481 21335
rect 6972 21304 7481 21332
rect 6972 21292 6978 21304
rect 7469 21301 7481 21304
rect 7515 21301 7527 21335
rect 7469 21295 7527 21301
rect 7558 21292 7564 21344
rect 7616 21292 7622 21344
rect 9766 21292 9772 21344
rect 9824 21332 9830 21344
rect 13722 21332 13728 21344
rect 9824 21304 13728 21332
rect 9824 21292 9830 21304
rect 13722 21292 13728 21304
rect 13780 21292 13786 21344
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 15565 21335 15623 21341
rect 15565 21332 15577 21335
rect 15528 21304 15577 21332
rect 15528 21292 15534 21304
rect 15565 21301 15577 21304
rect 15611 21301 15623 21335
rect 15672 21332 15700 21372
rect 18064 21332 18092 21440
rect 20257 21437 20269 21440
rect 20303 21437 20315 21471
rect 20364 21468 20392 21508
rect 20625 21505 20637 21539
rect 20671 21536 20683 21539
rect 22002 21536 22008 21548
rect 20671 21508 22008 21536
rect 20671 21505 20683 21508
rect 20625 21499 20683 21505
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 20714 21468 20720 21480
rect 20364 21440 20720 21468
rect 20257 21431 20315 21437
rect 20714 21428 20720 21440
rect 20772 21428 20778 21480
rect 20990 21428 20996 21480
rect 21048 21428 21054 21480
rect 22388 21468 22416 21576
rect 25314 21564 25320 21576
rect 25372 21564 25378 21616
rect 23106 21496 23112 21548
rect 23164 21496 23170 21548
rect 23382 21545 23388 21548
rect 23376 21499 23388 21545
rect 23382 21496 23388 21499
rect 23440 21496 23446 21548
rect 24486 21496 24492 21548
rect 24544 21536 24550 21548
rect 24949 21539 25007 21545
rect 24949 21536 24961 21539
rect 24544 21508 24961 21536
rect 24544 21496 24550 21508
rect 24949 21505 24961 21508
rect 24995 21505 25007 21539
rect 24949 21499 25007 21505
rect 26970 21496 26976 21548
rect 27028 21536 27034 21548
rect 28626 21536 28632 21548
rect 27028 21508 28632 21536
rect 27028 21496 27034 21508
rect 28626 21496 28632 21508
rect 28684 21496 28690 21548
rect 33318 21496 33324 21548
rect 33376 21496 33382 21548
rect 21100 21440 22416 21468
rect 22465 21471 22523 21477
rect 18138 21360 18144 21412
rect 18196 21400 18202 21412
rect 21100 21400 21128 21440
rect 22465 21437 22477 21471
rect 22511 21468 22523 21471
rect 22830 21468 22836 21480
rect 22511 21440 22836 21468
rect 22511 21437 22523 21440
rect 22465 21431 22523 21437
rect 22830 21428 22836 21440
rect 22888 21428 22894 21480
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24412 21440 25145 21468
rect 18196 21372 21128 21400
rect 21361 21403 21419 21409
rect 18196 21360 18202 21372
rect 21361 21369 21373 21403
rect 21407 21400 21419 21403
rect 21634 21400 21640 21412
rect 21407 21372 21640 21400
rect 21407 21369 21419 21372
rect 21361 21363 21419 21369
rect 21634 21360 21640 21372
rect 21692 21360 21698 21412
rect 15672 21304 18092 21332
rect 15565 21295 15623 21301
rect 20346 21292 20352 21344
rect 20404 21332 20410 21344
rect 20901 21335 20959 21341
rect 20901 21332 20913 21335
rect 20404 21304 20913 21332
rect 20404 21292 20410 21304
rect 20901 21301 20913 21304
rect 20947 21301 20959 21335
rect 20901 21295 20959 21301
rect 21450 21292 21456 21344
rect 21508 21292 21514 21344
rect 22922 21292 22928 21344
rect 22980 21332 22986 21344
rect 24412 21332 24440 21440
rect 25133 21437 25145 21440
rect 25179 21468 25191 21471
rect 28813 21471 28871 21477
rect 28813 21468 28825 21471
rect 25179 21440 28825 21468
rect 25179 21437 25191 21440
rect 25133 21431 25191 21437
rect 28813 21437 28825 21440
rect 28859 21468 28871 21471
rect 30834 21468 30840 21480
rect 28859 21440 30840 21468
rect 28859 21437 28871 21440
rect 28813 21431 28871 21437
rect 30834 21428 30840 21440
rect 30892 21428 30898 21480
rect 22980 21304 24440 21332
rect 22980 21292 22986 21304
rect 24486 21292 24492 21344
rect 24544 21292 24550 21344
rect 24578 21292 24584 21344
rect 24636 21292 24642 21344
rect 28261 21335 28319 21341
rect 28261 21301 28273 21335
rect 28307 21332 28319 21335
rect 29730 21332 29736 21344
rect 28307 21304 29736 21332
rect 28307 21301 28319 21304
rect 28261 21295 28319 21301
rect 29730 21292 29736 21304
rect 29788 21292 29794 21344
rect 31018 21292 31024 21344
rect 31076 21332 31082 21344
rect 31386 21332 31392 21344
rect 31076 21304 31392 21332
rect 31076 21292 31082 21304
rect 31386 21292 31392 21304
rect 31444 21292 31450 21344
rect 33137 21335 33195 21341
rect 33137 21301 33149 21335
rect 33183 21332 33195 21335
rect 33226 21332 33232 21344
rect 33183 21304 33232 21332
rect 33183 21301 33195 21304
rect 33137 21295 33195 21301
rect 33226 21292 33232 21304
rect 33284 21292 33290 21344
rect 1104 21242 36800 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 36800 21242
rect 1104 21168 36800 21190
rect 2682 21088 2688 21140
rect 2740 21128 2746 21140
rect 2740 21100 7880 21128
rect 2740 21088 2746 21100
rect 2792 21001 2820 21100
rect 6457 21063 6515 21069
rect 6457 21029 6469 21063
rect 6503 21060 6515 21063
rect 7653 21063 7711 21069
rect 7653 21060 7665 21063
rect 6503 21032 7665 21060
rect 6503 21029 6515 21032
rect 6457 21023 6515 21029
rect 7653 21029 7665 21032
rect 7699 21029 7711 21063
rect 7852 21060 7880 21100
rect 8662 21088 8668 21140
rect 8720 21128 8726 21140
rect 9858 21128 9864 21140
rect 8720 21100 9864 21128
rect 8720 21088 8726 21100
rect 9858 21088 9864 21100
rect 9916 21088 9922 21140
rect 9968 21100 14504 21128
rect 9674 21060 9680 21072
rect 7852 21032 9680 21060
rect 7653 21023 7711 21029
rect 9674 21020 9680 21032
rect 9732 21020 9738 21072
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20961 2835 20995
rect 2777 20955 2835 20961
rect 2976 20964 3924 20992
rect 2976 20936 3004 20964
rect 2593 20927 2651 20933
rect 2593 20893 2605 20927
rect 2639 20924 2651 20927
rect 2958 20924 2964 20936
rect 2639 20896 2964 20924
rect 2639 20893 2651 20896
rect 2593 20887 2651 20893
rect 2958 20884 2964 20896
rect 3016 20884 3022 20936
rect 3605 20927 3663 20933
rect 3605 20893 3617 20927
rect 3651 20924 3663 20927
rect 3896 20924 3924 20964
rect 3970 20952 3976 21004
rect 4028 20992 4034 21004
rect 4341 20995 4399 21001
rect 4341 20992 4353 20995
rect 4028 20964 4353 20992
rect 4028 20952 4034 20964
rect 4341 20961 4353 20964
rect 4387 20961 4399 20995
rect 4341 20955 4399 20961
rect 4614 20952 4620 21004
rect 4672 20952 4678 21004
rect 5258 20952 5264 21004
rect 5316 20952 5322 21004
rect 5350 20952 5356 21004
rect 5408 20992 5414 21004
rect 5537 20995 5595 21001
rect 5537 20992 5549 20995
rect 5408 20964 5549 20992
rect 5408 20952 5414 20964
rect 5537 20961 5549 20964
rect 5583 20961 5595 20995
rect 5537 20955 5595 20961
rect 5626 20952 5632 21004
rect 5684 21001 5690 21004
rect 5684 20995 5712 21001
rect 5700 20961 5712 20995
rect 5684 20955 5712 20961
rect 5684 20952 5690 20955
rect 7190 20952 7196 21004
rect 7248 20952 7254 21004
rect 9309 20995 9367 21001
rect 9309 20961 9321 20995
rect 9355 20992 9367 20995
rect 9582 20992 9588 21004
rect 9355 20964 9588 20992
rect 9355 20961 9367 20964
rect 9309 20955 9367 20961
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 9968 20992 9996 21100
rect 10870 21020 10876 21072
rect 10928 21020 10934 21072
rect 13725 21063 13783 21069
rect 11348 21032 12434 21060
rect 9784 20964 9996 20992
rect 10965 20995 11023 21001
rect 4062 20924 4068 20936
rect 3651 20896 3832 20924
rect 3896 20896 4068 20924
rect 3651 20893 3663 20896
rect 3605 20887 3663 20893
rect 2682 20816 2688 20868
rect 2740 20856 2746 20868
rect 2774 20856 2780 20868
rect 2740 20828 2780 20856
rect 2740 20816 2746 20828
rect 2774 20816 2780 20828
rect 2832 20816 2838 20868
rect 2038 20748 2044 20800
rect 2096 20788 2102 20800
rect 2225 20791 2283 20797
rect 2225 20788 2237 20791
rect 2096 20760 2237 20788
rect 2096 20748 2102 20760
rect 2225 20757 2237 20760
rect 2271 20757 2283 20791
rect 2225 20751 2283 20757
rect 3418 20748 3424 20800
rect 3476 20748 3482 20800
rect 3804 20797 3832 20896
rect 4062 20884 4068 20896
rect 4120 20924 4126 20936
rect 4801 20927 4859 20933
rect 4801 20924 4813 20927
rect 4120 20896 4813 20924
rect 4120 20884 4126 20896
rect 4801 20893 4813 20896
rect 4847 20893 4859 20927
rect 4801 20887 4859 20893
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 6914 20884 6920 20936
rect 6972 20884 6978 20936
rect 7006 20884 7012 20936
rect 7064 20884 7070 20936
rect 7285 20927 7343 20933
rect 7285 20893 7297 20927
rect 7331 20924 7343 20927
rect 7558 20924 7564 20936
rect 7331 20896 7564 20924
rect 7331 20893 7343 20896
rect 7285 20887 7343 20893
rect 7558 20884 7564 20896
rect 7616 20884 7622 20936
rect 8018 20884 8024 20936
rect 8076 20924 8082 20936
rect 9401 20927 9459 20933
rect 9401 20924 9413 20927
rect 8076 20896 9413 20924
rect 8076 20884 8082 20896
rect 9401 20893 9413 20896
rect 9447 20924 9459 20927
rect 9784 20924 9812 20964
rect 10965 20961 10977 20995
rect 11011 20992 11023 20995
rect 11238 20992 11244 21004
rect 11011 20964 11244 20992
rect 11011 20961 11023 20964
rect 10965 20955 11023 20961
rect 11238 20952 11244 20964
rect 11296 20952 11302 21004
rect 9447 20896 9812 20924
rect 9447 20893 9459 20896
rect 9401 20887 9459 20893
rect 9858 20884 9864 20936
rect 9916 20924 9922 20936
rect 11057 20927 11115 20933
rect 11057 20924 11069 20927
rect 9916 20896 11069 20924
rect 9916 20884 9922 20896
rect 11057 20893 11069 20896
rect 11103 20924 11115 20927
rect 11348 20924 11376 21032
rect 11422 20952 11428 21004
rect 11480 20952 11486 21004
rect 11514 20952 11520 21004
rect 11572 20992 11578 21004
rect 12406 20992 12434 21032
rect 13725 21029 13737 21063
rect 13771 21060 13783 21063
rect 14366 21060 14372 21072
rect 13771 21032 14372 21060
rect 13771 21029 13783 21032
rect 13725 21023 13783 21029
rect 14366 21020 14372 21032
rect 14424 21020 14430 21072
rect 14182 20992 14188 21004
rect 11572 20964 12296 20992
rect 12406 20964 14188 20992
rect 11572 20952 11578 20964
rect 11977 20927 12035 20933
rect 11977 20924 11989 20927
rect 11103 20896 11989 20924
rect 11103 20893 11115 20896
rect 11057 20887 11115 20893
rect 11977 20893 11989 20896
rect 12023 20893 12035 20927
rect 11977 20887 12035 20893
rect 12066 20884 12072 20936
rect 12124 20924 12130 20936
rect 12268 20933 12296 20964
rect 14182 20952 14188 20964
rect 14240 20952 14246 21004
rect 12161 20927 12219 20933
rect 12161 20924 12173 20927
rect 12124 20896 12173 20924
rect 12124 20884 12130 20896
rect 12161 20893 12173 20896
rect 12207 20893 12219 20927
rect 12161 20887 12219 20893
rect 12253 20927 12311 20933
rect 12253 20893 12265 20927
rect 12299 20924 12311 20927
rect 14274 20924 14280 20936
rect 12299 20896 14280 20924
rect 12299 20893 12311 20896
rect 12253 20887 12311 20893
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 14476 20924 14504 21100
rect 14550 21088 14556 21140
rect 14608 21128 14614 21140
rect 16301 21131 16359 21137
rect 14608 21100 15976 21128
rect 14608 21088 14614 21100
rect 14553 20995 14611 21001
rect 14553 20961 14565 20995
rect 14599 20992 14611 20995
rect 14599 20964 15056 20992
rect 14599 20961 14611 20964
rect 14553 20955 14611 20961
rect 14645 20927 14703 20933
rect 14645 20924 14657 20927
rect 14476 20896 14657 20924
rect 14645 20893 14657 20896
rect 14691 20893 14703 20927
rect 14645 20887 14703 20893
rect 4157 20859 4215 20865
rect 4157 20825 4169 20859
rect 4203 20856 4215 20859
rect 4430 20856 4436 20868
rect 4203 20828 4436 20856
rect 4203 20825 4215 20828
rect 4157 20819 4215 20825
rect 4430 20816 4436 20828
rect 4488 20856 4494 20868
rect 4488 20828 4844 20856
rect 4488 20816 4494 20828
rect 3789 20791 3847 20797
rect 3789 20757 3801 20791
rect 3835 20757 3847 20791
rect 3789 20751 3847 20757
rect 3878 20748 3884 20800
rect 3936 20788 3942 20800
rect 4249 20791 4307 20797
rect 4249 20788 4261 20791
rect 3936 20760 4261 20788
rect 3936 20748 3942 20760
rect 4249 20757 4261 20760
rect 4295 20788 4307 20791
rect 4614 20788 4620 20800
rect 4295 20760 4620 20788
rect 4295 20757 4307 20760
rect 4249 20751 4307 20757
rect 4614 20748 4620 20760
rect 4672 20748 4678 20800
rect 4816 20788 4844 20828
rect 7374 20816 7380 20868
rect 7432 20816 7438 20868
rect 8941 20859 8999 20865
rect 8941 20825 8953 20859
rect 8987 20856 8999 20859
rect 9306 20856 9312 20868
rect 8987 20828 9312 20856
rect 8987 20825 8999 20828
rect 8941 20819 8999 20825
rect 9306 20816 9312 20828
rect 9364 20856 9370 20868
rect 9766 20856 9772 20868
rect 9364 20828 9772 20856
rect 9364 20816 9370 20828
rect 9766 20816 9772 20828
rect 9824 20816 9830 20868
rect 10502 20816 10508 20868
rect 10560 20856 10566 20868
rect 11882 20856 11888 20868
rect 10560 20828 11888 20856
rect 10560 20816 10566 20828
rect 11882 20816 11888 20828
rect 11940 20816 11946 20868
rect 13446 20816 13452 20868
rect 13504 20856 13510 20868
rect 14550 20856 14556 20868
rect 13504 20828 14556 20856
rect 13504 20816 13510 20828
rect 14550 20816 14556 20828
rect 14608 20816 14614 20868
rect 14660 20856 14688 20887
rect 14918 20884 14924 20936
rect 14976 20884 14982 20936
rect 15028 20924 15056 20964
rect 15746 20924 15752 20936
rect 15028 20896 15752 20924
rect 15746 20884 15752 20896
rect 15804 20884 15810 20936
rect 15948 20924 15976 21100
rect 16301 21097 16313 21131
rect 16347 21128 16359 21131
rect 16850 21128 16856 21140
rect 16347 21100 16856 21128
rect 16347 21097 16359 21100
rect 16301 21091 16359 21097
rect 16850 21088 16856 21100
rect 16908 21088 16914 21140
rect 16942 21088 16948 21140
rect 17000 21128 17006 21140
rect 17313 21131 17371 21137
rect 17313 21128 17325 21131
rect 17000 21100 17325 21128
rect 17000 21088 17006 21100
rect 17313 21097 17325 21100
rect 17359 21097 17371 21131
rect 17313 21091 17371 21097
rect 17402 21088 17408 21140
rect 17460 21128 17466 21140
rect 17770 21128 17776 21140
rect 17460 21100 17776 21128
rect 17460 21088 17466 21100
rect 17770 21088 17776 21100
rect 17828 21088 17834 21140
rect 19702 21088 19708 21140
rect 19760 21088 19766 21140
rect 20346 21088 20352 21140
rect 20404 21088 20410 21140
rect 20990 21088 20996 21140
rect 21048 21128 21054 21140
rect 21048 21100 23336 21128
rect 21048 21088 21054 21100
rect 17126 21020 17132 21072
rect 17184 21020 17190 21072
rect 19426 21060 19432 21072
rect 17297 21032 19432 21060
rect 16761 20927 16819 20933
rect 16761 20924 16773 20927
rect 15948 20896 16773 20924
rect 16761 20893 16773 20896
rect 16807 20924 16819 20927
rect 17297 20924 17325 21032
rect 19426 21020 19432 21032
rect 19484 21020 19490 21072
rect 20714 21020 20720 21072
rect 20772 21060 20778 21072
rect 21174 21060 21180 21072
rect 20772 21032 21180 21060
rect 20772 21020 20778 21032
rect 21174 21020 21180 21032
rect 21232 21020 21238 21072
rect 17586 20952 17592 21004
rect 17644 20992 17650 21004
rect 17773 20995 17831 21001
rect 17773 20992 17785 20995
rect 17644 20964 17785 20992
rect 17644 20952 17650 20964
rect 17773 20961 17785 20964
rect 17819 20961 17831 20995
rect 17773 20955 17831 20961
rect 17862 20952 17868 21004
rect 17920 20952 17926 21004
rect 18509 20995 18567 21001
rect 18509 20961 18521 20995
rect 18555 20992 18567 20995
rect 18690 20992 18696 21004
rect 18555 20964 18696 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 18690 20952 18696 20964
rect 18748 20952 18754 21004
rect 20533 20995 20591 21001
rect 20533 20992 20545 20995
rect 20180 20964 20545 20992
rect 16807 20896 17325 20924
rect 16807 20893 16819 20896
rect 16761 20887 16819 20893
rect 17402 20884 17408 20936
rect 17460 20924 17466 20936
rect 17681 20927 17739 20933
rect 17681 20924 17693 20927
rect 17460 20896 17693 20924
rect 17460 20884 17466 20896
rect 17681 20893 17693 20896
rect 17727 20893 17739 20927
rect 18601 20927 18659 20933
rect 18601 20924 18613 20927
rect 17681 20887 17739 20893
rect 17788 20896 18613 20924
rect 15188 20859 15246 20865
rect 14660 20828 14964 20856
rect 5626 20788 5632 20800
rect 4816 20760 5632 20788
rect 5626 20748 5632 20760
rect 5684 20748 5690 20800
rect 6733 20791 6791 20797
rect 6733 20757 6745 20791
rect 6779 20788 6791 20791
rect 7282 20788 7288 20800
rect 6779 20760 7288 20788
rect 6779 20757 6791 20760
rect 6733 20751 6791 20757
rect 7282 20748 7288 20760
rect 7340 20748 7346 20800
rect 7837 20791 7895 20797
rect 7837 20757 7849 20791
rect 7883 20788 7895 20791
rect 8478 20788 8484 20800
rect 7883 20760 8484 20788
rect 7883 20757 7895 20760
rect 7837 20751 7895 20757
rect 8478 20748 8484 20760
rect 8536 20748 8542 20800
rect 9582 20748 9588 20800
rect 9640 20748 9646 20800
rect 11698 20748 11704 20800
rect 11756 20748 11762 20800
rect 11790 20748 11796 20800
rect 11848 20748 11854 20800
rect 13906 20748 13912 20800
rect 13964 20748 13970 20800
rect 14826 20748 14832 20800
rect 14884 20748 14890 20800
rect 14936 20788 14964 20828
rect 15188 20825 15200 20859
rect 15234 20856 15246 20859
rect 15286 20856 15292 20868
rect 15234 20828 15292 20856
rect 15234 20825 15246 20828
rect 15188 20819 15246 20825
rect 15286 20816 15292 20828
rect 15344 20816 15350 20868
rect 17788 20856 17816 20896
rect 18601 20893 18613 20896
rect 18647 20924 18659 20927
rect 19702 20924 19708 20936
rect 18647 20896 19708 20924
rect 18647 20893 18659 20896
rect 18601 20887 18659 20893
rect 19702 20884 19708 20896
rect 19760 20884 19766 20936
rect 19886 20884 19892 20936
rect 19944 20884 19950 20936
rect 20070 20884 20076 20936
rect 20128 20884 20134 20936
rect 20180 20933 20208 20964
rect 20533 20961 20545 20964
rect 20579 20961 20591 20995
rect 21450 20992 21456 21004
rect 20533 20955 20591 20961
rect 20640 20964 21456 20992
rect 20165 20927 20223 20933
rect 20165 20893 20177 20927
rect 20211 20893 20223 20927
rect 20165 20887 20223 20893
rect 20441 20927 20499 20933
rect 20441 20893 20453 20927
rect 20487 20924 20499 20927
rect 20640 20924 20668 20964
rect 21450 20952 21456 20964
rect 21508 20952 21514 21004
rect 23308 20992 23336 21100
rect 23382 21088 23388 21140
rect 23440 21088 23446 21140
rect 27062 21128 27068 21140
rect 24780 21100 27068 21128
rect 24780 21001 24808 21100
rect 27062 21088 27068 21100
rect 27120 21088 27126 21140
rect 27249 21131 27307 21137
rect 27249 21097 27261 21131
rect 27295 21128 27307 21131
rect 27893 21131 27951 21137
rect 27893 21128 27905 21131
rect 27295 21100 27905 21128
rect 27295 21097 27307 21100
rect 27249 21091 27307 21097
rect 27893 21097 27905 21100
rect 27939 21097 27951 21131
rect 27893 21091 27951 21097
rect 27982 21088 27988 21140
rect 28040 21088 28046 21140
rect 28626 21088 28632 21140
rect 28684 21128 28690 21140
rect 29365 21131 29423 21137
rect 29365 21128 29377 21131
rect 28684 21100 29377 21128
rect 28684 21088 28690 21100
rect 29365 21097 29377 21100
rect 29411 21097 29423 21131
rect 29365 21091 29423 21097
rect 31202 21088 31208 21140
rect 31260 21128 31266 21140
rect 31662 21128 31668 21140
rect 31260 21100 31668 21128
rect 31260 21088 31266 21100
rect 31662 21088 31668 21100
rect 31720 21088 31726 21140
rect 32030 21088 32036 21140
rect 32088 21128 32094 21140
rect 32309 21131 32367 21137
rect 32309 21128 32321 21131
rect 32088 21100 32321 21128
rect 32088 21088 32094 21100
rect 32309 21097 32321 21100
rect 32355 21097 32367 21131
rect 32309 21091 32367 21097
rect 25130 21020 25136 21072
rect 25188 21020 25194 21072
rect 27154 21060 27160 21072
rect 25700 21032 27160 21060
rect 25700 21001 25728 21032
rect 27154 21020 27160 21032
rect 27212 21020 27218 21072
rect 27709 21063 27767 21069
rect 27709 21029 27721 21063
rect 27755 21060 27767 21063
rect 28000 21060 28028 21088
rect 27755 21032 28028 21060
rect 30837 21063 30895 21069
rect 27755 21029 27767 21032
rect 27709 21023 27767 21029
rect 30837 21029 30849 21063
rect 30883 21060 30895 21063
rect 31018 21060 31024 21072
rect 30883 21032 31024 21060
rect 30883 21029 30895 21032
rect 30837 21023 30895 21029
rect 31018 21020 31024 21032
rect 31076 21020 31082 21072
rect 31389 21063 31447 21069
rect 31389 21029 31401 21063
rect 31435 21060 31447 21063
rect 31754 21060 31760 21072
rect 31435 21032 31760 21060
rect 31435 21029 31447 21032
rect 31389 21023 31447 21029
rect 31754 21020 31760 21032
rect 31812 21060 31818 21072
rect 32861 21063 32919 21069
rect 32861 21060 32873 21063
rect 31812 21032 32873 21060
rect 31812 21020 31818 21032
rect 32861 21029 32873 21032
rect 32907 21060 32919 21063
rect 33042 21060 33048 21072
rect 32907 21032 33048 21060
rect 32907 21029 32919 21032
rect 32861 21023 32919 21029
rect 33042 21020 33048 21032
rect 33100 21020 33106 21072
rect 24765 20995 24823 21001
rect 24765 20992 24777 20995
rect 23308 20964 24777 20992
rect 24765 20961 24777 20964
rect 24811 20961 24823 20995
rect 24765 20955 24823 20961
rect 25685 20995 25743 21001
rect 25685 20961 25697 20995
rect 25731 20961 25743 20995
rect 25685 20955 25743 20961
rect 25777 20995 25835 21001
rect 25777 20961 25789 20995
rect 25823 20992 25835 20995
rect 25958 20992 25964 21004
rect 25823 20964 25964 20992
rect 25823 20961 25835 20964
rect 25777 20955 25835 20961
rect 25958 20952 25964 20964
rect 26016 20992 26022 21004
rect 26421 20995 26479 21001
rect 26016 20964 26188 20992
rect 26016 20952 26022 20964
rect 20487 20896 20668 20924
rect 20717 20927 20775 20933
rect 20487 20893 20499 20896
rect 20441 20887 20499 20893
rect 20717 20893 20729 20927
rect 20763 20893 20775 20927
rect 20717 20887 20775 20893
rect 15396 20828 17816 20856
rect 15396 20788 15424 20828
rect 17954 20816 17960 20868
rect 18012 20856 18018 20868
rect 18785 20859 18843 20865
rect 18785 20856 18797 20859
rect 18012 20828 18797 20856
rect 18012 20816 18018 20828
rect 18785 20825 18797 20828
rect 18831 20825 18843 20859
rect 18785 20819 18843 20825
rect 19610 20816 19616 20868
rect 19668 20816 19674 20868
rect 20732 20856 20760 20887
rect 20806 20884 20812 20936
rect 20864 20924 20870 20936
rect 20901 20927 20959 20933
rect 20901 20924 20913 20927
rect 20864 20896 20913 20924
rect 20864 20884 20870 20896
rect 20901 20893 20913 20896
rect 20947 20893 20959 20927
rect 20901 20887 20959 20893
rect 20993 20927 21051 20933
rect 20993 20893 21005 20927
rect 21039 20924 21051 20927
rect 21174 20924 21180 20936
rect 21039 20896 21180 20924
rect 21039 20893 21051 20896
rect 20993 20887 21051 20893
rect 21174 20884 21180 20896
rect 21232 20884 21238 20936
rect 23569 20927 23627 20933
rect 23569 20893 23581 20927
rect 23615 20924 23627 20927
rect 24578 20924 24584 20936
rect 23615 20896 24584 20924
rect 23615 20893 23627 20896
rect 23569 20887 23627 20893
rect 24578 20884 24584 20896
rect 24636 20884 24642 20936
rect 26160 20924 26188 20964
rect 26421 20961 26433 20995
rect 26467 20992 26479 20995
rect 26602 20992 26608 21004
rect 26467 20964 26608 20992
rect 26467 20961 26479 20964
rect 26421 20955 26479 20961
rect 26602 20952 26608 20964
rect 26660 20952 26666 21004
rect 26697 20995 26755 21001
rect 26697 20961 26709 20995
rect 26743 20992 26755 20995
rect 26743 20964 27384 20992
rect 26743 20961 26755 20964
rect 26697 20955 26755 20961
rect 26326 20924 26332 20936
rect 26160 20896 26332 20924
rect 26326 20884 26332 20896
rect 26384 20924 26390 20936
rect 26513 20927 26571 20933
rect 26513 20924 26525 20927
rect 26384 20896 26525 20924
rect 26384 20884 26390 20896
rect 26513 20893 26525 20896
rect 26559 20893 26571 20927
rect 26513 20887 26571 20893
rect 26786 20884 26792 20936
rect 26844 20924 26850 20936
rect 27356 20933 27384 20964
rect 27798 20952 27804 21004
rect 27856 20992 27862 21004
rect 27985 20995 28043 21001
rect 27985 20992 27997 20995
rect 27856 20964 27997 20992
rect 27856 20952 27862 20964
rect 27985 20961 27997 20964
rect 28031 20961 28043 20995
rect 27985 20955 28043 20961
rect 30377 20995 30435 21001
rect 30377 20961 30389 20995
rect 30423 20992 30435 20995
rect 30742 20992 30748 21004
rect 30423 20964 30748 20992
rect 30423 20961 30435 20964
rect 30377 20955 30435 20961
rect 30742 20952 30748 20964
rect 30800 20952 30806 21004
rect 30926 20952 30932 21004
rect 30984 20992 30990 21004
rect 30984 20964 32720 20992
rect 30984 20952 30990 20964
rect 26973 20927 27031 20933
rect 26973 20924 26985 20927
rect 26844 20896 26985 20924
rect 26844 20884 26850 20896
rect 26973 20893 26985 20896
rect 27019 20893 27031 20927
rect 26973 20887 27031 20893
rect 27065 20927 27123 20933
rect 27065 20893 27077 20927
rect 27111 20893 27123 20927
rect 27065 20887 27123 20893
rect 27341 20927 27399 20933
rect 27341 20893 27353 20927
rect 27387 20893 27399 20927
rect 27341 20887 27399 20893
rect 24302 20856 24308 20868
rect 20732 20828 24308 20856
rect 14936 20760 15424 20788
rect 17221 20791 17279 20797
rect 17221 20757 17233 20791
rect 17267 20788 17279 20791
rect 17586 20788 17592 20800
rect 17267 20760 17592 20788
rect 17267 20757 17279 20760
rect 17221 20751 17279 20757
rect 17586 20748 17592 20760
rect 17644 20748 17650 20800
rect 17862 20748 17868 20800
rect 17920 20788 17926 20800
rect 18138 20788 18144 20800
rect 17920 20760 18144 20788
rect 17920 20748 17926 20760
rect 18138 20748 18144 20760
rect 18196 20748 18202 20800
rect 18414 20748 18420 20800
rect 18472 20788 18478 20800
rect 20732 20788 20760 20828
rect 24302 20816 24308 20828
rect 24360 20816 24366 20868
rect 24854 20816 24860 20868
rect 24912 20856 24918 20868
rect 25961 20859 26019 20865
rect 25961 20856 25973 20859
rect 24912 20828 25973 20856
rect 24912 20816 24918 20828
rect 25961 20825 25973 20828
rect 26007 20825 26019 20859
rect 25961 20819 26019 20825
rect 18472 20760 20760 20788
rect 18472 20748 18478 20760
rect 25222 20748 25228 20800
rect 25280 20748 25286 20800
rect 25314 20748 25320 20800
rect 25372 20788 25378 20800
rect 26053 20791 26111 20797
rect 26053 20788 26065 20791
rect 25372 20760 26065 20788
rect 25372 20748 25378 20760
rect 26053 20757 26065 20760
rect 26099 20788 26111 20791
rect 26142 20788 26148 20800
rect 26099 20760 26148 20788
rect 26099 20757 26111 20760
rect 26053 20751 26111 20757
rect 26142 20748 26148 20760
rect 26200 20748 26206 20800
rect 26510 20748 26516 20800
rect 26568 20788 26574 20800
rect 26789 20791 26847 20797
rect 26789 20788 26801 20791
rect 26568 20760 26801 20788
rect 26568 20748 26574 20760
rect 26789 20757 26801 20760
rect 26835 20757 26847 20791
rect 27080 20788 27108 20887
rect 29730 20884 29736 20936
rect 29788 20884 29794 20936
rect 30469 20927 30527 20933
rect 30469 20893 30481 20927
rect 30515 20924 30527 20927
rect 30558 20924 30564 20936
rect 30515 20896 30564 20924
rect 30515 20893 30527 20896
rect 30469 20887 30527 20893
rect 30558 20884 30564 20896
rect 30616 20924 30622 20936
rect 31202 20924 31208 20936
rect 30616 20896 31208 20924
rect 30616 20884 30622 20896
rect 31202 20884 31208 20896
rect 31260 20924 31266 20936
rect 31757 20927 31815 20933
rect 31757 20924 31769 20927
rect 31260 20896 31769 20924
rect 31260 20884 31266 20896
rect 31757 20893 31769 20896
rect 31803 20893 31815 20927
rect 31757 20887 31815 20893
rect 32122 20884 32128 20936
rect 32180 20884 32186 20936
rect 32692 20933 32720 20964
rect 33134 20952 33140 21004
rect 33192 20952 33198 21004
rect 32677 20927 32735 20933
rect 32677 20893 32689 20927
rect 32723 20893 32735 20927
rect 32677 20887 32735 20893
rect 27154 20816 27160 20868
rect 27212 20856 27218 20868
rect 27433 20859 27491 20865
rect 27433 20856 27445 20859
rect 27212 20828 27445 20856
rect 27212 20816 27218 20828
rect 27433 20825 27445 20828
rect 27479 20825 27491 20859
rect 27433 20819 27491 20825
rect 28252 20859 28310 20865
rect 28252 20825 28264 20859
rect 28298 20856 28310 20859
rect 31665 20859 31723 20865
rect 28298 20828 29592 20856
rect 28298 20825 28310 20828
rect 28252 20819 28310 20825
rect 28074 20788 28080 20800
rect 27080 20760 28080 20788
rect 26789 20751 26847 20757
rect 28074 20748 28080 20760
rect 28132 20748 28138 20800
rect 29564 20797 29592 20828
rect 31665 20825 31677 20859
rect 31711 20856 31723 20859
rect 32030 20856 32036 20868
rect 31711 20828 32036 20856
rect 31711 20825 31723 20828
rect 31665 20819 31723 20825
rect 32030 20816 32036 20828
rect 32088 20816 32094 20868
rect 32692 20856 32720 20887
rect 33226 20884 33232 20936
rect 33284 20924 33290 20936
rect 33393 20927 33451 20933
rect 33393 20924 33405 20927
rect 33284 20896 33405 20924
rect 33284 20884 33290 20896
rect 33393 20893 33405 20896
rect 33439 20893 33451 20927
rect 33393 20887 33451 20893
rect 36081 20859 36139 20865
rect 32692 20828 34560 20856
rect 29549 20791 29607 20797
rect 29549 20757 29561 20791
rect 29595 20757 29607 20791
rect 29549 20751 29607 20757
rect 30374 20748 30380 20800
rect 30432 20788 30438 20800
rect 31205 20791 31263 20797
rect 31205 20788 31217 20791
rect 30432 20760 31217 20788
rect 30432 20748 30438 20760
rect 31205 20757 31217 20760
rect 31251 20757 31263 20791
rect 31205 20751 31263 20757
rect 31294 20748 31300 20800
rect 31352 20788 31358 20800
rect 31573 20791 31631 20797
rect 31573 20788 31585 20791
rect 31352 20760 31585 20788
rect 31352 20748 31358 20760
rect 31573 20757 31585 20760
rect 31619 20757 31631 20791
rect 31573 20751 31631 20757
rect 31938 20748 31944 20800
rect 31996 20748 32002 20800
rect 34532 20797 34560 20828
rect 36081 20825 36093 20859
rect 36127 20856 36139 20859
rect 36262 20856 36268 20868
rect 36127 20828 36268 20856
rect 36127 20825 36139 20828
rect 36081 20819 36139 20825
rect 36262 20816 36268 20828
rect 36320 20816 36326 20868
rect 34517 20791 34575 20797
rect 34517 20757 34529 20791
rect 34563 20757 34575 20791
rect 34517 20751 34575 20757
rect 36354 20748 36360 20800
rect 36412 20748 36418 20800
rect 1104 20698 36800 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 36800 20698
rect 1104 20624 36800 20646
rect 2869 20587 2927 20593
rect 2869 20553 2881 20587
rect 2915 20584 2927 20587
rect 2958 20584 2964 20596
rect 2915 20556 2964 20584
rect 2915 20553 2927 20556
rect 2869 20547 2927 20553
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 4430 20544 4436 20596
rect 4488 20544 4494 20596
rect 7650 20544 7656 20596
rect 7708 20584 7714 20596
rect 8113 20587 8171 20593
rect 8113 20584 8125 20587
rect 7708 20556 8125 20584
rect 7708 20544 7714 20556
rect 8113 20553 8125 20556
rect 8159 20553 8171 20587
rect 8113 20547 8171 20553
rect 8754 20544 8760 20596
rect 8812 20544 8818 20596
rect 14461 20587 14519 20593
rect 14461 20553 14473 20587
rect 14507 20584 14519 20587
rect 15194 20584 15200 20596
rect 14507 20556 15200 20584
rect 14507 20553 14519 20556
rect 14461 20547 14519 20553
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 15286 20544 15292 20596
rect 15344 20544 15350 20596
rect 18325 20587 18383 20593
rect 18325 20553 18337 20587
rect 18371 20584 18383 20587
rect 18874 20584 18880 20596
rect 18371 20556 18880 20584
rect 18371 20553 18383 20556
rect 18325 20547 18383 20553
rect 18874 20544 18880 20556
rect 18932 20544 18938 20596
rect 19334 20584 19340 20596
rect 19306 20544 19340 20584
rect 19392 20544 19398 20596
rect 19426 20544 19432 20596
rect 19484 20544 19490 20596
rect 20070 20544 20076 20596
rect 20128 20584 20134 20596
rect 20625 20587 20683 20593
rect 20625 20584 20637 20587
rect 20128 20556 20637 20584
rect 20128 20544 20134 20556
rect 20625 20553 20637 20556
rect 20671 20553 20683 20587
rect 20625 20547 20683 20553
rect 22278 20544 22284 20596
rect 22336 20544 22342 20596
rect 25225 20587 25283 20593
rect 25225 20553 25237 20587
rect 25271 20584 25283 20587
rect 25866 20584 25872 20596
rect 25271 20556 25872 20584
rect 25271 20553 25283 20556
rect 25225 20547 25283 20553
rect 25866 20544 25872 20556
rect 25924 20544 25930 20596
rect 27154 20544 27160 20596
rect 27212 20584 27218 20596
rect 27709 20587 27767 20593
rect 27709 20584 27721 20587
rect 27212 20556 27721 20584
rect 27212 20544 27218 20556
rect 27709 20553 27721 20556
rect 27755 20553 27767 20587
rect 27709 20547 27767 20553
rect 28074 20544 28080 20596
rect 28132 20544 28138 20596
rect 28537 20587 28595 20593
rect 28537 20553 28549 20587
rect 28583 20584 28595 20587
rect 29270 20584 29276 20596
rect 28583 20556 29276 20584
rect 28583 20553 28595 20556
rect 28537 20547 28595 20553
rect 29270 20544 29276 20556
rect 29328 20544 29334 20596
rect 30650 20544 30656 20596
rect 30708 20544 30714 20596
rect 32122 20544 32128 20596
rect 32180 20584 32186 20596
rect 33505 20587 33563 20593
rect 33505 20584 33517 20587
rect 32180 20556 33517 20584
rect 32180 20544 32186 20556
rect 33505 20553 33517 20556
rect 33551 20553 33563 20587
rect 33505 20547 33563 20553
rect 3320 20519 3378 20525
rect 1504 20488 2774 20516
rect 1504 20460 1532 20488
rect 1486 20408 1492 20460
rect 1544 20408 1550 20460
rect 1762 20457 1768 20460
rect 1756 20411 1768 20457
rect 1762 20408 1768 20411
rect 1820 20408 1826 20460
rect 2746 20448 2774 20488
rect 3320 20485 3332 20519
rect 3366 20516 3378 20519
rect 3418 20516 3424 20528
rect 3366 20488 3424 20516
rect 3366 20485 3378 20488
rect 3320 20479 3378 20485
rect 3418 20476 3424 20488
rect 3476 20476 3482 20528
rect 11790 20516 11796 20528
rect 10980 20488 11796 20516
rect 3053 20451 3111 20457
rect 3053 20448 3065 20451
rect 2746 20420 3065 20448
rect 3053 20417 3065 20420
rect 3099 20417 3111 20451
rect 3053 20411 3111 20417
rect 7282 20408 7288 20460
rect 7340 20448 7346 20460
rect 7377 20451 7435 20457
rect 7377 20448 7389 20451
rect 7340 20420 7389 20448
rect 7340 20408 7346 20420
rect 7377 20417 7389 20420
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 8202 20408 8208 20460
rect 8260 20448 8266 20460
rect 8665 20451 8723 20457
rect 8665 20448 8677 20451
rect 8260 20420 8677 20448
rect 8260 20408 8266 20420
rect 8665 20417 8677 20420
rect 8711 20417 8723 20451
rect 8665 20411 8723 20417
rect 9306 20408 9312 20460
rect 9364 20408 9370 20460
rect 10870 20408 10876 20460
rect 10928 20408 10934 20460
rect 10980 20457 11008 20488
rect 11790 20476 11796 20488
rect 11848 20476 11854 20528
rect 11882 20476 11888 20528
rect 11940 20516 11946 20528
rect 19306 20516 19334 20544
rect 11940 20488 19334 20516
rect 19444 20516 19472 20544
rect 20165 20519 20223 20525
rect 20165 20516 20177 20519
rect 19444 20488 20177 20516
rect 11940 20476 11946 20488
rect 10965 20451 11023 20457
rect 10965 20417 10977 20451
rect 11011 20417 11023 20451
rect 10965 20411 11023 20417
rect 11238 20408 11244 20460
rect 11296 20408 11302 20460
rect 12710 20448 12716 20460
rect 11808 20420 12716 20448
rect 7101 20383 7159 20389
rect 7101 20349 7113 20383
rect 7147 20349 7159 20383
rect 7101 20343 7159 20349
rect 8941 20383 8999 20389
rect 8941 20349 8953 20383
rect 8987 20380 8999 20383
rect 10502 20380 10508 20392
rect 8987 20352 10508 20380
rect 8987 20349 8999 20352
rect 8941 20343 8999 20349
rect 7116 20244 7144 20343
rect 10502 20340 10508 20352
rect 10560 20340 10566 20392
rect 11149 20383 11207 20389
rect 11149 20349 11161 20383
rect 11195 20380 11207 20383
rect 11698 20380 11704 20392
rect 11195 20352 11704 20380
rect 11195 20349 11207 20352
rect 11149 20343 11207 20349
rect 11698 20340 11704 20352
rect 11756 20340 11762 20392
rect 11808 20312 11836 20420
rect 12710 20408 12716 20420
rect 12768 20408 12774 20460
rect 12989 20451 13047 20457
rect 12989 20417 13001 20451
rect 13035 20448 13047 20451
rect 13354 20448 13360 20460
rect 13035 20420 13360 20448
rect 13035 20417 13047 20420
rect 12989 20411 13047 20417
rect 13354 20408 13360 20420
rect 13412 20408 13418 20460
rect 14366 20408 14372 20460
rect 14424 20408 14430 20460
rect 14721 20448 14749 20488
rect 20165 20485 20177 20488
rect 20211 20485 20223 20519
rect 20165 20479 20223 20485
rect 21818 20476 21824 20528
rect 21876 20516 21882 20528
rect 22189 20519 22247 20525
rect 22189 20516 22201 20519
rect 21876 20488 22201 20516
rect 21876 20476 21882 20488
rect 22189 20485 22201 20488
rect 22235 20485 22247 20519
rect 25133 20519 25191 20525
rect 22189 20479 22247 20485
rect 23032 20488 25084 20516
rect 14660 20420 14749 20448
rect 14660 20389 14688 20420
rect 15470 20408 15476 20460
rect 15528 20408 15534 20460
rect 17402 20408 17408 20460
rect 17460 20408 17466 20460
rect 17497 20451 17555 20457
rect 17497 20417 17509 20451
rect 17543 20417 17555 20451
rect 17497 20411 17555 20417
rect 14645 20383 14703 20389
rect 14645 20349 14657 20383
rect 14691 20349 14703 20383
rect 14645 20343 14703 20349
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 17420 20380 17448 20408
rect 14792 20352 17448 20380
rect 14792 20340 14798 20352
rect 8036 20284 11836 20312
rect 8036 20244 8064 20284
rect 17126 20272 17132 20324
rect 17184 20312 17190 20324
rect 17512 20312 17540 20411
rect 17770 20408 17776 20460
rect 17828 20408 17834 20460
rect 18230 20408 18236 20460
rect 18288 20408 18294 20460
rect 19337 20451 19395 20457
rect 19337 20448 19349 20451
rect 18524 20420 19349 20448
rect 18524 20389 18552 20420
rect 19337 20417 19349 20420
rect 19383 20448 19395 20451
rect 19610 20448 19616 20460
rect 19383 20420 19616 20448
rect 19383 20417 19395 20420
rect 19337 20411 19395 20417
rect 19610 20408 19616 20420
rect 19668 20448 19674 20460
rect 23032 20448 23060 20488
rect 19668 20420 23060 20448
rect 23109 20451 23167 20457
rect 19668 20408 19674 20420
rect 23109 20417 23121 20451
rect 23155 20448 23167 20451
rect 23566 20448 23572 20460
rect 23155 20420 23572 20448
rect 23155 20417 23167 20420
rect 23109 20411 23167 20417
rect 18509 20383 18567 20389
rect 18509 20349 18521 20383
rect 18555 20349 18567 20383
rect 18509 20343 18567 20349
rect 18598 20340 18604 20392
rect 18656 20380 18662 20392
rect 18656 20352 21956 20380
rect 18656 20340 18662 20352
rect 17184 20284 17540 20312
rect 20533 20315 20591 20321
rect 17184 20272 17190 20284
rect 20533 20281 20545 20315
rect 20579 20312 20591 20315
rect 21174 20312 21180 20324
rect 20579 20284 21180 20312
rect 20579 20281 20591 20284
rect 20533 20275 20591 20281
rect 21174 20272 21180 20284
rect 21232 20272 21238 20324
rect 7116 20216 8064 20244
rect 8294 20204 8300 20256
rect 8352 20204 8358 20256
rect 9493 20247 9551 20253
rect 9493 20213 9505 20247
rect 9539 20244 9551 20247
rect 9674 20244 9680 20256
rect 9539 20216 9680 20244
rect 9539 20213 9551 20216
rect 9493 20207 9551 20213
rect 9674 20204 9680 20216
rect 9732 20244 9738 20256
rect 10410 20244 10416 20256
rect 9732 20216 10416 20244
rect 9732 20204 9738 20216
rect 10410 20204 10416 20216
rect 10468 20204 10474 20256
rect 10689 20247 10747 20253
rect 10689 20213 10701 20247
rect 10735 20244 10747 20247
rect 10778 20244 10784 20256
rect 10735 20216 10784 20244
rect 10735 20213 10747 20216
rect 10689 20207 10747 20213
rect 10778 20204 10784 20216
rect 10836 20204 10842 20256
rect 13722 20204 13728 20256
rect 13780 20204 13786 20256
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 14001 20247 14059 20253
rect 14001 20244 14013 20247
rect 13872 20216 14013 20244
rect 13872 20204 13878 20216
rect 14001 20213 14013 20216
rect 14047 20213 14059 20247
rect 14001 20207 14059 20213
rect 17221 20247 17279 20253
rect 17221 20213 17233 20247
rect 17267 20244 17279 20247
rect 17494 20244 17500 20256
rect 17267 20216 17500 20244
rect 17267 20213 17279 20216
rect 17221 20207 17279 20213
rect 17494 20204 17500 20216
rect 17552 20204 17558 20256
rect 17586 20204 17592 20256
rect 17644 20244 17650 20256
rect 17681 20247 17739 20253
rect 17681 20244 17693 20247
rect 17644 20216 17693 20244
rect 17644 20204 17650 20216
rect 17681 20213 17693 20216
rect 17727 20213 17739 20247
rect 17681 20207 17739 20213
rect 17862 20204 17868 20256
rect 17920 20204 17926 20256
rect 21358 20204 21364 20256
rect 21416 20244 21422 20256
rect 21821 20247 21879 20253
rect 21821 20244 21833 20247
rect 21416 20216 21833 20244
rect 21416 20204 21422 20216
rect 21821 20213 21833 20216
rect 21867 20213 21879 20247
rect 21928 20244 21956 20352
rect 22278 20340 22284 20392
rect 22336 20380 22342 20392
rect 22373 20383 22431 20389
rect 22373 20380 22385 20383
rect 22336 20352 22385 20380
rect 22336 20340 22342 20352
rect 22373 20349 22385 20352
rect 22419 20380 22431 20383
rect 22922 20380 22928 20392
rect 22419 20352 22928 20380
rect 22419 20349 22431 20352
rect 22373 20343 22431 20349
rect 22922 20340 22928 20352
rect 22980 20340 22986 20392
rect 23124 20244 23152 20411
rect 23566 20408 23572 20420
rect 23624 20448 23630 20460
rect 24210 20448 24216 20460
rect 23624 20420 24216 20448
rect 23624 20408 23630 20420
rect 24210 20408 24216 20420
rect 24268 20408 24274 20460
rect 24302 20408 24308 20460
rect 24360 20408 24366 20460
rect 24397 20451 24455 20457
rect 24397 20417 24409 20451
rect 24443 20417 24455 20451
rect 24397 20411 24455 20417
rect 24673 20451 24731 20457
rect 24673 20417 24685 20451
rect 24719 20448 24731 20451
rect 24854 20448 24860 20460
rect 24719 20420 24860 20448
rect 24719 20417 24731 20420
rect 24673 20411 24731 20417
rect 24412 20380 24440 20411
rect 24854 20408 24860 20420
rect 24912 20408 24918 20460
rect 25056 20380 25084 20488
rect 25133 20485 25145 20519
rect 25179 20516 25191 20519
rect 26234 20516 26240 20528
rect 25179 20488 26240 20516
rect 25179 20485 25191 20488
rect 25133 20479 25191 20485
rect 26234 20476 26240 20488
rect 26292 20476 26298 20528
rect 26326 20476 26332 20528
rect 26384 20476 26390 20528
rect 28445 20519 28503 20525
rect 28445 20485 28457 20519
rect 28491 20516 28503 20519
rect 29178 20516 29184 20528
rect 28491 20488 29184 20516
rect 28491 20485 28503 20488
rect 28445 20479 28503 20485
rect 29178 20476 29184 20488
rect 29236 20476 29242 20528
rect 30558 20476 30564 20528
rect 30616 20516 30622 20528
rect 30837 20519 30895 20525
rect 30837 20516 30849 20519
rect 30616 20488 30849 20516
rect 30616 20476 30622 20488
rect 30837 20485 30849 20488
rect 30883 20485 30895 20519
rect 30837 20479 30895 20485
rect 31481 20519 31539 20525
rect 31481 20485 31493 20519
rect 31527 20516 31539 20519
rect 32370 20519 32428 20525
rect 32370 20516 32382 20519
rect 31527 20488 32382 20516
rect 31527 20485 31539 20488
rect 31481 20479 31539 20485
rect 32370 20485 32382 20488
rect 32416 20485 32428 20519
rect 32370 20479 32428 20485
rect 26145 20451 26203 20457
rect 26145 20417 26157 20451
rect 26191 20417 26203 20451
rect 26145 20411 26203 20417
rect 27617 20451 27675 20457
rect 27617 20417 27629 20451
rect 27663 20448 27675 20451
rect 28997 20451 29055 20457
rect 28997 20448 29009 20451
rect 27663 20420 29009 20448
rect 27663 20417 27675 20420
rect 27617 20411 27675 20417
rect 28997 20417 29009 20420
rect 29043 20448 29055 20451
rect 30466 20448 30472 20460
rect 29043 20420 30472 20448
rect 29043 20417 29055 20420
rect 28997 20411 29055 20417
rect 25317 20383 25375 20389
rect 25317 20380 25329 20383
rect 24412 20352 24808 20380
rect 25056 20352 25329 20380
rect 23290 20272 23296 20324
rect 23348 20272 23354 20324
rect 24780 20321 24808 20352
rect 25317 20349 25329 20352
rect 25363 20380 25375 20383
rect 26160 20380 26188 20411
rect 30466 20408 30472 20420
rect 30524 20408 30530 20460
rect 30926 20448 30932 20460
rect 30668 20420 30932 20448
rect 28629 20383 28687 20389
rect 28629 20380 28641 20383
rect 25363 20352 28641 20380
rect 25363 20349 25375 20352
rect 25317 20343 25375 20349
rect 28629 20349 28641 20352
rect 28675 20380 28687 20383
rect 29181 20383 29239 20389
rect 29181 20380 29193 20383
rect 28675 20352 29193 20380
rect 28675 20349 28687 20352
rect 28629 20343 28687 20349
rect 29181 20349 29193 20352
rect 29227 20349 29239 20383
rect 29181 20343 29239 20349
rect 30377 20383 30435 20389
rect 30377 20349 30389 20383
rect 30423 20380 30435 20383
rect 30668 20380 30696 20420
rect 30926 20408 30932 20420
rect 30984 20408 30990 20460
rect 31662 20408 31668 20460
rect 31720 20408 31726 20460
rect 31846 20408 31852 20460
rect 31904 20408 31910 20460
rect 31941 20451 31999 20457
rect 31941 20417 31953 20451
rect 31987 20448 31999 20451
rect 32030 20448 32036 20460
rect 31987 20420 32036 20448
rect 31987 20417 31999 20420
rect 31941 20411 31999 20417
rect 32030 20408 32036 20420
rect 32088 20408 32094 20460
rect 32125 20451 32183 20457
rect 32125 20417 32137 20451
rect 32171 20448 32183 20451
rect 33134 20448 33140 20460
rect 32171 20420 33140 20448
rect 32171 20417 32183 20420
rect 32125 20411 32183 20417
rect 33134 20408 33140 20420
rect 33192 20408 33198 20460
rect 30423 20352 30696 20380
rect 30423 20349 30435 20352
rect 30377 20343 30435 20349
rect 30742 20340 30748 20392
rect 30800 20340 30806 20392
rect 24765 20315 24823 20321
rect 24765 20281 24777 20315
rect 24811 20281 24823 20315
rect 30760 20312 30788 20340
rect 32122 20312 32128 20324
rect 30760 20284 32128 20312
rect 24765 20275 24823 20281
rect 32122 20272 32128 20284
rect 32180 20272 32186 20324
rect 21928 20216 23152 20244
rect 21821 20207 21879 20213
rect 24118 20204 24124 20256
rect 24176 20204 24182 20256
rect 24581 20247 24639 20253
rect 24581 20213 24593 20247
rect 24627 20244 24639 20247
rect 25222 20244 25228 20256
rect 24627 20216 25228 20244
rect 24627 20213 24639 20216
rect 24581 20207 24639 20213
rect 25222 20204 25228 20216
rect 25280 20204 25286 20256
rect 30650 20204 30656 20256
rect 30708 20244 30714 20256
rect 31021 20247 31079 20253
rect 31021 20244 31033 20247
rect 30708 20216 31033 20244
rect 30708 20204 30714 20216
rect 31021 20213 31033 20216
rect 31067 20213 31079 20247
rect 31021 20207 31079 20213
rect 31846 20204 31852 20256
rect 31904 20244 31910 20256
rect 34790 20244 34796 20256
rect 31904 20216 34796 20244
rect 31904 20204 31910 20216
rect 34790 20204 34796 20216
rect 34848 20204 34854 20256
rect 1104 20154 36800 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 36800 20154
rect 1104 20080 36800 20102
rect 1762 20000 1768 20052
rect 1820 20040 1826 20052
rect 1857 20043 1915 20049
rect 1857 20040 1869 20043
rect 1820 20012 1869 20040
rect 1820 20000 1826 20012
rect 1857 20009 1869 20012
rect 1903 20009 1915 20043
rect 1857 20003 1915 20009
rect 6825 20043 6883 20049
rect 6825 20009 6837 20043
rect 6871 20040 6883 20043
rect 7190 20040 7196 20052
rect 6871 20012 7196 20040
rect 6871 20009 6883 20012
rect 6825 20003 6883 20009
rect 7190 20000 7196 20012
rect 7248 20000 7254 20052
rect 8478 20000 8484 20052
rect 8536 20000 8542 20052
rect 10870 20000 10876 20052
rect 10928 20040 10934 20052
rect 10965 20043 11023 20049
rect 10965 20040 10977 20043
rect 10928 20012 10977 20040
rect 10928 20000 10934 20012
rect 10965 20009 10977 20012
rect 11011 20009 11023 20043
rect 10965 20003 11023 20009
rect 13354 20000 13360 20052
rect 13412 20000 13418 20052
rect 13817 20043 13875 20049
rect 13817 20009 13829 20043
rect 13863 20040 13875 20043
rect 13906 20040 13912 20052
rect 13863 20012 13912 20040
rect 13863 20009 13875 20012
rect 13817 20003 13875 20009
rect 13906 20000 13912 20012
rect 13964 20000 13970 20052
rect 15028 20012 23520 20040
rect 6638 19932 6644 19984
rect 6696 19932 6702 19984
rect 7374 19932 7380 19984
rect 7432 19972 7438 19984
rect 10781 19975 10839 19981
rect 7432 19944 10548 19972
rect 7432 19932 7438 19944
rect 1578 19864 1584 19916
rect 1636 19904 1642 19916
rect 10520 19913 10548 19944
rect 10781 19941 10793 19975
rect 10827 19972 10839 19975
rect 11238 19972 11244 19984
rect 10827 19944 11244 19972
rect 10827 19941 10839 19944
rect 10781 19935 10839 19941
rect 11238 19932 11244 19944
rect 11296 19932 11302 19984
rect 10505 19907 10563 19913
rect 1636 19876 9812 19904
rect 1636 19864 1642 19876
rect 2038 19796 2044 19848
rect 2096 19796 2102 19848
rect 6365 19839 6423 19845
rect 6365 19805 6377 19839
rect 6411 19836 6423 19839
rect 7374 19836 7380 19848
rect 6411 19808 7380 19836
rect 6411 19805 6423 19808
rect 6365 19799 6423 19805
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 8205 19839 8263 19845
rect 8205 19805 8217 19839
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 8220 19768 8248 19799
rect 8294 19796 8300 19848
rect 8352 19796 8358 19848
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 9582 19836 9588 19848
rect 8619 19808 9588 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 9582 19796 9588 19808
rect 9640 19796 9646 19848
rect 9674 19768 9680 19780
rect 8220 19740 9680 19768
rect 9674 19728 9680 19740
rect 9732 19728 9738 19780
rect 4338 19660 4344 19712
rect 4396 19700 4402 19712
rect 4614 19700 4620 19712
rect 4396 19672 4620 19700
rect 4396 19660 4402 19672
rect 4614 19660 4620 19672
rect 4672 19700 4678 19712
rect 5902 19700 5908 19712
rect 4672 19672 5908 19700
rect 4672 19660 4678 19672
rect 5902 19660 5908 19672
rect 5960 19660 5966 19712
rect 8021 19703 8079 19709
rect 8021 19669 8033 19703
rect 8067 19700 8079 19703
rect 8110 19700 8116 19712
rect 8067 19672 8116 19700
rect 8067 19669 8079 19672
rect 8021 19663 8079 19669
rect 8110 19660 8116 19672
rect 8168 19660 8174 19712
rect 9784 19700 9812 19876
rect 10505 19873 10517 19907
rect 10551 19904 10563 19907
rect 13446 19904 13452 19916
rect 10551 19876 13452 19904
rect 10551 19873 10563 19876
rect 10505 19867 10563 19873
rect 13446 19864 13452 19876
rect 13504 19864 13510 19916
rect 14734 19904 14740 19916
rect 13556 19876 14740 19904
rect 10410 19796 10416 19848
rect 10468 19836 10474 19848
rect 13556 19845 13584 19876
rect 14734 19864 14740 19876
rect 14792 19864 14798 19916
rect 15028 19913 15056 20012
rect 16945 19975 17003 19981
rect 16945 19972 16957 19975
rect 16592 19944 16957 19972
rect 15013 19907 15071 19913
rect 15013 19873 15025 19907
rect 15059 19873 15071 19907
rect 15013 19867 15071 19873
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 16592 19913 16620 19944
rect 16945 19941 16957 19944
rect 16991 19941 17003 19975
rect 23492 19972 23520 20012
rect 23566 20000 23572 20052
rect 23624 20000 23630 20052
rect 32677 20043 32735 20049
rect 32677 20009 32689 20043
rect 32723 20040 32735 20043
rect 33318 20040 33324 20052
rect 32723 20012 33324 20040
rect 32723 20009 32735 20012
rect 32677 20003 32735 20009
rect 33318 20000 33324 20012
rect 33376 20000 33382 20052
rect 30834 19972 30840 19984
rect 23492 19944 30840 19972
rect 16945 19935 17003 19941
rect 30834 19932 30840 19944
rect 30892 19972 30898 19984
rect 30892 19944 34376 19972
rect 30892 19932 30898 19944
rect 16577 19907 16635 19913
rect 16577 19904 16589 19907
rect 15252 19876 16589 19904
rect 15252 19864 15258 19876
rect 16577 19873 16589 19876
rect 16623 19873 16635 19907
rect 20990 19904 20996 19916
rect 16577 19867 16635 19873
rect 16776 19876 20996 19904
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 10468 19808 13553 19836
rect 10468 19796 10474 19808
rect 13541 19805 13553 19808
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 13633 19839 13691 19845
rect 13633 19805 13645 19839
rect 13679 19836 13691 19839
rect 13814 19836 13820 19848
rect 13679 19808 13820 19836
rect 13679 19805 13691 19808
rect 13633 19799 13691 19805
rect 13814 19796 13820 19808
rect 13872 19796 13878 19848
rect 13909 19839 13967 19845
rect 13909 19805 13921 19839
rect 13955 19836 13967 19839
rect 14826 19836 14832 19848
rect 13955 19808 14832 19836
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 15102 19796 15108 19848
rect 15160 19836 15166 19848
rect 15289 19839 15347 19845
rect 15289 19836 15301 19839
rect 15160 19808 15301 19836
rect 15160 19796 15166 19808
rect 15289 19805 15301 19808
rect 15335 19805 15347 19839
rect 15289 19799 15347 19805
rect 16114 19796 16120 19848
rect 16172 19836 16178 19848
rect 16776 19845 16804 19876
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 21453 19907 21511 19913
rect 21453 19904 21465 19907
rect 21284 19876 21465 19904
rect 21284 19848 21312 19876
rect 21453 19873 21465 19876
rect 21499 19873 21511 19907
rect 23658 19904 23664 19916
rect 21453 19867 21511 19873
rect 22940 19876 23664 19904
rect 16393 19839 16451 19845
rect 16393 19836 16405 19839
rect 16172 19808 16405 19836
rect 16172 19796 16178 19808
rect 16393 19805 16405 19808
rect 16439 19805 16451 19839
rect 16393 19799 16451 19805
rect 16761 19839 16819 19845
rect 16761 19805 16773 19839
rect 16807 19805 16819 19839
rect 16761 19799 16819 19805
rect 21266 19796 21272 19848
rect 21324 19796 21330 19848
rect 22940 19845 22968 19876
rect 23658 19864 23664 19876
rect 23716 19864 23722 19916
rect 30926 19864 30932 19916
rect 30984 19904 30990 19916
rect 31662 19904 31668 19916
rect 30984 19876 31668 19904
rect 30984 19864 30990 19876
rect 31662 19864 31668 19876
rect 31720 19904 31726 19916
rect 32674 19904 32680 19916
rect 31720 19876 32680 19904
rect 31720 19864 31726 19876
rect 32674 19864 32680 19876
rect 32732 19904 32738 19916
rect 33229 19907 33287 19913
rect 33229 19904 33241 19907
rect 32732 19876 33241 19904
rect 32732 19864 32738 19876
rect 33229 19873 33241 19876
rect 33275 19873 33287 19907
rect 33229 19867 33287 19873
rect 21361 19844 21419 19845
rect 21358 19792 21364 19844
rect 21416 19832 21422 19844
rect 22925 19839 22983 19845
rect 21416 19804 21457 19832
rect 22925 19805 22937 19839
rect 22971 19805 22983 19839
rect 21416 19792 21422 19804
rect 22925 19799 22983 19805
rect 12434 19728 12440 19780
rect 12492 19768 12498 19780
rect 16022 19768 16028 19780
rect 12492 19740 16028 19768
rect 12492 19728 12498 19740
rect 16022 19728 16028 19740
rect 16080 19728 16086 19780
rect 19981 19771 20039 19777
rect 19981 19737 19993 19771
rect 20027 19768 20039 19771
rect 20990 19768 20996 19780
rect 20027 19740 20996 19768
rect 20027 19737 20039 19740
rect 19981 19731 20039 19737
rect 20990 19728 20996 19740
rect 21048 19728 21054 19780
rect 21542 19728 21548 19780
rect 21600 19768 21606 19780
rect 21698 19771 21756 19777
rect 21698 19768 21710 19771
rect 21600 19740 21710 19768
rect 21600 19728 21606 19740
rect 21698 19737 21710 19740
rect 21744 19737 21756 19771
rect 21698 19731 21756 19737
rect 22002 19728 22008 19780
rect 22060 19768 22066 19780
rect 22940 19768 22968 19799
rect 23382 19796 23388 19848
rect 23440 19796 23446 19848
rect 27985 19839 28043 19845
rect 27985 19805 27997 19839
rect 28031 19836 28043 19839
rect 28626 19836 28632 19848
rect 28031 19808 28632 19836
rect 28031 19805 28043 19808
rect 27985 19799 28043 19805
rect 28626 19796 28632 19808
rect 28684 19796 28690 19848
rect 29914 19796 29920 19848
rect 29972 19796 29978 19848
rect 33042 19796 33048 19848
rect 33100 19796 33106 19848
rect 34348 19845 34376 19944
rect 34333 19839 34391 19845
rect 34333 19805 34345 19839
rect 34379 19805 34391 19839
rect 34333 19799 34391 19805
rect 22060 19740 22968 19768
rect 34517 19771 34575 19777
rect 22060 19728 22066 19740
rect 34517 19737 34529 19771
rect 34563 19768 34575 19771
rect 34698 19768 34704 19780
rect 34563 19740 34704 19768
rect 34563 19737 34575 19740
rect 34517 19731 34575 19737
rect 34698 19728 34704 19740
rect 34756 19768 34762 19780
rect 34793 19771 34851 19777
rect 34793 19768 34805 19771
rect 34756 19740 34805 19768
rect 34756 19728 34762 19740
rect 34793 19737 34805 19740
rect 34839 19737 34851 19771
rect 34793 19731 34851 19737
rect 13722 19700 13728 19712
rect 9784 19672 13728 19700
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 15378 19660 15384 19712
rect 15436 19700 15442 19712
rect 15933 19703 15991 19709
rect 15933 19700 15945 19703
rect 15436 19672 15945 19700
rect 15436 19660 15442 19672
rect 15933 19669 15945 19672
rect 15979 19669 15991 19703
rect 15933 19663 15991 19669
rect 16298 19660 16304 19712
rect 16356 19660 16362 19712
rect 20070 19660 20076 19712
rect 20128 19660 20134 19712
rect 21177 19703 21235 19709
rect 21177 19669 21189 19703
rect 21223 19700 21235 19703
rect 21266 19700 21272 19712
rect 21223 19672 21272 19700
rect 21223 19669 21235 19672
rect 21177 19663 21235 19669
rect 21266 19660 21272 19672
rect 21324 19660 21330 19712
rect 21818 19660 21824 19712
rect 21876 19700 21882 19712
rect 22833 19703 22891 19709
rect 22833 19700 22845 19703
rect 21876 19672 22845 19700
rect 21876 19660 21882 19672
rect 22833 19669 22845 19672
rect 22879 19669 22891 19703
rect 22833 19663 22891 19669
rect 23106 19660 23112 19712
rect 23164 19660 23170 19712
rect 26326 19660 26332 19712
rect 26384 19700 26390 19712
rect 28169 19703 28227 19709
rect 28169 19700 28181 19703
rect 26384 19672 28181 19700
rect 26384 19660 26390 19672
rect 28169 19669 28181 19672
rect 28215 19669 28227 19703
rect 28169 19663 28227 19669
rect 29730 19660 29736 19712
rect 29788 19660 29794 19712
rect 33134 19660 33140 19712
rect 33192 19660 33198 19712
rect 34606 19660 34612 19712
rect 34664 19700 34670 19712
rect 34885 19703 34943 19709
rect 34885 19700 34897 19703
rect 34664 19672 34897 19700
rect 34664 19660 34670 19672
rect 34885 19669 34897 19672
rect 34931 19669 34943 19703
rect 34885 19663 34943 19669
rect 1104 19610 36800 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 36800 19610
rect 1104 19536 36800 19558
rect 12434 19496 12440 19508
rect 2746 19468 12440 19496
rect 1489 19431 1547 19437
rect 1489 19397 1501 19431
rect 1535 19428 1547 19431
rect 2746 19428 2774 19468
rect 12434 19456 12440 19468
rect 12492 19456 12498 19508
rect 12529 19499 12587 19505
rect 12529 19465 12541 19499
rect 12575 19496 12587 19499
rect 13078 19496 13084 19508
rect 12575 19468 13084 19496
rect 12575 19465 12587 19468
rect 12529 19459 12587 19465
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 14366 19456 14372 19508
rect 14424 19496 14430 19508
rect 14737 19499 14795 19505
rect 14737 19496 14749 19499
rect 14424 19468 14749 19496
rect 14424 19456 14430 19468
rect 14737 19465 14749 19468
rect 14783 19465 14795 19499
rect 14737 19459 14795 19465
rect 16022 19456 16028 19508
rect 16080 19496 16086 19508
rect 16206 19496 16212 19508
rect 16080 19468 16212 19496
rect 16080 19456 16086 19468
rect 16206 19456 16212 19468
rect 16264 19496 16270 19508
rect 19245 19499 19303 19505
rect 19245 19496 19257 19499
rect 16264 19468 19257 19496
rect 16264 19456 16270 19468
rect 19245 19465 19257 19468
rect 19291 19465 19303 19499
rect 19245 19459 19303 19465
rect 21266 19456 21272 19508
rect 21324 19496 21330 19508
rect 21542 19496 21548 19508
rect 21324 19468 21548 19496
rect 21324 19456 21330 19468
rect 21542 19456 21548 19468
rect 21600 19456 21606 19508
rect 22002 19456 22008 19508
rect 22060 19456 22066 19508
rect 25038 19456 25044 19508
rect 25096 19496 25102 19508
rect 25317 19499 25375 19505
rect 25317 19496 25329 19499
rect 25096 19468 25329 19496
rect 25096 19456 25102 19468
rect 25317 19465 25329 19468
rect 25363 19465 25375 19499
rect 25317 19459 25375 19465
rect 26050 19456 26056 19508
rect 26108 19456 26114 19508
rect 35434 19456 35440 19508
rect 35492 19496 35498 19508
rect 35529 19499 35587 19505
rect 35529 19496 35541 19499
rect 35492 19468 35541 19496
rect 35492 19456 35498 19468
rect 35529 19465 35541 19468
rect 35575 19465 35587 19499
rect 35529 19459 35587 19465
rect 1535 19400 2774 19428
rect 1535 19397 1547 19400
rect 1489 19391 1547 19397
rect 2958 19388 2964 19440
rect 3016 19428 3022 19440
rect 4157 19431 4215 19437
rect 4157 19428 4169 19431
rect 3016 19400 4169 19428
rect 3016 19388 3022 19400
rect 4157 19397 4169 19400
rect 4203 19397 4215 19431
rect 4157 19391 4215 19397
rect 4264 19400 4660 19428
rect 2409 19363 2467 19369
rect 2409 19329 2421 19363
rect 2455 19360 2467 19363
rect 2455 19332 2544 19360
rect 2455 19329 2467 19332
rect 2409 19323 2467 19329
rect 2516 19233 2544 19332
rect 2866 19320 2872 19372
rect 2924 19320 2930 19372
rect 3602 19320 3608 19372
rect 3660 19360 3666 19372
rect 3973 19363 4031 19369
rect 3973 19360 3985 19363
rect 3660 19332 3985 19360
rect 3660 19320 3666 19332
rect 3973 19329 3985 19332
rect 4019 19360 4031 19363
rect 4264 19360 4292 19400
rect 4632 19372 4660 19400
rect 14826 19388 14832 19440
rect 14884 19428 14890 19440
rect 20806 19428 20812 19440
rect 14884 19400 16988 19428
rect 14884 19388 14890 19400
rect 4019 19332 4292 19360
rect 4019 19329 4031 19332
rect 3973 19323 4031 19329
rect 4338 19320 4344 19372
rect 4396 19320 4402 19372
rect 4614 19320 4620 19372
rect 4672 19360 4678 19372
rect 8294 19369 8300 19372
rect 4709 19363 4767 19369
rect 4709 19360 4721 19363
rect 4672 19332 4721 19360
rect 4672 19320 4678 19332
rect 4709 19329 4721 19332
rect 4755 19329 4767 19363
rect 8288 19360 8300 19369
rect 8255 19332 8300 19360
rect 4709 19323 4767 19329
rect 8288 19323 8300 19332
rect 8294 19320 8300 19323
rect 8352 19320 8358 19372
rect 12437 19363 12495 19369
rect 12437 19329 12449 19363
rect 12483 19360 12495 19363
rect 12894 19360 12900 19372
rect 12483 19332 12900 19360
rect 12483 19329 12495 19332
rect 12437 19323 12495 19329
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 16960 19369 16988 19400
rect 19996 19400 20812 19428
rect 15289 19363 15347 19369
rect 15289 19329 15301 19363
rect 15335 19360 15347 19363
rect 16945 19363 17003 19369
rect 15335 19332 16712 19360
rect 15335 19329 15347 19332
rect 15289 19323 15347 19329
rect 2958 19252 2964 19304
rect 3016 19292 3022 19304
rect 3145 19295 3203 19301
rect 3145 19292 3157 19295
rect 3016 19264 3157 19292
rect 3016 19252 3022 19264
rect 3145 19261 3157 19264
rect 3191 19292 3203 19295
rect 3191 19264 7328 19292
rect 3191 19261 3203 19264
rect 3145 19255 3203 19261
rect 2501 19227 2559 19233
rect 2501 19193 2513 19227
rect 2547 19193 2559 19227
rect 4525 19227 4583 19233
rect 4525 19224 4537 19227
rect 2501 19187 2559 19193
rect 3620 19196 4537 19224
rect 934 19116 940 19168
rect 992 19156 998 19168
rect 1581 19159 1639 19165
rect 1581 19156 1593 19159
rect 992 19128 1593 19156
rect 992 19116 998 19128
rect 1581 19125 1593 19128
rect 1627 19125 1639 19159
rect 1581 19119 1639 19125
rect 2130 19116 2136 19168
rect 2188 19156 2194 19168
rect 2225 19159 2283 19165
rect 2225 19156 2237 19159
rect 2188 19128 2237 19156
rect 2188 19116 2194 19128
rect 2225 19125 2237 19128
rect 2271 19125 2283 19159
rect 2225 19119 2283 19125
rect 2682 19116 2688 19168
rect 2740 19156 2746 19168
rect 3620 19156 3648 19196
rect 4525 19193 4537 19196
rect 4571 19193 4583 19227
rect 4525 19187 4583 19193
rect 2740 19128 3648 19156
rect 2740 19116 2746 19128
rect 4706 19116 4712 19168
rect 4764 19156 4770 19168
rect 4801 19159 4859 19165
rect 4801 19156 4813 19159
rect 4764 19128 4813 19156
rect 4764 19116 4770 19128
rect 4801 19125 4813 19128
rect 4847 19125 4859 19159
rect 7300 19156 7328 19264
rect 8018 19252 8024 19304
rect 8076 19252 8082 19304
rect 9214 19252 9220 19304
rect 9272 19292 9278 19304
rect 12713 19295 12771 19301
rect 12713 19292 12725 19295
rect 9272 19264 12725 19292
rect 9272 19252 9278 19264
rect 12713 19261 12725 19264
rect 12759 19292 12771 19295
rect 12759 19264 13032 19292
rect 12759 19261 12771 19264
rect 12713 19255 12771 19261
rect 9030 19184 9036 19236
rect 9088 19224 9094 19236
rect 12618 19224 12624 19236
rect 9088 19196 12624 19224
rect 9088 19184 9094 19196
rect 12618 19184 12624 19196
rect 12676 19184 12682 19236
rect 9214 19156 9220 19168
rect 7300 19128 9220 19156
rect 4801 19119 4859 19125
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 9398 19116 9404 19168
rect 9456 19116 9462 19168
rect 9858 19116 9864 19168
rect 9916 19156 9922 19168
rect 10594 19156 10600 19168
rect 9916 19128 10600 19156
rect 9916 19116 9922 19128
rect 10594 19116 10600 19128
rect 10652 19156 10658 19168
rect 11974 19156 11980 19168
rect 10652 19128 11980 19156
rect 10652 19116 10658 19128
rect 11974 19116 11980 19128
rect 12032 19116 12038 19168
rect 12066 19116 12072 19168
rect 12124 19116 12130 19168
rect 13004 19156 13032 19264
rect 13078 19252 13084 19304
rect 13136 19252 13142 19304
rect 13446 19252 13452 19304
rect 13504 19292 13510 19304
rect 13541 19295 13599 19301
rect 13541 19292 13553 19295
rect 13504 19264 13553 19292
rect 13504 19252 13510 19264
rect 13541 19261 13553 19264
rect 13587 19261 13599 19295
rect 13541 19255 13599 19261
rect 13814 19252 13820 19304
rect 13872 19252 13878 19304
rect 13906 19252 13912 19304
rect 13964 19301 13970 19304
rect 13964 19295 13992 19301
rect 13980 19261 13992 19295
rect 13964 19255 13992 19261
rect 14093 19295 14151 19301
rect 14093 19261 14105 19295
rect 14139 19292 14151 19295
rect 14274 19292 14280 19304
rect 14139 19264 14280 19292
rect 14139 19261 14151 19264
rect 14093 19255 14151 19261
rect 13964 19252 13970 19255
rect 14274 19252 14280 19264
rect 14332 19252 14338 19304
rect 14642 19252 14648 19304
rect 14700 19292 14706 19304
rect 15013 19295 15071 19301
rect 15013 19292 15025 19295
rect 14700 19264 15025 19292
rect 14700 19252 14706 19264
rect 15013 19261 15025 19264
rect 15059 19292 15071 19295
rect 15102 19292 15108 19304
rect 15059 19264 15108 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 16684 19301 16712 19332
rect 16945 19329 16957 19363
rect 16991 19329 17003 19363
rect 16945 19323 17003 19329
rect 18138 19320 18144 19372
rect 18196 19360 18202 19372
rect 18233 19363 18291 19369
rect 18233 19360 18245 19363
rect 18196 19332 18245 19360
rect 18196 19320 18202 19332
rect 18233 19329 18245 19332
rect 18279 19329 18291 19363
rect 18233 19323 18291 19329
rect 18509 19363 18567 19369
rect 18509 19329 18521 19363
rect 18555 19360 18567 19363
rect 19886 19360 19892 19372
rect 18555 19332 19892 19360
rect 18555 19329 18567 19332
rect 18509 19323 18567 19329
rect 19886 19320 19892 19332
rect 19944 19320 19950 19372
rect 19996 19369 20024 19400
rect 20806 19388 20812 19400
rect 20864 19388 20870 19440
rect 20990 19388 20996 19440
rect 21048 19428 21054 19440
rect 24762 19428 24768 19440
rect 21048 19400 21956 19428
rect 21048 19388 21054 19400
rect 19981 19363 20039 19369
rect 19981 19329 19993 19363
rect 20027 19329 20039 19363
rect 19981 19323 20039 19329
rect 20070 19320 20076 19372
rect 20128 19360 20134 19372
rect 20128 19332 20944 19360
rect 20128 19320 20134 19332
rect 16669 19295 16727 19301
rect 16669 19261 16681 19295
rect 16715 19292 16727 19295
rect 16758 19292 16764 19304
rect 16715 19264 16764 19292
rect 16715 19261 16727 19264
rect 16669 19255 16727 19261
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 17034 19252 17040 19304
rect 17092 19292 17098 19304
rect 17402 19292 17408 19304
rect 17092 19264 17408 19292
rect 17092 19252 17098 19264
rect 17402 19252 17408 19264
rect 17460 19252 17466 19304
rect 20916 19292 20944 19332
rect 21542 19320 21548 19372
rect 21600 19360 21606 19372
rect 21821 19363 21879 19369
rect 21821 19360 21833 19363
rect 21600 19332 21833 19360
rect 21600 19320 21606 19332
rect 21821 19329 21833 19332
rect 21867 19329 21879 19363
rect 21928 19360 21956 19400
rect 23308 19400 24768 19428
rect 23308 19360 23336 19400
rect 24762 19388 24768 19400
rect 24820 19428 24826 19440
rect 26326 19428 26332 19440
rect 24820 19400 26332 19428
rect 24820 19388 24826 19400
rect 26326 19388 26332 19400
rect 26384 19388 26390 19440
rect 29730 19437 29736 19440
rect 29724 19428 29736 19437
rect 29691 19400 29736 19428
rect 29724 19391 29736 19400
rect 29730 19388 29736 19391
rect 29788 19388 29794 19440
rect 33229 19431 33287 19437
rect 33229 19397 33241 19431
rect 33275 19428 33287 19431
rect 34606 19428 34612 19440
rect 33275 19400 34612 19428
rect 33275 19397 33287 19400
rect 33229 19391 33287 19397
rect 34606 19388 34612 19400
rect 34664 19388 34670 19440
rect 21928 19332 23336 19360
rect 21821 19323 21879 19329
rect 23382 19320 23388 19372
rect 23440 19320 23446 19372
rect 24854 19320 24860 19372
rect 24912 19360 24918 19372
rect 25406 19360 25412 19372
rect 24912 19332 25412 19360
rect 24912 19320 24918 19332
rect 25406 19320 25412 19332
rect 25464 19320 25470 19372
rect 25866 19320 25872 19372
rect 25924 19320 25930 19372
rect 26970 19320 26976 19372
rect 27028 19360 27034 19372
rect 27338 19360 27344 19372
rect 27028 19332 27344 19360
rect 27028 19320 27034 19332
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 29457 19363 29515 19369
rect 29457 19329 29469 19363
rect 29503 19360 29515 19363
rect 29546 19360 29552 19372
rect 29503 19332 29552 19360
rect 29503 19329 29515 19332
rect 29457 19323 29515 19329
rect 29546 19320 29552 19332
rect 29604 19360 29610 19372
rect 29604 19332 30512 19360
rect 29604 19320 29610 19332
rect 21726 19292 21732 19304
rect 20916 19264 21732 19292
rect 21726 19252 21732 19264
rect 21784 19252 21790 19304
rect 23290 19292 23296 19304
rect 21928 19264 23296 19292
rect 19334 19184 19340 19236
rect 19392 19224 19398 19236
rect 21818 19224 21824 19236
rect 19392 19196 21824 19224
rect 19392 19184 19398 19196
rect 21818 19184 21824 19196
rect 21876 19184 21882 19236
rect 15194 19156 15200 19168
rect 13004 19128 15200 19156
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 17586 19116 17592 19168
rect 17644 19156 17650 19168
rect 18046 19156 18052 19168
rect 17644 19128 18052 19156
rect 17644 19116 17650 19128
rect 18046 19116 18052 19128
rect 18104 19156 18110 19168
rect 20070 19156 20076 19168
rect 18104 19128 20076 19156
rect 18104 19116 18110 19128
rect 20070 19116 20076 19128
rect 20128 19116 20134 19168
rect 20162 19116 20168 19168
rect 20220 19116 20226 19168
rect 20254 19116 20260 19168
rect 20312 19156 20318 19168
rect 21928 19156 21956 19264
rect 23290 19252 23296 19264
rect 23348 19292 23354 19304
rect 25593 19295 25651 19301
rect 23348 19264 25452 19292
rect 23348 19252 23354 19264
rect 25424 19224 25452 19264
rect 25593 19261 25605 19295
rect 25639 19292 25651 19295
rect 25682 19292 25688 19304
rect 25639 19264 25688 19292
rect 25639 19261 25651 19264
rect 25593 19255 25651 19261
rect 25682 19252 25688 19264
rect 25740 19292 25746 19304
rect 27062 19292 27068 19304
rect 25740 19264 27068 19292
rect 25740 19252 25746 19264
rect 27062 19252 27068 19264
rect 27120 19252 27126 19304
rect 27157 19295 27215 19301
rect 27157 19261 27169 19295
rect 27203 19292 27215 19295
rect 27522 19292 27528 19304
rect 27203 19264 27528 19292
rect 27203 19261 27215 19264
rect 27157 19255 27215 19261
rect 27522 19252 27528 19264
rect 27580 19252 27586 19304
rect 28074 19301 28080 19304
rect 27893 19295 27951 19301
rect 27893 19292 27905 19295
rect 27724 19264 27905 19292
rect 27617 19227 27675 19233
rect 27617 19224 27629 19227
rect 22066 19196 25360 19224
rect 25424 19196 27629 19224
rect 22066 19168 22094 19196
rect 20312 19128 21956 19156
rect 20312 19116 20318 19128
rect 22002 19116 22008 19168
rect 22060 19128 22094 19168
rect 22060 19116 22066 19128
rect 23658 19116 23664 19168
rect 23716 19116 23722 19168
rect 24946 19116 24952 19168
rect 25004 19116 25010 19168
rect 25332 19156 25360 19196
rect 27617 19193 27629 19196
rect 27663 19193 27675 19227
rect 27617 19187 27675 19193
rect 25590 19156 25596 19168
rect 25332 19128 25596 19156
rect 25590 19116 25596 19128
rect 25648 19116 25654 19168
rect 26418 19116 26424 19168
rect 26476 19116 26482 19168
rect 27724 19156 27752 19264
rect 27893 19261 27905 19264
rect 27939 19261 27951 19295
rect 27893 19255 27951 19261
rect 28031 19295 28080 19301
rect 28031 19261 28043 19295
rect 28077 19261 28080 19295
rect 28031 19255 28080 19261
rect 28074 19252 28080 19255
rect 28132 19252 28138 19304
rect 28179 19295 28237 19301
rect 28179 19261 28191 19295
rect 28225 19292 28237 19295
rect 28534 19292 28540 19304
rect 28225 19264 28540 19292
rect 28225 19261 28237 19264
rect 28179 19255 28237 19261
rect 28534 19252 28540 19264
rect 28592 19252 28598 19304
rect 28810 19252 28816 19304
rect 28868 19252 28874 19304
rect 30484 19292 30512 19332
rect 34146 19320 34152 19372
rect 34204 19320 34210 19372
rect 34416 19363 34474 19369
rect 34416 19329 34428 19363
rect 34462 19360 34474 19363
rect 35342 19360 35348 19372
rect 34462 19332 35348 19360
rect 34462 19329 34474 19332
rect 34416 19323 34474 19329
rect 35342 19320 35348 19332
rect 35400 19320 35406 19372
rect 32398 19292 32404 19304
rect 30484 19264 32404 19292
rect 32398 19252 32404 19264
rect 32456 19292 32462 19304
rect 33413 19295 33471 19301
rect 33413 19292 33425 19295
rect 32456 19264 33425 19292
rect 32456 19252 32462 19264
rect 33413 19261 33425 19264
rect 33459 19261 33471 19295
rect 33413 19255 33471 19261
rect 28258 19156 28264 19168
rect 27724 19128 28264 19156
rect 28258 19116 28264 19128
rect 28316 19116 28322 19168
rect 28350 19116 28356 19168
rect 28408 19156 28414 19168
rect 30374 19156 30380 19168
rect 28408 19128 30380 19156
rect 28408 19116 28414 19128
rect 30374 19116 30380 19128
rect 30432 19116 30438 19168
rect 30834 19116 30840 19168
rect 30892 19116 30898 19168
rect 1104 19066 36800 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 36800 19066
rect 1104 18992 36800 19014
rect 2866 18912 2872 18964
rect 2924 18952 2930 18964
rect 3237 18955 3295 18961
rect 3237 18952 3249 18955
rect 2924 18924 3249 18952
rect 2924 18912 2930 18924
rect 3237 18921 3249 18924
rect 3283 18921 3295 18955
rect 5258 18952 5264 18964
rect 3237 18915 3295 18921
rect 5000 18924 5264 18952
rect 3252 18816 3280 18915
rect 4062 18816 4068 18828
rect 3252 18788 4068 18816
rect 4062 18776 4068 18788
rect 4120 18816 4126 18828
rect 5000 18825 5028 18924
rect 5258 18912 5264 18924
rect 5316 18952 5322 18964
rect 6181 18955 6239 18961
rect 5316 18924 5948 18952
rect 5316 18912 5322 18924
rect 5920 18884 5948 18924
rect 6181 18921 6193 18955
rect 6227 18952 6239 18955
rect 6638 18952 6644 18964
rect 6227 18924 6644 18952
rect 6227 18921 6239 18924
rect 6181 18915 6239 18921
rect 6638 18912 6644 18924
rect 6696 18912 6702 18964
rect 8018 18912 8024 18964
rect 8076 18952 8082 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 8076 18924 8125 18952
rect 8076 18912 8082 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8113 18915 8171 18921
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 8941 18955 8999 18961
rect 8941 18952 8953 18955
rect 8352 18924 8953 18952
rect 8352 18912 8358 18924
rect 8941 18921 8953 18924
rect 8987 18921 8999 18955
rect 8941 18915 8999 18921
rect 11238 18912 11244 18964
rect 11296 18912 11302 18964
rect 11348 18924 12848 18952
rect 5920 18856 10088 18884
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 4120 18788 4353 18816
rect 4120 18776 4126 18788
rect 4341 18785 4353 18788
rect 4387 18785 4399 18819
rect 4341 18779 4399 18785
rect 4985 18819 5043 18825
rect 4985 18785 4997 18819
rect 5031 18785 5043 18819
rect 4985 18779 5043 18785
rect 7558 18776 7564 18828
rect 7616 18816 7622 18828
rect 7926 18816 7932 18828
rect 7616 18788 7932 18816
rect 7616 18776 7622 18788
rect 7926 18776 7932 18788
rect 7984 18776 7990 18828
rect 9030 18776 9036 18828
rect 9088 18776 9094 18828
rect 9398 18776 9404 18828
rect 9456 18776 9462 18828
rect 9585 18819 9643 18825
rect 9585 18785 9597 18819
rect 9631 18816 9643 18819
rect 9674 18816 9680 18828
rect 9631 18788 9680 18816
rect 9631 18785 9643 18788
rect 9585 18779 9643 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 10060 18825 10088 18856
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18816 10103 18819
rect 11348 18816 11376 18924
rect 12820 18884 12848 18924
rect 12894 18912 12900 18964
rect 12952 18912 12958 18964
rect 16209 18955 16267 18961
rect 16209 18921 16221 18955
rect 16255 18952 16267 18955
rect 16298 18952 16304 18964
rect 16255 18924 16304 18952
rect 16255 18921 16267 18924
rect 16209 18915 16267 18921
rect 16298 18912 16304 18924
rect 16356 18952 16362 18964
rect 16356 18924 16436 18952
rect 16356 18912 16362 18924
rect 13170 18884 13176 18896
rect 12820 18856 13176 18884
rect 13170 18844 13176 18856
rect 13228 18844 13234 18896
rect 10091 18788 11376 18816
rect 10091 18785 10103 18788
rect 10045 18779 10103 18785
rect 14826 18776 14832 18828
rect 14884 18776 14890 18828
rect 16408 18825 16436 18924
rect 18230 18912 18236 18964
rect 18288 18912 18294 18964
rect 18800 18924 21404 18952
rect 16482 18844 16488 18896
rect 16540 18884 16546 18896
rect 16540 18856 17172 18884
rect 16540 18844 16546 18856
rect 16393 18819 16451 18825
rect 16393 18785 16405 18819
rect 16439 18785 16451 18819
rect 16393 18779 16451 18785
rect 17034 18776 17040 18828
rect 17092 18776 17098 18828
rect 17144 18816 17172 18856
rect 17144 18788 17356 18816
rect 1486 18708 1492 18760
rect 1544 18748 1550 18760
rect 2130 18757 2136 18760
rect 1857 18751 1915 18757
rect 1857 18748 1869 18751
rect 1544 18720 1869 18748
rect 1544 18708 1550 18720
rect 1857 18717 1869 18720
rect 1903 18717 1915 18751
rect 2124 18748 2136 18757
rect 2091 18720 2136 18748
rect 1857 18711 1915 18717
rect 2124 18711 2136 18720
rect 2130 18708 2136 18711
rect 2188 18708 2194 18760
rect 4522 18708 4528 18760
rect 4580 18708 4586 18760
rect 5258 18708 5264 18760
rect 5316 18708 5322 18760
rect 5442 18757 5448 18760
rect 5399 18751 5448 18757
rect 5399 18717 5411 18751
rect 5445 18717 5448 18751
rect 5399 18711 5448 18717
rect 5442 18708 5448 18711
rect 5500 18708 5506 18760
rect 5534 18708 5540 18760
rect 5592 18708 5598 18760
rect 6178 18708 6184 18760
rect 6236 18748 6242 18760
rect 9048 18748 9076 18776
rect 6236 18720 9076 18748
rect 6236 18708 6242 18720
rect 9122 18708 9128 18760
rect 9180 18708 9186 18760
rect 9214 18708 9220 18760
rect 9272 18708 9278 18760
rect 10318 18708 10324 18760
rect 10376 18708 10382 18760
rect 10502 18757 10508 18760
rect 10459 18751 10508 18757
rect 10459 18717 10471 18751
rect 10505 18717 10508 18751
rect 10459 18711 10508 18717
rect 10502 18708 10508 18711
rect 10560 18708 10566 18760
rect 10594 18708 10600 18760
rect 10652 18708 10658 18760
rect 11514 18708 11520 18760
rect 11572 18708 11578 18760
rect 13630 18748 13636 18760
rect 11624 18720 13636 18748
rect 7926 18640 7932 18692
rect 7984 18680 7990 18692
rect 8021 18683 8079 18689
rect 8021 18680 8033 18683
rect 7984 18652 8033 18680
rect 7984 18640 7990 18652
rect 8021 18649 8033 18652
rect 8067 18649 8079 18683
rect 8021 18643 8079 18649
rect 8941 18683 8999 18689
rect 8941 18649 8953 18683
rect 8987 18680 8999 18683
rect 9030 18680 9036 18692
rect 8987 18652 9036 18680
rect 8987 18649 8999 18652
rect 8941 18643 8999 18649
rect 9030 18640 9036 18652
rect 9088 18640 9094 18692
rect 5534 18572 5540 18624
rect 5592 18612 5598 18624
rect 5810 18612 5816 18624
rect 5592 18584 5816 18612
rect 5592 18572 5598 18584
rect 5810 18572 5816 18584
rect 5868 18612 5874 18624
rect 10594 18612 10600 18624
rect 5868 18584 10600 18612
rect 5868 18572 5874 18584
rect 10594 18572 10600 18584
rect 10652 18612 10658 18624
rect 11624 18612 11652 18720
rect 13630 18708 13636 18720
rect 13688 18708 13694 18760
rect 16574 18708 16580 18760
rect 16632 18708 16638 18760
rect 17328 18757 17356 18788
rect 17313 18751 17371 18757
rect 17313 18717 17325 18751
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17402 18708 17408 18760
rect 17460 18757 17466 18760
rect 17460 18751 17488 18757
rect 17476 18717 17488 18751
rect 17460 18711 17488 18717
rect 17460 18708 17466 18711
rect 17586 18708 17592 18760
rect 17644 18708 17650 18760
rect 11784 18683 11842 18689
rect 11784 18649 11796 18683
rect 11830 18680 11842 18683
rect 11882 18680 11888 18692
rect 11830 18652 11888 18680
rect 11830 18649 11842 18652
rect 11784 18643 11842 18649
rect 11882 18640 11888 18652
rect 11940 18640 11946 18692
rect 11974 18640 11980 18692
rect 12032 18680 12038 18692
rect 14274 18680 14280 18692
rect 12032 18652 14280 18680
rect 12032 18640 12038 18652
rect 14274 18640 14280 18652
rect 14332 18640 14338 18692
rect 15096 18683 15154 18689
rect 15096 18649 15108 18683
rect 15142 18680 15154 18683
rect 15194 18680 15200 18692
rect 15142 18652 15200 18680
rect 15142 18649 15154 18652
rect 15096 18643 15154 18649
rect 15194 18640 15200 18652
rect 15252 18640 15258 18692
rect 10652 18584 11652 18612
rect 10652 18572 10658 18584
rect 11698 18572 11704 18624
rect 11756 18612 11762 18624
rect 18800 18612 18828 18924
rect 18874 18844 18880 18896
rect 18932 18884 18938 18896
rect 20254 18884 20260 18896
rect 18932 18856 20260 18884
rect 18932 18844 18938 18856
rect 20254 18844 20260 18856
rect 20312 18844 20318 18896
rect 21376 18884 21404 18924
rect 21450 18912 21456 18964
rect 21508 18912 21514 18964
rect 22005 18955 22063 18961
rect 22005 18952 22017 18955
rect 21928 18924 22017 18952
rect 21928 18884 21956 18924
rect 22005 18921 22017 18924
rect 22051 18952 22063 18955
rect 24210 18952 24216 18964
rect 22051 18924 24216 18952
rect 22051 18921 22063 18924
rect 22005 18915 22063 18921
rect 24210 18912 24216 18924
rect 24268 18912 24274 18964
rect 26234 18912 26240 18964
rect 26292 18912 26298 18964
rect 27172 18924 28948 18952
rect 21376 18856 21956 18884
rect 23842 18844 23848 18896
rect 23900 18884 23906 18896
rect 27172 18893 27200 18924
rect 27157 18887 27215 18893
rect 23900 18856 25176 18884
rect 23900 18844 23906 18856
rect 20346 18776 20352 18828
rect 20404 18816 20410 18828
rect 20650 18819 20708 18825
rect 20650 18816 20662 18819
rect 20404 18788 20662 18816
rect 20404 18776 20410 18788
rect 20650 18785 20662 18788
rect 20696 18785 20708 18819
rect 20650 18779 20708 18785
rect 20806 18776 20812 18828
rect 20864 18816 20870 18828
rect 23106 18816 23112 18828
rect 20864 18788 23112 18816
rect 20864 18776 20870 18788
rect 23106 18776 23112 18788
rect 23164 18776 23170 18828
rect 25038 18776 25044 18828
rect 25096 18776 25102 18828
rect 25148 18816 25176 18856
rect 27157 18853 27169 18887
rect 27203 18853 27215 18887
rect 27157 18847 27215 18853
rect 25434 18819 25492 18825
rect 25434 18816 25446 18819
rect 25148 18788 25446 18816
rect 25434 18785 25446 18788
rect 25480 18785 25492 18819
rect 25434 18779 25492 18785
rect 25590 18776 25596 18828
rect 25648 18816 25654 18828
rect 27172 18816 27200 18847
rect 27890 18816 27896 18828
rect 25648 18788 27200 18816
rect 27264 18788 27896 18816
rect 25648 18776 25654 18788
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19392 18720 19625 18748
rect 19392 18708 19398 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 19702 18708 19708 18760
rect 19760 18748 19766 18760
rect 19797 18751 19855 18757
rect 19797 18748 19809 18751
rect 19760 18720 19809 18748
rect 19760 18708 19766 18720
rect 19797 18717 19809 18720
rect 19843 18717 19855 18751
rect 19797 18711 19855 18717
rect 20530 18708 20536 18760
rect 20588 18708 20594 18760
rect 21542 18708 21548 18760
rect 21600 18748 21606 18760
rect 21821 18751 21879 18757
rect 21821 18748 21833 18751
rect 21600 18720 21833 18748
rect 21600 18708 21606 18720
rect 21821 18717 21833 18720
rect 21867 18717 21879 18751
rect 21821 18711 21879 18717
rect 23566 18708 23572 18760
rect 23624 18748 23630 18760
rect 24397 18751 24455 18757
rect 24397 18748 24409 18751
rect 23624 18720 24409 18748
rect 23624 18708 23630 18720
rect 24397 18717 24409 18720
rect 24443 18748 24455 18751
rect 24486 18748 24492 18760
rect 24443 18720 24492 18748
rect 24443 18717 24455 18720
rect 24397 18711 24455 18717
rect 24486 18708 24492 18720
rect 24544 18708 24550 18760
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18748 24639 18751
rect 24762 18748 24768 18760
rect 24627 18720 24768 18748
rect 24627 18717 24639 18720
rect 24581 18711 24639 18717
rect 23198 18640 23204 18692
rect 23256 18680 23262 18692
rect 24596 18680 24624 18711
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 25314 18708 25320 18760
rect 25372 18708 25378 18760
rect 26970 18708 26976 18760
rect 27028 18708 27034 18760
rect 23256 18652 24624 18680
rect 23256 18640 23262 18652
rect 26142 18640 26148 18692
rect 26200 18680 26206 18692
rect 27264 18680 27292 18788
rect 27890 18776 27896 18788
rect 27948 18816 27954 18828
rect 27985 18819 28043 18825
rect 27985 18816 27997 18819
rect 27948 18788 27997 18816
rect 27948 18776 27954 18788
rect 27985 18785 27997 18788
rect 28031 18785 28043 18819
rect 27985 18779 28043 18785
rect 28074 18776 28080 18828
rect 28132 18816 28138 18828
rect 28537 18819 28595 18825
rect 28132 18788 28396 18816
rect 28132 18776 28138 18788
rect 28368 18760 28396 18788
rect 28537 18785 28549 18819
rect 28583 18816 28595 18819
rect 28920 18816 28948 18924
rect 29178 18912 29184 18964
rect 29236 18912 29242 18964
rect 29825 18955 29883 18961
rect 29825 18921 29837 18955
rect 29871 18952 29883 18955
rect 29914 18952 29920 18964
rect 29871 18924 29920 18952
rect 29871 18921 29883 18924
rect 29825 18915 29883 18921
rect 29914 18912 29920 18924
rect 29972 18912 29978 18964
rect 30466 18912 30472 18964
rect 30524 18952 30530 18964
rect 33781 18955 33839 18961
rect 33781 18952 33793 18955
rect 30524 18924 33793 18952
rect 30524 18912 30530 18924
rect 33781 18921 33793 18924
rect 33827 18921 33839 18955
rect 33781 18915 33839 18921
rect 28583 18788 28948 18816
rect 28583 18785 28595 18788
rect 28537 18779 28595 18785
rect 30374 18776 30380 18828
rect 30432 18776 30438 18828
rect 32398 18776 32404 18828
rect 32456 18776 32462 18828
rect 34146 18776 34152 18828
rect 34204 18816 34210 18828
rect 34977 18819 35035 18825
rect 34977 18816 34989 18819
rect 34204 18788 34989 18816
rect 34204 18776 34210 18788
rect 34977 18785 34989 18788
rect 35023 18785 35035 18819
rect 34977 18779 35035 18785
rect 27338 18708 27344 18760
rect 27396 18708 27402 18760
rect 27522 18708 27528 18760
rect 27580 18708 27586 18760
rect 28258 18708 28264 18760
rect 28316 18708 28322 18760
rect 28350 18708 28356 18760
rect 28408 18757 28414 18760
rect 28408 18751 28436 18757
rect 28424 18717 28436 18751
rect 28408 18711 28436 18717
rect 28408 18708 28414 18711
rect 29822 18708 29828 18760
rect 29880 18748 29886 18760
rect 30193 18751 30251 18757
rect 30193 18748 30205 18751
rect 29880 18720 30205 18748
rect 29880 18708 29886 18720
rect 30193 18717 30205 18720
rect 30239 18717 30251 18751
rect 30193 18711 30251 18717
rect 30285 18751 30343 18757
rect 30285 18717 30297 18751
rect 30331 18748 30343 18751
rect 30834 18748 30840 18760
rect 30331 18720 30840 18748
rect 30331 18717 30343 18720
rect 30285 18711 30343 18717
rect 26200 18652 27292 18680
rect 26200 18640 26206 18652
rect 11756 18584 18828 18612
rect 11756 18572 11762 18584
rect 20254 18572 20260 18624
rect 20312 18612 20318 18624
rect 20530 18612 20536 18624
rect 20312 18584 20536 18612
rect 20312 18572 20318 18584
rect 20530 18572 20536 18584
rect 20588 18572 20594 18624
rect 23934 18572 23940 18624
rect 23992 18612 23998 18624
rect 25314 18612 25320 18624
rect 23992 18584 25320 18612
rect 23992 18572 23998 18584
rect 25314 18572 25320 18584
rect 25372 18572 25378 18624
rect 27540 18612 27568 18708
rect 30300 18612 30328 18711
rect 30834 18708 30840 18720
rect 30892 18708 30898 18760
rect 30929 18751 30987 18757
rect 30929 18717 30941 18751
rect 30975 18748 30987 18751
rect 31570 18748 31576 18760
rect 30975 18720 31576 18748
rect 30975 18717 30987 18720
rect 30929 18711 30987 18717
rect 31570 18708 31576 18720
rect 31628 18708 31634 18760
rect 34606 18708 34612 18760
rect 34664 18748 34670 18760
rect 34701 18751 34759 18757
rect 34701 18748 34713 18751
rect 34664 18720 34713 18748
rect 34664 18708 34670 18720
rect 34701 18717 34713 18720
rect 34747 18717 34759 18751
rect 34701 18711 34759 18717
rect 31202 18689 31208 18692
rect 31196 18643 31208 18689
rect 31202 18640 31208 18643
rect 31260 18640 31266 18692
rect 32214 18640 32220 18692
rect 32272 18680 32278 18692
rect 32646 18683 32704 18689
rect 32646 18680 32658 18683
rect 32272 18652 32658 18680
rect 32272 18640 32278 18652
rect 32646 18649 32658 18652
rect 32692 18649 32704 18683
rect 32646 18643 32704 18649
rect 27540 18584 30328 18612
rect 31018 18572 31024 18624
rect 31076 18612 31082 18624
rect 32309 18615 32367 18621
rect 32309 18612 32321 18615
rect 31076 18584 32321 18612
rect 31076 18572 31082 18584
rect 32309 18581 32321 18584
rect 32355 18581 32367 18615
rect 32309 18575 32367 18581
rect 1104 18522 36800 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 36800 18522
rect 1104 18448 36800 18470
rect 4982 18368 4988 18420
rect 5040 18408 5046 18420
rect 5626 18408 5632 18420
rect 5040 18380 5632 18408
rect 5040 18368 5046 18380
rect 5626 18368 5632 18380
rect 5684 18368 5690 18420
rect 6181 18411 6239 18417
rect 6181 18377 6193 18411
rect 6227 18408 6239 18411
rect 6362 18408 6368 18420
rect 6227 18380 6368 18408
rect 6227 18377 6239 18380
rect 6181 18371 6239 18377
rect 6362 18368 6368 18380
rect 6420 18368 6426 18420
rect 7190 18408 7196 18420
rect 6564 18380 7196 18408
rect 2685 18343 2743 18349
rect 2685 18309 2697 18343
rect 2731 18340 2743 18343
rect 2866 18340 2872 18352
rect 2731 18312 2872 18340
rect 2731 18309 2743 18312
rect 2685 18303 2743 18309
rect 2866 18300 2872 18312
rect 2924 18300 2930 18352
rect 6086 18300 6092 18352
rect 6144 18340 6150 18352
rect 6564 18340 6592 18380
rect 7190 18368 7196 18380
rect 7248 18408 7254 18420
rect 7248 18380 8156 18408
rect 7248 18368 7254 18380
rect 6144 18312 6592 18340
rect 8128 18340 8156 18380
rect 8202 18368 8208 18420
rect 8260 18368 8266 18420
rect 9030 18368 9036 18420
rect 9088 18368 9094 18420
rect 9122 18368 9128 18420
rect 9180 18408 9186 18420
rect 10502 18408 10508 18420
rect 9180 18380 10508 18408
rect 9180 18368 9186 18380
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 11146 18368 11152 18420
rect 11204 18408 11210 18420
rect 11333 18411 11391 18417
rect 11333 18408 11345 18411
rect 11204 18380 11345 18408
rect 11204 18368 11210 18380
rect 11333 18377 11345 18380
rect 11379 18377 11391 18411
rect 11333 18371 11391 18377
rect 11882 18368 11888 18420
rect 11940 18368 11946 18420
rect 13998 18368 14004 18420
rect 14056 18408 14062 18420
rect 14737 18411 14795 18417
rect 14737 18408 14749 18411
rect 14056 18380 14749 18408
rect 14056 18368 14062 18380
rect 14737 18377 14749 18380
rect 14783 18377 14795 18411
rect 14737 18371 14795 18377
rect 15194 18368 15200 18420
rect 15252 18368 15258 18420
rect 16482 18368 16488 18420
rect 16540 18408 16546 18420
rect 17586 18408 17592 18420
rect 16540 18380 17592 18408
rect 16540 18368 16546 18380
rect 17586 18368 17592 18380
rect 17644 18368 17650 18420
rect 18506 18368 18512 18420
rect 18564 18368 18570 18420
rect 18616 18380 21036 18408
rect 8846 18340 8852 18352
rect 8128 18312 8852 18340
rect 6144 18300 6150 18312
rect 8846 18300 8852 18312
rect 8904 18300 8910 18352
rect 9214 18340 9220 18352
rect 8956 18312 9220 18340
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 4341 18275 4399 18281
rect 4341 18272 4353 18275
rect 4120 18244 4353 18272
rect 4120 18232 4126 18244
rect 4341 18241 4353 18244
rect 4387 18241 4399 18275
rect 4341 18235 4399 18241
rect 4522 18232 4528 18284
rect 4580 18232 4586 18284
rect 8956 18281 8984 18312
rect 9214 18300 9220 18312
rect 9272 18300 9278 18352
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18241 8999 18275
rect 8941 18235 8999 18241
rect 9125 18275 9183 18281
rect 9125 18241 9137 18275
rect 9171 18272 9183 18275
rect 9398 18272 9404 18284
rect 9171 18244 9404 18272
rect 9171 18241 9183 18244
rect 9125 18235 9183 18241
rect 9398 18232 9404 18244
rect 9456 18272 9462 18284
rect 9493 18275 9551 18281
rect 9493 18272 9505 18275
rect 9456 18244 9505 18272
rect 9456 18232 9462 18244
rect 9493 18241 9505 18244
rect 9539 18241 9551 18275
rect 9858 18272 9864 18284
rect 9493 18235 9551 18241
rect 9600 18244 9864 18272
rect 2682 18164 2688 18216
rect 2740 18204 2746 18216
rect 2777 18207 2835 18213
rect 2777 18204 2789 18207
rect 2740 18176 2789 18204
rect 2740 18164 2746 18176
rect 2777 18173 2789 18176
rect 2823 18173 2835 18207
rect 2777 18167 2835 18173
rect 2958 18164 2964 18216
rect 3016 18164 3022 18216
rect 4540 18204 4568 18232
rect 5074 18204 5080 18216
rect 4540 18176 5080 18204
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 5258 18164 5264 18216
rect 5316 18164 5322 18216
rect 5442 18213 5448 18216
rect 5399 18207 5448 18213
rect 5399 18173 5411 18207
rect 5445 18173 5448 18207
rect 5399 18167 5448 18173
rect 5442 18164 5448 18167
rect 5500 18164 5506 18216
rect 5537 18207 5595 18213
rect 5537 18173 5549 18207
rect 5583 18204 5595 18207
rect 6086 18204 6092 18216
rect 5583 18176 6092 18204
rect 5583 18173 5595 18176
rect 5537 18167 5595 18173
rect 6086 18164 6092 18176
rect 6144 18164 6150 18216
rect 6362 18164 6368 18216
rect 6420 18164 6426 18216
rect 6546 18164 6552 18216
rect 6604 18164 6610 18216
rect 6914 18164 6920 18216
rect 6972 18204 6978 18216
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 6972 18176 7297 18204
rect 6972 18164 6978 18176
rect 7285 18173 7297 18176
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 7374 18164 7380 18216
rect 7432 18213 7438 18216
rect 7432 18207 7460 18213
rect 7448 18173 7460 18207
rect 7432 18167 7460 18173
rect 7561 18207 7619 18213
rect 7561 18173 7573 18207
rect 7607 18204 7619 18207
rect 9600 18204 9628 18244
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 10410 18232 10416 18284
rect 10468 18232 10474 18284
rect 10502 18232 10508 18284
rect 10560 18281 10566 18284
rect 10560 18275 10588 18281
rect 10576 18241 10588 18275
rect 10560 18235 10588 18241
rect 10560 18232 10566 18235
rect 10686 18232 10692 18284
rect 10744 18232 10750 18284
rect 12066 18232 12072 18284
rect 12124 18232 12130 18284
rect 12894 18232 12900 18284
rect 12952 18232 12958 18284
rect 13078 18232 13084 18284
rect 13136 18232 13142 18284
rect 13814 18232 13820 18284
rect 13872 18232 13878 18284
rect 13906 18232 13912 18284
rect 13964 18281 13970 18284
rect 13964 18275 13992 18281
rect 13980 18241 13992 18275
rect 13964 18235 13992 18241
rect 13964 18232 13970 18235
rect 15378 18232 15384 18284
rect 15436 18232 15442 18284
rect 16298 18232 16304 18284
rect 16356 18272 16362 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16356 18244 16681 18272
rect 16356 18232 16362 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 17586 18232 17592 18284
rect 17644 18232 17650 18284
rect 17862 18232 17868 18284
rect 17920 18232 17926 18284
rect 18616 18281 18644 18380
rect 21008 18340 21036 18380
rect 21174 18368 21180 18420
rect 21232 18368 21238 18420
rect 21634 18368 21640 18420
rect 21692 18408 21698 18420
rect 22189 18411 22247 18417
rect 22189 18408 22201 18411
rect 21692 18380 22201 18408
rect 21692 18368 21698 18380
rect 22189 18377 22201 18380
rect 22235 18377 22247 18411
rect 22189 18371 22247 18377
rect 24857 18411 24915 18417
rect 24857 18377 24869 18411
rect 24903 18408 24915 18411
rect 25130 18408 25136 18420
rect 24903 18380 25136 18408
rect 24903 18377 24915 18380
rect 24857 18371 24915 18377
rect 25130 18368 25136 18380
rect 25188 18368 25194 18420
rect 25406 18368 25412 18420
rect 25464 18408 25470 18420
rect 26329 18411 26387 18417
rect 26329 18408 26341 18411
rect 25464 18380 26341 18408
rect 25464 18368 25470 18380
rect 26329 18377 26341 18380
rect 26375 18377 26387 18411
rect 26329 18371 26387 18377
rect 28442 18368 28448 18420
rect 28500 18408 28506 18420
rect 28629 18411 28687 18417
rect 28629 18408 28641 18411
rect 28500 18380 28641 18408
rect 28500 18368 28506 18380
rect 28629 18377 28641 18380
rect 28675 18377 28687 18411
rect 28629 18371 28687 18377
rect 31202 18368 31208 18420
rect 31260 18368 31266 18420
rect 32214 18368 32220 18420
rect 32272 18368 32278 18420
rect 32398 18368 32404 18420
rect 32456 18368 32462 18420
rect 35342 18368 35348 18420
rect 35400 18368 35406 18420
rect 27985 18343 28043 18349
rect 21008 18312 22508 18340
rect 18601 18275 18659 18281
rect 18601 18241 18613 18275
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 19334 18232 19340 18284
rect 19392 18232 19398 18284
rect 20254 18232 20260 18284
rect 20312 18232 20318 18284
rect 20530 18232 20536 18284
rect 20588 18232 20594 18284
rect 7607 18176 9628 18204
rect 7607 18173 7619 18176
rect 7561 18167 7619 18173
rect 7432 18164 7438 18167
rect 9674 18164 9680 18216
rect 9732 18164 9738 18216
rect 13170 18164 13176 18216
rect 13228 18204 13234 18216
rect 13924 18204 13952 18232
rect 13228 18176 13952 18204
rect 14093 18207 14151 18213
rect 13228 18164 13234 18176
rect 14093 18173 14105 18207
rect 14139 18204 14151 18207
rect 14458 18204 14464 18216
rect 14139 18176 14464 18204
rect 14139 18173 14151 18176
rect 14093 18167 14151 18173
rect 14458 18164 14464 18176
rect 14516 18164 14522 18216
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 16850 18204 16856 18216
rect 16632 18176 16856 18204
rect 16632 18164 16638 18176
rect 16850 18164 16856 18176
rect 16908 18164 16914 18216
rect 17402 18164 17408 18216
rect 17460 18204 17466 18216
rect 17706 18207 17764 18213
rect 17706 18204 17718 18207
rect 17460 18176 17718 18204
rect 17460 18164 17466 18176
rect 17706 18173 17718 18176
rect 17752 18173 17764 18207
rect 17880 18204 17908 18232
rect 19426 18204 19432 18216
rect 17880 18176 19432 18204
rect 17706 18167 17764 18173
rect 19426 18164 19432 18176
rect 19484 18164 19490 18216
rect 19521 18207 19579 18213
rect 19521 18173 19533 18207
rect 19567 18204 19579 18207
rect 19702 18204 19708 18216
rect 19567 18176 19708 18204
rect 19567 18173 19579 18176
rect 19521 18167 19579 18173
rect 19702 18164 19708 18176
rect 19760 18204 19766 18216
rect 19760 18176 20116 18204
rect 19760 18164 19766 18176
rect 4982 18096 4988 18148
rect 5040 18096 5046 18148
rect 7006 18096 7012 18148
rect 7064 18096 7070 18148
rect 10134 18096 10140 18148
rect 10192 18096 10198 18148
rect 13541 18139 13599 18145
rect 13541 18136 13553 18139
rect 12406 18108 13553 18136
rect 2038 18028 2044 18080
rect 2096 18068 2102 18080
rect 2317 18071 2375 18077
rect 2317 18068 2329 18071
rect 2096 18040 2329 18068
rect 2096 18028 2102 18040
rect 2317 18037 2329 18040
rect 2363 18037 2375 18071
rect 2317 18031 2375 18037
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 12406 18068 12434 18108
rect 13541 18105 13553 18108
rect 13587 18136 13599 18139
rect 13630 18136 13636 18148
rect 13587 18108 13636 18136
rect 13587 18105 13599 18108
rect 13541 18099 13599 18105
rect 13630 18096 13636 18108
rect 13688 18096 13694 18148
rect 4856 18040 12434 18068
rect 4856 18028 4862 18040
rect 12618 18028 12624 18080
rect 12676 18068 12682 18080
rect 14476 18068 14504 18164
rect 17313 18139 17371 18145
rect 17313 18105 17325 18139
rect 17359 18105 17371 18139
rect 18874 18136 18880 18148
rect 17313 18099 17371 18105
rect 18248 18108 18880 18136
rect 12676 18040 14504 18068
rect 12676 18028 12682 18040
rect 14550 18028 14556 18080
rect 14608 18068 14614 18080
rect 17328 18068 17356 18099
rect 18248 18068 18276 18108
rect 18874 18096 18880 18108
rect 18932 18096 18938 18148
rect 19978 18096 19984 18148
rect 20036 18096 20042 18148
rect 14608 18040 18276 18068
rect 14608 18028 14614 18040
rect 18782 18028 18788 18080
rect 18840 18028 18846 18080
rect 20088 18068 20116 18176
rect 20346 18164 20352 18216
rect 20404 18213 20410 18216
rect 20404 18207 20432 18213
rect 20420 18173 20432 18207
rect 22094 18204 22100 18216
rect 20404 18167 20432 18173
rect 20916 18176 22100 18204
rect 20404 18164 20410 18167
rect 20916 18068 20944 18176
rect 22094 18164 22100 18176
rect 22152 18204 22158 18216
rect 22480 18213 22508 18312
rect 27985 18309 27997 18343
rect 28031 18340 28043 18343
rect 28031 18309 28053 18340
rect 27985 18303 28053 18309
rect 22922 18232 22928 18284
rect 22980 18232 22986 18284
rect 23198 18232 23204 18284
rect 23256 18232 23262 18284
rect 23934 18232 23940 18284
rect 23992 18232 23998 18284
rect 24210 18232 24216 18284
rect 24268 18232 24274 18284
rect 25038 18232 25044 18284
rect 25096 18272 25102 18284
rect 25205 18275 25263 18281
rect 25205 18272 25217 18275
rect 25096 18244 25217 18272
rect 25096 18232 25102 18244
rect 25205 18241 25217 18244
rect 25251 18241 25263 18275
rect 25205 18235 25263 18241
rect 25958 18232 25964 18284
rect 26016 18272 26022 18284
rect 27249 18275 27307 18281
rect 27249 18272 27261 18275
rect 26016 18244 27261 18272
rect 26016 18232 26022 18244
rect 27249 18241 27261 18244
rect 27295 18241 27307 18275
rect 27249 18235 27307 18241
rect 22281 18207 22339 18213
rect 22281 18204 22293 18207
rect 22152 18176 22293 18204
rect 22152 18164 22158 18176
rect 22281 18173 22293 18176
rect 22327 18173 22339 18207
rect 22281 18167 22339 18173
rect 22465 18207 22523 18213
rect 22465 18173 22477 18207
rect 22511 18204 22523 18207
rect 23017 18207 23075 18213
rect 22511 18176 22968 18204
rect 22511 18173 22523 18176
rect 22465 18167 22523 18173
rect 20088 18040 20944 18068
rect 21818 18028 21824 18080
rect 21876 18028 21882 18080
rect 22738 18028 22744 18080
rect 22796 18028 22802 18080
rect 22940 18068 22968 18176
rect 23017 18173 23029 18207
rect 23063 18204 23075 18207
rect 23566 18204 23572 18216
rect 23063 18176 23572 18204
rect 23063 18173 23075 18176
rect 23017 18167 23075 18173
rect 23566 18164 23572 18176
rect 23624 18164 23630 18216
rect 23658 18164 23664 18216
rect 23716 18164 23722 18216
rect 23750 18164 23756 18216
rect 23808 18204 23814 18216
rect 23952 18204 23980 18232
rect 23808 18176 23980 18204
rect 23808 18164 23814 18176
rect 24026 18164 24032 18216
rect 24084 18213 24090 18216
rect 24084 18207 24112 18213
rect 24100 18173 24112 18207
rect 24084 18167 24112 18173
rect 24084 18164 24090 18167
rect 24854 18164 24860 18216
rect 24912 18204 24918 18216
rect 24949 18207 25007 18213
rect 24949 18204 24961 18207
rect 24912 18176 24961 18204
rect 24912 18164 24918 18176
rect 24949 18173 24961 18176
rect 24995 18173 25007 18207
rect 24949 18167 25007 18173
rect 26878 18164 26884 18216
rect 26936 18204 26942 18216
rect 26973 18207 27031 18213
rect 26973 18204 26985 18207
rect 26936 18176 26985 18204
rect 26936 18164 26942 18176
rect 26973 18173 26985 18176
rect 27019 18173 27031 18207
rect 28025 18204 28053 18303
rect 28534 18300 28540 18352
rect 28592 18340 28598 18352
rect 30745 18343 30803 18349
rect 28592 18312 28994 18340
rect 28592 18300 28598 18312
rect 28966 18272 28994 18312
rect 30745 18309 30757 18343
rect 30791 18340 30803 18343
rect 31294 18340 31300 18352
rect 30791 18312 31300 18340
rect 30791 18309 30803 18312
rect 30745 18303 30803 18309
rect 31294 18300 31300 18312
rect 31352 18300 31358 18352
rect 32416 18340 32444 18368
rect 34698 18340 34704 18352
rect 32416 18312 33088 18340
rect 30374 18272 30380 18284
rect 28966 18244 30380 18272
rect 30374 18232 30380 18244
rect 30432 18232 30438 18284
rect 30484 18244 31064 18272
rect 28626 18204 28632 18216
rect 28025 18176 28632 18204
rect 26973 18167 27031 18173
rect 25682 18068 25688 18080
rect 22940 18040 25688 18068
rect 25682 18028 25688 18040
rect 25740 18028 25746 18080
rect 26988 18068 27016 18167
rect 28626 18164 28632 18176
rect 28684 18164 28690 18216
rect 30484 18204 30512 18244
rect 28736 18176 30512 18204
rect 27890 18096 27896 18148
rect 27948 18136 27954 18148
rect 28169 18139 28227 18145
rect 28169 18136 28181 18139
rect 27948 18108 28181 18136
rect 27948 18096 27954 18108
rect 28169 18105 28181 18108
rect 28215 18105 28227 18139
rect 28736 18136 28764 18176
rect 30558 18164 30564 18216
rect 30616 18204 30622 18216
rect 30837 18207 30895 18213
rect 30837 18204 30849 18207
rect 30616 18176 30849 18204
rect 30616 18164 30622 18176
rect 30837 18173 30849 18176
rect 30883 18173 30895 18207
rect 30837 18167 30895 18173
rect 30926 18164 30932 18216
rect 30984 18164 30990 18216
rect 31036 18204 31064 18244
rect 31386 18232 31392 18284
rect 31444 18232 31450 18284
rect 32398 18232 32404 18284
rect 32456 18232 32462 18284
rect 33060 18281 33088 18312
rect 33152 18312 34704 18340
rect 33045 18275 33103 18281
rect 33045 18241 33057 18275
rect 33091 18241 33103 18275
rect 33045 18235 33103 18241
rect 33152 18204 33180 18312
rect 34698 18300 34704 18312
rect 34756 18300 34762 18352
rect 33318 18281 33324 18284
rect 33312 18235 33324 18281
rect 33318 18232 33324 18235
rect 33376 18232 33382 18284
rect 35161 18275 35219 18281
rect 35161 18241 35173 18275
rect 35207 18272 35219 18275
rect 35434 18272 35440 18284
rect 35207 18244 35440 18272
rect 35207 18241 35219 18244
rect 35161 18235 35219 18241
rect 35434 18232 35440 18244
rect 35492 18232 35498 18284
rect 31036 18176 33180 18204
rect 34514 18164 34520 18216
rect 34572 18204 34578 18216
rect 34701 18207 34759 18213
rect 34701 18204 34713 18207
rect 34572 18176 34713 18204
rect 34572 18164 34578 18176
rect 34701 18173 34713 18176
rect 34747 18173 34759 18207
rect 34701 18167 34759 18173
rect 34790 18164 34796 18216
rect 34848 18204 34854 18216
rect 35069 18207 35127 18213
rect 35069 18204 35081 18207
rect 34848 18176 35081 18204
rect 34848 18164 34854 18176
rect 35069 18173 35081 18176
rect 35115 18173 35127 18207
rect 35069 18167 35127 18173
rect 28169 18099 28227 18105
rect 28552 18108 28764 18136
rect 30377 18139 30435 18145
rect 28552 18068 28580 18108
rect 30377 18105 30389 18139
rect 30423 18136 30435 18139
rect 31386 18136 31392 18148
rect 30423 18108 31392 18136
rect 30423 18105 30435 18108
rect 30377 18099 30435 18105
rect 31386 18096 31392 18108
rect 31444 18096 31450 18148
rect 31726 18108 32352 18136
rect 26988 18040 28580 18068
rect 28626 18028 28632 18080
rect 28684 18068 28690 18080
rect 31726 18068 31754 18108
rect 28684 18040 31754 18068
rect 32324 18068 32352 18108
rect 34425 18071 34483 18077
rect 34425 18068 34437 18071
rect 32324 18040 34437 18068
rect 28684 18028 28690 18040
rect 34425 18037 34437 18040
rect 34471 18037 34483 18071
rect 34425 18031 34483 18037
rect 34698 18028 34704 18080
rect 34756 18068 34762 18080
rect 35342 18068 35348 18080
rect 34756 18040 35348 18068
rect 34756 18028 34762 18040
rect 35342 18028 35348 18040
rect 35400 18028 35406 18080
rect 1104 17978 36800 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 36800 17978
rect 1104 17904 36800 17926
rect 5074 17824 5080 17876
rect 5132 17864 5138 17876
rect 5169 17867 5227 17873
rect 5169 17864 5181 17867
rect 5132 17836 5181 17864
rect 5132 17824 5138 17836
rect 5169 17833 5181 17836
rect 5215 17864 5227 17867
rect 5258 17864 5264 17876
rect 5215 17836 5264 17864
rect 5215 17833 5227 17836
rect 5169 17827 5227 17833
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 5368 17836 7604 17864
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17660 1455 17663
rect 1486 17660 1492 17672
rect 1443 17632 1492 17660
rect 1443 17629 1455 17632
rect 1397 17623 1455 17629
rect 1486 17620 1492 17632
rect 1544 17660 1550 17672
rect 2774 17660 2780 17672
rect 1544 17632 2780 17660
rect 1544 17620 1550 17632
rect 2774 17620 2780 17632
rect 2832 17660 2838 17672
rect 3789 17663 3847 17669
rect 3789 17660 3801 17663
rect 2832 17632 3801 17660
rect 2832 17620 2838 17632
rect 3789 17629 3801 17632
rect 3835 17660 3847 17663
rect 5368 17660 5396 17836
rect 5626 17756 5632 17808
rect 5684 17796 5690 17808
rect 6638 17796 6644 17808
rect 5684 17768 6644 17796
rect 5684 17756 5690 17768
rect 6638 17756 6644 17768
rect 6696 17756 6702 17808
rect 7576 17796 7604 17836
rect 7742 17824 7748 17876
rect 7800 17864 7806 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 7800 17836 7849 17864
rect 7800 17824 7806 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 7837 17827 7895 17833
rect 9490 17824 9496 17876
rect 9548 17864 9554 17876
rect 9677 17867 9735 17873
rect 9677 17864 9689 17867
rect 9548 17836 9689 17864
rect 9548 17824 9554 17836
rect 9677 17833 9689 17836
rect 9723 17833 9735 17867
rect 10183 17867 10241 17873
rect 10183 17864 10195 17867
rect 9677 17827 9735 17833
rect 9784 17836 10195 17864
rect 8018 17796 8024 17808
rect 7576 17768 8024 17796
rect 8018 17756 8024 17768
rect 8076 17756 8082 17808
rect 9784 17796 9812 17836
rect 10183 17833 10195 17836
rect 10229 17833 10241 17867
rect 10183 17827 10241 17833
rect 10410 17824 10416 17876
rect 10468 17864 10474 17876
rect 14642 17864 14648 17876
rect 10468 17836 14648 17864
rect 10468 17824 10474 17836
rect 14642 17824 14648 17836
rect 14700 17824 14706 17876
rect 22094 17824 22100 17876
rect 22152 17824 22158 17876
rect 23842 17824 23848 17876
rect 23900 17824 23906 17876
rect 24949 17867 25007 17873
rect 24949 17833 24961 17867
rect 24995 17864 25007 17867
rect 25038 17864 25044 17876
rect 24995 17836 25044 17864
rect 24995 17833 25007 17836
rect 24949 17827 25007 17833
rect 25038 17824 25044 17836
rect 25096 17824 25102 17876
rect 25130 17824 25136 17876
rect 25188 17864 25194 17876
rect 25188 17836 28120 17864
rect 25188 17824 25194 17836
rect 9508 17768 9812 17796
rect 27341 17799 27399 17805
rect 5997 17731 6055 17737
rect 5997 17697 6009 17731
rect 6043 17728 6055 17731
rect 6362 17728 6368 17740
rect 6043 17700 6368 17728
rect 6043 17697 6055 17700
rect 5997 17691 6055 17697
rect 3835 17632 5396 17660
rect 3835 17629 3847 17632
rect 3789 17623 3847 17629
rect 1664 17595 1722 17601
rect 1664 17561 1676 17595
rect 1710 17592 1722 17595
rect 1854 17592 1860 17604
rect 1710 17564 1860 17592
rect 1710 17561 1722 17564
rect 1664 17555 1722 17561
rect 1854 17552 1860 17564
rect 1912 17552 1918 17604
rect 4062 17601 4068 17604
rect 4056 17555 4068 17601
rect 4062 17552 4068 17555
rect 4120 17552 4126 17604
rect 2777 17527 2835 17533
rect 2777 17493 2789 17527
rect 2823 17524 2835 17527
rect 2866 17524 2872 17536
rect 2823 17496 2872 17524
rect 2823 17493 2835 17496
rect 2777 17487 2835 17493
rect 2866 17484 2872 17496
rect 2924 17524 2930 17536
rect 6012 17524 6040 17691
rect 6362 17688 6368 17700
rect 6420 17688 6426 17740
rect 6914 17688 6920 17740
rect 6972 17688 6978 17740
rect 7374 17728 7380 17740
rect 7024 17700 7380 17728
rect 7024 17672 7052 17700
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 6181 17663 6239 17669
rect 6181 17629 6193 17663
rect 6227 17629 6239 17663
rect 6181 17623 6239 17629
rect 2924 17496 6040 17524
rect 6196 17524 6224 17623
rect 7006 17620 7012 17672
rect 7064 17669 7070 17672
rect 7064 17663 7092 17669
rect 7080 17629 7092 17663
rect 7064 17623 7092 17629
rect 7064 17620 7070 17623
rect 7190 17620 7196 17672
rect 7248 17620 7254 17672
rect 7926 17620 7932 17672
rect 7984 17660 7990 17672
rect 9508 17669 9536 17768
rect 27341 17765 27353 17799
rect 27387 17765 27399 17799
rect 27341 17759 27399 17765
rect 9861 17731 9919 17737
rect 9861 17697 9873 17731
rect 9907 17728 9919 17731
rect 10965 17731 11023 17737
rect 10965 17728 10977 17731
rect 9907 17700 10977 17728
rect 9907 17697 9919 17700
rect 9861 17691 9919 17697
rect 10965 17697 10977 17700
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 13078 17688 13084 17740
rect 13136 17728 13142 17740
rect 14550 17728 14556 17740
rect 13136 17700 14556 17728
rect 13136 17688 13142 17700
rect 14550 17688 14556 17700
rect 14608 17688 14614 17740
rect 14645 17731 14703 17737
rect 14645 17697 14657 17731
rect 14691 17728 14703 17731
rect 17589 17731 17647 17737
rect 17589 17728 17601 17731
rect 14691 17700 17601 17728
rect 14691 17697 14703 17700
rect 14645 17691 14703 17697
rect 17589 17697 17601 17700
rect 17635 17728 17647 17731
rect 18782 17728 18788 17740
rect 17635 17700 18788 17728
rect 17635 17697 17647 17700
rect 17589 17691 17647 17697
rect 9493 17663 9551 17669
rect 9493 17660 9505 17663
rect 7984 17632 9505 17660
rect 7984 17620 7990 17632
rect 9493 17629 9505 17632
rect 9539 17629 9551 17663
rect 9493 17623 9551 17629
rect 9582 17620 9588 17672
rect 9640 17620 9646 17672
rect 9953 17663 10011 17669
rect 9953 17629 9965 17663
rect 9999 17660 10011 17663
rect 10410 17660 10416 17672
rect 9999 17632 10416 17660
rect 9999 17629 10011 17632
rect 9953 17623 10011 17629
rect 10410 17620 10416 17632
rect 10468 17620 10474 17672
rect 10870 17620 10876 17672
rect 10928 17620 10934 17672
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17660 11115 17663
rect 14660 17660 14688 17691
rect 18782 17688 18788 17700
rect 18840 17688 18846 17740
rect 11103 17632 14688 17660
rect 11103 17629 11115 17632
rect 11057 17623 11115 17629
rect 9600 17592 9628 17620
rect 11072 17592 11100 17623
rect 17310 17620 17316 17672
rect 17368 17660 17374 17672
rect 17405 17663 17463 17669
rect 17405 17660 17417 17663
rect 17368 17632 17417 17660
rect 17368 17620 17374 17632
rect 17405 17629 17417 17632
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 18874 17620 18880 17672
rect 18932 17660 18938 17672
rect 18969 17663 19027 17669
rect 18969 17660 18981 17663
rect 18932 17632 18981 17660
rect 18932 17620 18938 17632
rect 18969 17629 18981 17632
rect 19015 17629 19027 17663
rect 18969 17623 19027 17629
rect 19242 17620 19248 17672
rect 19300 17620 19306 17672
rect 20717 17663 20775 17669
rect 20717 17629 20729 17663
rect 20763 17660 20775 17663
rect 20806 17660 20812 17672
rect 20763 17632 20812 17660
rect 20763 17629 20775 17632
rect 20717 17623 20775 17629
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 22738 17669 22744 17672
rect 22465 17663 22523 17669
rect 22465 17629 22477 17663
rect 22511 17629 22523 17663
rect 22732 17660 22744 17669
rect 22699 17632 22744 17660
rect 22465 17623 22523 17629
rect 22732 17623 22744 17632
rect 9600 17564 11100 17592
rect 13538 17552 13544 17604
rect 13596 17592 13602 17604
rect 14461 17595 14519 17601
rect 14461 17592 14473 17595
rect 13596 17564 14473 17592
rect 13596 17552 13602 17564
rect 14461 17561 14473 17564
rect 14507 17561 14519 17595
rect 14461 17555 14519 17561
rect 16850 17552 16856 17604
rect 16908 17592 16914 17604
rect 20990 17601 20996 17604
rect 19490 17595 19548 17601
rect 19490 17592 19502 17595
rect 16908 17564 17540 17592
rect 16908 17552 16914 17564
rect 6546 17524 6552 17536
rect 6196 17496 6552 17524
rect 2924 17484 2930 17496
rect 6546 17484 6552 17496
rect 6604 17524 6610 17536
rect 6822 17524 6828 17536
rect 6604 17496 6828 17524
rect 6604 17484 6610 17496
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 9306 17484 9312 17536
rect 9364 17484 9370 17536
rect 9861 17527 9919 17533
rect 9861 17493 9873 17527
rect 9907 17524 9919 17527
rect 9950 17524 9956 17536
rect 9907 17496 9956 17524
rect 9907 17493 9919 17496
rect 9861 17487 9919 17493
rect 9950 17484 9956 17496
rect 10008 17484 10014 17536
rect 13446 17484 13452 17536
rect 13504 17524 13510 17536
rect 14093 17527 14151 17533
rect 14093 17524 14105 17527
rect 13504 17496 14105 17524
rect 13504 17484 13510 17496
rect 14093 17493 14105 17496
rect 14139 17493 14151 17527
rect 14093 17487 14151 17493
rect 17034 17484 17040 17536
rect 17092 17484 17098 17536
rect 17512 17533 17540 17564
rect 18800 17564 19502 17592
rect 17497 17527 17555 17533
rect 17497 17493 17509 17527
rect 17543 17524 17555 17527
rect 17586 17524 17592 17536
rect 17543 17496 17592 17524
rect 17543 17493 17555 17496
rect 17497 17487 17555 17493
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 18800 17533 18828 17564
rect 19490 17561 19502 17564
rect 19536 17561 19548 17595
rect 19490 17555 19548 17561
rect 20984 17555 20996 17601
rect 20990 17552 20996 17555
rect 21048 17552 21054 17604
rect 22480 17592 22508 17623
rect 22738 17620 22744 17623
rect 22796 17620 22802 17672
rect 24946 17620 24952 17672
rect 25004 17660 25010 17672
rect 25133 17663 25191 17669
rect 25133 17660 25145 17663
rect 25004 17632 25145 17660
rect 25004 17620 25010 17632
rect 25133 17629 25145 17632
rect 25179 17629 25191 17663
rect 25133 17623 25191 17629
rect 25866 17620 25872 17672
rect 25924 17620 25930 17672
rect 25961 17663 26019 17669
rect 25961 17629 25973 17663
rect 26007 17629 26019 17663
rect 27356 17660 27384 17759
rect 28092 17737 28120 17836
rect 30466 17824 30472 17876
rect 30524 17864 30530 17876
rect 30929 17867 30987 17873
rect 30929 17864 30941 17867
rect 30524 17836 30941 17864
rect 30524 17824 30530 17836
rect 30929 17833 30941 17836
rect 30975 17833 30987 17867
rect 30929 17827 30987 17833
rect 33318 17824 33324 17876
rect 33376 17864 33382 17876
rect 33505 17867 33563 17873
rect 33505 17864 33517 17867
rect 33376 17836 33517 17864
rect 33376 17824 33382 17836
rect 33505 17833 33517 17836
rect 33551 17833 33563 17867
rect 33505 17827 33563 17833
rect 28077 17731 28135 17737
rect 28077 17697 28089 17731
rect 28123 17728 28135 17731
rect 28123 17700 28488 17728
rect 28123 17697 28135 17700
rect 28077 17691 28135 17697
rect 27801 17663 27859 17669
rect 27801 17660 27813 17663
rect 27356 17632 27813 17660
rect 25961 17623 26019 17629
rect 27801 17629 27813 17632
rect 27847 17660 27859 17663
rect 28350 17660 28356 17672
rect 27847 17632 28356 17660
rect 27847 17629 27859 17632
rect 27801 17623 27859 17629
rect 22646 17592 22652 17604
rect 22480 17564 22652 17592
rect 22646 17552 22652 17564
rect 22704 17592 22710 17604
rect 24854 17592 24860 17604
rect 22704 17564 24860 17592
rect 22704 17552 22710 17564
rect 24854 17552 24860 17564
rect 24912 17592 24918 17604
rect 25976 17592 26004 17623
rect 28350 17620 28356 17632
rect 28408 17620 28414 17672
rect 28460 17660 28488 17700
rect 29178 17688 29184 17740
rect 29236 17728 29242 17740
rect 29546 17728 29552 17740
rect 29236 17700 29552 17728
rect 29236 17688 29242 17700
rect 29546 17688 29552 17700
rect 29604 17688 29610 17740
rect 30650 17660 30656 17672
rect 28460 17632 30656 17660
rect 30650 17620 30656 17632
rect 30708 17620 30714 17672
rect 33594 17620 33600 17672
rect 33652 17660 33658 17672
rect 33689 17663 33747 17669
rect 33689 17660 33701 17663
rect 33652 17632 33701 17660
rect 33652 17620 33658 17632
rect 33689 17629 33701 17632
rect 33735 17629 33747 17663
rect 33689 17623 33747 17629
rect 26234 17601 26240 17604
rect 24912 17564 26004 17592
rect 24912 17552 24918 17564
rect 18785 17527 18843 17533
rect 18785 17493 18797 17527
rect 18831 17493 18843 17527
rect 18785 17487 18843 17493
rect 20622 17484 20628 17536
rect 20680 17484 20686 17536
rect 25700 17533 25728 17564
rect 26228 17555 26240 17601
rect 26234 17552 26240 17555
rect 26292 17552 26298 17604
rect 26418 17552 26424 17604
rect 26476 17592 26482 17604
rect 26476 17564 27476 17592
rect 26476 17552 26482 17564
rect 27448 17533 27476 17564
rect 29454 17552 29460 17604
rect 29512 17592 29518 17604
rect 29794 17595 29852 17601
rect 29794 17592 29806 17595
rect 29512 17564 29806 17592
rect 29512 17552 29518 17564
rect 29794 17561 29806 17564
rect 29840 17561 29852 17595
rect 29794 17555 29852 17561
rect 25685 17527 25743 17533
rect 25685 17493 25697 17527
rect 25731 17493 25743 17527
rect 25685 17487 25743 17493
rect 27433 17527 27491 17533
rect 27433 17493 27445 17527
rect 27479 17493 27491 17527
rect 27433 17487 27491 17493
rect 27893 17527 27951 17533
rect 27893 17493 27905 17527
rect 27939 17524 27951 17527
rect 28166 17524 28172 17536
rect 27939 17496 28172 17524
rect 27939 17493 27951 17496
rect 27893 17487 27951 17493
rect 28166 17484 28172 17496
rect 28224 17524 28230 17536
rect 30190 17524 30196 17536
rect 28224 17496 30196 17524
rect 28224 17484 28230 17496
rect 30190 17484 30196 17496
rect 30248 17484 30254 17536
rect 1104 17434 36800 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 36800 17434
rect 1104 17360 36800 17382
rect 1854 17280 1860 17332
rect 1912 17280 1918 17332
rect 3973 17323 4031 17329
rect 3973 17289 3985 17323
rect 4019 17320 4031 17323
rect 4062 17320 4068 17332
rect 4019 17292 4068 17320
rect 4019 17289 4031 17292
rect 3973 17283 4031 17289
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4433 17323 4491 17329
rect 4433 17289 4445 17323
rect 4479 17289 4491 17323
rect 4433 17283 4491 17289
rect 2038 17144 2044 17196
rect 2096 17144 2102 17196
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17184 4215 17187
rect 4448 17184 4476 17283
rect 4706 17280 4712 17332
rect 4764 17320 4770 17332
rect 4801 17323 4859 17329
rect 4801 17320 4813 17323
rect 4764 17292 4813 17320
rect 4764 17280 4770 17292
rect 4801 17289 4813 17292
rect 4847 17289 4859 17323
rect 4801 17283 4859 17289
rect 4893 17323 4951 17329
rect 4893 17289 4905 17323
rect 4939 17320 4951 17323
rect 5258 17320 5264 17332
rect 4939 17292 5264 17320
rect 4939 17289 4951 17292
rect 4893 17283 4951 17289
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 6089 17323 6147 17329
rect 6089 17289 6101 17323
rect 6135 17320 6147 17323
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 6135 17292 6837 17320
rect 6135 17289 6147 17292
rect 6089 17283 6147 17289
rect 6825 17289 6837 17292
rect 6871 17320 6883 17323
rect 7098 17320 7104 17332
rect 6871 17292 7104 17320
rect 6871 17289 6883 17292
rect 6825 17283 6883 17289
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 9674 17280 9680 17332
rect 9732 17320 9738 17332
rect 10870 17320 10876 17332
rect 9732 17292 10876 17320
rect 9732 17280 9738 17292
rect 10870 17280 10876 17292
rect 10928 17320 10934 17332
rect 11057 17323 11115 17329
rect 11057 17320 11069 17323
rect 10928 17292 11069 17320
rect 10928 17280 10934 17292
rect 11057 17289 11069 17292
rect 11103 17289 11115 17323
rect 11057 17283 11115 17289
rect 12897 17323 12955 17329
rect 12897 17289 12909 17323
rect 12943 17320 12955 17323
rect 13170 17320 13176 17332
rect 12943 17292 13176 17320
rect 12943 17289 12955 17292
rect 12897 17283 12955 17289
rect 13170 17280 13176 17292
rect 13228 17280 13234 17332
rect 13265 17323 13323 17329
rect 13265 17289 13277 17323
rect 13311 17289 13323 17323
rect 13265 17283 13323 17289
rect 9582 17252 9588 17264
rect 4203 17156 4476 17184
rect 5092 17224 9588 17252
rect 4203 17153 4215 17156
rect 4157 17147 4215 17153
rect 5092 17125 5120 17224
rect 5994 17144 6000 17196
rect 6052 17144 6058 17196
rect 7024 17125 7052 17224
rect 9582 17212 9588 17224
rect 9640 17212 9646 17264
rect 13280 17252 13308 17283
rect 14550 17280 14556 17332
rect 14608 17320 14614 17332
rect 14921 17323 14979 17329
rect 14921 17320 14933 17323
rect 14608 17292 14933 17320
rect 14608 17280 14614 17292
rect 14921 17289 14933 17292
rect 14967 17289 14979 17323
rect 14921 17283 14979 17289
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 18049 17323 18107 17329
rect 18049 17320 18061 17323
rect 17644 17292 18061 17320
rect 17644 17280 17650 17292
rect 18049 17289 18061 17292
rect 18095 17289 18107 17323
rect 18049 17283 18107 17289
rect 18874 17280 18880 17332
rect 18932 17280 18938 17332
rect 19245 17323 19303 17329
rect 19245 17289 19257 17323
rect 19291 17320 19303 17323
rect 20346 17320 20352 17332
rect 19291 17292 20352 17320
rect 19291 17289 19303 17292
rect 19245 17283 19303 17289
rect 20346 17280 20352 17292
rect 20404 17320 20410 17332
rect 20622 17320 20628 17332
rect 20404 17292 20628 17320
rect 20404 17280 20410 17292
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 20990 17280 20996 17332
rect 21048 17280 21054 17332
rect 22833 17323 22891 17329
rect 22833 17289 22845 17323
rect 22879 17320 22891 17323
rect 22922 17320 22928 17332
rect 22879 17292 22928 17320
rect 22879 17289 22891 17292
rect 22833 17283 22891 17289
rect 22922 17280 22928 17292
rect 22980 17280 22986 17332
rect 23201 17323 23259 17329
rect 23201 17289 23213 17323
rect 23247 17320 23259 17323
rect 23842 17320 23848 17332
rect 23247 17292 23848 17320
rect 23247 17289 23259 17292
rect 23201 17283 23259 17289
rect 23842 17280 23848 17292
rect 23900 17280 23906 17332
rect 26234 17280 26240 17332
rect 26292 17280 26298 17332
rect 27065 17323 27123 17329
rect 27065 17289 27077 17323
rect 27111 17289 27123 17323
rect 27065 17283 27123 17289
rect 13786 17255 13844 17261
rect 13786 17252 13798 17255
rect 13280 17224 13798 17252
rect 13786 17221 13798 17224
rect 13832 17221 13844 17255
rect 23293 17255 23351 17261
rect 13786 17215 13844 17221
rect 16224 17224 22094 17252
rect 9950 17193 9956 17196
rect 9944 17184 9956 17193
rect 9911 17156 9956 17184
rect 9944 17147 9956 17156
rect 9950 17144 9956 17147
rect 10008 17144 10014 17196
rect 11514 17144 11520 17196
rect 11572 17144 11578 17196
rect 11790 17193 11796 17196
rect 11784 17147 11796 17193
rect 11790 17144 11796 17147
rect 11848 17144 11854 17196
rect 13446 17144 13452 17196
rect 13504 17144 13510 17196
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17184 13599 17187
rect 14826 17184 14832 17196
rect 13587 17156 14832 17184
rect 13587 17153 13599 17156
rect 13541 17147 13599 17153
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17085 5135 17119
rect 6917 17119 6975 17125
rect 6917 17116 6929 17119
rect 5077 17079 5135 17085
rect 6840 17088 6929 17116
rect 6840 17060 6868 17088
rect 6917 17085 6929 17088
rect 6963 17085 6975 17119
rect 6917 17079 6975 17085
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17085 7067 17119
rect 7009 17079 7067 17085
rect 8846 17076 8852 17128
rect 8904 17116 8910 17128
rect 9306 17116 9312 17128
rect 8904 17088 9312 17116
rect 8904 17076 8910 17088
rect 9306 17076 9312 17088
rect 9364 17116 9370 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 9364 17088 9689 17116
rect 9364 17076 9370 17088
rect 9677 17085 9689 17088
rect 9723 17085 9735 17119
rect 9677 17079 9735 17085
rect 5258 17008 5264 17060
rect 5316 17048 5322 17060
rect 5316 17020 6684 17048
rect 5316 17008 5322 17020
rect 6457 16983 6515 16989
rect 6457 16949 6469 16983
rect 6503 16980 6515 16983
rect 6546 16980 6552 16992
rect 6503 16952 6552 16980
rect 6503 16949 6515 16952
rect 6457 16943 6515 16949
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 6656 16980 6684 17020
rect 6822 17008 6828 17060
rect 6880 17008 6886 17060
rect 8386 16980 8392 16992
rect 6656 16952 8392 16980
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 11514 16940 11520 16992
rect 11572 16980 11578 16992
rect 12526 16980 12532 16992
rect 11572 16952 12532 16980
rect 11572 16940 11578 16952
rect 12526 16940 12532 16952
rect 12584 16980 12590 16992
rect 13556 16980 13584 17147
rect 14826 17144 14832 17156
rect 14884 17144 14890 17196
rect 16224 17193 16252 17224
rect 16209 17187 16267 17193
rect 16209 17153 16221 17187
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 16632 17156 16681 17184
rect 16632 17144 16638 17156
rect 16669 17153 16681 17156
rect 16715 17184 16727 17187
rect 16758 17184 16764 17196
rect 16715 17156 16764 17184
rect 16715 17153 16727 17156
rect 16669 17147 16727 17153
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 16936 17187 16994 17193
rect 16936 17153 16948 17187
rect 16982 17184 16994 17187
rect 17218 17184 17224 17196
rect 16982 17156 17224 17184
rect 16982 17153 16994 17156
rect 16936 17147 16994 17153
rect 17218 17144 17224 17156
rect 17276 17144 17282 17196
rect 19444 17125 19472 17224
rect 21177 17187 21235 17193
rect 21177 17153 21189 17187
rect 21223 17184 21235 17187
rect 21818 17184 21824 17196
rect 21223 17156 21824 17184
rect 21223 17153 21235 17156
rect 21177 17147 21235 17153
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 19337 17119 19395 17125
rect 19337 17085 19349 17119
rect 19383 17085 19395 17119
rect 19337 17079 19395 17085
rect 19429 17119 19487 17125
rect 19429 17085 19441 17119
rect 19475 17085 19487 17119
rect 22066 17116 22094 17224
rect 23293 17221 23305 17255
rect 23339 17252 23351 17255
rect 23658 17252 23664 17264
rect 23339 17224 23664 17252
rect 23339 17221 23351 17224
rect 23293 17215 23351 17221
rect 23658 17212 23664 17224
rect 23716 17252 23722 17264
rect 24670 17252 24676 17264
rect 23716 17224 24676 17252
rect 23716 17212 23722 17224
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 27080 17252 27108 17283
rect 28258 17280 28264 17332
rect 28316 17320 28322 17332
rect 28721 17323 28779 17329
rect 28721 17320 28733 17323
rect 28316 17292 28733 17320
rect 28316 17280 28322 17292
rect 28721 17289 28733 17292
rect 28767 17289 28779 17323
rect 28721 17283 28779 17289
rect 29454 17280 29460 17332
rect 29512 17280 29518 17332
rect 32125 17323 32183 17329
rect 32125 17289 32137 17323
rect 32171 17320 32183 17323
rect 32398 17320 32404 17332
rect 32171 17292 32404 17320
rect 32171 17289 32183 17292
rect 32125 17283 32183 17289
rect 32398 17280 32404 17292
rect 32456 17280 32462 17332
rect 33594 17280 33600 17332
rect 33652 17280 33658 17332
rect 27586 17255 27644 17261
rect 27586 17252 27598 17255
rect 27080 17224 27598 17252
rect 27586 17221 27598 17224
rect 27632 17221 27644 17255
rect 27586 17215 27644 17221
rect 27706 17212 27712 17264
rect 27764 17212 27770 17264
rect 26418 17144 26424 17196
rect 26476 17144 26482 17196
rect 27249 17187 27307 17193
rect 27249 17153 27261 17187
rect 27295 17184 27307 17187
rect 27724 17184 27752 17212
rect 27295 17156 27752 17184
rect 27295 17153 27307 17156
rect 27249 17147 27307 17153
rect 29638 17144 29644 17196
rect 29696 17144 29702 17196
rect 32490 17144 32496 17196
rect 32548 17144 32554 17196
rect 33965 17187 34023 17193
rect 33965 17153 33977 17187
rect 34011 17184 34023 17187
rect 34422 17184 34428 17196
rect 34011 17156 34428 17184
rect 34011 17153 34023 17156
rect 33965 17147 34023 17153
rect 34422 17144 34428 17156
rect 34480 17144 34486 17196
rect 36446 17144 36452 17196
rect 36504 17144 36510 17196
rect 23385 17119 23443 17125
rect 23385 17116 23397 17119
rect 22066 17088 23397 17116
rect 19429 17079 19487 17085
rect 23385 17085 23397 17088
rect 23431 17116 23443 17119
rect 25130 17116 25136 17128
rect 23431 17088 25136 17116
rect 23431 17085 23443 17088
rect 23385 17079 23443 17085
rect 18230 17008 18236 17060
rect 18288 17048 18294 17060
rect 19352 17048 19380 17079
rect 25130 17076 25136 17088
rect 25188 17076 25194 17128
rect 27341 17119 27399 17125
rect 27341 17085 27353 17119
rect 27387 17085 27399 17119
rect 27341 17079 27399 17085
rect 32585 17119 32643 17125
rect 32585 17085 32597 17119
rect 32631 17116 32643 17119
rect 32674 17116 32680 17128
rect 32631 17088 32680 17116
rect 32631 17085 32643 17088
rect 32585 17079 32643 17085
rect 19794 17048 19800 17060
rect 18288 17020 19800 17048
rect 18288 17008 18294 17020
rect 19794 17008 19800 17020
rect 19852 17008 19858 17060
rect 12584 16952 13584 16980
rect 12584 16940 12590 16952
rect 16390 16940 16396 16992
rect 16448 16940 16454 16992
rect 27356 16980 27384 17079
rect 32674 17076 32680 17088
rect 32732 17076 32738 17128
rect 32769 17119 32827 17125
rect 32769 17085 32781 17119
rect 32815 17085 32827 17119
rect 32769 17079 32827 17085
rect 30282 17008 30288 17060
rect 30340 17048 30346 17060
rect 32784 17048 32812 17079
rect 34054 17076 34060 17128
rect 34112 17076 34118 17128
rect 34241 17119 34299 17125
rect 34241 17085 34253 17119
rect 34287 17116 34299 17119
rect 34330 17116 34336 17128
rect 34287 17088 34336 17116
rect 34287 17085 34299 17088
rect 34241 17079 34299 17085
rect 34256 17048 34284 17079
rect 34330 17076 34336 17088
rect 34388 17076 34394 17128
rect 30340 17020 34284 17048
rect 30340 17008 30346 17020
rect 29178 16980 29184 16992
rect 27356 16952 29184 16980
rect 29178 16940 29184 16952
rect 29236 16940 29242 16992
rect 36170 16940 36176 16992
rect 36228 16980 36234 16992
rect 36265 16983 36323 16989
rect 36265 16980 36277 16983
rect 36228 16952 36277 16980
rect 36228 16940 36234 16952
rect 36265 16949 36277 16952
rect 36311 16949 36323 16983
rect 36265 16943 36323 16949
rect 1104 16890 36800 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 36800 16890
rect 1104 16816 36800 16838
rect 8846 16776 8852 16788
rect 5920 16748 8852 16776
rect 4706 16708 4712 16720
rect 4264 16680 4712 16708
rect 4264 16649 4292 16680
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 4249 16643 4307 16649
rect 4249 16609 4261 16643
rect 4295 16609 4307 16643
rect 4249 16603 4307 16609
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 5258 16640 5264 16652
rect 4479 16612 5264 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 5258 16600 5264 16612
rect 5316 16600 5322 16652
rect 5920 16649 5948 16748
rect 7392 16649 7420 16748
rect 8846 16736 8852 16748
rect 8904 16736 8910 16788
rect 11790 16736 11796 16788
rect 11848 16736 11854 16788
rect 16390 16776 16396 16788
rect 14568 16748 16396 16776
rect 8757 16711 8815 16717
rect 8757 16677 8769 16711
rect 8803 16708 8815 16711
rect 9122 16708 9128 16720
rect 8803 16680 9128 16708
rect 8803 16677 8815 16680
rect 8757 16671 8815 16677
rect 9122 16668 9128 16680
rect 9180 16668 9186 16720
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16609 5963 16643
rect 5905 16603 5963 16609
rect 7377 16643 7435 16649
rect 7377 16609 7389 16643
rect 7423 16609 7435 16643
rect 12713 16643 12771 16649
rect 12713 16640 12725 16643
rect 7377 16603 7435 16609
rect 8956 16612 12725 16640
rect 4798 16532 4804 16584
rect 4856 16532 4862 16584
rect 8386 16532 8392 16584
rect 8444 16572 8450 16584
rect 8956 16581 8984 16612
rect 12713 16609 12725 16612
rect 12759 16640 12771 16643
rect 14568 16640 14596 16748
rect 16390 16736 16396 16748
rect 16448 16736 16454 16788
rect 17218 16736 17224 16788
rect 17276 16736 17282 16788
rect 24872 16748 25820 16776
rect 12759 16612 14596 16640
rect 12759 16609 12771 16612
rect 12713 16603 12771 16609
rect 14826 16600 14832 16652
rect 14884 16640 14890 16652
rect 14921 16643 14979 16649
rect 14921 16640 14933 16643
rect 14884 16612 14933 16640
rect 14884 16600 14890 16612
rect 14921 16609 14933 16612
rect 14967 16609 14979 16643
rect 14921 16603 14979 16609
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 16448 16612 16957 16640
rect 16448 16600 16454 16612
rect 16945 16609 16957 16612
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 22186 16600 22192 16652
rect 22244 16640 22250 16652
rect 23658 16640 23664 16652
rect 22244 16612 23664 16640
rect 22244 16600 22250 16612
rect 23658 16600 23664 16612
rect 23716 16640 23722 16652
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 23716 16612 23765 16640
rect 23716 16600 23722 16612
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 23934 16600 23940 16652
rect 23992 16640 23998 16652
rect 24872 16640 24900 16748
rect 25792 16708 25820 16748
rect 27706 16736 27712 16788
rect 27764 16736 27770 16788
rect 29638 16736 29644 16788
rect 29696 16776 29702 16788
rect 29733 16779 29791 16785
rect 29733 16776 29745 16779
rect 29696 16748 29745 16776
rect 29696 16736 29702 16748
rect 29733 16745 29745 16748
rect 29779 16745 29791 16779
rect 31938 16776 31944 16788
rect 29733 16739 29791 16745
rect 29840 16748 31944 16776
rect 25792 16680 28396 16708
rect 23992 16612 24900 16640
rect 23992 16600 23998 16612
rect 27798 16600 27804 16652
rect 27856 16640 27862 16652
rect 28166 16640 28172 16652
rect 27856 16612 28172 16640
rect 27856 16600 27862 16612
rect 28166 16600 28172 16612
rect 28224 16600 28230 16652
rect 28368 16649 28396 16680
rect 28353 16643 28411 16649
rect 28353 16609 28365 16643
rect 28399 16640 28411 16643
rect 29840 16640 29868 16748
rect 31938 16736 31944 16748
rect 31996 16736 32002 16788
rect 32490 16736 32496 16788
rect 32548 16776 32554 16788
rect 32953 16779 33011 16785
rect 32953 16776 32965 16779
rect 32548 16748 32965 16776
rect 32548 16736 32554 16748
rect 32953 16745 32965 16748
rect 32999 16745 33011 16779
rect 34146 16776 34152 16788
rect 32953 16739 33011 16745
rect 33152 16748 34152 16776
rect 30098 16668 30104 16720
rect 30156 16708 30162 16720
rect 30156 16680 31064 16708
rect 30156 16668 30162 16680
rect 28399 16612 29868 16640
rect 28399 16609 28411 16612
rect 28353 16603 28411 16609
rect 30282 16600 30288 16652
rect 30340 16600 30346 16652
rect 31036 16649 31064 16680
rect 31021 16643 31079 16649
rect 31021 16609 31033 16643
rect 31067 16609 31079 16643
rect 31021 16603 31079 16609
rect 31110 16600 31116 16652
rect 31168 16600 31174 16652
rect 31570 16600 31576 16652
rect 31628 16640 31634 16652
rect 33152 16649 33180 16748
rect 34146 16736 34152 16748
rect 34204 16736 34210 16788
rect 34422 16736 34428 16788
rect 34480 16776 34486 16788
rect 34517 16779 34575 16785
rect 34517 16776 34529 16779
rect 34480 16748 34529 16776
rect 34480 16736 34486 16748
rect 34517 16745 34529 16748
rect 34563 16745 34575 16779
rect 34517 16739 34575 16745
rect 33137 16643 33195 16649
rect 33137 16640 33149 16643
rect 31628 16612 31708 16640
rect 31628 16600 31634 16612
rect 8941 16575 8999 16581
rect 8941 16572 8953 16575
rect 8444 16544 8953 16572
rect 8444 16532 8450 16544
rect 8941 16541 8953 16544
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 9122 16532 9128 16584
rect 9180 16532 9186 16584
rect 11977 16575 12035 16581
rect 11977 16541 11989 16575
rect 12023 16572 12035 16575
rect 12437 16575 12495 16581
rect 12023 16544 12112 16572
rect 12023 16541 12035 16544
rect 11977 16535 12035 16541
rect 5442 16504 5448 16516
rect 4172 16476 5448 16504
rect 4172 16448 4200 16476
rect 5442 16464 5448 16476
rect 5500 16464 5506 16516
rect 6172 16507 6230 16513
rect 6172 16473 6184 16507
rect 6218 16504 6230 16507
rect 6362 16504 6368 16516
rect 6218 16476 6368 16504
rect 6218 16473 6230 16476
rect 6172 16467 6230 16473
rect 6362 16464 6368 16476
rect 6420 16464 6426 16516
rect 7644 16507 7702 16513
rect 7644 16473 7656 16507
rect 7690 16504 7702 16507
rect 8018 16504 8024 16516
rect 7690 16476 8024 16504
rect 7690 16473 7702 16476
rect 7644 16467 7702 16473
rect 8018 16464 8024 16476
rect 8076 16464 8082 16516
rect 3050 16396 3056 16448
rect 3108 16436 3114 16448
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 3108 16408 3801 16436
rect 3108 16396 3114 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 4154 16396 4160 16448
rect 4212 16396 4218 16448
rect 4614 16396 4620 16448
rect 4672 16396 4678 16448
rect 6822 16396 6828 16448
rect 6880 16436 6886 16448
rect 7285 16439 7343 16445
rect 7285 16436 7297 16439
rect 6880 16408 7297 16436
rect 6880 16396 6886 16408
rect 7285 16405 7297 16408
rect 7331 16405 7343 16439
rect 7285 16399 7343 16405
rect 9030 16396 9036 16448
rect 9088 16396 9094 16448
rect 12084 16445 12112 16544
rect 12437 16541 12449 16575
rect 12483 16572 12495 16575
rect 13170 16572 13176 16584
rect 12483 16544 13176 16572
rect 12483 16541 12495 16544
rect 12437 16535 12495 16541
rect 13170 16532 13176 16544
rect 13228 16532 13234 16584
rect 17034 16532 17040 16584
rect 17092 16572 17098 16584
rect 17405 16575 17463 16581
rect 17405 16572 17417 16575
rect 17092 16544 17417 16572
rect 17092 16532 17098 16544
rect 17405 16541 17417 16544
rect 17451 16541 17463 16575
rect 17405 16535 17463 16541
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 24854 16572 24860 16584
rect 20864 16544 24860 16572
rect 20864 16532 20870 16544
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 28077 16575 28135 16581
rect 28077 16541 28089 16575
rect 28123 16572 28135 16575
rect 28258 16572 28264 16584
rect 28123 16544 28264 16572
rect 28123 16541 28135 16544
rect 28077 16535 28135 16541
rect 28258 16532 28264 16544
rect 28316 16532 28322 16584
rect 29546 16532 29552 16584
rect 29604 16572 29610 16584
rect 30300 16572 30328 16600
rect 29604 16544 30328 16572
rect 31680 16572 31708 16612
rect 32600 16612 33149 16640
rect 32600 16572 32628 16612
rect 33137 16609 33149 16612
rect 33183 16609 33195 16643
rect 33137 16603 33195 16609
rect 31680 16544 32628 16572
rect 29604 16532 29610 16544
rect 33778 16532 33784 16584
rect 33836 16572 33842 16584
rect 34885 16575 34943 16581
rect 34885 16572 34897 16575
rect 33836 16544 34897 16572
rect 33836 16532 33842 16544
rect 34885 16541 34897 16544
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 15188 16507 15246 16513
rect 15188 16473 15200 16507
rect 15234 16504 15246 16507
rect 15286 16504 15292 16516
rect 15234 16476 15292 16504
rect 15234 16473 15246 16476
rect 15188 16467 15246 16473
rect 15286 16464 15292 16476
rect 15344 16464 15350 16516
rect 16761 16507 16819 16513
rect 16761 16504 16773 16507
rect 16316 16476 16773 16504
rect 12069 16439 12127 16445
rect 12069 16405 12081 16439
rect 12115 16405 12127 16439
rect 12069 16399 12127 16405
rect 12529 16439 12587 16445
rect 12529 16405 12541 16439
rect 12575 16436 12587 16439
rect 13354 16436 13360 16448
rect 12575 16408 13360 16436
rect 12575 16405 12587 16408
rect 12529 16399 12587 16405
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 16316 16445 16344 16476
rect 16761 16473 16773 16476
rect 16807 16504 16819 16507
rect 17310 16504 17316 16516
rect 16807 16476 17316 16504
rect 16807 16473 16819 16476
rect 16761 16467 16819 16473
rect 17310 16464 17316 16476
rect 17368 16464 17374 16516
rect 23658 16464 23664 16516
rect 23716 16464 23722 16516
rect 25124 16507 25182 16513
rect 25124 16473 25136 16507
rect 25170 16504 25182 16507
rect 26326 16504 26332 16516
rect 25170 16476 26332 16504
rect 25170 16473 25182 16476
rect 25124 16467 25182 16473
rect 26326 16464 26332 16476
rect 26384 16464 26390 16516
rect 30190 16464 30196 16516
rect 30248 16504 30254 16516
rect 31846 16513 31852 16516
rect 30929 16507 30987 16513
rect 30929 16504 30941 16507
rect 30248 16476 30941 16504
rect 30248 16464 30254 16476
rect 30929 16473 30941 16476
rect 30975 16473 30987 16507
rect 30929 16467 30987 16473
rect 31840 16467 31852 16513
rect 31846 16464 31852 16467
rect 31904 16464 31910 16516
rect 33404 16507 33462 16513
rect 33404 16473 33416 16507
rect 33450 16504 33462 16507
rect 33450 16476 34744 16504
rect 33450 16473 33462 16476
rect 33404 16467 33462 16473
rect 16301 16439 16359 16445
rect 16301 16405 16313 16439
rect 16347 16405 16359 16439
rect 16301 16399 16359 16405
rect 16390 16396 16396 16448
rect 16448 16396 16454 16448
rect 16853 16439 16911 16445
rect 16853 16405 16865 16439
rect 16899 16436 16911 16439
rect 16942 16436 16948 16448
rect 16899 16408 16948 16436
rect 16899 16405 16911 16408
rect 16853 16399 16911 16405
rect 16942 16396 16948 16408
rect 17000 16396 17006 16448
rect 22830 16396 22836 16448
rect 22888 16436 22894 16448
rect 23293 16439 23351 16445
rect 23293 16436 23305 16439
rect 22888 16408 23305 16436
rect 22888 16396 22894 16408
rect 23293 16405 23305 16408
rect 23339 16405 23351 16439
rect 23293 16399 23351 16405
rect 26050 16396 26056 16448
rect 26108 16436 26114 16448
rect 26237 16439 26295 16445
rect 26237 16436 26249 16439
rect 26108 16408 26249 16436
rect 26108 16396 26114 16408
rect 26237 16405 26249 16408
rect 26283 16405 26295 16439
rect 26237 16399 26295 16405
rect 30098 16396 30104 16448
rect 30156 16396 30162 16448
rect 30558 16396 30564 16448
rect 30616 16396 30622 16448
rect 34716 16445 34744 16476
rect 34701 16439 34759 16445
rect 34701 16405 34713 16439
rect 34747 16405 34759 16439
rect 34701 16399 34759 16405
rect 1104 16346 36800 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 36800 16346
rect 1104 16272 36800 16294
rect 3789 16235 3847 16241
rect 3789 16201 3801 16235
rect 3835 16232 3847 16235
rect 4154 16232 4160 16244
rect 3835 16204 4160 16232
rect 3835 16201 3847 16204
rect 3789 16195 3847 16201
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 6362 16192 6368 16244
rect 6420 16192 6426 16244
rect 7834 16192 7840 16244
rect 7892 16232 7898 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 7892 16204 8217 16232
rect 7892 16192 7898 16204
rect 8205 16201 8217 16204
rect 8251 16232 8263 16235
rect 9214 16232 9220 16244
rect 8251 16204 9220 16232
rect 8251 16201 8263 16204
rect 8205 16195 8263 16201
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 10229 16235 10287 16241
rect 10229 16201 10241 16235
rect 10275 16232 10287 16235
rect 10318 16232 10324 16244
rect 10275 16204 10324 16232
rect 10275 16201 10287 16204
rect 10229 16195 10287 16201
rect 10318 16192 10324 16204
rect 10376 16192 10382 16244
rect 12253 16235 12311 16241
rect 12253 16201 12265 16235
rect 12299 16232 12311 16235
rect 12299 16204 12434 16232
rect 12299 16201 12311 16204
rect 12253 16195 12311 16201
rect 2774 16164 2780 16176
rect 2424 16136 2780 16164
rect 1397 16099 1455 16105
rect 1397 16065 1409 16099
rect 1443 16096 1455 16099
rect 1854 16096 1860 16108
rect 1443 16068 1860 16096
rect 1443 16065 1455 16068
rect 1397 16059 1455 16065
rect 1854 16056 1860 16068
rect 1912 16056 1918 16108
rect 2424 16105 2452 16136
rect 2774 16124 2780 16136
rect 2832 16164 2838 16176
rect 4614 16173 4620 16176
rect 4608 16164 4620 16173
rect 2832 16136 4384 16164
rect 4575 16136 4620 16164
rect 2832 16124 2838 16136
rect 2682 16105 2688 16108
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16065 2467 16099
rect 2409 16059 2467 16065
rect 2676 16059 2688 16105
rect 2682 16056 2688 16059
rect 2740 16056 2746 16108
rect 4356 16105 4384 16136
rect 4608 16127 4620 16136
rect 4614 16124 4620 16127
rect 4672 16124 4678 16176
rect 8021 16167 8079 16173
rect 8021 16133 8033 16167
rect 8067 16164 8079 16167
rect 9030 16164 9036 16176
rect 8067 16136 9036 16164
rect 8067 16133 8079 16136
rect 8021 16127 8079 16133
rect 9030 16124 9036 16136
rect 9088 16124 9094 16176
rect 10336 16164 10364 16192
rect 12406 16164 12434 16204
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 13909 16235 13967 16241
rect 13909 16232 13921 16235
rect 13872 16204 13921 16232
rect 13872 16192 13878 16204
rect 13909 16201 13921 16204
rect 13955 16201 13967 16235
rect 13909 16195 13967 16201
rect 15286 16192 15292 16244
rect 15344 16192 15350 16244
rect 19610 16192 19616 16244
rect 19668 16232 19674 16244
rect 19797 16235 19855 16241
rect 19797 16232 19809 16235
rect 19668 16204 19809 16232
rect 19668 16192 19674 16204
rect 19797 16201 19809 16204
rect 19843 16232 19855 16235
rect 20254 16232 20260 16244
rect 19843 16204 20260 16232
rect 19843 16201 19855 16204
rect 19797 16195 19855 16201
rect 20254 16192 20260 16204
rect 20312 16192 20318 16244
rect 21542 16192 21548 16244
rect 21600 16192 21606 16244
rect 22649 16235 22707 16241
rect 22649 16201 22661 16235
rect 22695 16201 22707 16235
rect 22649 16195 22707 16201
rect 12774 16167 12832 16173
rect 12774 16164 12786 16167
rect 10336 16136 10548 16164
rect 12406 16136 12786 16164
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 8297 16099 8355 16105
rect 8297 16065 8309 16099
rect 8343 16096 8355 16099
rect 8386 16096 8392 16108
rect 8343 16068 8392 16096
rect 8343 16065 8355 16068
rect 8297 16059 8355 16065
rect 8386 16056 8392 16068
rect 8444 16056 8450 16108
rect 8846 16056 8852 16108
rect 8904 16056 8910 16108
rect 9122 16105 9128 16108
rect 9116 16096 9128 16105
rect 9083 16068 9128 16096
rect 9116 16059 9128 16068
rect 9122 16056 9128 16059
rect 9180 16056 9186 16108
rect 10226 16056 10232 16108
rect 10284 16096 10290 16108
rect 10520 16105 10548 16136
rect 12774 16133 12786 16136
rect 12820 16133 12832 16167
rect 19242 16164 19248 16176
rect 12774 16127 12832 16133
rect 18432 16136 19248 16164
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 10284 16068 10333 16096
rect 10284 16056 10290 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 10505 16099 10563 16105
rect 10505 16065 10517 16099
rect 10551 16065 10563 16099
rect 10505 16059 10563 16065
rect 12434 16056 12440 16108
rect 12492 16056 12498 16108
rect 12526 16056 12532 16108
rect 12584 16056 12590 16108
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16096 15531 16099
rect 16390 16096 16396 16108
rect 15519 16068 16396 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 17586 16056 17592 16108
rect 17644 16056 17650 16108
rect 18432 16105 18460 16136
rect 19242 16124 19248 16136
rect 19300 16164 19306 16176
rect 22664 16164 22692 16195
rect 23750 16192 23756 16244
rect 23808 16232 23814 16244
rect 24305 16235 24363 16241
rect 24305 16232 24317 16235
rect 23808 16204 24317 16232
rect 23808 16192 23814 16204
rect 24305 16201 24317 16204
rect 24351 16201 24363 16235
rect 24305 16195 24363 16201
rect 24854 16192 24860 16244
rect 24912 16232 24918 16244
rect 25777 16235 25835 16241
rect 25777 16232 25789 16235
rect 24912 16204 25789 16232
rect 24912 16192 24918 16204
rect 25777 16201 25789 16204
rect 25823 16201 25835 16235
rect 25777 16195 25835 16201
rect 25866 16192 25872 16244
rect 25924 16192 25930 16244
rect 26326 16192 26332 16244
rect 26384 16192 26390 16244
rect 28905 16235 28963 16241
rect 28905 16201 28917 16235
rect 28951 16201 28963 16235
rect 28905 16195 28963 16201
rect 23170 16167 23228 16173
rect 23170 16164 23182 16167
rect 19300 16136 20029 16164
rect 22664 16136 23182 16164
rect 19300 16124 19306 16136
rect 18690 16105 18696 16108
rect 18417 16099 18475 16105
rect 18417 16065 18429 16099
rect 18463 16065 18475 16099
rect 18417 16059 18475 16065
rect 18684 16059 18696 16105
rect 18690 16056 18696 16059
rect 18748 16056 18754 16108
rect 20001 16028 20029 16136
rect 23170 16133 23182 16136
rect 23216 16133 23228 16167
rect 23170 16127 23228 16133
rect 25685 16167 25743 16173
rect 25685 16133 25697 16167
rect 25731 16164 25743 16167
rect 25884 16164 25912 16192
rect 26142 16164 26148 16176
rect 25731 16136 26148 16164
rect 25731 16133 25743 16136
rect 25685 16127 25743 16133
rect 26142 16124 26148 16136
rect 26200 16124 26206 16176
rect 28920 16164 28948 16195
rect 30098 16192 30104 16244
rect 30156 16232 30162 16244
rect 30561 16235 30619 16241
rect 30561 16232 30573 16235
rect 30156 16204 30573 16232
rect 30156 16192 30162 16204
rect 30561 16201 30573 16204
rect 30607 16201 30619 16235
rect 30561 16195 30619 16201
rect 31757 16235 31815 16241
rect 31757 16201 31769 16235
rect 31803 16232 31815 16235
rect 31846 16232 31852 16244
rect 31803 16204 31852 16232
rect 31803 16201 31815 16204
rect 31757 16195 31815 16201
rect 31846 16192 31852 16204
rect 31904 16192 31910 16244
rect 32125 16235 32183 16241
rect 32125 16201 32137 16235
rect 32171 16201 32183 16235
rect 32125 16195 32183 16201
rect 29426 16167 29484 16173
rect 29426 16164 29438 16167
rect 28920 16136 29438 16164
rect 29426 16133 29438 16136
rect 29472 16133 29484 16167
rect 29426 16127 29484 16133
rect 20070 16056 20076 16108
rect 20128 16096 20134 16108
rect 20421 16099 20479 16105
rect 20421 16096 20433 16099
rect 20128 16068 20433 16096
rect 20128 16056 20134 16068
rect 20421 16065 20433 16068
rect 20467 16065 20479 16099
rect 20421 16059 20479 16065
rect 22830 16056 22836 16108
rect 22888 16056 22894 16108
rect 25866 16056 25872 16108
rect 25924 16096 25930 16108
rect 25961 16099 26019 16105
rect 25961 16096 25973 16099
rect 25924 16068 25973 16096
rect 25924 16056 25930 16068
rect 25961 16065 25973 16068
rect 26007 16065 26019 16099
rect 25961 16059 26019 16065
rect 26513 16099 26571 16105
rect 26513 16065 26525 16099
rect 26559 16096 26571 16099
rect 26970 16096 26976 16108
rect 26559 16068 26976 16096
rect 26559 16065 26571 16068
rect 26513 16059 26571 16065
rect 26970 16056 26976 16068
rect 27028 16056 27034 16108
rect 29089 16099 29147 16105
rect 29089 16065 29101 16099
rect 29135 16096 29147 16099
rect 29730 16096 29736 16108
rect 29135 16068 29736 16096
rect 29135 16065 29147 16068
rect 29089 16059 29147 16065
rect 29730 16056 29736 16068
rect 29788 16056 29794 16108
rect 31941 16099 31999 16105
rect 31941 16065 31953 16099
rect 31987 16096 31999 16099
rect 32140 16096 32168 16195
rect 32490 16192 32496 16244
rect 32548 16192 32554 16244
rect 32582 16192 32588 16244
rect 32640 16232 32646 16244
rect 32953 16235 33011 16241
rect 32953 16232 32965 16235
rect 32640 16204 32965 16232
rect 32640 16192 32646 16204
rect 32953 16201 32965 16204
rect 32999 16201 33011 16235
rect 32953 16195 33011 16201
rect 33778 16192 33784 16244
rect 33836 16192 33842 16244
rect 34149 16235 34207 16241
rect 34149 16201 34161 16235
rect 34195 16232 34207 16235
rect 34422 16232 34428 16244
rect 34195 16204 34428 16232
rect 34195 16201 34207 16204
rect 34149 16195 34207 16201
rect 34422 16192 34428 16204
rect 34480 16192 34486 16244
rect 33413 16167 33471 16173
rect 33413 16133 33425 16167
rect 33459 16164 33471 16167
rect 33502 16164 33508 16176
rect 33459 16136 33508 16164
rect 33459 16133 33471 16136
rect 33413 16127 33471 16133
rect 33502 16124 33508 16136
rect 33560 16124 33566 16176
rect 34054 16124 34060 16176
rect 34112 16164 34118 16176
rect 34241 16167 34299 16173
rect 34241 16164 34253 16167
rect 34112 16136 34253 16164
rect 34112 16124 34118 16136
rect 34241 16133 34253 16136
rect 34287 16133 34299 16167
rect 34241 16127 34299 16133
rect 33321 16099 33379 16105
rect 33321 16096 33333 16099
rect 31987 16068 32168 16096
rect 32600 16068 33333 16096
rect 31987 16065 31999 16068
rect 31941 16059 31999 16065
rect 32600 16040 32628 16068
rect 33321 16065 33333 16068
rect 33367 16065 33379 16099
rect 33321 16059 33379 16065
rect 20165 16031 20223 16037
rect 20165 16028 20177 16031
rect 20001 16000 20177 16028
rect 20165 15997 20177 16000
rect 20211 15997 20223 16031
rect 20165 15991 20223 15997
rect 8018 15920 8024 15972
rect 8076 15920 8082 15972
rect 934 15852 940 15904
rect 992 15892 998 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 992 15864 1593 15892
rect 992 15852 998 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 1581 15855 1639 15861
rect 5718 15852 5724 15904
rect 5776 15892 5782 15904
rect 7006 15892 7012 15904
rect 5776 15864 7012 15892
rect 5776 15852 5782 15864
rect 7006 15852 7012 15864
rect 7064 15852 7070 15904
rect 10318 15852 10324 15904
rect 10376 15852 10382 15904
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 12710 15892 12716 15904
rect 10560 15864 12716 15892
rect 10560 15852 10566 15864
rect 12710 15852 12716 15864
rect 12768 15892 12774 15904
rect 15470 15892 15476 15904
rect 12768 15864 15476 15892
rect 12768 15852 12774 15864
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 16758 15852 16764 15904
rect 16816 15892 16822 15904
rect 17773 15895 17831 15901
rect 17773 15892 17785 15895
rect 16816 15864 17785 15892
rect 16816 15852 16822 15864
rect 17773 15861 17785 15864
rect 17819 15861 17831 15895
rect 20180 15892 20208 15991
rect 22646 15988 22652 16040
rect 22704 16028 22710 16040
rect 22925 16031 22983 16037
rect 22925 16028 22937 16031
rect 22704 16000 22937 16028
rect 22704 15988 22710 16000
rect 22925 15997 22937 16000
rect 22971 15997 22983 16031
rect 22925 15991 22983 15997
rect 29178 15988 29184 16040
rect 29236 15988 29242 16040
rect 32582 15988 32588 16040
rect 32640 15988 32646 16040
rect 32674 15988 32680 16040
rect 32732 15988 32738 16040
rect 33597 16031 33655 16037
rect 33597 15997 33609 16031
rect 33643 16028 33655 16031
rect 33686 16028 33692 16040
rect 33643 16000 33692 16028
rect 33643 15997 33655 16000
rect 33597 15991 33655 15997
rect 33612 15960 33640 15991
rect 33686 15988 33692 16000
rect 33744 15988 33750 16040
rect 34330 15988 34336 16040
rect 34388 15988 34394 16040
rect 31726 15932 33640 15960
rect 20806 15892 20812 15904
rect 20180 15864 20812 15892
rect 17773 15855 17831 15861
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 25406 15852 25412 15904
rect 25464 15892 25470 15904
rect 26145 15895 26203 15901
rect 26145 15892 26157 15895
rect 25464 15864 26157 15892
rect 25464 15852 25470 15864
rect 26145 15861 26157 15864
rect 26191 15861 26203 15895
rect 26145 15855 26203 15861
rect 28442 15852 28448 15904
rect 28500 15892 28506 15904
rect 31110 15892 31116 15904
rect 28500 15864 31116 15892
rect 28500 15852 28506 15864
rect 31110 15852 31116 15864
rect 31168 15892 31174 15904
rect 31726 15892 31754 15932
rect 31168 15864 31754 15892
rect 31168 15852 31174 15864
rect 1104 15802 36800 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 36800 15802
rect 1104 15728 36800 15750
rect 2682 15648 2688 15700
rect 2740 15688 2746 15700
rect 2869 15691 2927 15697
rect 2869 15688 2881 15691
rect 2740 15660 2881 15688
rect 2740 15648 2746 15660
rect 2869 15657 2881 15660
rect 2915 15657 2927 15691
rect 2869 15651 2927 15657
rect 4798 15648 4804 15700
rect 4856 15648 4862 15700
rect 9033 15691 9091 15697
rect 9033 15657 9045 15691
rect 9079 15688 9091 15691
rect 9122 15688 9128 15700
rect 9079 15660 9128 15688
rect 9079 15657 9091 15660
rect 9033 15651 9091 15657
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 12897 15691 12955 15697
rect 12897 15688 12909 15691
rect 12492 15660 12909 15688
rect 12492 15648 12498 15660
rect 12897 15657 12909 15660
rect 12943 15657 12955 15691
rect 12897 15651 12955 15657
rect 18690 15648 18696 15700
rect 18748 15648 18754 15700
rect 20070 15648 20076 15700
rect 20128 15648 20134 15700
rect 22097 15691 22155 15697
rect 20548 15660 21772 15688
rect 16117 15623 16175 15629
rect 16117 15589 16129 15623
rect 16163 15620 16175 15623
rect 16850 15620 16856 15632
rect 16163 15592 16856 15620
rect 16163 15589 16175 15592
rect 16117 15583 16175 15589
rect 16850 15580 16856 15592
rect 16908 15580 16914 15632
rect 20548 15620 20576 15660
rect 20714 15620 20720 15632
rect 19812 15592 20576 15620
rect 20640 15592 20720 15620
rect 5258 15512 5264 15564
rect 5316 15552 5322 15564
rect 5353 15555 5411 15561
rect 5353 15552 5365 15555
rect 5316 15524 5365 15552
rect 5316 15512 5322 15524
rect 5353 15521 5365 15524
rect 5399 15521 5411 15555
rect 10318 15552 10324 15564
rect 5353 15515 5411 15521
rect 9048 15524 10324 15552
rect 3050 15444 3056 15496
rect 3108 15444 3114 15496
rect 5169 15487 5227 15493
rect 5169 15453 5181 15487
rect 5215 15484 5227 15487
rect 5718 15484 5724 15496
rect 5215 15456 5724 15484
rect 5215 15453 5227 15456
rect 5169 15447 5227 15453
rect 5718 15444 5724 15456
rect 5776 15444 5782 15496
rect 9048 15493 9076 15524
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 13541 15555 13599 15561
rect 13541 15552 13553 15555
rect 12406 15524 13553 15552
rect 9033 15487 9091 15493
rect 9033 15453 9045 15487
rect 9079 15453 9091 15487
rect 9033 15447 9091 15453
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15484 9367 15487
rect 10226 15484 10232 15496
rect 9355 15456 10232 15484
rect 9355 15453 9367 15456
rect 9309 15447 9367 15453
rect 7742 15376 7748 15428
rect 7800 15416 7806 15428
rect 9324 15416 9352 15447
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 10502 15444 10508 15496
rect 10560 15444 10566 15496
rect 10778 15444 10784 15496
rect 10836 15444 10842 15496
rect 7800 15388 9352 15416
rect 10244 15416 10272 15444
rect 12406 15416 12434 15524
rect 13541 15521 13553 15524
rect 13587 15552 13599 15555
rect 16758 15552 16764 15564
rect 13587 15524 16764 15552
rect 13587 15521 13599 15524
rect 13541 15515 13599 15521
rect 16758 15512 16764 15524
rect 16816 15512 16822 15564
rect 17586 15512 17592 15564
rect 17644 15552 17650 15564
rect 19812 15561 19840 15592
rect 19797 15555 19855 15561
rect 19797 15552 19809 15555
rect 17644 15524 19809 15552
rect 17644 15512 17650 15524
rect 19797 15521 19809 15524
rect 19843 15521 19855 15555
rect 19797 15515 19855 15521
rect 13265 15487 13323 15493
rect 13265 15453 13277 15487
rect 13311 15484 13323 15487
rect 13814 15484 13820 15496
rect 13311 15456 13820 15484
rect 13311 15453 13323 15456
rect 13265 15447 13323 15453
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15484 18935 15487
rect 18923 15456 19288 15484
rect 18923 15453 18935 15456
rect 18877 15447 18935 15453
rect 10244 15388 12434 15416
rect 7800 15376 7806 15388
rect 13354 15376 13360 15428
rect 13412 15416 13418 15428
rect 18966 15416 18972 15428
rect 13412 15388 18972 15416
rect 13412 15376 13418 15388
rect 18966 15376 18972 15388
rect 19024 15376 19030 15428
rect 5261 15351 5319 15357
rect 5261 15317 5273 15351
rect 5307 15348 5319 15351
rect 5994 15348 6000 15360
rect 5307 15320 6000 15348
rect 5307 15317 5319 15320
rect 5261 15311 5319 15317
rect 5994 15308 6000 15320
rect 6052 15348 6058 15360
rect 6638 15348 6644 15360
rect 6052 15320 6644 15348
rect 6052 15308 6058 15320
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 9214 15308 9220 15360
rect 9272 15308 9278 15360
rect 11517 15351 11575 15357
rect 11517 15317 11529 15351
rect 11563 15348 11575 15351
rect 12158 15348 12164 15360
rect 11563 15320 12164 15348
rect 11563 15317 11575 15320
rect 11517 15311 11575 15317
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 16482 15308 16488 15360
rect 16540 15308 16546 15360
rect 16577 15351 16635 15357
rect 16577 15317 16589 15351
rect 16623 15348 16635 15351
rect 16942 15348 16948 15360
rect 16623 15320 16948 15348
rect 16623 15317 16635 15320
rect 16577 15311 16635 15317
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 19260 15357 19288 15456
rect 19610 15444 19616 15496
rect 19668 15444 19674 15496
rect 20254 15444 20260 15496
rect 20312 15444 20318 15496
rect 20640 15493 20668 15592
rect 20714 15580 20720 15592
rect 20772 15580 20778 15632
rect 21744 15552 21772 15660
rect 22097 15657 22109 15691
rect 22143 15688 22155 15691
rect 22554 15688 22560 15700
rect 22143 15660 22560 15688
rect 22143 15657 22155 15660
rect 22097 15651 22155 15657
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 23382 15648 23388 15700
rect 23440 15688 23446 15700
rect 23661 15691 23719 15697
rect 23661 15688 23673 15691
rect 23440 15660 23673 15688
rect 23440 15648 23446 15660
rect 23661 15657 23673 15660
rect 23707 15657 23719 15691
rect 23661 15651 23719 15657
rect 26970 15648 26976 15700
rect 27028 15648 27034 15700
rect 28813 15691 28871 15697
rect 28813 15688 28825 15691
rect 27540 15660 28825 15688
rect 21744 15524 22416 15552
rect 20625 15487 20683 15493
rect 20625 15453 20637 15487
rect 20671 15453 20683 15487
rect 20625 15447 20683 15453
rect 20717 15487 20775 15493
rect 20717 15453 20729 15487
rect 20763 15484 20775 15487
rect 20806 15484 20812 15496
rect 20763 15456 20812 15484
rect 20763 15453 20775 15456
rect 20717 15447 20775 15453
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 22281 15487 22339 15493
rect 22281 15484 22293 15487
rect 22152 15456 22293 15484
rect 22152 15444 22158 15456
rect 22281 15453 22293 15456
rect 22327 15453 22339 15487
rect 22388 15484 22416 15524
rect 27246 15512 27252 15564
rect 27304 15552 27310 15564
rect 27540 15561 27568 15660
rect 28813 15657 28825 15660
rect 28859 15688 28871 15691
rect 29546 15688 29552 15700
rect 28859 15660 29552 15688
rect 28859 15657 28871 15660
rect 28813 15651 28871 15657
rect 29546 15648 29552 15660
rect 29604 15648 29610 15700
rect 29730 15648 29736 15700
rect 29788 15648 29794 15700
rect 27801 15623 27859 15629
rect 27801 15589 27813 15623
rect 27847 15620 27859 15623
rect 33410 15620 33416 15632
rect 27847 15592 33416 15620
rect 27847 15589 27859 15592
rect 27801 15583 27859 15589
rect 33410 15580 33416 15592
rect 33468 15580 33474 15632
rect 27525 15555 27583 15561
rect 27525 15552 27537 15555
rect 27304 15524 27537 15552
rect 27304 15512 27310 15524
rect 27525 15521 27537 15524
rect 27571 15521 27583 15555
rect 27525 15515 27583 15521
rect 28442 15512 28448 15564
rect 28500 15512 28506 15564
rect 30190 15512 30196 15564
rect 30248 15512 30254 15564
rect 30285 15555 30343 15561
rect 30285 15521 30297 15555
rect 30331 15552 30343 15555
rect 32674 15552 32680 15564
rect 30331 15524 32680 15552
rect 30331 15521 30343 15524
rect 30285 15515 30343 15521
rect 23934 15484 23940 15496
rect 22388 15456 23940 15484
rect 22281 15447 22339 15453
rect 23934 15444 23940 15456
rect 23992 15444 23998 15496
rect 24486 15444 24492 15496
rect 24544 15484 24550 15496
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 24544 15456 24593 15484
rect 24544 15444 24550 15456
rect 24581 15453 24593 15456
rect 24627 15484 24639 15487
rect 26142 15484 26148 15496
rect 24627 15456 26148 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 26142 15444 26148 15456
rect 26200 15444 26206 15496
rect 27341 15487 27399 15493
rect 27341 15453 27353 15487
rect 27387 15484 27399 15487
rect 27430 15484 27436 15496
rect 27387 15456 27436 15484
rect 27387 15453 27399 15456
rect 27341 15447 27399 15453
rect 27430 15444 27436 15456
rect 27488 15444 27494 15496
rect 19705 15419 19763 15425
rect 19705 15385 19717 15419
rect 19751 15416 19763 15419
rect 19794 15416 19800 15428
rect 19751 15388 19800 15416
rect 19751 15385 19763 15388
rect 19705 15379 19763 15385
rect 19794 15376 19800 15388
rect 19852 15376 19858 15428
rect 20962 15419 21020 15425
rect 20962 15416 20974 15419
rect 20456 15388 20974 15416
rect 20456 15357 20484 15388
rect 20962 15385 20974 15388
rect 21008 15385 21020 15419
rect 20962 15379 21020 15385
rect 22370 15376 22376 15428
rect 22428 15416 22434 15428
rect 22526 15419 22584 15425
rect 22526 15416 22538 15419
rect 22428 15388 22538 15416
rect 22428 15376 22434 15388
rect 22526 15385 22538 15388
rect 22572 15385 22584 15419
rect 22526 15379 22584 15385
rect 24848 15419 24906 15425
rect 24848 15385 24860 15419
rect 24894 15416 24906 15419
rect 25130 15416 25136 15428
rect 24894 15388 25136 15416
rect 24894 15385 24906 15388
rect 24848 15379 24906 15385
rect 25130 15376 25136 15388
rect 25188 15376 25194 15428
rect 28460 15416 28488 15512
rect 28626 15444 28632 15496
rect 28684 15444 28690 15496
rect 30098 15444 30104 15496
rect 30156 15444 30162 15496
rect 30300 15484 30328 15515
rect 32674 15512 32680 15524
rect 32732 15512 32738 15564
rect 30208 15456 30328 15484
rect 25240 15388 28488 15416
rect 28644 15416 28672 15444
rect 30208 15416 30236 15456
rect 28644 15388 30236 15416
rect 19245 15351 19303 15357
rect 19245 15317 19257 15351
rect 19291 15317 19303 15351
rect 19245 15311 19303 15317
rect 20441 15351 20499 15357
rect 20441 15317 20453 15351
rect 20487 15317 20499 15351
rect 20441 15311 20499 15317
rect 24394 15308 24400 15360
rect 24452 15348 24458 15360
rect 25240 15348 25268 15388
rect 24452 15320 25268 15348
rect 24452 15308 24458 15320
rect 25866 15308 25872 15360
rect 25924 15348 25930 15360
rect 25961 15351 26019 15357
rect 25961 15348 25973 15351
rect 25924 15320 25973 15348
rect 25924 15308 25930 15320
rect 25961 15317 25973 15320
rect 26007 15317 26019 15351
rect 25961 15311 26019 15317
rect 27433 15351 27491 15357
rect 27433 15317 27445 15351
rect 27479 15348 27491 15351
rect 27522 15348 27528 15360
rect 27479 15320 27528 15348
rect 27479 15317 27491 15320
rect 27433 15311 27491 15317
rect 27522 15308 27528 15320
rect 27580 15348 27586 15360
rect 28169 15351 28227 15357
rect 28169 15348 28181 15351
rect 27580 15320 28181 15348
rect 27580 15308 27586 15320
rect 28169 15317 28181 15320
rect 28215 15317 28227 15351
rect 28169 15311 28227 15317
rect 28258 15308 28264 15360
rect 28316 15308 28322 15360
rect 1104 15258 36800 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 36800 15258
rect 1104 15184 36800 15206
rect 6365 15147 6423 15153
rect 6365 15113 6377 15147
rect 6411 15113 6423 15147
rect 6365 15107 6423 15113
rect 6733 15147 6791 15153
rect 6733 15113 6745 15147
rect 6779 15144 6791 15147
rect 6914 15144 6920 15156
rect 6779 15116 6920 15144
rect 6779 15113 6791 15116
rect 6733 15107 6791 15113
rect 4433 15079 4491 15085
rect 4433 15045 4445 15079
rect 4479 15076 4491 15079
rect 4614 15076 4620 15088
rect 4479 15048 4620 15076
rect 4479 15045 4491 15048
rect 4433 15039 4491 15045
rect 4614 15036 4620 15048
rect 4672 15076 4678 15088
rect 5350 15076 5356 15088
rect 4672 15048 5356 15076
rect 4672 15036 4678 15048
rect 5350 15036 5356 15048
rect 5408 15036 5414 15088
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 4798 15008 4804 15020
rect 4571 14980 4804 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 4798 14968 4804 14980
rect 4856 14968 4862 15020
rect 5537 15011 5595 15017
rect 5537 14977 5549 15011
rect 5583 15008 5595 15011
rect 6380 15008 6408 15107
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 16482 15104 16488 15156
rect 16540 15104 16546 15156
rect 16669 15147 16727 15153
rect 16669 15113 16681 15147
rect 16715 15113 16727 15147
rect 16669 15107 16727 15113
rect 10502 15076 10508 15088
rect 7852 15048 10508 15076
rect 7852 15017 7880 15048
rect 10502 15036 10508 15048
rect 10560 15036 10566 15088
rect 15194 15076 15200 15088
rect 13832 15048 15200 15076
rect 5583 14980 6408 15008
rect 7837 15011 7895 15017
rect 5583 14977 5595 14980
rect 5537 14971 5595 14977
rect 7837 14977 7849 15011
rect 7883 14977 7895 15011
rect 7837 14971 7895 14977
rect 8110 14968 8116 15020
rect 8168 14968 8174 15020
rect 13832 15017 13860 15048
rect 15194 15036 15200 15048
rect 15252 15036 15258 15088
rect 15372 15079 15430 15085
rect 15372 15045 15384 15079
rect 15418 15076 15430 15079
rect 16684 15076 16712 15107
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 24118 15144 24124 15156
rect 18472 15116 24124 15144
rect 18472 15104 18478 15116
rect 24118 15104 24124 15116
rect 24176 15104 24182 15156
rect 25130 15104 25136 15156
rect 25188 15104 25194 15156
rect 27246 15144 27252 15156
rect 25332 15116 27252 15144
rect 15418 15048 16712 15076
rect 15418 15045 15430 15048
rect 15372 15039 15430 15045
rect 17218 15036 17224 15088
rect 17276 15076 17282 15088
rect 23014 15076 23020 15088
rect 17276 15048 23020 15076
rect 17276 15036 17282 15048
rect 23014 15036 23020 15048
rect 23072 15036 23078 15088
rect 13817 15011 13875 15017
rect 13817 14977 13829 15011
rect 13863 14977 13875 15011
rect 13817 14971 13875 14977
rect 14090 14968 14096 15020
rect 14148 14968 14154 15020
rect 15105 15011 15163 15017
rect 15105 14977 15117 15011
rect 15151 15008 15163 15011
rect 16298 15008 16304 15020
rect 15151 14980 16304 15008
rect 15151 14977 15163 14980
rect 15105 14971 15163 14977
rect 16298 14968 16304 14980
rect 16356 15008 16362 15020
rect 16574 15008 16580 15020
rect 16356 14980 16580 15008
rect 16356 14968 16362 14980
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 16850 14968 16856 15020
rect 16908 14968 16914 15020
rect 17494 14968 17500 15020
rect 17552 15008 17558 15020
rect 17589 15011 17647 15017
rect 17589 15008 17601 15011
rect 17552 14980 17601 15008
rect 17552 14968 17558 14980
rect 17589 14977 17601 14980
rect 17635 14977 17647 15011
rect 17589 14971 17647 14977
rect 22278 14968 22284 15020
rect 22336 15008 22342 15020
rect 25332 15017 25360 15116
rect 27246 15104 27252 15116
rect 27304 15104 27310 15156
rect 33597 15147 33655 15153
rect 33597 15113 33609 15147
rect 33643 15144 33655 15147
rect 34054 15144 34060 15156
rect 33643 15116 34060 15144
rect 33643 15113 33655 15116
rect 33597 15107 33655 15113
rect 34054 15104 34060 15116
rect 34112 15104 34118 15156
rect 25501 15079 25559 15085
rect 25501 15045 25513 15079
rect 25547 15076 25559 15079
rect 25682 15076 25688 15088
rect 25547 15048 25688 15076
rect 25547 15045 25559 15048
rect 25501 15039 25559 15045
rect 25682 15036 25688 15048
rect 25740 15036 25746 15088
rect 28626 15076 28632 15088
rect 27356 15048 28632 15076
rect 22557 15011 22615 15017
rect 22557 15008 22569 15011
rect 22336 14980 22569 15008
rect 22336 14968 22342 14980
rect 22557 14977 22569 14980
rect 22603 14977 22615 15011
rect 22557 14971 22615 14977
rect 25317 15011 25375 15017
rect 25317 14977 25329 15011
rect 25363 14977 25375 15011
rect 25317 14971 25375 14977
rect 25406 14968 25412 15020
rect 25464 15008 25470 15020
rect 25593 15011 25651 15017
rect 25593 15008 25605 15011
rect 25464 14980 25605 15008
rect 25464 14968 25470 14980
rect 25593 14977 25605 14980
rect 25639 14977 25651 15011
rect 25593 14971 25651 14977
rect 4709 14943 4767 14949
rect 4709 14909 4721 14943
rect 4755 14909 4767 14943
rect 4709 14903 4767 14909
rect 4724 14872 4752 14903
rect 6638 14900 6644 14952
rect 6696 14940 6702 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6696 14912 6837 14940
rect 6696 14900 6702 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14940 6975 14943
rect 7742 14940 7748 14952
rect 6963 14912 7748 14940
rect 6963 14909 6975 14912
rect 6917 14903 6975 14909
rect 6932 14872 6960 14903
rect 7742 14900 7748 14912
rect 7800 14900 7806 14952
rect 17310 14900 17316 14952
rect 17368 14900 17374 14952
rect 24854 14900 24860 14952
rect 24912 14940 24918 14952
rect 27356 14940 27384 15048
rect 27430 14968 27436 15020
rect 27488 14968 27494 15020
rect 24912 14912 27384 14940
rect 24912 14900 24918 14912
rect 27522 14900 27528 14952
rect 27580 14900 27586 14952
rect 27632 14949 27660 15048
rect 28626 15036 28632 15048
rect 28684 15036 28690 15088
rect 30742 14968 30748 15020
rect 30800 15008 30806 15020
rect 31849 15011 31907 15017
rect 31849 15008 31861 15011
rect 30800 14980 31861 15008
rect 30800 14968 30806 14980
rect 31849 14977 31861 14980
rect 31895 14977 31907 15011
rect 31849 14971 31907 14977
rect 34238 14968 34244 15020
rect 34296 15008 34302 15020
rect 36170 15008 36176 15020
rect 34296 14980 36176 15008
rect 34296 14968 34302 14980
rect 36170 14968 36176 14980
rect 36228 14968 36234 15020
rect 27617 14943 27675 14949
rect 27617 14909 27629 14943
rect 27663 14909 27675 14943
rect 27617 14903 27675 14909
rect 33410 14900 33416 14952
rect 33468 14940 33474 14952
rect 33689 14943 33747 14949
rect 33689 14940 33701 14943
rect 33468 14912 33701 14940
rect 33468 14900 33474 14912
rect 33689 14909 33701 14912
rect 33735 14909 33747 14943
rect 33689 14903 33747 14909
rect 33781 14943 33839 14949
rect 33781 14909 33793 14943
rect 33827 14909 33839 14943
rect 33781 14903 33839 14909
rect 27982 14872 27988 14884
rect 4724 14844 6960 14872
rect 22066 14844 27988 14872
rect 3970 14764 3976 14816
rect 4028 14804 4034 14816
rect 4065 14807 4123 14813
rect 4065 14804 4077 14807
rect 4028 14776 4077 14804
rect 4028 14764 4034 14776
rect 4065 14773 4077 14776
rect 4111 14773 4123 14807
rect 4065 14767 4123 14773
rect 5350 14764 5356 14816
rect 5408 14764 5414 14816
rect 8849 14807 8907 14813
rect 8849 14773 8861 14807
rect 8895 14804 8907 14807
rect 9858 14804 9864 14816
rect 8895 14776 9864 14804
rect 8895 14773 8907 14776
rect 8849 14767 8907 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 14826 14764 14832 14816
rect 14884 14764 14890 14816
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18325 14807 18383 14813
rect 18325 14804 18337 14807
rect 18012 14776 18337 14804
rect 18012 14764 18018 14776
rect 18325 14773 18337 14776
rect 18371 14804 18383 14807
rect 22066 14804 22094 14844
rect 27982 14832 27988 14844
rect 28040 14832 28046 14884
rect 30282 14832 30288 14884
rect 30340 14872 30346 14884
rect 33796 14872 33824 14903
rect 30340 14844 33824 14872
rect 30340 14832 30346 14844
rect 18371 14776 22094 14804
rect 18371 14773 18383 14776
rect 18325 14767 18383 14773
rect 22370 14764 22376 14816
rect 22428 14764 22434 14816
rect 27065 14807 27123 14813
rect 27065 14773 27077 14807
rect 27111 14804 27123 14807
rect 27154 14804 27160 14816
rect 27111 14776 27160 14804
rect 27111 14773 27123 14776
rect 27065 14767 27123 14773
rect 27154 14764 27160 14776
rect 27212 14764 27218 14816
rect 31665 14807 31723 14813
rect 31665 14773 31677 14807
rect 31711 14804 31723 14807
rect 31846 14804 31852 14816
rect 31711 14776 31852 14804
rect 31711 14773 31723 14776
rect 31665 14767 31723 14773
rect 31846 14764 31852 14776
rect 31904 14764 31910 14816
rect 33226 14764 33232 14816
rect 33284 14764 33290 14816
rect 33318 14764 33324 14816
rect 33376 14804 33382 14816
rect 34057 14807 34115 14813
rect 34057 14804 34069 14807
rect 33376 14776 34069 14804
rect 33376 14764 33382 14776
rect 34057 14773 34069 14776
rect 34103 14773 34115 14807
rect 34057 14767 34115 14773
rect 1104 14714 36800 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 36800 14714
rect 1104 14640 36800 14662
rect 6457 14603 6515 14609
rect 6457 14569 6469 14603
rect 6503 14600 6515 14603
rect 6914 14600 6920 14612
rect 6503 14572 6920 14600
rect 6503 14569 6515 14572
rect 6457 14563 6515 14569
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 9858 14560 9864 14612
rect 9916 14560 9922 14612
rect 17218 14600 17224 14612
rect 9968 14572 17224 14600
rect 9968 14532 9996 14572
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 19245 14603 19303 14609
rect 19245 14569 19257 14603
rect 19291 14600 19303 14603
rect 20254 14600 20260 14612
rect 19291 14572 20260 14600
rect 19291 14569 19303 14572
rect 19245 14563 19303 14569
rect 20254 14560 20260 14572
rect 20312 14560 20318 14612
rect 22278 14560 22284 14612
rect 22336 14560 22342 14612
rect 27430 14560 27436 14612
rect 27488 14600 27494 14612
rect 27893 14603 27951 14609
rect 27893 14600 27905 14603
rect 27488 14572 27905 14600
rect 27488 14560 27494 14572
rect 27893 14569 27905 14572
rect 27939 14569 27951 14603
rect 27893 14563 27951 14569
rect 27982 14560 27988 14612
rect 28040 14600 28046 14612
rect 28040 14572 36216 14600
rect 28040 14560 28046 14572
rect 9692 14504 9996 14532
rect 3970 14356 3976 14408
rect 4028 14356 4034 14408
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 5350 14405 5356 14408
rect 5077 14399 5135 14405
rect 5077 14396 5089 14399
rect 4764 14368 5089 14396
rect 4764 14356 4770 14368
rect 5077 14365 5089 14368
rect 5123 14365 5135 14399
rect 5344 14396 5356 14405
rect 5311 14368 5356 14396
rect 5077 14359 5135 14365
rect 5344 14359 5356 14368
rect 5092 14328 5120 14359
rect 5350 14356 5356 14359
rect 5408 14356 5414 14408
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 7101 14399 7159 14405
rect 7101 14396 7113 14399
rect 6880 14368 7113 14396
rect 6880 14356 6886 14368
rect 7101 14365 7113 14368
rect 7147 14365 7159 14399
rect 7101 14359 7159 14365
rect 7377 14399 7435 14405
rect 7377 14365 7389 14399
rect 7423 14396 7435 14399
rect 9692 14396 9720 14504
rect 11698 14492 11704 14544
rect 11756 14492 11762 14544
rect 17310 14492 17316 14544
rect 17368 14532 17374 14544
rect 18138 14532 18144 14544
rect 17368 14504 18144 14532
rect 17368 14492 17374 14504
rect 18138 14492 18144 14504
rect 18196 14532 18202 14544
rect 18196 14504 19932 14532
rect 18196 14492 18202 14504
rect 10229 14467 10287 14473
rect 10229 14433 10241 14467
rect 10275 14464 10287 14467
rect 10275 14436 10548 14464
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 7423 14368 9720 14396
rect 7423 14365 7435 14368
rect 7377 14359 7435 14365
rect 9766 14356 9772 14408
rect 9824 14356 9830 14408
rect 10520 14405 10548 14436
rect 10962 14424 10968 14476
rect 11020 14464 11026 14476
rect 13906 14464 13912 14476
rect 11020 14436 13912 14464
rect 11020 14424 11026 14436
rect 13906 14424 13912 14436
rect 13964 14424 13970 14476
rect 19518 14424 19524 14476
rect 19576 14464 19582 14476
rect 19705 14467 19763 14473
rect 19705 14464 19717 14467
rect 19576 14436 19717 14464
rect 19576 14424 19582 14436
rect 19705 14433 19717 14436
rect 19751 14433 19763 14467
rect 19705 14427 19763 14433
rect 19797 14467 19855 14473
rect 19797 14433 19809 14467
rect 19843 14433 19855 14467
rect 19797 14427 19855 14433
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 10686 14356 10692 14408
rect 10744 14356 10750 14408
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 10836 14368 11928 14396
rect 10836 14356 10842 14368
rect 7926 14328 7932 14340
rect 5092 14300 7932 14328
rect 7926 14288 7932 14300
rect 7984 14288 7990 14340
rect 11425 14331 11483 14337
rect 11425 14297 11437 14331
rect 11471 14328 11483 14331
rect 11514 14328 11520 14340
rect 11471 14300 11520 14328
rect 11471 14297 11483 14300
rect 11425 14291 11483 14297
rect 11514 14288 11520 14300
rect 11572 14288 11578 14340
rect 11900 14328 11928 14368
rect 12066 14356 12072 14408
rect 12124 14356 12130 14408
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14365 12219 14399
rect 12161 14359 12219 14365
rect 13633 14399 13691 14405
rect 13633 14365 13645 14399
rect 13679 14396 13691 14399
rect 13722 14396 13728 14408
rect 13679 14368 13728 14396
rect 13679 14365 13691 14368
rect 13633 14359 13691 14365
rect 12176 14328 12204 14359
rect 13722 14356 13728 14368
rect 13780 14396 13786 14408
rect 13780 14368 13952 14396
rect 13780 14356 13786 14368
rect 12526 14328 12532 14340
rect 11900 14300 12532 14328
rect 12526 14288 12532 14300
rect 12584 14288 12590 14340
rect 13924 14328 13952 14368
rect 14090 14356 14096 14408
rect 14148 14396 14154 14408
rect 14826 14396 14832 14408
rect 14148 14368 14832 14396
rect 14148 14356 14154 14368
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 15470 14356 15476 14408
rect 15528 14356 15534 14408
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14396 15807 14399
rect 18414 14396 18420 14408
rect 15795 14368 18420 14396
rect 15795 14365 15807 14368
rect 15749 14359 15807 14365
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 18506 14356 18512 14408
rect 18564 14356 18570 14408
rect 14277 14331 14335 14337
rect 14277 14328 14289 14331
rect 13924 14300 14289 14328
rect 14277 14297 14289 14300
rect 14323 14297 14335 14331
rect 14277 14291 14335 14297
rect 17770 14288 17776 14340
rect 17828 14328 17834 14340
rect 19812 14328 19840 14427
rect 19904 14396 19932 14504
rect 19978 14492 19984 14544
rect 20036 14532 20042 14544
rect 25406 14532 25412 14544
rect 20036 14504 25412 14532
rect 20036 14492 20042 14504
rect 25406 14492 25412 14504
rect 25464 14492 25470 14544
rect 30190 14492 30196 14544
rect 30248 14532 30254 14544
rect 30561 14535 30619 14541
rect 30561 14532 30573 14535
rect 30248 14504 30573 14532
rect 30248 14492 30254 14504
rect 30561 14501 30573 14504
rect 30607 14501 30619 14535
rect 30561 14495 30619 14501
rect 30742 14492 30748 14544
rect 30800 14492 30806 14544
rect 34054 14492 34060 14544
rect 34112 14532 34118 14544
rect 34333 14535 34391 14541
rect 34333 14532 34345 14535
rect 34112 14504 34345 14532
rect 34112 14492 34118 14504
rect 34333 14501 34345 14504
rect 34379 14501 34391 14535
rect 34333 14495 34391 14501
rect 20990 14424 20996 14476
rect 21048 14424 21054 14476
rect 21358 14424 21364 14476
rect 21416 14464 21422 14476
rect 22925 14467 22983 14473
rect 22925 14464 22937 14467
rect 21416 14436 22937 14464
rect 21416 14424 21422 14436
rect 22925 14433 22937 14436
rect 22971 14464 22983 14467
rect 23014 14464 23020 14476
rect 22971 14436 23020 14464
rect 22971 14433 22983 14436
rect 22925 14427 22983 14433
rect 23014 14424 23020 14436
rect 23072 14424 23078 14476
rect 26142 14424 26148 14476
rect 26200 14464 26206 14476
rect 26513 14467 26571 14473
rect 26513 14464 26525 14467
rect 26200 14436 26525 14464
rect 26200 14424 26206 14436
rect 26513 14433 26525 14436
rect 26559 14433 26571 14467
rect 26513 14427 26571 14433
rect 28166 14424 28172 14476
rect 28224 14464 28230 14476
rect 29549 14467 29607 14473
rect 29549 14464 29561 14467
rect 28224 14436 29561 14464
rect 28224 14424 28230 14436
rect 29549 14433 29561 14436
rect 29595 14433 29607 14467
rect 29549 14427 29607 14433
rect 30282 14424 30288 14476
rect 30340 14464 30346 14476
rect 31297 14467 31355 14473
rect 31297 14464 31309 14467
rect 30340 14436 31309 14464
rect 30340 14424 30346 14436
rect 31297 14433 31309 14436
rect 31343 14433 31355 14467
rect 31297 14427 31355 14433
rect 32858 14424 32864 14476
rect 32916 14464 32922 14476
rect 33318 14464 33324 14476
rect 32916 14436 33324 14464
rect 32916 14424 32922 14436
rect 33318 14424 33324 14436
rect 33376 14424 33382 14476
rect 25406 14396 25412 14408
rect 19904 14368 25412 14396
rect 25406 14356 25412 14368
rect 25464 14356 25470 14408
rect 25685 14399 25743 14405
rect 25685 14365 25697 14399
rect 25731 14396 25743 14399
rect 26418 14396 26424 14408
rect 25731 14368 26424 14396
rect 25731 14365 25743 14368
rect 25685 14359 25743 14365
rect 26418 14356 26424 14368
rect 26476 14356 26482 14408
rect 29362 14356 29368 14408
rect 29420 14356 29426 14408
rect 29825 14399 29883 14405
rect 29825 14365 29837 14399
rect 29871 14365 29883 14399
rect 29825 14359 29883 14365
rect 31573 14399 31631 14405
rect 31573 14365 31585 14399
rect 31619 14396 31631 14399
rect 31619 14368 31754 14396
rect 31619 14365 31631 14368
rect 31573 14359 31631 14365
rect 21358 14328 21364 14340
rect 17828 14300 21364 14328
rect 17828 14288 17834 14300
rect 21358 14288 21364 14300
rect 21416 14288 21422 14340
rect 22738 14288 22744 14340
rect 22796 14288 22802 14340
rect 24486 14288 24492 14340
rect 24544 14288 24550 14340
rect 26780 14331 26838 14337
rect 26780 14297 26792 14331
rect 26826 14328 26838 14331
rect 26970 14328 26976 14340
rect 26826 14300 26976 14328
rect 26826 14297 26838 14300
rect 26780 14291 26838 14297
rect 26970 14288 26976 14300
rect 27028 14288 27034 14340
rect 29840 14328 29868 14359
rect 29196 14300 29868 14328
rect 31113 14331 31171 14337
rect 3786 14220 3792 14272
rect 3844 14220 3850 14272
rect 8113 14263 8171 14269
rect 8113 14229 8125 14263
rect 8159 14260 8171 14263
rect 8202 14260 8208 14272
rect 8159 14232 8208 14260
rect 8159 14229 8171 14232
rect 8113 14223 8171 14229
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 10689 14263 10747 14269
rect 10689 14229 10701 14263
rect 10735 14260 10747 14263
rect 11790 14260 11796 14272
rect 10735 14232 11796 14260
rect 10735 14229 10747 14232
rect 10689 14223 10747 14229
rect 11790 14220 11796 14232
rect 11848 14220 11854 14272
rect 11882 14220 11888 14272
rect 11940 14220 11946 14272
rect 12342 14220 12348 14272
rect 12400 14220 12406 14272
rect 13262 14220 13268 14272
rect 13320 14260 13326 14272
rect 13722 14260 13728 14272
rect 13320 14232 13728 14260
rect 13320 14220 13326 14232
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 14461 14263 14519 14269
rect 14461 14229 14473 14263
rect 14507 14260 14519 14263
rect 14550 14260 14556 14272
rect 14507 14232 14556 14260
rect 14507 14229 14519 14232
rect 14461 14223 14519 14229
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 16482 14220 16488 14272
rect 16540 14220 16546 14272
rect 18325 14263 18383 14269
rect 18325 14229 18337 14263
rect 18371 14260 18383 14263
rect 18598 14260 18604 14272
rect 18371 14232 18604 14260
rect 18371 14229 18383 14232
rect 18325 14223 18383 14229
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 19610 14220 19616 14272
rect 19668 14220 19674 14272
rect 20438 14220 20444 14272
rect 20496 14220 20502 14272
rect 20806 14220 20812 14272
rect 20864 14220 20870 14272
rect 20901 14263 20959 14269
rect 20901 14229 20913 14263
rect 20947 14260 20959 14263
rect 21174 14260 21180 14272
rect 20947 14232 21180 14260
rect 20947 14229 20959 14232
rect 20901 14223 20959 14229
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 22646 14220 22652 14272
rect 22704 14220 22710 14272
rect 24118 14220 24124 14272
rect 24176 14260 24182 14272
rect 24581 14263 24639 14269
rect 24581 14260 24593 14263
rect 24176 14232 24593 14260
rect 24176 14220 24182 14232
rect 24581 14229 24593 14232
rect 24627 14229 24639 14263
rect 24581 14223 24639 14229
rect 26418 14220 26424 14272
rect 26476 14220 26482 14272
rect 29196 14269 29224 14300
rect 31113 14297 31125 14331
rect 31159 14328 31171 14331
rect 31726 14328 31754 14368
rect 31846 14356 31852 14408
rect 31904 14356 31910 14408
rect 33226 14356 33232 14408
rect 33284 14356 33290 14408
rect 36188 14405 36216 14572
rect 33597 14399 33655 14405
rect 33597 14365 33609 14399
rect 33643 14365 33655 14399
rect 33597 14359 33655 14365
rect 36173 14399 36231 14405
rect 36173 14365 36185 14399
rect 36219 14365 36231 14399
rect 36173 14359 36231 14365
rect 32858 14328 32864 14340
rect 31159 14300 31432 14328
rect 31726 14300 32864 14328
rect 31159 14297 31171 14300
rect 31113 14291 31171 14297
rect 29181 14263 29239 14269
rect 29181 14229 29193 14263
rect 29227 14229 29239 14263
rect 29181 14223 29239 14229
rect 29270 14220 29276 14272
rect 29328 14260 29334 14272
rect 30006 14260 30012 14272
rect 29328 14232 30012 14260
rect 29328 14220 29334 14232
rect 30006 14220 30012 14232
rect 30064 14220 30070 14272
rect 31202 14220 31208 14272
rect 31260 14220 31266 14272
rect 31404 14260 31432 14300
rect 32858 14288 32864 14300
rect 32916 14288 32922 14340
rect 33612 14328 33640 14359
rect 33060 14300 33640 14328
rect 32582 14260 32588 14272
rect 31404 14232 32588 14260
rect 32582 14220 32588 14232
rect 32640 14220 32646 14272
rect 33060 14269 33088 14300
rect 33045 14263 33103 14269
rect 33045 14229 33057 14263
rect 33091 14229 33103 14263
rect 33045 14223 33103 14229
rect 36354 14220 36360 14272
rect 36412 14220 36418 14272
rect 1104 14170 36800 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 36800 14170
rect 1104 14096 36800 14118
rect 4525 14059 4583 14065
rect 4525 14025 4537 14059
rect 4571 14056 4583 14059
rect 4614 14056 4620 14068
rect 4571 14028 4620 14056
rect 4571 14025 4583 14028
rect 4525 14019 4583 14025
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 7929 14059 7987 14065
rect 7929 14025 7941 14059
rect 7975 14025 7987 14059
rect 7929 14019 7987 14025
rect 10597 14059 10655 14065
rect 10597 14025 10609 14059
rect 10643 14056 10655 14059
rect 10686 14056 10692 14068
rect 10643 14028 10692 14056
rect 10643 14025 10655 14028
rect 10597 14019 10655 14025
rect 3412 13991 3470 13997
rect 3412 13957 3424 13991
rect 3458 13988 3470 13991
rect 3786 13988 3792 14000
rect 3458 13960 3792 13988
rect 3458 13957 3470 13960
rect 3412 13951 3470 13957
rect 3786 13948 3792 13960
rect 3844 13948 3850 14000
rect 6730 13948 6736 14000
rect 6788 13988 6794 14000
rect 6788 13960 7236 13988
rect 6788 13948 6794 13960
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 4706 13920 4712 13932
rect 3191 13892 4712 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 6822 13880 6828 13932
rect 6880 13920 6886 13932
rect 7208 13929 7236 13960
rect 6917 13923 6975 13929
rect 6917 13920 6929 13923
rect 6880 13892 6929 13920
rect 6880 13880 6886 13892
rect 6917 13889 6929 13892
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 7193 13923 7251 13929
rect 7193 13889 7205 13923
rect 7239 13889 7251 13923
rect 7944 13920 7972 14019
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 10962 14016 10968 14068
rect 11020 14056 11026 14068
rect 11149 14059 11207 14065
rect 11149 14056 11161 14059
rect 11020 14028 11161 14056
rect 11020 14016 11026 14028
rect 11149 14025 11161 14028
rect 11195 14025 11207 14059
rect 12066 14056 12072 14068
rect 11149 14019 11207 14025
rect 11256 14028 12072 14056
rect 9766 13988 9772 14000
rect 8404 13960 9772 13988
rect 8404 13929 8432 13960
rect 9766 13948 9772 13960
rect 9824 13948 9830 14000
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 7944 13892 8401 13920
rect 7193 13883 7251 13889
rect 8389 13889 8401 13892
rect 8435 13889 8447 13923
rect 8389 13883 8447 13889
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13889 8631 13923
rect 8573 13883 8631 13889
rect 9309 13923 9367 13929
rect 9309 13889 9321 13923
rect 9355 13920 9367 13923
rect 9858 13920 9864 13932
rect 9355 13892 9864 13920
rect 9355 13889 9367 13892
rect 9309 13883 9367 13889
rect 8588 13852 8616 13883
rect 9858 13880 9864 13892
rect 9916 13920 9922 13932
rect 10137 13923 10195 13929
rect 10137 13920 10149 13923
rect 9916 13892 10149 13920
rect 9916 13880 9922 13892
rect 10137 13889 10149 13892
rect 10183 13920 10195 13923
rect 10226 13920 10232 13932
rect 10183 13892 10232 13920
rect 10183 13889 10195 13892
rect 10137 13883 10195 13889
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13920 10747 13923
rect 11256 13920 11284 14028
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 14090 14056 14096 14068
rect 13096 14028 14096 14056
rect 12526 13948 12532 14000
rect 12584 13948 12590 14000
rect 10735 13892 11284 13920
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 8588 13824 9505 13852
rect 9493 13821 9505 13824
rect 9539 13852 9551 13855
rect 10704 13852 10732 13883
rect 11606 13880 11612 13932
rect 11664 13920 11670 13932
rect 12161 13923 12219 13929
rect 12161 13920 12173 13923
rect 11664 13892 12173 13920
rect 11664 13880 11670 13892
rect 12161 13889 12173 13892
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12342 13880 12348 13932
rect 12400 13880 12406 13932
rect 13096 13929 13124 14028
rect 13170 13948 13176 14000
rect 13228 13948 13234 14000
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 12912 13892 13093 13920
rect 9539 13824 10732 13852
rect 9539 13821 9551 13824
rect 9493 13815 9551 13821
rect 11514 13812 11520 13864
rect 11572 13812 11578 13864
rect 11698 13812 11704 13864
rect 11756 13812 11762 13864
rect 11790 13812 11796 13864
rect 11848 13852 11854 13864
rect 11885 13855 11943 13861
rect 11885 13852 11897 13855
rect 11848 13824 11897 13852
rect 11848 13812 11854 13824
rect 11885 13821 11897 13824
rect 11931 13821 11943 13855
rect 12912 13852 12940 13892
rect 13081 13889 13093 13892
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13262 13880 13268 13932
rect 13320 13880 13326 13932
rect 13556 13929 13584 14028
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 19337 14059 19395 14065
rect 15528 14028 18368 14056
rect 15528 14016 15534 14028
rect 14182 13988 14188 14000
rect 14016 13960 14188 13988
rect 13722 13929 13728 13932
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13706 13923 13728 13929
rect 13706 13889 13718 13923
rect 13706 13883 13728 13889
rect 13722 13880 13728 13883
rect 13780 13880 13786 13932
rect 13817 13923 13875 13929
rect 13817 13889 13829 13923
rect 13863 13889 13875 13923
rect 13817 13883 13875 13889
rect 11885 13815 11943 13821
rect 11992 13824 12940 13852
rect 12989 13855 13047 13861
rect 10594 13784 10600 13796
rect 7576 13756 10600 13784
rect 2314 13676 2320 13728
rect 2372 13716 2378 13728
rect 7576 13716 7604 13756
rect 10594 13744 10600 13756
rect 10652 13744 10658 13796
rect 10778 13784 10784 13796
rect 10704 13756 10784 13784
rect 2372 13688 7604 13716
rect 2372 13676 2378 13688
rect 8386 13676 8392 13728
rect 8444 13716 8450 13728
rect 8481 13719 8539 13725
rect 8481 13716 8493 13719
rect 8444 13688 8493 13716
rect 8444 13676 8450 13688
rect 8481 13685 8493 13688
rect 8527 13685 8539 13719
rect 8481 13679 8539 13685
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 10229 13719 10287 13725
rect 10229 13716 10241 13719
rect 9824 13688 10241 13716
rect 9824 13676 9830 13688
rect 10229 13685 10241 13688
rect 10275 13716 10287 13719
rect 10704 13716 10732 13756
rect 10778 13744 10784 13756
rect 10836 13784 10842 13796
rect 10965 13787 11023 13793
rect 10965 13784 10977 13787
rect 10836 13756 10977 13784
rect 10836 13744 10842 13756
rect 10965 13753 10977 13756
rect 11011 13753 11023 13787
rect 11716 13784 11744 13812
rect 11992 13784 12020 13824
rect 12989 13821 13001 13855
rect 13035 13852 13047 13855
rect 13832 13852 13860 13883
rect 13906 13880 13912 13932
rect 13964 13880 13970 13932
rect 14016 13929 14044 13960
rect 14182 13948 14188 13960
rect 14240 13988 14246 14000
rect 18340 13988 18368 14028
rect 19337 14025 19349 14059
rect 19383 14056 19395 14059
rect 19610 14056 19616 14068
rect 19383 14028 19616 14056
rect 19383 14025 19395 14028
rect 19337 14019 19395 14025
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 19978 14056 19984 14068
rect 19720 14028 19984 14056
rect 19720 13988 19748 14028
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 21361 14059 21419 14065
rect 21361 14056 21373 14059
rect 20864 14028 21373 14056
rect 20864 14016 20870 14028
rect 21361 14025 21373 14028
rect 21407 14025 21419 14059
rect 21361 14019 21419 14025
rect 22646 14016 22652 14068
rect 22704 14056 22710 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 22704 14028 23397 14056
rect 22704 14016 22710 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 23845 14059 23903 14065
rect 23845 14025 23857 14059
rect 23891 14025 23903 14059
rect 23845 14019 23903 14025
rect 21266 13988 21272 14000
rect 14240 13960 14780 13988
rect 18340 13960 19748 13988
rect 19996 13960 21272 13988
rect 14240 13948 14246 13960
rect 14001 13923 14059 13929
rect 14001 13889 14013 13923
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 14090 13880 14096 13932
rect 14148 13920 14154 13932
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 14148 13892 14289 13920
rect 14148 13880 14154 13892
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13889 14519 13923
rect 14461 13883 14519 13889
rect 14476 13852 14504 13883
rect 14550 13880 14556 13932
rect 14608 13880 14614 13932
rect 14752 13929 14780 13960
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 16298 13880 16304 13932
rect 16356 13920 16362 13932
rect 17957 13923 18015 13929
rect 17957 13920 17969 13923
rect 16356 13892 17969 13920
rect 16356 13880 16362 13892
rect 17957 13889 17969 13892
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 18224 13923 18282 13929
rect 18224 13889 18236 13923
rect 18270 13920 18282 13923
rect 18598 13920 18604 13932
rect 18270 13892 18604 13920
rect 18270 13889 18282 13892
rect 18224 13883 18282 13889
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 19996 13929 20024 13960
rect 21266 13948 21272 13960
rect 21324 13988 21330 14000
rect 21542 13988 21548 14000
rect 21324 13960 21548 13988
rect 21324 13948 21330 13960
rect 21542 13948 21548 13960
rect 21600 13948 21606 14000
rect 22278 13997 22284 14000
rect 22272 13988 22284 13997
rect 22239 13960 22284 13988
rect 22272 13951 22284 13960
rect 22278 13948 22284 13951
rect 22336 13948 22342 14000
rect 23860 13988 23888 14019
rect 25406 14016 25412 14068
rect 25464 14056 25470 14068
rect 25685 14059 25743 14065
rect 25685 14056 25697 14059
rect 25464 14028 25697 14056
rect 25464 14016 25470 14028
rect 25685 14025 25697 14028
rect 25731 14025 25743 14059
rect 25685 14019 25743 14025
rect 26970 14016 26976 14068
rect 27028 14016 27034 14068
rect 29362 14016 29368 14068
rect 29420 14056 29426 14068
rect 29549 14059 29607 14065
rect 29549 14056 29561 14059
rect 29420 14028 29561 14056
rect 29420 14016 29426 14028
rect 29549 14025 29561 14028
rect 29595 14025 29607 14059
rect 29549 14019 29607 14025
rect 29917 14059 29975 14065
rect 29917 14025 29929 14059
rect 29963 14056 29975 14059
rect 30190 14056 30196 14068
rect 29963 14028 30196 14056
rect 29963 14025 29975 14028
rect 29917 14019 29975 14025
rect 30190 14016 30196 14028
rect 30248 14016 30254 14068
rect 30561 14059 30619 14065
rect 30561 14025 30573 14059
rect 30607 14025 30619 14059
rect 30561 14019 30619 14025
rect 24366 13991 24424 13997
rect 24366 13988 24378 13991
rect 23860 13960 24378 13988
rect 24366 13957 24378 13960
rect 24412 13957 24424 13991
rect 24366 13951 24424 13957
rect 28166 13948 28172 14000
rect 28224 13988 28230 14000
rect 30576 13988 30604 14019
rect 33134 14016 33140 14068
rect 33192 14016 33198 14068
rect 33505 14059 33563 14065
rect 33505 14025 33517 14059
rect 33551 14056 33563 14059
rect 34054 14056 34060 14068
rect 33551 14028 34060 14056
rect 33551 14025 33563 14028
rect 33505 14019 33563 14025
rect 34054 14016 34060 14028
rect 34112 14016 34118 14068
rect 28224 13960 29408 13988
rect 30576 13960 31156 13988
rect 28224 13948 28230 13960
rect 20254 13929 20260 13932
rect 19981 13923 20039 13929
rect 19981 13889 19993 13923
rect 20027 13889 20039 13923
rect 19981 13883 20039 13889
rect 20248 13883 20260 13929
rect 20254 13880 20260 13883
rect 20312 13880 20318 13932
rect 21637 13923 21695 13929
rect 21637 13889 21649 13923
rect 21683 13889 21695 13923
rect 21637 13883 21695 13889
rect 22112 13892 23060 13920
rect 13035 13824 14504 13852
rect 14921 13855 14979 13861
rect 13035 13821 13047 13824
rect 12989 13815 13047 13821
rect 14921 13821 14933 13855
rect 14967 13852 14979 13855
rect 15194 13852 15200 13864
rect 14967 13824 15200 13852
rect 14967 13821 14979 13824
rect 14921 13815 14979 13821
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 21652 13852 21680 13883
rect 21818 13852 21824 13864
rect 21652 13824 21824 13852
rect 21818 13812 21824 13824
rect 21876 13812 21882 13864
rect 22002 13852 22008 13864
rect 21963 13824 22008 13852
rect 22002 13812 22008 13824
rect 22060 13852 22066 13864
rect 22112 13852 22140 13892
rect 22060 13824 22140 13852
rect 23032 13852 23060 13892
rect 24026 13880 24032 13932
rect 24084 13880 24090 13932
rect 24118 13880 24124 13932
rect 24176 13880 24182 13932
rect 24210 13880 24216 13932
rect 24268 13920 24274 13932
rect 24268 13892 25820 13920
rect 24268 13880 24274 13892
rect 24136 13852 24164 13880
rect 23032 13824 24164 13852
rect 25792 13852 25820 13892
rect 25866 13880 25872 13932
rect 25924 13880 25930 13932
rect 27154 13880 27160 13932
rect 27212 13880 27218 13932
rect 28442 13880 28448 13932
rect 28500 13880 28506 13932
rect 29270 13880 29276 13932
rect 29328 13880 29334 13932
rect 29380 13920 29408 13960
rect 29380 13892 30420 13920
rect 25792 13824 28120 13852
rect 22060 13812 22066 13824
rect 10965 13747 11023 13753
rect 11072 13756 11284 13784
rect 11716 13756 12020 13784
rect 10275 13688 10732 13716
rect 10275 13685 10287 13688
rect 10229 13679 10287 13685
rect 10870 13676 10876 13728
rect 10928 13716 10934 13728
rect 11072 13716 11100 13756
rect 10928 13688 11100 13716
rect 11256 13716 11284 13756
rect 12066 13744 12072 13796
rect 12124 13784 12130 13796
rect 12342 13784 12348 13796
rect 12124 13756 12348 13784
rect 12124 13744 12130 13756
rect 12342 13744 12348 13756
rect 12400 13784 12406 13796
rect 12805 13787 12863 13793
rect 12805 13784 12817 13787
rect 12400 13756 12817 13784
rect 12400 13744 12406 13756
rect 12805 13753 12817 13756
rect 12851 13753 12863 13787
rect 17954 13784 17960 13796
rect 12805 13747 12863 13753
rect 13280 13756 17960 13784
rect 13280 13716 13308 13756
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 25498 13744 25504 13796
rect 25556 13744 25562 13796
rect 11256 13688 13308 13716
rect 13357 13719 13415 13725
rect 10928 13676 10934 13688
rect 13357 13685 13369 13719
rect 13403 13716 13415 13719
rect 13906 13716 13912 13728
rect 13403 13688 13912 13716
rect 13403 13685 13415 13688
rect 13357 13679 13415 13685
rect 13906 13676 13912 13688
rect 13964 13676 13970 13728
rect 13998 13676 14004 13728
rect 14056 13716 14062 13728
rect 14277 13719 14335 13725
rect 14277 13716 14289 13719
rect 14056 13688 14289 13716
rect 14056 13676 14062 13688
rect 14277 13685 14289 13688
rect 14323 13685 14335 13719
rect 14277 13679 14335 13685
rect 21453 13719 21511 13725
rect 21453 13685 21465 13719
rect 21499 13716 21511 13719
rect 22278 13716 22284 13728
rect 21499 13688 22284 13716
rect 21499 13685 21511 13688
rect 21453 13679 21511 13685
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 23842 13676 23848 13728
rect 23900 13716 23906 13728
rect 27982 13716 27988 13728
rect 23900 13688 27988 13716
rect 23900 13676 23906 13688
rect 27982 13676 27988 13688
rect 28040 13676 28046 13728
rect 28092 13716 28120 13824
rect 28166 13812 28172 13864
rect 28224 13812 28230 13864
rect 30009 13855 30067 13861
rect 30009 13852 30021 13855
rect 28828 13824 30021 13852
rect 28534 13716 28540 13728
rect 28092 13688 28540 13716
rect 28534 13676 28540 13688
rect 28592 13716 28598 13728
rect 28828 13716 28856 13824
rect 28592 13688 28856 13716
rect 29840 13716 29868 13824
rect 30009 13821 30021 13824
rect 30055 13821 30067 13855
rect 30009 13815 30067 13821
rect 30101 13855 30159 13861
rect 30101 13821 30113 13855
rect 30147 13852 30159 13855
rect 30282 13852 30288 13864
rect 30147 13824 30288 13852
rect 30147 13821 30159 13824
rect 30101 13815 30159 13821
rect 29914 13744 29920 13796
rect 29972 13784 29978 13796
rect 30116 13784 30144 13815
rect 30282 13812 30288 13824
rect 30340 13812 30346 13864
rect 30392 13852 30420 13892
rect 30742 13880 30748 13932
rect 30800 13880 30806 13932
rect 31128 13929 31156 13960
rect 31113 13923 31171 13929
rect 31113 13889 31125 13923
rect 31159 13889 31171 13923
rect 31113 13883 31171 13889
rect 31938 13880 31944 13932
rect 31996 13920 32002 13932
rect 33502 13920 33508 13932
rect 31996 13892 33508 13920
rect 31996 13880 32002 13892
rect 33502 13880 33508 13892
rect 33560 13880 33566 13932
rect 30837 13855 30895 13861
rect 30837 13852 30849 13855
rect 30392 13824 30849 13852
rect 30837 13821 30849 13824
rect 30883 13821 30895 13855
rect 30837 13815 30895 13821
rect 29972 13756 30144 13784
rect 29972 13744 29978 13756
rect 30650 13716 30656 13728
rect 29840 13688 30656 13716
rect 28592 13676 28598 13688
rect 30650 13676 30656 13688
rect 30708 13676 30714 13728
rect 30852 13716 30880 13815
rect 33594 13812 33600 13864
rect 33652 13812 33658 13864
rect 33686 13812 33692 13864
rect 33744 13812 33750 13864
rect 32950 13716 32956 13728
rect 30852 13688 32956 13716
rect 32950 13676 32956 13688
rect 33008 13676 33014 13728
rect 1104 13626 36800 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 36800 13626
rect 1104 13552 36800 13574
rect 5920 13484 9352 13512
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13308 4491 13311
rect 4614 13308 4620 13320
rect 4479 13280 4620 13308
rect 4479 13277 4491 13280
rect 4433 13271 4491 13277
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 5920 13308 5948 13484
rect 7190 13404 7196 13456
rect 7248 13444 7254 13456
rect 8113 13447 8171 13453
rect 8113 13444 8125 13447
rect 7248 13416 8125 13444
rect 7248 13404 7254 13416
rect 8113 13413 8125 13416
rect 8159 13413 8171 13447
rect 9324 13444 9352 13484
rect 9398 13472 9404 13524
rect 9456 13512 9462 13524
rect 16393 13515 16451 13521
rect 16393 13512 16405 13515
rect 9456 13484 16405 13512
rect 9456 13472 9462 13484
rect 16393 13481 16405 13484
rect 16439 13481 16451 13515
rect 16666 13512 16672 13524
rect 16393 13475 16451 13481
rect 16500 13484 16672 13512
rect 10042 13444 10048 13456
rect 9324 13416 10048 13444
rect 8113 13407 8171 13413
rect 10042 13404 10048 13416
rect 10100 13404 10106 13456
rect 10321 13447 10379 13453
rect 10321 13413 10333 13447
rect 10367 13444 10379 13447
rect 10962 13444 10968 13456
rect 10367 13416 10968 13444
rect 10367 13413 10379 13416
rect 10321 13407 10379 13413
rect 10962 13404 10968 13416
rect 11020 13404 11026 13456
rect 16500 13444 16528 13484
rect 16666 13472 16672 13484
rect 16724 13472 16730 13524
rect 17678 13472 17684 13524
rect 17736 13512 17742 13524
rect 17865 13515 17923 13521
rect 17865 13512 17877 13515
rect 17736 13484 17877 13512
rect 17736 13472 17742 13484
rect 17865 13481 17877 13484
rect 17911 13481 17923 13515
rect 17865 13475 17923 13481
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 18564 13484 19257 13512
rect 18564 13472 18570 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 20254 13472 20260 13524
rect 20312 13472 20318 13524
rect 20714 13472 20720 13524
rect 20772 13472 20778 13524
rect 21818 13472 21824 13524
rect 21876 13512 21882 13524
rect 22281 13515 22339 13521
rect 22281 13512 22293 13515
rect 21876 13484 22293 13512
rect 21876 13472 21882 13484
rect 22281 13481 22293 13484
rect 22327 13481 22339 13515
rect 22281 13475 22339 13481
rect 24026 13472 24032 13524
rect 24084 13512 24090 13524
rect 24397 13515 24455 13521
rect 24397 13512 24409 13515
rect 24084 13484 24409 13512
rect 24084 13472 24090 13484
rect 24397 13481 24409 13484
rect 24443 13481 24455 13515
rect 24397 13475 24455 13481
rect 28442 13472 28448 13524
rect 28500 13512 28506 13524
rect 28905 13515 28963 13521
rect 28905 13512 28917 13515
rect 28500 13484 28917 13512
rect 28500 13472 28506 13484
rect 28905 13481 28917 13484
rect 28951 13481 28963 13515
rect 28905 13475 28963 13481
rect 30742 13472 30748 13524
rect 30800 13512 30806 13524
rect 30929 13515 30987 13521
rect 30929 13512 30941 13515
rect 30800 13484 30941 13512
rect 30800 13472 30806 13484
rect 30929 13481 30941 13484
rect 30975 13481 30987 13515
rect 30929 13475 30987 13481
rect 23842 13444 23848 13456
rect 16224 13416 16528 13444
rect 17512 13416 23848 13444
rect 6638 13336 6644 13388
rect 6696 13376 6702 13388
rect 10505 13379 10563 13385
rect 6696 13348 10364 13376
rect 6696 13336 6702 13348
rect 4755 13280 5948 13308
rect 5997 13311 6055 13317
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 5997 13277 6009 13311
rect 6043 13277 6055 13311
rect 5997 13271 6055 13277
rect 6012 13240 6040 13271
rect 6270 13268 6276 13320
rect 6328 13268 6334 13320
rect 8386 13268 8392 13320
rect 8444 13268 8450 13320
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10336 13308 10364 13348
rect 10505 13345 10517 13379
rect 10551 13376 10563 13379
rect 10686 13376 10692 13388
rect 10551 13348 10692 13376
rect 10551 13345 10563 13348
rect 10505 13339 10563 13345
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 11701 13379 11759 13385
rect 11701 13345 11713 13379
rect 11747 13376 11759 13379
rect 11790 13376 11796 13388
rect 11747 13348 11796 13376
rect 11747 13345 11759 13348
rect 11701 13339 11759 13345
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 11977 13379 12035 13385
rect 11977 13345 11989 13379
rect 12023 13376 12035 13379
rect 13078 13376 13084 13388
rect 12023 13348 13084 13376
rect 12023 13345 12035 13348
rect 11977 13339 12035 13345
rect 13078 13336 13084 13348
rect 13136 13336 13142 13388
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 15381 13379 15439 13385
rect 15381 13376 15393 13379
rect 15344 13348 15393 13376
rect 15344 13336 15350 13348
rect 15381 13345 15393 13348
rect 15427 13345 15439 13379
rect 15381 13339 15439 13345
rect 11054 13308 11060 13320
rect 10336 13280 11060 13308
rect 10229 13271 10287 13277
rect 6822 13240 6828 13252
rect 6012 13212 6828 13240
rect 6822 13200 6828 13212
rect 6880 13200 6886 13252
rect 8113 13243 8171 13249
rect 8113 13209 8125 13243
rect 8159 13240 8171 13243
rect 8846 13240 8852 13252
rect 8159 13212 8852 13240
rect 8159 13209 8171 13212
rect 8113 13203 8171 13209
rect 8846 13200 8852 13212
rect 8904 13200 8910 13252
rect 10244 13240 10272 13271
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 11609 13311 11667 13317
rect 11609 13277 11621 13311
rect 11655 13308 11667 13311
rect 11882 13308 11888 13320
rect 11655 13280 11888 13308
rect 11655 13277 11667 13280
rect 11609 13271 11667 13277
rect 11624 13240 11652 13271
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13308 15715 13311
rect 16224 13308 16252 13416
rect 16298 13336 16304 13388
rect 16356 13376 16362 13388
rect 16485 13379 16543 13385
rect 16485 13376 16497 13379
rect 16356 13348 16497 13376
rect 16356 13336 16362 13348
rect 16485 13345 16497 13348
rect 16531 13345 16543 13379
rect 16485 13339 16543 13345
rect 17512 13308 17540 13416
rect 23842 13404 23848 13416
rect 23900 13404 23906 13456
rect 28077 13447 28135 13453
rect 23952 13416 25636 13444
rect 18417 13379 18475 13385
rect 18417 13345 18429 13379
rect 18463 13376 18475 13379
rect 19058 13376 19064 13388
rect 18463 13348 19064 13376
rect 18463 13345 18475 13348
rect 18417 13339 18475 13345
rect 19058 13336 19064 13348
rect 19116 13336 19122 13388
rect 19518 13336 19524 13388
rect 19576 13376 19582 13388
rect 19705 13379 19763 13385
rect 19705 13376 19717 13379
rect 19576 13348 19717 13376
rect 19576 13336 19582 13348
rect 19705 13345 19717 13348
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 19797 13379 19855 13385
rect 19797 13345 19809 13379
rect 19843 13345 19855 13379
rect 19797 13339 19855 13345
rect 15703 13280 16252 13308
rect 16592 13280 17540 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 10244 13212 11652 13240
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 16592 13240 16620 13280
rect 17586 13268 17592 13320
rect 17644 13308 17650 13320
rect 17644 13280 19564 13308
rect 17644 13268 17650 13280
rect 16758 13249 16764 13252
rect 14976 13212 16620 13240
rect 14976 13200 14982 13212
rect 16752 13203 16764 13249
rect 16758 13200 16764 13203
rect 16816 13200 16822 13252
rect 18046 13200 18052 13252
rect 18104 13240 18110 13252
rect 18141 13243 18199 13249
rect 18141 13240 18153 13243
rect 18104 13212 18153 13240
rect 18104 13200 18110 13212
rect 18141 13209 18153 13212
rect 18187 13209 18199 13243
rect 19536 13240 19564 13280
rect 19610 13268 19616 13320
rect 19668 13268 19674 13320
rect 19812 13240 19840 13339
rect 21174 13336 21180 13388
rect 21232 13336 21238 13388
rect 21358 13336 21364 13388
rect 21416 13336 21422 13388
rect 22922 13376 22928 13388
rect 21468 13348 22928 13376
rect 20438 13268 20444 13320
rect 20496 13268 20502 13320
rect 20806 13268 20812 13320
rect 20864 13308 20870 13320
rect 21085 13311 21143 13317
rect 21085 13308 21097 13311
rect 20864 13280 21097 13308
rect 20864 13268 20870 13280
rect 21085 13277 21097 13280
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 20990 13240 20996 13252
rect 19536 13212 20996 13240
rect 18141 13203 18199 13209
rect 20990 13200 20996 13212
rect 21048 13240 21054 13252
rect 21468 13240 21496 13348
rect 22922 13336 22928 13348
rect 22980 13336 22986 13388
rect 22646 13268 22652 13320
rect 22704 13268 22710 13320
rect 22738 13268 22744 13320
rect 22796 13268 22802 13320
rect 23952 13240 23980 13416
rect 24026 13336 24032 13388
rect 24084 13376 24090 13388
rect 24949 13379 25007 13385
rect 24949 13376 24961 13379
rect 24084 13348 24961 13376
rect 24084 13336 24090 13348
rect 24949 13345 24961 13348
rect 24995 13345 25007 13379
rect 24949 13339 25007 13345
rect 25498 13336 25504 13388
rect 25556 13336 25562 13388
rect 24857 13311 24915 13317
rect 24857 13277 24869 13311
rect 24903 13308 24915 13311
rect 25516 13308 25544 13336
rect 24903 13280 25544 13308
rect 25608 13308 25636 13416
rect 26344 13416 27384 13444
rect 26344 13388 26372 13416
rect 26326 13336 26332 13388
rect 26384 13336 26390 13388
rect 27356 13376 27384 13416
rect 28077 13413 28089 13447
rect 28123 13444 28135 13447
rect 29086 13444 29092 13456
rect 28123 13416 29092 13444
rect 28123 13413 28135 13416
rect 28077 13407 28135 13413
rect 29086 13404 29092 13416
rect 29144 13404 29150 13456
rect 31128 13416 31524 13444
rect 28629 13379 28687 13385
rect 28629 13376 28641 13379
rect 26436 13348 27292 13376
rect 27356 13348 28641 13376
rect 26436 13308 26464 13348
rect 25608 13280 26464 13308
rect 24903 13277 24915 13280
rect 24857 13271 24915 13277
rect 27154 13268 27160 13320
rect 27212 13268 27218 13320
rect 27264 13308 27292 13348
rect 28629 13345 28641 13348
rect 28675 13376 28687 13379
rect 31128 13376 31156 13416
rect 31496 13385 31524 13416
rect 28675 13348 31156 13376
rect 31481 13379 31539 13385
rect 28675 13345 28687 13348
rect 28629 13339 28687 13345
rect 31481 13345 31493 13379
rect 31527 13376 31539 13379
rect 32030 13376 32036 13388
rect 31527 13348 32036 13376
rect 31527 13345 31539 13348
rect 31481 13339 31539 13345
rect 32030 13336 32036 13348
rect 32088 13336 32094 13388
rect 32950 13336 32956 13388
rect 33008 13376 33014 13388
rect 33321 13379 33379 13385
rect 33321 13376 33333 13379
rect 33008 13348 33333 13376
rect 33008 13336 33014 13348
rect 33321 13345 33333 13348
rect 33367 13345 33379 13379
rect 33321 13339 33379 13345
rect 28994 13308 29000 13320
rect 27264 13280 29000 13308
rect 28994 13268 29000 13280
rect 29052 13268 29058 13320
rect 29086 13268 29092 13320
rect 29144 13268 29150 13320
rect 32858 13268 32864 13320
rect 32916 13308 32922 13320
rect 33045 13311 33103 13317
rect 33045 13308 33057 13311
rect 32916 13280 33057 13308
rect 32916 13268 32922 13280
rect 33045 13277 33057 13280
rect 33091 13277 33103 13311
rect 33045 13271 33103 13277
rect 21048 13212 21496 13240
rect 21551 13212 23980 13240
rect 21048 13200 21054 13212
rect 5442 13132 5448 13184
rect 5500 13132 5506 13184
rect 7009 13175 7067 13181
rect 7009 13141 7021 13175
rect 7055 13172 7067 13175
rect 7374 13172 7380 13184
rect 7055 13144 7380 13172
rect 7055 13141 7067 13144
rect 7009 13135 7067 13141
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 8294 13132 8300 13184
rect 8352 13132 8358 13184
rect 10410 13132 10416 13184
rect 10468 13172 10474 13184
rect 10505 13175 10563 13181
rect 10505 13172 10517 13175
rect 10468 13144 10517 13172
rect 10468 13132 10474 13144
rect 10505 13141 10517 13144
rect 10551 13141 10563 13175
rect 10505 13135 10563 13141
rect 10594 13132 10600 13184
rect 10652 13172 10658 13184
rect 15010 13172 15016 13184
rect 10652 13144 15016 13172
rect 10652 13132 10658 13144
rect 15010 13132 15016 13144
rect 15068 13132 15074 13184
rect 15286 13132 15292 13184
rect 15344 13172 15350 13184
rect 16390 13172 16396 13184
rect 15344 13144 16396 13172
rect 15344 13132 15350 13144
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 19058 13132 19064 13184
rect 19116 13172 19122 13184
rect 21551 13172 21579 13212
rect 24302 13200 24308 13252
rect 24360 13240 24366 13252
rect 30561 13243 30619 13249
rect 30561 13240 30573 13243
rect 24360 13212 30573 13240
rect 24360 13200 24366 13212
rect 30561 13209 30573 13212
rect 30607 13240 30619 13243
rect 31297 13243 31355 13249
rect 31297 13240 31309 13243
rect 30607 13212 31309 13240
rect 30607 13209 30619 13212
rect 30561 13203 30619 13209
rect 31297 13209 31309 13212
rect 31343 13240 31355 13243
rect 31938 13240 31944 13252
rect 31343 13212 31944 13240
rect 31343 13209 31355 13212
rect 31297 13203 31355 13209
rect 31938 13200 31944 13212
rect 31996 13200 32002 13252
rect 19116 13144 21579 13172
rect 19116 13132 19122 13144
rect 22094 13132 22100 13184
rect 22152 13172 22158 13184
rect 22738 13172 22744 13184
rect 22152 13144 22744 13172
rect 22152 13132 22158 13144
rect 22738 13132 22744 13144
rect 22796 13172 22802 13184
rect 23382 13172 23388 13184
rect 22796 13144 23388 13172
rect 22796 13132 22802 13144
rect 23382 13132 23388 13144
rect 23440 13132 23446 13184
rect 24762 13132 24768 13184
rect 24820 13132 24826 13184
rect 25590 13132 25596 13184
rect 25648 13172 25654 13184
rect 25777 13175 25835 13181
rect 25777 13172 25789 13175
rect 25648 13144 25789 13172
rect 25648 13132 25654 13144
rect 25777 13141 25789 13144
rect 25823 13141 25835 13175
rect 25777 13135 25835 13141
rect 26142 13132 26148 13184
rect 26200 13132 26206 13184
rect 26234 13132 26240 13184
rect 26292 13132 26298 13184
rect 26973 13175 27031 13181
rect 26973 13141 26985 13175
rect 27019 13172 27031 13175
rect 27246 13172 27252 13184
rect 27019 13144 27252 13172
rect 27019 13141 27031 13144
rect 26973 13135 27031 13141
rect 27246 13132 27252 13144
rect 27304 13132 27310 13184
rect 27982 13132 27988 13184
rect 28040 13172 28046 13184
rect 28442 13172 28448 13184
rect 28040 13144 28448 13172
rect 28040 13132 28046 13144
rect 28442 13132 28448 13144
rect 28500 13132 28506 13184
rect 28534 13132 28540 13184
rect 28592 13132 28598 13184
rect 28994 13132 29000 13184
rect 29052 13172 29058 13184
rect 30098 13172 30104 13184
rect 29052 13144 30104 13172
rect 29052 13132 29058 13144
rect 30098 13132 30104 13144
rect 30156 13132 30162 13184
rect 31110 13132 31116 13184
rect 31168 13172 31174 13184
rect 31389 13175 31447 13181
rect 31389 13172 31401 13175
rect 31168 13144 31401 13172
rect 31168 13132 31174 13144
rect 31389 13141 31401 13144
rect 31435 13141 31447 13175
rect 31389 13135 31447 13141
rect 1104 13082 36800 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 36800 13082
rect 1104 13008 36800 13030
rect 7561 12971 7619 12977
rect 7561 12937 7573 12971
rect 7607 12968 7619 12971
rect 7742 12968 7748 12980
rect 7607 12940 7748 12968
rect 7607 12937 7619 12940
rect 7561 12931 7619 12937
rect 7742 12928 7748 12940
rect 7800 12968 7806 12980
rect 8665 12971 8723 12977
rect 8665 12968 8677 12971
rect 7800 12940 8677 12968
rect 7800 12928 7806 12940
rect 8665 12937 8677 12940
rect 8711 12937 8723 12971
rect 8665 12931 8723 12937
rect 8757 12971 8815 12977
rect 8757 12937 8769 12971
rect 8803 12937 8815 12971
rect 8757 12931 8815 12937
rect 5350 12860 5356 12912
rect 5408 12900 5414 12912
rect 8772 12900 8800 12931
rect 8846 12928 8852 12980
rect 8904 12928 8910 12980
rect 13633 12971 13691 12977
rect 13633 12937 13645 12971
rect 13679 12968 13691 12971
rect 13817 12971 13875 12977
rect 13817 12968 13829 12971
rect 13679 12940 13829 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 13817 12937 13829 12940
rect 13863 12937 13875 12971
rect 16669 12971 16727 12977
rect 13817 12931 13875 12937
rect 14108 12940 15884 12968
rect 9766 12900 9772 12912
rect 5408 12872 8708 12900
rect 8772 12872 9772 12900
rect 5408 12860 5414 12872
rect 1489 12835 1547 12841
rect 1489 12801 1501 12835
rect 1535 12832 1547 12835
rect 4985 12835 5043 12841
rect 4985 12832 4997 12835
rect 1535 12804 4997 12832
rect 1535 12801 1547 12804
rect 1489 12795 1547 12801
rect 4985 12801 4997 12804
rect 5031 12832 5043 12835
rect 5261 12835 5319 12841
rect 5031 12804 5212 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5184 12696 5212 12804
rect 5261 12801 5273 12835
rect 5307 12832 5319 12835
rect 5442 12832 5448 12844
rect 5307 12804 5448 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 6822 12832 6828 12844
rect 6687 12804 6828 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7374 12832 7380 12844
rect 7156 12804 7380 12832
rect 7156 12792 7162 12804
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 7607 12804 7972 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 5629 12767 5687 12773
rect 5629 12733 5641 12767
rect 5675 12764 5687 12767
rect 5902 12764 5908 12776
rect 5675 12736 5908 12764
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 6362 12724 6368 12776
rect 6420 12724 6426 12776
rect 7650 12724 7656 12776
rect 7708 12724 7714 12776
rect 7944 12773 7972 12804
rect 8570 12792 8576 12844
rect 8628 12792 8634 12844
rect 8680 12832 8708 12872
rect 9766 12860 9772 12872
rect 9824 12860 9830 12912
rect 14108 12900 14136 12940
rect 10980 12872 14136 12900
rect 15105 12903 15163 12909
rect 8680 12804 9076 12832
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12764 7987 12767
rect 8018 12764 8024 12776
rect 7975 12736 8024 12764
rect 7975 12733 7987 12736
rect 7929 12727 7987 12733
rect 8018 12724 8024 12736
rect 8076 12724 8082 12776
rect 8938 12724 8944 12776
rect 8996 12724 9002 12776
rect 9048 12764 9076 12804
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9398 12832 9404 12844
rect 9180 12804 9404 12832
rect 9180 12792 9186 12804
rect 9398 12792 9404 12804
rect 9456 12792 9462 12844
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 10870 12832 10876 12844
rect 9631 12804 10876 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 10980 12764 11008 12872
rect 15105 12869 15117 12903
rect 15151 12900 15163 12903
rect 15378 12900 15384 12912
rect 15151 12872 15384 12900
rect 15151 12869 15163 12872
rect 15105 12863 15163 12869
rect 15378 12860 15384 12872
rect 15436 12860 15442 12912
rect 15856 12909 15884 12940
rect 16669 12937 16681 12971
rect 16715 12968 16727 12971
rect 16758 12968 16764 12980
rect 16715 12940 16764 12968
rect 16715 12937 16727 12940
rect 16669 12931 16727 12937
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 21174 12928 21180 12980
rect 21232 12968 21238 12980
rect 24578 12968 24584 12980
rect 21232 12940 24584 12968
rect 21232 12928 21238 12940
rect 24578 12928 24584 12940
rect 24636 12968 24642 12980
rect 24762 12968 24768 12980
rect 24636 12940 24768 12968
rect 24636 12928 24642 12940
rect 24762 12928 24768 12940
rect 24820 12928 24826 12980
rect 25409 12971 25467 12977
rect 25409 12937 25421 12971
rect 25455 12968 25467 12971
rect 28258 12968 28264 12980
rect 25455 12940 25820 12968
rect 25455 12937 25467 12940
rect 25409 12931 25467 12937
rect 15841 12903 15899 12909
rect 15841 12869 15853 12903
rect 15887 12869 15899 12903
rect 25792 12900 25820 12940
rect 26804 12940 28264 12968
rect 25792 12872 26004 12900
rect 15841 12863 15899 12869
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 13265 12835 13323 12841
rect 13265 12832 13277 12835
rect 11112 12804 13277 12832
rect 11112 12792 11118 12804
rect 13265 12801 13277 12804
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 13449 12835 13507 12841
rect 13449 12801 13461 12835
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 9048 12736 11008 12764
rect 12158 12696 12164 12708
rect 5184 12668 12164 12696
rect 12158 12656 12164 12668
rect 12216 12656 12222 12708
rect 13464 12696 13492 12795
rect 13722 12792 13728 12844
rect 13780 12792 13786 12844
rect 13906 12792 13912 12844
rect 13964 12832 13970 12844
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13964 12804 14197 12832
rect 13964 12792 13970 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 14918 12792 14924 12844
rect 14976 12792 14982 12844
rect 15010 12792 15016 12844
rect 15068 12832 15074 12844
rect 15197 12835 15255 12841
rect 15197 12832 15209 12835
rect 15068 12804 15209 12832
rect 15068 12792 15074 12804
rect 15197 12801 15209 12804
rect 15243 12801 15255 12835
rect 15197 12795 15255 12801
rect 15286 12792 15292 12844
rect 15344 12792 15350 12844
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12801 15623 12835
rect 15565 12795 15623 12801
rect 13998 12724 14004 12776
rect 14056 12724 14062 12776
rect 14090 12724 14096 12776
rect 14148 12724 14154 12776
rect 14274 12724 14280 12776
rect 14332 12724 14338 12776
rect 15580 12764 15608 12795
rect 15746 12792 15752 12844
rect 15804 12792 15810 12844
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12832 15991 12835
rect 16114 12832 16120 12844
rect 15979 12804 16120 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 16114 12792 16120 12804
rect 16172 12792 16178 12844
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 18322 12792 18328 12844
rect 18380 12832 18386 12844
rect 24302 12832 24308 12844
rect 18380 12804 24308 12832
rect 18380 12792 18386 12804
rect 24302 12792 24308 12804
rect 24360 12792 24366 12844
rect 25590 12792 25596 12844
rect 25648 12792 25654 12844
rect 25976 12841 26004 12872
rect 25961 12835 26019 12841
rect 25961 12801 25973 12835
rect 26007 12801 26019 12835
rect 25961 12795 26019 12801
rect 26142 12792 26148 12844
rect 26200 12832 26206 12844
rect 26804 12841 26832 12940
rect 28258 12928 28264 12940
rect 28316 12928 28322 12980
rect 28442 12928 28448 12980
rect 28500 12968 28506 12980
rect 29270 12968 29276 12980
rect 28500 12940 29276 12968
rect 28500 12928 28506 12940
rect 29270 12928 29276 12940
rect 29328 12928 29334 12980
rect 29638 12928 29644 12980
rect 29696 12968 29702 12980
rect 30285 12971 30343 12977
rect 30285 12968 30297 12971
rect 29696 12940 30297 12968
rect 29696 12928 29702 12940
rect 30285 12937 30297 12940
rect 30331 12937 30343 12971
rect 30285 12931 30343 12937
rect 32769 12971 32827 12977
rect 32769 12937 32781 12971
rect 32815 12937 32827 12971
rect 32769 12931 32827 12937
rect 28166 12900 28172 12912
rect 26988 12872 28172 12900
rect 26789 12835 26847 12841
rect 26789 12832 26801 12835
rect 26200 12804 26801 12832
rect 26200 12792 26206 12804
rect 26789 12801 26801 12804
rect 26835 12801 26847 12835
rect 26789 12795 26847 12801
rect 17126 12764 17132 12776
rect 15580 12736 17132 12764
rect 17126 12724 17132 12736
rect 17184 12764 17190 12776
rect 18233 12767 18291 12773
rect 17184 12736 18184 12764
rect 17184 12724 17190 12736
rect 15473 12699 15531 12705
rect 15473 12696 15485 12699
rect 13464 12668 15485 12696
rect 15473 12665 15485 12668
rect 15519 12665 15531 12699
rect 15473 12659 15531 12665
rect 15746 12656 15752 12708
rect 15804 12696 15810 12708
rect 18156 12696 18184 12736
rect 18233 12733 18245 12767
rect 18279 12764 18291 12767
rect 18414 12764 18420 12776
rect 18279 12736 18420 12764
rect 18279 12733 18291 12736
rect 18233 12727 18291 12733
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 25406 12764 25412 12776
rect 18524 12736 25412 12764
rect 18524 12696 18552 12736
rect 25406 12724 25412 12736
rect 25464 12724 25470 12776
rect 26988 12773 27016 12872
rect 28166 12860 28172 12872
rect 28224 12860 28230 12912
rect 32784 12900 32812 12931
rect 33318 12928 33324 12980
rect 33376 12968 33382 12980
rect 33594 12968 33600 12980
rect 33376 12940 33600 12968
rect 33376 12928 33382 12940
rect 33594 12928 33600 12940
rect 33652 12968 33658 12980
rect 34057 12971 34115 12977
rect 34057 12968 34069 12971
rect 33652 12940 34069 12968
rect 33652 12928 33658 12940
rect 34057 12937 34069 12940
rect 34103 12937 34115 12971
rect 34057 12931 34115 12937
rect 35986 12928 35992 12980
rect 36044 12928 36050 12980
rect 32784 12872 33364 12900
rect 27246 12792 27252 12844
rect 27304 12792 27310 12844
rect 29178 12841 29184 12844
rect 29172 12795 29184 12841
rect 29178 12792 29184 12795
rect 29236 12792 29242 12844
rect 32950 12792 32956 12844
rect 33008 12792 33014 12844
rect 33042 12792 33048 12844
rect 33100 12792 33106 12844
rect 33336 12841 33364 12872
rect 33321 12835 33379 12841
rect 33321 12801 33333 12835
rect 33367 12801 33379 12835
rect 33321 12795 33379 12801
rect 34698 12792 34704 12844
rect 34756 12832 34762 12844
rect 34865 12835 34923 12841
rect 34865 12832 34877 12835
rect 34756 12804 34877 12832
rect 34756 12792 34762 12804
rect 34865 12801 34877 12804
rect 34911 12801 34923 12835
rect 34865 12795 34923 12801
rect 25685 12767 25743 12773
rect 25685 12733 25697 12767
rect 25731 12733 25743 12767
rect 25685 12727 25743 12733
rect 26973 12767 27031 12773
rect 26973 12733 26985 12767
rect 27019 12733 27031 12767
rect 26973 12727 27031 12733
rect 28905 12767 28963 12773
rect 28905 12733 28917 12767
rect 28951 12733 28963 12767
rect 28905 12727 28963 12733
rect 34609 12767 34667 12773
rect 34609 12733 34621 12767
rect 34655 12733 34667 12767
rect 34609 12727 34667 12733
rect 15804 12668 17356 12696
rect 18156 12668 18552 12696
rect 15804 12656 15810 12668
rect 1578 12588 1584 12640
rect 1636 12588 1642 12640
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 13998 12628 14004 12640
rect 8352 12600 14004 12628
rect 8352 12588 8358 12600
rect 13998 12588 14004 12600
rect 14056 12588 14062 12640
rect 15654 12588 15660 12640
rect 15712 12628 15718 12640
rect 16117 12631 16175 12637
rect 16117 12628 16129 12631
rect 15712 12600 16129 12628
rect 15712 12588 15718 12600
rect 16117 12597 16129 12600
rect 16163 12597 16175 12631
rect 17328 12628 17356 12668
rect 18598 12656 18604 12708
rect 18656 12656 18662 12708
rect 18693 12631 18751 12637
rect 18693 12628 18705 12631
rect 17328 12600 18705 12628
rect 16117 12591 16175 12597
rect 18693 12597 18705 12600
rect 18739 12628 18751 12631
rect 18874 12628 18880 12640
rect 18739 12600 18880 12628
rect 18739 12597 18751 12600
rect 18693 12591 18751 12597
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 22738 12588 22744 12640
rect 22796 12628 22802 12640
rect 24210 12628 24216 12640
rect 22796 12600 24216 12628
rect 22796 12588 22802 12600
rect 24210 12588 24216 12600
rect 24268 12588 24274 12640
rect 25700 12628 25728 12727
rect 26988 12628 27016 12727
rect 25700 12600 27016 12628
rect 27614 12588 27620 12640
rect 27672 12628 27678 12640
rect 27982 12628 27988 12640
rect 27672 12600 27988 12628
rect 27672 12588 27678 12600
rect 27982 12588 27988 12600
rect 28040 12588 28046 12640
rect 28920 12628 28948 12727
rect 30208 12668 31754 12696
rect 30208 12628 30236 12668
rect 28920 12600 30236 12628
rect 31726 12628 31754 12668
rect 34624 12640 34652 12727
rect 34606 12628 34612 12640
rect 31726 12600 34612 12628
rect 34606 12588 34612 12600
rect 34664 12588 34670 12640
rect 1104 12538 36800 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 36800 12538
rect 1104 12464 36800 12486
rect 8938 12384 8944 12436
rect 8996 12424 9002 12436
rect 9217 12427 9275 12433
rect 9217 12424 9229 12427
rect 8996 12396 9229 12424
rect 8996 12384 9002 12396
rect 9217 12393 9229 12396
rect 9263 12393 9275 12427
rect 9217 12387 9275 12393
rect 9493 12427 9551 12433
rect 9493 12393 9505 12427
rect 9539 12424 9551 12427
rect 11422 12424 11428 12436
rect 9539 12396 11428 12424
rect 9539 12393 9551 12396
rect 9493 12387 9551 12393
rect 7742 12248 7748 12300
rect 7800 12248 7806 12300
rect 9232 12288 9260 12387
rect 11422 12384 11428 12396
rect 11480 12424 11486 12436
rect 11606 12424 11612 12436
rect 11480 12396 11612 12424
rect 11480 12384 11486 12396
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 12529 12427 12587 12433
rect 12529 12393 12541 12427
rect 12575 12393 12587 12427
rect 12529 12387 12587 12393
rect 9582 12316 9588 12368
rect 9640 12316 9646 12368
rect 10318 12356 10324 12368
rect 10152 12328 10324 12356
rect 10152 12297 10180 12328
rect 10318 12316 10324 12328
rect 10376 12316 10382 12368
rect 11149 12359 11207 12365
rect 11149 12325 11161 12359
rect 11195 12356 11207 12359
rect 12544 12356 12572 12387
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 18877 12427 18935 12433
rect 18877 12424 18889 12427
rect 17000 12396 18889 12424
rect 17000 12384 17006 12396
rect 18877 12393 18889 12396
rect 18923 12393 18935 12427
rect 18877 12387 18935 12393
rect 19242 12384 19248 12436
rect 19300 12424 19306 12436
rect 21082 12424 21088 12436
rect 19300 12396 21088 12424
rect 19300 12384 19306 12396
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 21192 12396 22876 12424
rect 21192 12356 21220 12396
rect 11195 12328 12572 12356
rect 19076 12328 21220 12356
rect 22848 12356 22876 12396
rect 22922 12384 22928 12436
rect 22980 12384 22986 12436
rect 25777 12427 25835 12433
rect 25777 12424 25789 12427
rect 24044 12396 25789 12424
rect 24044 12368 24072 12396
rect 25777 12393 25789 12396
rect 25823 12393 25835 12427
rect 25777 12387 25835 12393
rect 27065 12427 27123 12433
rect 27065 12393 27077 12427
rect 27111 12424 27123 12427
rect 27154 12424 27160 12436
rect 27111 12396 27160 12424
rect 27111 12393 27123 12396
rect 27065 12387 27123 12393
rect 27154 12384 27160 12396
rect 27212 12384 27218 12436
rect 29178 12384 29184 12436
rect 29236 12384 29242 12436
rect 29270 12384 29276 12436
rect 29328 12424 29334 12436
rect 29914 12424 29920 12436
rect 29328 12396 29920 12424
rect 29328 12384 29334 12396
rect 29914 12384 29920 12396
rect 29972 12384 29978 12436
rect 30006 12384 30012 12436
rect 30064 12424 30070 12436
rect 30064 12396 31892 12424
rect 30064 12384 30070 12396
rect 24026 12356 24032 12368
rect 22848 12328 24032 12356
rect 11195 12325 11207 12328
rect 11149 12319 11207 12325
rect 9677 12291 9735 12297
rect 9677 12288 9689 12291
rect 9232 12260 9689 12288
rect 9677 12257 9689 12260
rect 9723 12288 9735 12291
rect 10137 12291 10195 12297
rect 9723 12260 9996 12288
rect 9723 12257 9735 12260
rect 9677 12251 9735 12257
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12220 4675 12223
rect 5718 12220 5724 12232
rect 4663 12192 5724 12220
rect 4663 12189 4675 12192
rect 4617 12183 4675 12189
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 5997 12223 6055 12229
rect 5997 12189 6009 12223
rect 6043 12220 6055 12223
rect 6822 12220 6828 12232
rect 6043 12192 6828 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 4706 12112 4712 12164
rect 4764 12152 4770 12164
rect 6012 12152 6040 12183
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7374 12220 7380 12232
rect 7156 12192 7380 12220
rect 7156 12180 7162 12192
rect 7374 12180 7380 12192
rect 7432 12180 7438 12232
rect 7469 12223 7527 12229
rect 7469 12189 7481 12223
rect 7515 12220 7527 12223
rect 7558 12220 7564 12232
rect 7515 12192 7564 12220
rect 7515 12189 7527 12192
rect 7469 12183 7527 12189
rect 7558 12180 7564 12192
rect 7616 12220 7622 12232
rect 7929 12223 7987 12229
rect 7929 12220 7941 12223
rect 7616 12192 7941 12220
rect 7616 12180 7622 12192
rect 7929 12189 7941 12192
rect 7975 12220 7987 12223
rect 8570 12220 8576 12232
rect 7975 12192 8576 12220
rect 7975 12189 7987 12192
rect 7929 12183 7987 12189
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 4764 12124 6040 12152
rect 4764 12112 4770 12124
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 7285 12155 7343 12161
rect 7285 12152 7297 12155
rect 6972 12124 7297 12152
rect 6972 12112 6978 12124
rect 7285 12121 7297 12124
rect 7331 12152 7343 12155
rect 7834 12152 7840 12164
rect 7331 12124 7840 12152
rect 7331 12121 7343 12124
rect 7285 12115 7343 12121
rect 7834 12112 7840 12124
rect 7892 12112 7898 12164
rect 8202 12112 8208 12164
rect 8260 12152 8266 12164
rect 9324 12152 9352 12183
rect 8260 12124 9352 12152
rect 9416 12152 9444 12183
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 9968 12229 9996 12260
rect 10137 12257 10149 12291
rect 10183 12257 10195 12291
rect 10137 12251 10195 12257
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12288 10287 12291
rect 10870 12288 10876 12300
rect 10275 12260 10876 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 10152 12152 10180 12251
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 11072 12260 11560 12288
rect 10502 12180 10508 12232
rect 10560 12180 10566 12232
rect 10520 12152 10548 12180
rect 9416 12124 10180 12152
rect 10244 12124 10548 12152
rect 8260 12112 8266 12124
rect 4985 12087 5043 12093
rect 4985 12053 4997 12087
rect 5031 12084 5043 12087
rect 5350 12084 5356 12096
rect 5031 12056 5356 12084
rect 5031 12053 5043 12056
rect 4985 12047 5043 12053
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 8113 12087 8171 12093
rect 8113 12053 8125 12087
rect 8159 12084 8171 12087
rect 8938 12084 8944 12096
rect 8159 12056 8944 12084
rect 8159 12053 8171 12056
rect 8113 12047 8171 12053
rect 8938 12044 8944 12056
rect 8996 12044 9002 12096
rect 9324 12084 9352 12124
rect 10244 12084 10272 12124
rect 9324 12056 10272 12084
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 11072 12084 11100 12260
rect 11422 12180 11428 12232
rect 11480 12180 11486 12232
rect 11532 12229 11560 12260
rect 11790 12248 11796 12300
rect 11848 12248 11854 12300
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12288 12219 12291
rect 12544 12288 12756 12296
rect 12207 12268 16620 12288
rect 12207 12260 12572 12268
rect 12728 12260 16620 12268
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12189 11575 12223
rect 11517 12183 11575 12189
rect 12391 12223 12449 12229
rect 12391 12189 12403 12223
rect 12437 12189 12449 12223
rect 12391 12183 12449 12189
rect 11149 12155 11207 12161
rect 11149 12121 11161 12155
rect 11195 12152 11207 12155
rect 11793 12155 11851 12161
rect 11793 12152 11805 12155
rect 11195 12124 11805 12152
rect 11195 12121 11207 12124
rect 11149 12115 11207 12121
rect 11793 12121 11805 12124
rect 11839 12121 11851 12155
rect 11793 12115 11851 12121
rect 11882 12112 11888 12164
rect 11940 12152 11946 12164
rect 12406 12152 12434 12183
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 15105 12223 15163 12229
rect 15105 12189 15117 12223
rect 15151 12189 15163 12223
rect 15105 12183 15163 12189
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12220 15347 12223
rect 15378 12220 15384 12232
rect 15335 12192 15384 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 11940 12124 12434 12152
rect 11940 12112 11946 12124
rect 11333 12087 11391 12093
rect 11333 12084 11345 12087
rect 10376 12056 11345 12084
rect 10376 12044 10382 12056
rect 11333 12053 11345 12056
rect 11379 12053 11391 12087
rect 12406 12084 12434 12124
rect 12526 12112 12532 12164
rect 12584 12152 12590 12164
rect 13446 12152 13452 12164
rect 12584 12124 13452 12152
rect 12584 12112 12590 12124
rect 13446 12112 13452 12124
rect 13504 12152 13510 12164
rect 14090 12152 14096 12164
rect 13504 12124 14096 12152
rect 13504 12112 13510 12124
rect 14090 12112 14096 12124
rect 14148 12112 14154 12164
rect 15120 12152 15148 12183
rect 15378 12180 15384 12192
rect 15436 12220 15442 12232
rect 15746 12220 15752 12232
rect 15436 12192 15752 12220
rect 15436 12180 15442 12192
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 16114 12180 16120 12232
rect 16172 12180 16178 12232
rect 16592 12220 16620 12260
rect 18598 12248 18604 12300
rect 18656 12288 18662 12300
rect 19076 12288 19104 12328
rect 24026 12316 24032 12328
rect 24084 12316 24090 12368
rect 24118 12316 24124 12368
rect 24176 12316 24182 12368
rect 27264 12328 30328 12356
rect 18656 12260 19104 12288
rect 19904 12260 21220 12288
rect 18656 12248 18662 12260
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 16592 12192 18245 12220
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 18322 12180 18328 12232
rect 18380 12180 18386 12232
rect 18698 12223 18756 12229
rect 18698 12220 18710 12223
rect 18432 12192 18710 12220
rect 15933 12155 15991 12161
rect 15933 12152 15945 12155
rect 15120 12124 15945 12152
rect 15304 12096 15332 12124
rect 15933 12121 15945 12124
rect 15979 12152 15991 12155
rect 16132 12152 16160 12180
rect 17954 12152 17960 12164
rect 15979 12124 17960 12152
rect 15979 12121 15991 12124
rect 15933 12115 15991 12121
rect 17954 12112 17960 12124
rect 18012 12112 18018 12164
rect 18141 12155 18199 12161
rect 18141 12121 18153 12155
rect 18187 12152 18199 12155
rect 18432 12152 18460 12192
rect 18698 12189 18710 12192
rect 18744 12220 18756 12223
rect 18966 12220 18972 12232
rect 18744 12192 18972 12220
rect 18744 12189 18756 12192
rect 18698 12183 18756 12189
rect 18966 12180 18972 12192
rect 19024 12180 19030 12232
rect 19518 12180 19524 12232
rect 19576 12180 19582 12232
rect 19669 12223 19727 12229
rect 19669 12189 19681 12223
rect 19715 12220 19727 12223
rect 19904 12220 19932 12260
rect 19715 12192 19932 12220
rect 19715 12189 19727 12192
rect 19669 12183 19727 12189
rect 19978 12180 19984 12232
rect 20036 12229 20042 12232
rect 20036 12220 20044 12229
rect 21192 12220 21220 12260
rect 21266 12248 21272 12300
rect 21324 12248 21330 12300
rect 23661 12291 23719 12297
rect 23661 12257 23673 12291
rect 23707 12288 23719 12291
rect 24136 12288 24164 12316
rect 24397 12291 24455 12297
rect 24397 12288 24409 12291
rect 23707 12260 24072 12288
rect 24136 12260 24409 12288
rect 23707 12257 23719 12260
rect 23661 12251 23719 12257
rect 21910 12220 21916 12232
rect 20036 12192 20081 12220
rect 21192 12192 21916 12220
rect 20036 12183 20044 12192
rect 20036 12180 20042 12183
rect 21910 12180 21916 12192
rect 21968 12180 21974 12232
rect 22002 12180 22008 12232
rect 22060 12220 22066 12232
rect 22462 12220 22468 12232
rect 22060 12192 22468 12220
rect 22060 12180 22066 12192
rect 22462 12180 22468 12192
rect 22520 12180 22526 12232
rect 22738 12180 22744 12232
rect 22796 12180 22802 12232
rect 23106 12180 23112 12232
rect 23164 12220 23170 12232
rect 23845 12223 23903 12229
rect 23845 12220 23857 12223
rect 23164 12192 23857 12220
rect 23164 12180 23170 12192
rect 23845 12189 23857 12192
rect 23891 12189 23903 12223
rect 23845 12183 23903 12189
rect 23937 12223 23995 12229
rect 23937 12189 23949 12223
rect 23983 12189 23995 12223
rect 23937 12183 23995 12189
rect 18187 12124 18460 12152
rect 18187 12121 18199 12124
rect 18141 12115 18199 12121
rect 18506 12112 18512 12164
rect 18564 12112 18570 12164
rect 18601 12155 18659 12161
rect 18601 12121 18613 12155
rect 18647 12152 18659 12155
rect 19150 12152 19156 12164
rect 18647 12124 19156 12152
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 19150 12112 19156 12124
rect 19208 12112 19214 12164
rect 19797 12155 19855 12161
rect 19797 12121 19809 12155
rect 19843 12121 19855 12155
rect 19797 12115 19855 12121
rect 13722 12084 13728 12096
rect 12406 12056 13728 12084
rect 11333 12047 11391 12053
rect 13722 12044 13728 12056
rect 13780 12084 13786 12096
rect 14918 12084 14924 12096
rect 13780 12056 14924 12084
rect 13780 12044 13786 12056
rect 14918 12044 14924 12056
rect 14976 12084 14982 12096
rect 15105 12087 15163 12093
rect 15105 12084 15117 12087
rect 14976 12056 15117 12084
rect 14976 12044 14982 12056
rect 15105 12053 15117 12056
rect 15151 12053 15163 12087
rect 15105 12047 15163 12053
rect 15286 12044 15292 12096
rect 15344 12044 15350 12096
rect 16114 12044 16120 12096
rect 16172 12044 16178 12096
rect 18524 12084 18552 12112
rect 19702 12084 19708 12096
rect 18524 12056 19708 12084
rect 19702 12044 19708 12056
rect 19760 12084 19766 12096
rect 19812 12084 19840 12115
rect 19886 12112 19892 12164
rect 19944 12112 19950 12164
rect 21536 12155 21594 12161
rect 21536 12121 21548 12155
rect 21582 12152 21594 12155
rect 21818 12152 21824 12164
rect 21582 12124 21824 12152
rect 21582 12121 21594 12124
rect 21536 12115 21594 12121
rect 21818 12112 21824 12124
rect 21876 12112 21882 12164
rect 22066 12124 23704 12152
rect 19760 12056 19840 12084
rect 20165 12087 20223 12093
rect 19760 12044 19766 12056
rect 20165 12053 20177 12087
rect 20211 12084 20223 12087
rect 22066 12084 22094 12124
rect 20211 12056 22094 12084
rect 20211 12053 20223 12056
rect 20165 12047 20223 12053
rect 22646 12044 22652 12096
rect 22704 12044 22710 12096
rect 23676 12084 23704 12124
rect 23750 12112 23756 12164
rect 23808 12152 23814 12164
rect 23952 12152 23980 12183
rect 23808 12124 23980 12152
rect 24044 12152 24072 12260
rect 24397 12257 24409 12260
rect 24443 12257 24455 12291
rect 24397 12251 24455 12257
rect 24118 12180 24124 12232
rect 24176 12180 24182 12232
rect 24210 12180 24216 12232
rect 24268 12180 24274 12232
rect 27264 12220 27292 12328
rect 27709 12291 27767 12297
rect 27709 12257 27721 12291
rect 27755 12288 27767 12291
rect 29270 12288 29276 12300
rect 27755 12260 29276 12288
rect 27755 12257 27767 12260
rect 27709 12251 27767 12257
rect 29270 12248 29276 12260
rect 29328 12248 29334 12300
rect 29546 12248 29552 12300
rect 29604 12288 29610 12300
rect 30009 12291 30067 12297
rect 30009 12288 30021 12291
rect 29604 12260 30021 12288
rect 29604 12248 29610 12260
rect 30009 12257 30021 12260
rect 30055 12257 30067 12291
rect 30009 12251 30067 12257
rect 30098 12248 30104 12300
rect 30156 12248 30162 12300
rect 30300 12288 30328 12328
rect 30650 12316 30656 12368
rect 30708 12356 30714 12368
rect 31570 12356 31576 12368
rect 30708 12328 31576 12356
rect 30708 12316 30714 12328
rect 31570 12316 31576 12328
rect 31628 12316 31634 12368
rect 31864 12356 31892 12396
rect 32030 12384 32036 12436
rect 32088 12424 32094 12436
rect 32088 12396 32352 12424
rect 32088 12384 32094 12396
rect 32324 12356 32352 12396
rect 32950 12384 32956 12436
rect 33008 12384 33014 12436
rect 34698 12384 34704 12436
rect 34756 12384 34762 12436
rect 31864 12328 32260 12356
rect 32324 12328 33548 12356
rect 30926 12288 30932 12300
rect 30300 12260 30932 12288
rect 30926 12248 30932 12260
rect 30984 12248 30990 12300
rect 32232 12288 32260 12328
rect 33318 12288 33324 12300
rect 31481 12261 31539 12267
rect 24320 12192 27292 12220
rect 27433 12223 27491 12229
rect 24320 12152 24348 12192
rect 27433 12189 27445 12223
rect 27479 12220 27491 12223
rect 27982 12220 27988 12232
rect 27479 12192 27988 12220
rect 27479 12189 27491 12192
rect 27433 12183 27491 12189
rect 27982 12180 27988 12192
rect 28040 12180 28046 12232
rect 29365 12223 29423 12229
rect 29365 12189 29377 12223
rect 29411 12220 29423 12223
rect 29411 12192 29592 12220
rect 29411 12189 29423 12192
rect 29365 12183 29423 12189
rect 24044 12124 24348 12152
rect 23808 12112 23814 12124
rect 24394 12112 24400 12164
rect 24452 12152 24458 12164
rect 24642 12155 24700 12161
rect 24642 12152 24654 12155
rect 24452 12124 24654 12152
rect 24452 12112 24458 12124
rect 24642 12121 24654 12124
rect 24688 12121 24700 12155
rect 27798 12152 27804 12164
rect 24642 12115 24700 12121
rect 24964 12124 27804 12152
rect 24964 12084 24992 12124
rect 27798 12112 27804 12124
rect 27856 12112 27862 12164
rect 23676 12056 24992 12084
rect 26234 12044 26240 12096
rect 26292 12084 26298 12096
rect 27525 12087 27583 12093
rect 27525 12084 27537 12087
rect 26292 12056 27537 12084
rect 26292 12044 26298 12056
rect 27525 12053 27537 12056
rect 27571 12084 27583 12087
rect 27982 12084 27988 12096
rect 27571 12056 27988 12084
rect 27571 12053 27583 12056
rect 27525 12047 27583 12053
rect 27982 12044 27988 12056
rect 28040 12044 28046 12096
rect 29564 12093 29592 12192
rect 29638 12180 29644 12232
rect 29696 12220 29702 12232
rect 31110 12220 31116 12232
rect 29696 12192 31116 12220
rect 29696 12180 29702 12192
rect 31110 12180 31116 12192
rect 31168 12220 31174 12232
rect 31205 12223 31263 12229
rect 31205 12220 31217 12223
rect 31168 12192 31217 12220
rect 31168 12180 31174 12192
rect 31205 12189 31217 12192
rect 31251 12189 31263 12223
rect 31205 12183 31263 12189
rect 31294 12180 31300 12232
rect 31352 12180 31358 12232
rect 31481 12227 31493 12261
rect 31527 12227 31539 12261
rect 32232 12260 33324 12288
rect 33318 12248 33324 12260
rect 33376 12248 33382 12300
rect 33410 12248 33416 12300
rect 33468 12248 33474 12300
rect 33520 12297 33548 12328
rect 33505 12291 33563 12297
rect 33505 12257 33517 12291
rect 33551 12257 33563 12291
rect 33505 12251 33563 12257
rect 31481 12221 31539 12227
rect 31496 12152 31524 12221
rect 31570 12180 31576 12232
rect 31628 12216 31634 12232
rect 31941 12223 31999 12229
rect 31941 12220 31953 12223
rect 31680 12216 31953 12220
rect 31628 12192 31953 12216
rect 31628 12188 31708 12192
rect 31941 12189 31953 12192
rect 31987 12189 31999 12223
rect 31628 12180 31634 12188
rect 31941 12183 31999 12189
rect 32122 12180 32128 12232
rect 32180 12180 32186 12232
rect 33336 12161 33364 12248
rect 34882 12180 34888 12232
rect 34940 12180 34946 12232
rect 35161 12223 35219 12229
rect 35161 12189 35173 12223
rect 35207 12220 35219 12223
rect 35986 12220 35992 12232
rect 35207 12192 35992 12220
rect 35207 12189 35219 12192
rect 35161 12183 35219 12189
rect 35986 12180 35992 12192
rect 36044 12180 36050 12232
rect 33321 12155 33379 12161
rect 31496 12124 31984 12152
rect 31956 12096 31984 12124
rect 33321 12121 33333 12155
rect 33367 12121 33379 12155
rect 33321 12115 33379 12121
rect 29549 12087 29607 12093
rect 29549 12053 29561 12087
rect 29595 12053 29607 12087
rect 29549 12047 29607 12053
rect 29914 12044 29920 12096
rect 29972 12044 29978 12096
rect 30282 12044 30288 12096
rect 30340 12084 30346 12096
rect 31481 12087 31539 12093
rect 31481 12084 31493 12087
rect 30340 12056 31493 12084
rect 30340 12044 30346 12056
rect 31481 12053 31493 12056
rect 31527 12053 31539 12087
rect 31481 12047 31539 12053
rect 31938 12044 31944 12096
rect 31996 12044 32002 12096
rect 32030 12044 32036 12096
rect 32088 12044 32094 12096
rect 34790 12044 34796 12096
rect 34848 12084 34854 12096
rect 35069 12087 35127 12093
rect 35069 12084 35081 12087
rect 34848 12056 35081 12084
rect 34848 12044 34854 12056
rect 35069 12053 35081 12056
rect 35115 12053 35127 12087
rect 35069 12047 35127 12053
rect 1104 11994 36800 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 36800 11994
rect 1104 11920 36800 11942
rect 7193 11883 7251 11889
rect 7193 11849 7205 11883
rect 7239 11880 7251 11883
rect 7742 11880 7748 11892
rect 7239 11852 7748 11880
rect 7239 11849 7251 11852
rect 7193 11843 7251 11849
rect 7742 11840 7748 11852
rect 7800 11880 7806 11892
rect 7800 11852 8331 11880
rect 7800 11840 7806 11852
rect 4614 11812 4620 11824
rect 3896 11784 4620 11812
rect 3896 11753 3924 11784
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 7558 11772 7564 11824
rect 7616 11772 7622 11824
rect 7653 11815 7711 11821
rect 7653 11781 7665 11815
rect 7699 11812 7711 11815
rect 8202 11812 8208 11824
rect 7699 11784 8208 11812
rect 7699 11781 7711 11784
rect 7653 11775 7711 11781
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 3881 11747 3939 11753
rect 3881 11713 3893 11747
rect 3927 11713 3939 11747
rect 3881 11707 3939 11713
rect 4154 11704 4160 11756
rect 4212 11704 4218 11756
rect 6914 11704 6920 11756
rect 6972 11704 6978 11756
rect 7009 11747 7067 11753
rect 7009 11713 7021 11747
rect 7055 11744 7067 11747
rect 7374 11744 7380 11756
rect 7055 11716 7380 11744
rect 7055 11713 7067 11716
rect 7009 11707 7067 11713
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11744 7527 11747
rect 7515 11716 7696 11744
rect 7515 11713 7527 11716
rect 7469 11707 7527 11713
rect 7668 11608 7696 11716
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 7837 11747 7895 11753
rect 7837 11744 7849 11747
rect 7800 11716 7849 11744
rect 7800 11704 7806 11716
rect 7837 11713 7849 11716
rect 7883 11713 7895 11747
rect 7837 11707 7895 11713
rect 7926 11704 7932 11756
rect 7984 11704 7990 11756
rect 8303 11744 8331 11852
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 11698 11880 11704 11892
rect 8444 11852 11704 11880
rect 8444 11840 8450 11852
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 11793 11883 11851 11889
rect 11793 11849 11805 11883
rect 11839 11880 11851 11883
rect 12250 11880 12256 11892
rect 11839 11852 12256 11880
rect 11839 11849 11851 11852
rect 11793 11843 11851 11849
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 12400 11840 12434 11880
rect 12618 11840 12624 11892
rect 12676 11880 12682 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 12676 11852 12725 11880
rect 12676 11840 12682 11852
rect 12713 11849 12725 11852
rect 12759 11849 12771 11883
rect 12713 11843 12771 11849
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 12860 11852 14044 11880
rect 12860 11840 12866 11852
rect 9122 11772 9128 11824
rect 9180 11812 9186 11824
rect 9309 11815 9367 11821
rect 9309 11812 9321 11815
rect 9180 11784 9321 11812
rect 9180 11772 9186 11784
rect 9309 11781 9321 11784
rect 9355 11781 9367 11815
rect 9309 11775 9367 11781
rect 12069 11815 12127 11821
rect 12069 11781 12081 11815
rect 12115 11812 12127 11815
rect 12406 11812 12434 11840
rect 12115 11784 13216 11812
rect 12115 11781 12127 11784
rect 12069 11775 12127 11781
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 8303 11716 8493 11744
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 10410 11704 10416 11756
rect 10468 11704 10474 11756
rect 10502 11704 10508 11756
rect 10560 11744 10566 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 10560 11716 11713 11744
rect 10560 11704 10566 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 8202 11636 8208 11688
rect 8260 11636 8266 11688
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 8570 11676 8576 11688
rect 8435 11648 8576 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 8312 11608 8340 11639
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 10318 11636 10324 11688
rect 10376 11636 10382 11688
rect 9122 11608 9128 11620
rect 7668 11580 9128 11608
rect 9122 11568 9128 11580
rect 9180 11568 9186 11620
rect 9677 11611 9735 11617
rect 9677 11577 9689 11611
rect 9723 11608 9735 11611
rect 10520 11608 10548 11704
rect 11716 11676 11744 11707
rect 12176 11676 12204 11707
rect 11716 11648 12204 11676
rect 12360 11676 12388 11707
rect 12434 11704 12440 11756
rect 12492 11704 12498 11756
rect 12526 11704 12532 11756
rect 12584 11704 12590 11756
rect 13078 11704 13084 11756
rect 13136 11704 13142 11756
rect 13188 11744 13216 11784
rect 14016 11753 14044 11852
rect 14274 11840 14280 11892
rect 14332 11880 14338 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 14332 11852 14381 11880
rect 14332 11840 14338 11852
rect 14369 11849 14381 11852
rect 14415 11849 14427 11883
rect 14369 11843 14427 11849
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 18012 11852 18368 11880
rect 18012 11840 18018 11852
rect 15289 11815 15347 11821
rect 15289 11781 15301 11815
rect 15335 11812 15347 11815
rect 18141 11815 18199 11821
rect 15335 11784 16160 11812
rect 15335 11781 15347 11784
rect 15289 11775 15347 11781
rect 16132 11756 16160 11784
rect 18141 11781 18153 11815
rect 18187 11812 18199 11815
rect 18230 11812 18236 11824
rect 18187 11784 18236 11812
rect 18187 11781 18199 11784
rect 18141 11775 18199 11781
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 18340 11812 18368 11852
rect 18506 11840 18512 11892
rect 18564 11880 18570 11892
rect 18969 11883 19027 11889
rect 18969 11880 18981 11883
rect 18564 11852 18981 11880
rect 18564 11840 18570 11852
rect 18969 11849 18981 11852
rect 19015 11849 19027 11883
rect 18969 11843 19027 11849
rect 19058 11840 19064 11892
rect 19116 11880 19122 11892
rect 20073 11883 20131 11889
rect 20073 11880 20085 11883
rect 19116 11852 20085 11880
rect 19116 11840 19122 11852
rect 20073 11849 20085 11852
rect 20119 11849 20131 11883
rect 20073 11843 20131 11849
rect 21818 11840 21824 11892
rect 21876 11840 21882 11892
rect 21910 11840 21916 11892
rect 21968 11880 21974 11892
rect 22094 11880 22100 11892
rect 21968 11852 22100 11880
rect 21968 11840 21974 11852
rect 22094 11840 22100 11852
rect 22152 11840 22158 11892
rect 23750 11840 23756 11892
rect 23808 11880 23814 11892
rect 24489 11883 24547 11889
rect 24489 11880 24501 11883
rect 23808 11852 24501 11880
rect 23808 11840 23814 11852
rect 24489 11849 24501 11852
rect 24535 11849 24547 11883
rect 34882 11880 34888 11892
rect 24489 11843 24547 11849
rect 28966 11852 34888 11880
rect 18690 11812 18696 11824
rect 18340 11784 18696 11812
rect 18690 11772 18696 11784
rect 18748 11772 18754 11824
rect 18874 11772 18880 11824
rect 18932 11772 18938 11824
rect 24213 11815 24271 11821
rect 19592 11784 23612 11812
rect 13817 11747 13875 11753
rect 13817 11744 13829 11747
rect 13188 11716 13829 11744
rect 13817 11713 13829 11716
rect 13863 11713 13875 11747
rect 13817 11707 13875 11713
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 14090 11704 14096 11756
rect 14148 11704 14154 11756
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 15473 11747 15531 11753
rect 15473 11713 15485 11747
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 12802 11676 12808 11688
rect 12360 11648 12808 11676
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 13265 11679 13323 11685
rect 13265 11645 13277 11679
rect 13311 11676 13323 11679
rect 13906 11676 13912 11688
rect 13311 11648 13912 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 14200 11676 14228 11707
rect 14016 11648 14228 11676
rect 9723 11580 10548 11608
rect 9723 11577 9735 11580
rect 9677 11571 9735 11577
rect 11330 11568 11336 11620
rect 11388 11608 11394 11620
rect 11885 11611 11943 11617
rect 11885 11608 11897 11611
rect 11388 11580 11897 11608
rect 11388 11568 11394 11580
rect 11885 11577 11897 11580
rect 11931 11608 11943 11611
rect 12434 11608 12440 11620
rect 11931 11580 12440 11608
rect 11931 11577 11943 11580
rect 11885 11571 11943 11577
rect 12434 11568 12440 11580
rect 12492 11568 12498 11620
rect 13725 11611 13783 11617
rect 13725 11577 13737 11611
rect 13771 11608 13783 11611
rect 14016 11608 14044 11648
rect 15488 11608 15516 11707
rect 15562 11704 15568 11756
rect 15620 11704 15626 11756
rect 16114 11704 16120 11756
rect 16172 11744 16178 11756
rect 17037 11747 17095 11753
rect 17037 11744 17049 11747
rect 16172 11716 17049 11744
rect 16172 11704 16178 11716
rect 17037 11713 17049 11716
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 17402 11704 17408 11756
rect 17460 11704 17466 11756
rect 17954 11704 17960 11756
rect 18012 11704 18018 11756
rect 18598 11744 18604 11756
rect 18248 11716 18604 11744
rect 18248 11685 18276 11716
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 19242 11704 19248 11756
rect 19300 11744 19306 11756
rect 19592 11753 19620 11784
rect 19429 11747 19487 11753
rect 19429 11744 19441 11747
rect 19300 11716 19441 11744
rect 19300 11704 19306 11716
rect 19429 11713 19441 11716
rect 19475 11713 19487 11747
rect 19429 11707 19487 11713
rect 19577 11747 19635 11753
rect 19577 11713 19589 11747
rect 19623 11713 19635 11747
rect 19577 11707 19635 11713
rect 19702 11704 19708 11756
rect 19760 11704 19766 11756
rect 19794 11704 19800 11756
rect 19852 11704 19858 11756
rect 19978 11753 19984 11756
rect 19935 11747 19984 11753
rect 19935 11713 19947 11747
rect 19981 11713 19984 11747
rect 19935 11707 19984 11713
rect 19978 11704 19984 11707
rect 20036 11744 20042 11756
rect 20438 11744 20444 11756
rect 20036 11716 20444 11744
rect 20036 11704 20042 11716
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 22005 11747 22063 11753
rect 22005 11713 22017 11747
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 18414 11636 18420 11688
rect 18472 11676 18478 11688
rect 22020 11676 22048 11707
rect 22278 11704 22284 11756
rect 22336 11704 22342 11756
rect 22465 11747 22523 11753
rect 22465 11713 22477 11747
rect 22511 11744 22523 11747
rect 22646 11744 22652 11756
rect 22511 11716 22652 11744
rect 22511 11713 22523 11716
rect 22465 11707 22523 11713
rect 22646 11704 22652 11716
rect 22704 11704 22710 11756
rect 23014 11704 23020 11756
rect 23072 11704 23078 11756
rect 22557 11679 22615 11685
rect 22557 11676 22569 11679
rect 18472 11648 19937 11676
rect 22020 11648 22569 11676
rect 18472 11636 18478 11648
rect 18524 11617 18552 11648
rect 13771 11580 14044 11608
rect 14108 11580 15516 11608
rect 18509 11611 18567 11617
rect 13771 11577 13783 11580
rect 13725 11571 13783 11577
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 4893 11543 4951 11549
rect 4893 11540 4905 11543
rect 4672 11512 4905 11540
rect 4672 11500 4678 11512
rect 4893 11509 4905 11512
rect 4939 11509 4951 11543
rect 4893 11503 4951 11509
rect 7282 11500 7288 11552
rect 7340 11500 7346 11552
rect 8018 11500 8024 11552
rect 8076 11500 8082 11552
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 9456 11512 9781 11540
rect 9456 11500 9462 11512
rect 9769 11509 9781 11512
rect 9815 11509 9827 11543
rect 9769 11503 9827 11509
rect 10781 11543 10839 11549
rect 10781 11509 10793 11543
rect 10827 11540 10839 11543
rect 11606 11540 11612 11552
rect 10827 11512 11612 11540
rect 10827 11509 10839 11512
rect 10781 11503 10839 11509
rect 11606 11500 11612 11512
rect 11664 11500 11670 11552
rect 11974 11500 11980 11552
rect 12032 11500 12038 11552
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 14108 11540 14136 11580
rect 18509 11577 18521 11611
rect 18555 11577 18567 11611
rect 19518 11608 19524 11620
rect 18509 11571 18567 11577
rect 18616 11580 19524 11608
rect 12124 11512 14136 11540
rect 15289 11543 15347 11549
rect 12124 11500 12130 11512
rect 15289 11509 15301 11543
rect 15335 11540 15347 11543
rect 18616 11540 18644 11580
rect 19518 11568 19524 11580
rect 19576 11568 19582 11620
rect 19909 11608 19937 11648
rect 22557 11645 22569 11648
rect 22603 11645 22615 11679
rect 22557 11639 22615 11645
rect 22664 11608 22692 11704
rect 22741 11679 22799 11685
rect 22741 11645 22753 11679
rect 22787 11645 22799 11679
rect 22741 11639 22799 11645
rect 19909 11580 22692 11608
rect 22756 11608 22784 11639
rect 22830 11636 22836 11688
rect 22888 11636 22894 11688
rect 22922 11636 22928 11688
rect 22980 11636 22986 11688
rect 23014 11608 23020 11620
rect 22756 11580 23020 11608
rect 23014 11568 23020 11580
rect 23072 11568 23078 11620
rect 15335 11512 18644 11540
rect 15335 11509 15347 11512
rect 15289 11503 15347 11509
rect 18690 11500 18696 11552
rect 18748 11500 18754 11552
rect 18966 11500 18972 11552
rect 19024 11540 19030 11552
rect 19978 11540 19984 11552
rect 19024 11512 19984 11540
rect 19024 11500 19030 11512
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 23584 11540 23612 11784
rect 24213 11781 24225 11815
rect 24259 11812 24271 11815
rect 24394 11812 24400 11824
rect 24259 11784 24400 11812
rect 24259 11781 24271 11784
rect 24213 11775 24271 11781
rect 24394 11772 24400 11784
rect 24452 11772 24458 11824
rect 23750 11704 23756 11756
rect 23808 11704 23814 11756
rect 23842 11704 23848 11756
rect 23900 11704 23906 11756
rect 24026 11704 24032 11756
rect 24084 11744 24090 11756
rect 24305 11747 24363 11753
rect 24084 11734 24256 11744
rect 24305 11734 24317 11747
rect 24084 11716 24317 11734
rect 24084 11704 24090 11716
rect 24228 11713 24317 11716
rect 24351 11713 24363 11747
rect 24228 11707 24363 11713
rect 24228 11706 24348 11707
rect 24578 11704 24584 11756
rect 24636 11704 24642 11756
rect 24118 11636 24124 11688
rect 24176 11676 24182 11688
rect 28966 11676 28994 11852
rect 34882 11840 34888 11852
rect 34940 11840 34946 11892
rect 31294 11812 31300 11824
rect 30484 11784 31300 11812
rect 30282 11704 30288 11756
rect 30340 11704 30346 11756
rect 30484 11753 30512 11784
rect 31294 11772 31300 11784
rect 31352 11812 31358 11824
rect 31352 11784 31616 11812
rect 31352 11772 31358 11784
rect 30469 11747 30527 11753
rect 30469 11713 30481 11747
rect 30515 11713 30527 11747
rect 30469 11707 30527 11713
rect 30650 11704 30656 11756
rect 30708 11744 30714 11756
rect 31588 11753 31616 11784
rect 31754 11772 31760 11824
rect 31812 11812 31818 11824
rect 31812 11784 33272 11812
rect 31812 11772 31818 11784
rect 30929 11747 30987 11753
rect 30929 11744 30941 11747
rect 30708 11716 30941 11744
rect 30708 11704 30714 11716
rect 30929 11713 30941 11716
rect 30975 11713 30987 11747
rect 30929 11707 30987 11713
rect 31573 11747 31631 11753
rect 31573 11713 31585 11747
rect 31619 11713 31631 11747
rect 31573 11707 31631 11713
rect 31662 11704 31668 11756
rect 31720 11704 31726 11756
rect 32217 11747 32275 11753
rect 32217 11713 32229 11747
rect 32263 11713 32275 11747
rect 32217 11707 32275 11713
rect 24176 11648 28994 11676
rect 31205 11679 31263 11685
rect 24176 11636 24182 11648
rect 31205 11645 31217 11679
rect 31251 11676 31263 11679
rect 31386 11676 31392 11688
rect 31251 11648 31392 11676
rect 31251 11645 31263 11648
rect 31205 11639 31263 11645
rect 31386 11636 31392 11648
rect 31444 11636 31450 11688
rect 31680 11676 31708 11704
rect 31496 11648 31708 11676
rect 24029 11611 24087 11617
rect 24029 11577 24041 11611
rect 24075 11608 24087 11611
rect 24305 11611 24363 11617
rect 24305 11608 24317 11611
rect 24075 11580 24317 11608
rect 24075 11577 24087 11580
rect 24029 11571 24087 11577
rect 24305 11577 24317 11580
rect 24351 11577 24363 11611
rect 24305 11571 24363 11577
rect 30374 11568 30380 11620
rect 30432 11608 30438 11620
rect 31496 11608 31524 11648
rect 31754 11636 31760 11688
rect 31812 11636 31818 11688
rect 32122 11636 32128 11688
rect 32180 11676 32186 11688
rect 32232 11676 32260 11707
rect 33134 11704 33140 11756
rect 33192 11704 33198 11756
rect 33244 11753 33272 11784
rect 33229 11747 33287 11753
rect 33229 11713 33241 11747
rect 33275 11744 33287 11747
rect 33689 11747 33747 11753
rect 33689 11744 33701 11747
rect 33275 11716 33701 11744
rect 33275 11713 33287 11716
rect 33229 11707 33287 11713
rect 33689 11713 33701 11716
rect 33735 11713 33747 11747
rect 33689 11707 33747 11713
rect 34606 11704 34612 11756
rect 34664 11744 34670 11756
rect 34977 11747 35035 11753
rect 34977 11744 34989 11747
rect 34664 11716 34989 11744
rect 34664 11704 34670 11716
rect 34977 11713 34989 11716
rect 35023 11713 35035 11747
rect 34977 11707 35035 11713
rect 35244 11747 35302 11753
rect 35244 11713 35256 11747
rect 35290 11744 35302 11747
rect 36262 11744 36268 11756
rect 35290 11716 36268 11744
rect 35290 11713 35302 11716
rect 35244 11707 35302 11713
rect 36262 11704 36268 11716
rect 36320 11704 36326 11756
rect 32180 11648 33456 11676
rect 32180 11636 32186 11648
rect 30432 11580 31524 11608
rect 30432 11568 30438 11580
rect 31570 11568 31576 11620
rect 31628 11608 31634 11620
rect 31665 11611 31723 11617
rect 31665 11608 31677 11611
rect 31628 11580 31677 11608
rect 31628 11568 31634 11580
rect 31665 11577 31677 11580
rect 31711 11577 31723 11611
rect 31665 11571 31723 11577
rect 31938 11568 31944 11620
rect 31996 11608 32002 11620
rect 33321 11611 33379 11617
rect 33321 11608 33333 11611
rect 31996 11580 33333 11608
rect 31996 11568 32002 11580
rect 33321 11577 33333 11580
rect 33367 11577 33379 11611
rect 33428 11608 33456 11648
rect 33502 11636 33508 11688
rect 33560 11636 33566 11688
rect 33428 11580 34008 11608
rect 33321 11571 33379 11577
rect 29914 11540 29920 11552
rect 23584 11512 29920 11540
rect 29914 11500 29920 11512
rect 29972 11500 29978 11552
rect 30285 11543 30343 11549
rect 30285 11509 30297 11543
rect 30331 11540 30343 11543
rect 31018 11540 31024 11552
rect 30331 11512 31024 11540
rect 30331 11509 30343 11512
rect 30285 11503 30343 11509
rect 31018 11500 31024 11512
rect 31076 11500 31082 11552
rect 32214 11500 32220 11552
rect 32272 11540 32278 11552
rect 32309 11543 32367 11549
rect 32309 11540 32321 11543
rect 32272 11512 32321 11540
rect 32272 11500 32278 11512
rect 32309 11509 32321 11512
rect 32355 11509 32367 11543
rect 32309 11503 32367 11509
rect 33594 11500 33600 11552
rect 33652 11540 33658 11552
rect 33873 11543 33931 11549
rect 33873 11540 33885 11543
rect 33652 11512 33885 11540
rect 33652 11500 33658 11512
rect 33873 11509 33885 11512
rect 33919 11509 33931 11543
rect 33980 11540 34008 11580
rect 36357 11543 36415 11549
rect 36357 11540 36369 11543
rect 33980 11512 36369 11540
rect 33873 11503 33931 11509
rect 36357 11509 36369 11512
rect 36403 11509 36415 11543
rect 36357 11503 36415 11509
rect 1104 11450 36800 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 36800 11450
rect 1104 11376 36800 11398
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11336 7251 11339
rect 7282 11336 7288 11348
rect 7239 11308 7288 11336
rect 7239 11305 7251 11308
rect 7193 11299 7251 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 12066 11336 12072 11348
rect 7607 11308 12072 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 12253 11339 12311 11345
rect 12253 11305 12265 11339
rect 12299 11336 12311 11339
rect 12526 11336 12532 11348
rect 12299 11308 12532 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 16761 11339 16819 11345
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 16850 11336 16856 11348
rect 16807 11308 16856 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 19797 11339 19855 11345
rect 19797 11336 19809 11339
rect 18012 11308 19809 11336
rect 18012 11296 18018 11308
rect 19797 11305 19809 11308
rect 19843 11305 19855 11339
rect 19797 11299 19855 11305
rect 22278 11296 22284 11348
rect 22336 11296 22342 11348
rect 22465 11339 22523 11345
rect 22465 11305 22477 11339
rect 22511 11336 22523 11339
rect 22738 11336 22744 11348
rect 22511 11308 22744 11336
rect 22511 11305 22523 11308
rect 22465 11299 22523 11305
rect 22738 11296 22744 11308
rect 22796 11296 22802 11348
rect 23477 11339 23535 11345
rect 23477 11305 23489 11339
rect 23523 11336 23535 11339
rect 23750 11336 23756 11348
rect 23523 11308 23756 11336
rect 23523 11305 23535 11308
rect 23477 11299 23535 11305
rect 23750 11296 23756 11308
rect 23808 11296 23814 11348
rect 24118 11296 24124 11348
rect 24176 11336 24182 11348
rect 29270 11336 29276 11348
rect 24176 11308 29276 11336
rect 24176 11296 24182 11308
rect 29270 11296 29276 11308
rect 29328 11296 29334 11348
rect 31294 11296 31300 11348
rect 31352 11296 31358 11348
rect 31386 11296 31392 11348
rect 31444 11336 31450 11348
rect 33134 11336 33140 11348
rect 31444 11308 33140 11336
rect 31444 11296 31450 11308
rect 33134 11296 33140 11308
rect 33192 11296 33198 11348
rect 36262 11296 36268 11348
rect 36320 11296 36326 11348
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 9401 11271 9459 11277
rect 9401 11268 9413 11271
rect 9088 11240 9413 11268
rect 9088 11228 9094 11240
rect 9401 11237 9413 11240
rect 9447 11237 9459 11271
rect 11790 11268 11796 11280
rect 9401 11231 9459 11237
rect 9508 11240 11796 11268
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 9508 11200 9536 11240
rect 11790 11228 11796 11240
rect 11848 11228 11854 11280
rect 14277 11271 14335 11277
rect 14277 11237 14289 11271
rect 14323 11268 14335 11271
rect 19242 11268 19248 11280
rect 14323 11240 19248 11268
rect 14323 11237 14335 11240
rect 14277 11231 14335 11237
rect 19242 11228 19248 11240
rect 19300 11228 19306 11280
rect 19978 11268 19984 11280
rect 19444 11240 19984 11268
rect 11330 11200 11336 11212
rect 7423 11172 9536 11200
rect 9600 11172 11336 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7190 11132 7196 11144
rect 7147 11104 7196 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 5718 10956 5724 11008
rect 5776 10996 5782 11008
rect 7392 10996 7420 11163
rect 7466 11092 7472 11144
rect 7524 11092 7530 11144
rect 9398 11092 9404 11144
rect 9456 11092 9462 11144
rect 9600 11132 9628 11172
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 11606 11160 11612 11212
rect 11664 11160 11670 11212
rect 16850 11160 16856 11212
rect 16908 11200 16914 11212
rect 17405 11203 17463 11209
rect 17405 11200 17417 11203
rect 16908 11172 17417 11200
rect 16908 11160 16914 11172
rect 17405 11169 17417 11172
rect 17451 11200 17463 11203
rect 17770 11200 17776 11212
rect 17451 11172 17776 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 17770 11160 17776 11172
rect 17828 11160 17834 11212
rect 18598 11160 18604 11212
rect 18656 11200 18662 11212
rect 19444 11200 19472 11240
rect 19978 11228 19984 11240
rect 20036 11228 20042 11280
rect 25038 11228 25044 11280
rect 25096 11268 25102 11280
rect 25682 11268 25688 11280
rect 25096 11240 25688 11268
rect 25096 11228 25102 11240
rect 25682 11228 25688 11240
rect 25740 11268 25746 11280
rect 34790 11268 34796 11280
rect 25740 11240 34796 11268
rect 25740 11228 25746 11240
rect 34790 11228 34796 11240
rect 34848 11228 34854 11280
rect 18656 11172 19472 11200
rect 18656 11160 18662 11172
rect 9508 11104 9628 11132
rect 9677 11135 9735 11141
rect 7834 11024 7840 11076
rect 7892 11064 7898 11076
rect 9508 11064 9536 11104
rect 9677 11101 9689 11135
rect 9723 11132 9735 11135
rect 10318 11132 10324 11144
rect 9723 11104 10324 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 11790 11092 11796 11144
rect 11848 11092 11854 11144
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 14553 11135 14611 11141
rect 14553 11132 14565 11135
rect 12860 11104 14565 11132
rect 12860 11092 12866 11104
rect 14553 11101 14565 11104
rect 14599 11101 14611 11135
rect 14553 11095 14611 11101
rect 14642 11092 14648 11144
rect 14700 11092 14706 11144
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 7892 11036 9536 11064
rect 9585 11067 9643 11073
rect 7892 11024 7898 11036
rect 9585 11033 9597 11067
rect 9631 11064 9643 11067
rect 10410 11064 10416 11076
rect 9631 11036 10416 11064
rect 9631 11033 9643 11036
rect 9585 11027 9643 11033
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 14090 11024 14096 11076
rect 14148 11064 14154 11076
rect 14752 11064 14780 11095
rect 14918 11092 14924 11144
rect 14976 11092 14982 11144
rect 15194 11092 15200 11144
rect 15252 11092 15258 11144
rect 18708 11141 18736 11172
rect 18509 11135 18567 11141
rect 18509 11132 18521 11135
rect 17512 11104 18521 11132
rect 14148 11036 14780 11064
rect 14148 11024 14154 11036
rect 17512 11008 17540 11104
rect 18509 11101 18521 11104
rect 18555 11101 18567 11135
rect 18509 11095 18567 11101
rect 18693 11135 18751 11141
rect 18693 11101 18705 11135
rect 18739 11101 18751 11135
rect 18693 11095 18751 11101
rect 18782 11092 18788 11144
rect 18840 11092 18846 11144
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11132 18935 11135
rect 18966 11132 18972 11144
rect 18923 11104 18972 11132
rect 18923 11101 18935 11104
rect 18877 11095 18935 11101
rect 18966 11092 18972 11104
rect 19024 11132 19030 11144
rect 19444 11141 19472 11172
rect 19521 11203 19579 11209
rect 19521 11169 19533 11203
rect 19567 11200 19579 11203
rect 21085 11203 21143 11209
rect 19567 11172 20760 11200
rect 19567 11169 19579 11172
rect 19521 11163 19579 11169
rect 19429 11135 19487 11141
rect 19024 11104 19380 11132
rect 19024 11092 19030 11104
rect 19242 11024 19248 11076
rect 19300 11024 19306 11076
rect 5776 10968 7420 10996
rect 5776 10956 5782 10968
rect 15010 10956 15016 11008
rect 15068 10956 15074 11008
rect 17126 10956 17132 11008
rect 17184 10956 17190 11008
rect 17221 10999 17279 11005
rect 17221 10965 17233 10999
rect 17267 10996 17279 10999
rect 17494 10996 17500 11008
rect 17267 10968 17500 10996
rect 17267 10965 17279 10968
rect 17221 10959 17279 10965
rect 17494 10956 17500 10968
rect 17552 10956 17558 11008
rect 19058 10956 19064 11008
rect 19116 10956 19122 11008
rect 19352 10996 19380 11104
rect 19429 11101 19441 11135
rect 19475 11101 19487 11135
rect 19889 11135 19947 11141
rect 19429 11095 19487 11101
rect 19618 11113 19676 11119
rect 19618 11079 19630 11113
rect 19664 11079 19676 11113
rect 19889 11101 19901 11135
rect 19935 11101 19947 11135
rect 19889 11095 19947 11101
rect 19518 11024 19524 11076
rect 19576 11024 19582 11076
rect 19618 11073 19676 11079
rect 19628 10996 19656 11073
rect 19904 11064 19932 11095
rect 19978 11092 19984 11144
rect 20036 11092 20042 11144
rect 20254 11092 20260 11144
rect 20312 11092 20318 11144
rect 20438 11092 20444 11144
rect 20496 11092 20502 11144
rect 20732 11141 20760 11172
rect 21085 11169 21097 11203
rect 21131 11200 21143 11203
rect 22186 11200 22192 11212
rect 21131 11172 22192 11200
rect 21131 11169 21143 11172
rect 21085 11163 21143 11169
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 23014 11160 23020 11212
rect 23072 11200 23078 11212
rect 24578 11200 24584 11212
rect 23072 11172 24584 11200
rect 23072 11160 23078 11172
rect 24578 11160 24584 11172
rect 24636 11160 24642 11212
rect 28813 11203 28871 11209
rect 28276 11172 28672 11200
rect 20717 11135 20775 11141
rect 20717 11101 20729 11135
rect 20763 11101 20775 11135
rect 20717 11095 20775 11101
rect 20806 11092 20812 11144
rect 20864 11132 20870 11144
rect 20901 11135 20959 11141
rect 20901 11132 20913 11135
rect 20864 11104 20913 11132
rect 20864 11092 20870 11104
rect 20901 11101 20913 11104
rect 20947 11101 20959 11135
rect 22922 11132 22928 11144
rect 20901 11095 20959 11101
rect 22112 11104 22928 11132
rect 22112 11076 22140 11104
rect 22922 11092 22928 11104
rect 22980 11132 22986 11144
rect 23109 11135 23167 11141
rect 23109 11132 23121 11135
rect 22980 11104 23121 11132
rect 22980 11092 22986 11104
rect 23109 11101 23121 11104
rect 23155 11101 23167 11135
rect 23109 11095 23167 11101
rect 23293 11135 23351 11141
rect 23293 11101 23305 11135
rect 23339 11101 23351 11135
rect 23293 11095 23351 11101
rect 26329 11135 26387 11141
rect 26329 11101 26341 11135
rect 26375 11132 26387 11135
rect 26878 11132 26884 11144
rect 26375 11104 26884 11132
rect 26375 11101 26387 11104
rect 26329 11095 26387 11101
rect 21174 11064 21180 11076
rect 19904 11036 20116 11064
rect 19352 10968 19656 10996
rect 20088 10996 20116 11036
rect 20272 11036 21180 11064
rect 20272 10996 20300 11036
rect 21174 11024 21180 11036
rect 21232 11024 21238 11076
rect 22094 11024 22100 11076
rect 22152 11024 22158 11076
rect 22830 11064 22836 11076
rect 22388 11036 22836 11064
rect 22388 11008 22416 11036
rect 22830 11024 22836 11036
rect 22888 11064 22894 11076
rect 23308 11064 23336 11095
rect 26878 11092 26884 11104
rect 26936 11092 26942 11144
rect 27982 11092 27988 11144
rect 28040 11132 28046 11144
rect 28077 11135 28135 11141
rect 28077 11132 28089 11135
rect 28040 11104 28089 11132
rect 28040 11092 28046 11104
rect 28077 11101 28089 11104
rect 28123 11101 28135 11135
rect 28077 11095 28135 11101
rect 22888 11036 23336 11064
rect 22888 11024 22894 11036
rect 25406 11024 25412 11076
rect 25464 11064 25470 11076
rect 26513 11067 26571 11073
rect 26513 11064 26525 11067
rect 25464 11036 26525 11064
rect 25464 11024 25470 11036
rect 26513 11033 26525 11036
rect 26559 11033 26571 11067
rect 28092 11064 28120 11095
rect 28166 11092 28172 11144
rect 28224 11132 28230 11144
rect 28276 11141 28304 11172
rect 28644 11141 28672 11172
rect 28813 11169 28825 11203
rect 28859 11200 28871 11203
rect 31478 11200 31484 11212
rect 28859 11172 31484 11200
rect 28859 11169 28871 11172
rect 28813 11163 28871 11169
rect 31478 11160 31484 11172
rect 31536 11200 31542 11212
rect 31662 11200 31668 11212
rect 31536 11172 31668 11200
rect 31536 11160 31542 11172
rect 31662 11160 31668 11172
rect 31720 11200 31726 11212
rect 31720 11160 31754 11200
rect 28261 11135 28319 11141
rect 28261 11132 28273 11135
rect 28224 11104 28273 11132
rect 28224 11092 28230 11104
rect 28261 11101 28273 11104
rect 28307 11101 28319 11135
rect 28261 11095 28319 11101
rect 28537 11135 28595 11141
rect 28537 11101 28549 11135
rect 28583 11101 28595 11135
rect 28537 11095 28595 11101
rect 28629 11135 28687 11141
rect 28629 11101 28641 11135
rect 28675 11132 28687 11135
rect 28718 11132 28724 11144
rect 28675 11104 28724 11132
rect 28675 11101 28687 11104
rect 28629 11095 28687 11101
rect 28552 11064 28580 11095
rect 28718 11092 28724 11104
rect 28776 11092 28782 11144
rect 31021 11135 31079 11141
rect 31021 11101 31033 11135
rect 31067 11101 31079 11135
rect 31021 11095 31079 11101
rect 31113 11135 31171 11141
rect 31113 11101 31125 11135
rect 31159 11132 31171 11135
rect 31386 11132 31392 11144
rect 31159 11104 31392 11132
rect 31159 11101 31171 11104
rect 31113 11095 31171 11101
rect 28092 11036 28580 11064
rect 31036 11064 31064 11095
rect 31386 11092 31392 11104
rect 31444 11092 31450 11144
rect 31726 11132 31754 11160
rect 31849 11135 31907 11141
rect 31849 11132 31861 11135
rect 31726 11104 31861 11132
rect 31849 11101 31861 11104
rect 31895 11101 31907 11135
rect 31849 11095 31907 11101
rect 31938 11092 31944 11144
rect 31996 11092 32002 11144
rect 32030 11092 32036 11144
rect 32088 11092 32094 11144
rect 32214 11092 32220 11144
rect 32272 11092 32278 11144
rect 35253 11135 35311 11141
rect 35253 11101 35265 11135
rect 35299 11132 35311 11135
rect 35342 11132 35348 11144
rect 35299 11104 35348 11132
rect 35299 11101 35311 11104
rect 35253 11095 35311 11101
rect 35342 11092 35348 11104
rect 35400 11092 35406 11144
rect 36446 11092 36452 11144
rect 36504 11092 36510 11144
rect 31294 11064 31300 11076
rect 31036 11036 31300 11064
rect 26513 11027 26571 11033
rect 31294 11024 31300 11036
rect 31352 11064 31358 11076
rect 32122 11064 32128 11076
rect 31352 11036 32128 11064
rect 31352 11024 31358 11036
rect 32122 11024 32128 11036
rect 32180 11024 32186 11076
rect 20088 10968 20300 10996
rect 22281 10999 22339 11005
rect 22281 10965 22293 10999
rect 22327 10996 22339 10999
rect 22370 10996 22376 11008
rect 22327 10968 22376 10996
rect 22327 10965 22339 10968
rect 22281 10959 22339 10965
rect 22370 10956 22376 10968
rect 22428 10956 22434 11008
rect 24302 10956 24308 11008
rect 24360 10996 24366 11008
rect 26326 10996 26332 11008
rect 24360 10968 26332 10996
rect 24360 10956 24366 10968
rect 26326 10956 26332 10968
rect 26384 10956 26390 11008
rect 28445 10999 28503 11005
rect 28445 10965 28457 10999
rect 28491 10996 28503 10999
rect 28534 10996 28540 11008
rect 28491 10968 28540 10996
rect 28491 10965 28503 10968
rect 28445 10959 28503 10965
rect 28534 10956 28540 10968
rect 28592 10956 28598 11008
rect 28626 10956 28632 11008
rect 28684 10996 28690 11008
rect 28813 10999 28871 11005
rect 28813 10996 28825 10999
rect 28684 10968 28825 10996
rect 28684 10956 28690 10968
rect 28813 10965 28825 10968
rect 28859 10965 28871 10999
rect 28813 10959 28871 10965
rect 28994 10956 29000 11008
rect 29052 10996 29058 11008
rect 34514 10996 34520 11008
rect 29052 10968 34520 10996
rect 29052 10956 29058 10968
rect 34514 10956 34520 10968
rect 34572 10956 34578 11008
rect 34698 10956 34704 11008
rect 34756 10996 34762 11008
rect 35069 10999 35127 11005
rect 35069 10996 35081 10999
rect 34756 10968 35081 10996
rect 34756 10956 34762 10968
rect 35069 10965 35081 10968
rect 35115 10965 35127 10999
rect 35069 10959 35127 10965
rect 1104 10906 36800 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 36800 10906
rect 1104 10832 36800 10854
rect 7466 10752 7472 10804
rect 7524 10752 7530 10804
rect 9214 10752 9220 10804
rect 9272 10792 9278 10804
rect 10229 10795 10287 10801
rect 10229 10792 10241 10795
rect 9272 10764 10241 10792
rect 9272 10752 9278 10764
rect 10229 10761 10241 10764
rect 10275 10761 10287 10795
rect 10229 10755 10287 10761
rect 14090 10752 14096 10804
rect 14148 10752 14154 10804
rect 14461 10795 14519 10801
rect 14461 10761 14473 10795
rect 14507 10792 14519 10795
rect 14642 10792 14648 10804
rect 14507 10764 14648 10792
rect 14507 10761 14519 10764
rect 14461 10755 14519 10761
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 14829 10795 14887 10801
rect 14829 10761 14841 10795
rect 14875 10792 14887 10795
rect 15010 10792 15016 10804
rect 14875 10764 15016 10792
rect 14875 10761 14887 10764
rect 14829 10755 14887 10761
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 16301 10795 16359 10801
rect 16301 10761 16313 10795
rect 16347 10761 16359 10795
rect 16301 10755 16359 10761
rect 5997 10727 6055 10733
rect 5997 10724 6009 10727
rect 5184 10696 6009 10724
rect 4982 10616 4988 10668
rect 5040 10616 5046 10668
rect 5074 10616 5080 10668
rect 5132 10616 5138 10668
rect 5184 10665 5212 10696
rect 5997 10693 6009 10696
rect 6043 10693 6055 10727
rect 8018 10724 8024 10736
rect 5997 10687 6055 10693
rect 7208 10696 8024 10724
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 5534 10616 5540 10668
rect 5592 10616 5598 10668
rect 5718 10616 5724 10668
rect 5776 10616 5782 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10588 5411 10591
rect 5828 10588 5856 10619
rect 5902 10616 5908 10668
rect 5960 10616 5966 10668
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7208 10665 7236 10696
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 13630 10724 13636 10736
rect 12406 10696 13636 10724
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 6972 10628 7205 10656
rect 6972 10616 6978 10628
rect 7193 10625 7205 10628
rect 7239 10625 7251 10659
rect 7193 10619 7251 10625
rect 7282 10616 7288 10668
rect 7340 10616 7346 10668
rect 10318 10616 10324 10668
rect 10376 10616 10382 10668
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 12406 10656 12434 10696
rect 13630 10684 13636 10696
rect 13688 10684 13694 10736
rect 16316 10724 16344 10755
rect 16390 10752 16396 10804
rect 16448 10792 16454 10804
rect 16448 10764 17080 10792
rect 16448 10752 16454 10764
rect 16914 10727 16972 10733
rect 16914 10724 16926 10727
rect 16316 10696 16926 10724
rect 16914 10693 16926 10696
rect 16960 10693 16972 10727
rect 17052 10724 17080 10764
rect 17126 10752 17132 10804
rect 17184 10792 17190 10804
rect 18049 10795 18107 10801
rect 18049 10792 18061 10795
rect 17184 10764 18061 10792
rect 17184 10752 17190 10764
rect 18049 10761 18061 10764
rect 18095 10761 18107 10795
rect 18049 10755 18107 10761
rect 24765 10795 24823 10801
rect 24765 10761 24777 10795
rect 24811 10792 24823 10795
rect 24811 10764 27844 10792
rect 24811 10761 24823 10764
rect 24765 10755 24823 10761
rect 21266 10724 21272 10736
rect 17052 10696 21272 10724
rect 16914 10687 16972 10693
rect 21266 10684 21272 10696
rect 21324 10684 21330 10736
rect 24857 10727 24915 10733
rect 24857 10693 24869 10727
rect 24903 10724 24915 10727
rect 25654 10727 25712 10733
rect 25654 10724 25666 10727
rect 24903 10696 25666 10724
rect 24903 10693 24915 10696
rect 24857 10687 24915 10693
rect 25654 10693 25666 10696
rect 25700 10693 25712 10727
rect 27816 10724 27844 10764
rect 27890 10752 27896 10804
rect 27948 10792 27954 10804
rect 28629 10795 28687 10801
rect 28629 10792 28641 10795
rect 27948 10764 28641 10792
rect 27948 10752 27954 10764
rect 28629 10761 28641 10764
rect 28675 10761 28687 10795
rect 28629 10755 28687 10761
rect 28810 10752 28816 10804
rect 28868 10792 28874 10804
rect 28868 10764 29316 10792
rect 28868 10752 28874 10764
rect 28994 10724 29000 10736
rect 27816 10696 29000 10724
rect 25654 10687 25712 10693
rect 28994 10684 29000 10696
rect 29052 10684 29058 10736
rect 29288 10733 29316 10764
rect 31478 10752 31484 10804
rect 31536 10752 31542 10804
rect 34238 10792 34244 10804
rect 31726 10764 34244 10792
rect 29273 10727 29331 10733
rect 29273 10693 29285 10727
rect 29319 10693 29331 10727
rect 29273 10687 29331 10693
rect 29362 10684 29368 10736
rect 29420 10724 29426 10736
rect 31726 10724 31754 10764
rect 34238 10752 34244 10764
rect 34296 10752 34302 10804
rect 35894 10792 35900 10804
rect 34624 10764 35900 10792
rect 33226 10724 33232 10736
rect 29420 10696 31754 10724
rect 32140 10696 33232 10724
rect 29420 10684 29426 10696
rect 10689 10619 10747 10625
rect 10796 10628 12434 10656
rect 5399 10560 5856 10588
rect 7469 10591 7527 10597
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 7558 10588 7564 10600
rect 7515 10560 7564 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 7558 10548 7564 10560
rect 7616 10588 7622 10600
rect 7926 10588 7932 10600
rect 7616 10560 7932 10588
rect 7616 10548 7622 10560
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 10704 10588 10732 10619
rect 8128 10560 10732 10588
rect 5813 10523 5871 10529
rect 5813 10489 5825 10523
rect 5859 10520 5871 10523
rect 8128 10520 8156 10560
rect 5859 10492 8156 10520
rect 5859 10489 5871 10492
rect 5813 10483 5871 10489
rect 6362 10412 6368 10464
rect 6420 10452 6426 10464
rect 10796 10452 10824 10628
rect 13538 10616 13544 10668
rect 13596 10656 13602 10668
rect 13725 10659 13783 10665
rect 13725 10656 13737 10659
rect 13596 10628 13737 10656
rect 13596 10616 13602 10628
rect 13725 10625 13737 10628
rect 13771 10625 13783 10659
rect 13725 10619 13783 10625
rect 14642 10616 14648 10668
rect 14700 10656 14706 10668
rect 16485 10659 16543 10665
rect 14700 10628 15056 10656
rect 14700 10616 14706 10628
rect 10962 10548 10968 10600
rect 11020 10548 11026 10600
rect 11974 10548 11980 10600
rect 12032 10588 12038 10600
rect 13262 10588 13268 10600
rect 12032 10560 13268 10588
rect 12032 10548 12038 10560
rect 13262 10548 13268 10560
rect 13320 10588 13326 10600
rect 13817 10591 13875 10597
rect 13817 10588 13829 10591
rect 13320 10560 13829 10588
rect 13320 10548 13326 10560
rect 13817 10557 13829 10560
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 14918 10548 14924 10600
rect 14976 10548 14982 10600
rect 15028 10597 15056 10628
rect 16485 10625 16497 10659
rect 16531 10656 16543 10659
rect 16758 10656 16764 10668
rect 16531 10628 16764 10656
rect 16531 10625 16543 10628
rect 16485 10619 16543 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 20622 10616 20628 10668
rect 20680 10656 20686 10668
rect 21545 10659 21603 10665
rect 21545 10656 21557 10659
rect 20680 10628 21557 10656
rect 20680 10616 20686 10628
rect 21545 10625 21557 10628
rect 21591 10625 21603 10659
rect 21545 10619 21603 10625
rect 21910 10616 21916 10668
rect 21968 10656 21974 10668
rect 22278 10656 22284 10668
rect 21968 10628 22284 10656
rect 21968 10616 21974 10628
rect 22278 10616 22284 10628
rect 22336 10616 22342 10668
rect 23934 10616 23940 10668
rect 23992 10656 23998 10668
rect 24210 10656 24216 10668
rect 23992 10628 24216 10656
rect 23992 10616 23998 10628
rect 24210 10616 24216 10628
rect 24268 10656 24274 10668
rect 24397 10659 24455 10665
rect 24397 10656 24409 10659
rect 24268 10628 24409 10656
rect 24268 10616 24274 10628
rect 24397 10625 24409 10628
rect 24443 10625 24455 10659
rect 24397 10619 24455 10625
rect 25038 10616 25044 10668
rect 25096 10616 25102 10668
rect 25225 10659 25283 10665
rect 25225 10625 25237 10659
rect 25271 10656 25283 10659
rect 27617 10659 27675 10665
rect 25271 10628 27568 10656
rect 25271 10625 25283 10628
rect 25225 10619 25283 10625
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 16669 10591 16727 10597
rect 16669 10557 16681 10591
rect 16715 10557 16727 10591
rect 16669 10551 16727 10557
rect 12342 10480 12348 10532
rect 12400 10520 12406 10532
rect 16684 10520 16712 10551
rect 21358 10548 21364 10600
rect 21416 10548 21422 10600
rect 24489 10591 24547 10597
rect 24489 10557 24501 10591
rect 24535 10588 24547 10591
rect 25130 10588 25136 10600
rect 24535 10560 25136 10588
rect 24535 10557 24547 10560
rect 24489 10551 24547 10557
rect 25130 10548 25136 10560
rect 25188 10588 25194 10600
rect 25317 10591 25375 10597
rect 25317 10588 25329 10591
rect 25188 10560 25329 10588
rect 25188 10548 25194 10560
rect 25317 10557 25329 10560
rect 25363 10557 25375 10591
rect 25317 10551 25375 10557
rect 25406 10548 25412 10600
rect 25464 10548 25470 10600
rect 27540 10588 27568 10628
rect 27617 10625 27629 10659
rect 27663 10656 27675 10659
rect 27893 10659 27951 10665
rect 27663 10628 27844 10656
rect 27663 10625 27675 10628
rect 27617 10619 27675 10625
rect 27706 10588 27712 10600
rect 27540 10560 27712 10588
rect 27706 10548 27712 10560
rect 27764 10548 27770 10600
rect 27816 10588 27844 10628
rect 27893 10625 27905 10659
rect 27939 10656 27951 10659
rect 28166 10656 28172 10668
rect 27939 10628 28172 10656
rect 27939 10625 27951 10628
rect 27893 10619 27951 10625
rect 28166 10616 28172 10628
rect 28224 10616 28230 10668
rect 28261 10659 28319 10665
rect 28261 10625 28273 10659
rect 28307 10625 28319 10659
rect 28261 10619 28319 10625
rect 28445 10659 28503 10665
rect 28445 10625 28457 10659
rect 28491 10656 28503 10659
rect 28626 10656 28632 10668
rect 28491 10628 28632 10656
rect 28491 10625 28503 10628
rect 28445 10619 28503 10625
rect 27982 10588 27988 10600
rect 27816 10560 27988 10588
rect 27982 10548 27988 10560
rect 28040 10548 28046 10600
rect 12400 10492 16712 10520
rect 12400 10480 12406 10492
rect 6420 10424 10824 10452
rect 6420 10412 6426 10424
rect 13446 10412 13452 10464
rect 13504 10452 13510 10464
rect 13725 10455 13783 10461
rect 13725 10452 13737 10455
rect 13504 10424 13737 10452
rect 13504 10412 13510 10424
rect 13725 10421 13737 10424
rect 13771 10452 13783 10455
rect 13814 10452 13820 10464
rect 13771 10424 13820 10452
rect 13771 10421 13783 10424
rect 13725 10415 13783 10421
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 16684 10452 16712 10492
rect 19242 10480 19248 10532
rect 19300 10520 19306 10532
rect 21266 10520 21272 10532
rect 19300 10492 21272 10520
rect 19300 10480 19306 10492
rect 21266 10480 21272 10492
rect 21324 10480 21330 10532
rect 17770 10452 17776 10464
rect 16684 10424 17776 10452
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 21376 10461 21404 10548
rect 24762 10480 24768 10532
rect 24820 10520 24826 10532
rect 25038 10520 25044 10532
rect 24820 10492 25044 10520
rect 24820 10480 24826 10492
rect 25038 10480 25044 10492
rect 25096 10520 25102 10532
rect 25424 10520 25452 10548
rect 25096 10492 25452 10520
rect 25096 10480 25102 10492
rect 27614 10480 27620 10532
rect 27672 10520 27678 10532
rect 27893 10523 27951 10529
rect 27893 10520 27905 10523
rect 27672 10492 27905 10520
rect 27672 10480 27678 10492
rect 27893 10489 27905 10492
rect 27939 10520 27951 10523
rect 28276 10520 28304 10619
rect 28626 10616 28632 10628
rect 28684 10616 28690 10668
rect 28810 10616 28816 10668
rect 28868 10616 28874 10668
rect 28905 10659 28963 10665
rect 28905 10625 28917 10659
rect 28951 10625 28963 10659
rect 28905 10619 28963 10625
rect 29181 10659 29239 10665
rect 29181 10625 29193 10659
rect 29227 10656 29239 10659
rect 29638 10656 29644 10668
rect 29227 10628 29644 10656
rect 29227 10625 29239 10628
rect 29181 10619 29239 10625
rect 28534 10548 28540 10600
rect 28592 10588 28598 10600
rect 28920 10588 28948 10619
rect 29638 10616 29644 10628
rect 29696 10616 29702 10668
rect 31294 10616 31300 10668
rect 31352 10616 31358 10668
rect 31386 10616 31392 10668
rect 31444 10616 31450 10668
rect 31662 10616 31668 10668
rect 31720 10656 31726 10668
rect 32140 10656 32168 10696
rect 33226 10684 33232 10696
rect 33284 10684 33290 10736
rect 33962 10724 33968 10736
rect 33428 10696 33968 10724
rect 33428 10668 33456 10696
rect 33962 10684 33968 10696
rect 34020 10684 34026 10736
rect 34517 10727 34575 10733
rect 34517 10724 34529 10727
rect 34164 10696 34529 10724
rect 34164 10668 34192 10696
rect 34517 10693 34529 10696
rect 34563 10693 34575 10727
rect 34517 10687 34575 10693
rect 31720 10628 32168 10656
rect 31720 10616 31726 10628
rect 32214 10616 32220 10668
rect 32272 10616 32278 10668
rect 32677 10659 32735 10665
rect 32677 10625 32689 10659
rect 32723 10625 32735 10659
rect 32677 10619 32735 10625
rect 29457 10591 29515 10597
rect 29457 10588 29469 10591
rect 28592 10560 29469 10588
rect 28592 10548 28598 10560
rect 29457 10557 29469 10560
rect 29503 10557 29515 10591
rect 29457 10551 29515 10557
rect 31018 10548 31024 10600
rect 31076 10588 31082 10600
rect 31757 10591 31815 10597
rect 31757 10588 31769 10591
rect 31076 10560 31769 10588
rect 31076 10548 31082 10560
rect 31757 10557 31769 10560
rect 31803 10557 31815 10591
rect 31757 10551 31815 10557
rect 31938 10548 31944 10600
rect 31996 10548 32002 10600
rect 32030 10548 32036 10600
rect 32088 10588 32094 10600
rect 32692 10588 32720 10619
rect 32858 10616 32864 10668
rect 32916 10656 32922 10668
rect 33045 10659 33103 10665
rect 33045 10656 33057 10659
rect 32916 10628 33057 10656
rect 32916 10616 32922 10628
rect 33045 10625 33057 10628
rect 33091 10656 33103 10659
rect 33410 10656 33416 10668
rect 33091 10628 33416 10656
rect 33091 10625 33103 10628
rect 33045 10619 33103 10625
rect 33410 10616 33416 10628
rect 33468 10616 33474 10668
rect 33594 10616 33600 10668
rect 33652 10616 33658 10668
rect 33778 10616 33784 10668
rect 33836 10616 33842 10668
rect 34057 10659 34115 10665
rect 34057 10625 34069 10659
rect 34103 10656 34115 10659
rect 34146 10656 34152 10668
rect 34103 10628 34152 10656
rect 34103 10625 34115 10628
rect 34057 10619 34115 10625
rect 34146 10616 34152 10628
rect 34204 10616 34210 10668
rect 34241 10659 34299 10665
rect 34241 10625 34253 10659
rect 34287 10656 34299 10659
rect 34624 10656 34652 10764
rect 35894 10752 35900 10764
rect 35952 10792 35958 10804
rect 36354 10792 36360 10804
rect 35952 10764 36360 10792
rect 35952 10752 35958 10764
rect 36354 10752 36360 10764
rect 36412 10752 36418 10804
rect 34287 10628 34652 10656
rect 34287 10625 34299 10628
rect 34241 10619 34299 10625
rect 34790 10616 34796 10668
rect 34848 10656 34854 10668
rect 35233 10659 35291 10665
rect 35233 10656 35245 10659
rect 34848 10628 35245 10656
rect 34848 10616 34854 10628
rect 35233 10625 35245 10628
rect 35279 10625 35291 10659
rect 35233 10619 35291 10625
rect 32088 10560 32720 10588
rect 32088 10548 32094 10560
rect 28902 10520 28908 10532
rect 27939 10492 28212 10520
rect 28276 10492 28908 10520
rect 27939 10489 27951 10492
rect 27893 10483 27951 10489
rect 21361 10455 21419 10461
rect 21361 10421 21373 10455
rect 21407 10421 21419 10455
rect 21361 10415 21419 10421
rect 21818 10412 21824 10464
rect 21876 10452 21882 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21876 10424 22017 10452
rect 21876 10412 21882 10424
rect 22005 10421 22017 10424
rect 22051 10452 22063 10455
rect 23290 10452 23296 10464
rect 22051 10424 23296 10452
rect 22051 10421 22063 10424
rect 22005 10415 22063 10421
rect 23290 10412 23296 10424
rect 23348 10452 23354 10464
rect 23842 10452 23848 10464
rect 23348 10424 23848 10452
rect 23348 10412 23354 10424
rect 23842 10412 23848 10424
rect 23900 10452 23906 10464
rect 24581 10455 24639 10461
rect 24581 10452 24593 10455
rect 23900 10424 24593 10452
rect 23900 10412 23906 10424
rect 24581 10421 24593 10424
rect 24627 10452 24639 10455
rect 24670 10452 24676 10464
rect 24627 10424 24676 10452
rect 24627 10421 24639 10424
rect 24581 10415 24639 10421
rect 24670 10412 24676 10424
rect 24728 10412 24734 10464
rect 26789 10455 26847 10461
rect 26789 10421 26801 10455
rect 26835 10452 26847 10455
rect 27154 10452 27160 10464
rect 26835 10424 27160 10452
rect 26835 10421 26847 10424
rect 26789 10415 26847 10421
rect 27154 10412 27160 10424
rect 27212 10412 27218 10464
rect 27798 10412 27804 10464
rect 27856 10452 27862 10464
rect 28077 10455 28135 10461
rect 28077 10452 28089 10455
rect 27856 10424 28089 10452
rect 27856 10412 27862 10424
rect 28077 10421 28089 10424
rect 28123 10421 28135 10455
rect 28184 10452 28212 10492
rect 28902 10480 28908 10492
rect 28960 10520 28966 10532
rect 29549 10523 29607 10529
rect 28960 10492 29215 10520
rect 28960 10480 28966 10492
rect 28810 10452 28816 10464
rect 28184 10424 28816 10452
rect 28077 10415 28135 10421
rect 28810 10412 28816 10424
rect 28868 10412 28874 10464
rect 29086 10412 29092 10464
rect 29144 10412 29150 10464
rect 29187 10452 29215 10492
rect 29549 10489 29561 10523
rect 29595 10520 29607 10523
rect 30282 10520 30288 10532
rect 29595 10492 30288 10520
rect 29595 10489 29607 10492
rect 29549 10483 29607 10489
rect 30282 10480 30288 10492
rect 30340 10480 30346 10532
rect 32309 10523 32367 10529
rect 32309 10520 32321 10523
rect 31726 10492 32321 10520
rect 29457 10455 29515 10461
rect 29457 10452 29469 10455
rect 29187 10424 29469 10452
rect 29457 10421 29469 10424
rect 29503 10421 29515 10455
rect 29457 10415 29515 10421
rect 30098 10412 30104 10464
rect 30156 10452 30162 10464
rect 31726 10452 31754 10492
rect 32309 10489 32321 10492
rect 32355 10489 32367 10523
rect 32309 10483 32367 10489
rect 32692 10464 32720 10560
rect 32769 10591 32827 10597
rect 32769 10557 32781 10591
rect 32815 10557 32827 10591
rect 32769 10551 32827 10557
rect 32784 10520 32812 10551
rect 32950 10548 32956 10600
rect 33008 10548 33014 10600
rect 33226 10548 33232 10600
rect 33284 10588 33290 10600
rect 33870 10588 33876 10600
rect 33284 10560 33876 10588
rect 33284 10548 33290 10560
rect 33870 10548 33876 10560
rect 33928 10548 33934 10600
rect 34698 10548 34704 10600
rect 34756 10588 34762 10600
rect 34977 10591 35035 10597
rect 34977 10588 34989 10591
rect 34756 10560 34989 10588
rect 34756 10548 34762 10560
rect 34977 10557 34989 10560
rect 35023 10557 35035 10591
rect 34977 10551 35035 10557
rect 33134 10520 33140 10532
rect 32784 10492 33140 10520
rect 33134 10480 33140 10492
rect 33192 10520 33198 10532
rect 33502 10520 33508 10532
rect 33192 10492 33508 10520
rect 33192 10480 33198 10492
rect 33502 10480 33508 10492
rect 33560 10480 33566 10532
rect 30156 10424 31754 10452
rect 30156 10412 30162 10424
rect 31846 10412 31852 10464
rect 31904 10412 31910 10464
rect 32674 10412 32680 10464
rect 32732 10452 32738 10464
rect 33594 10452 33600 10464
rect 32732 10424 33600 10452
rect 32732 10412 32738 10424
rect 33594 10412 33600 10424
rect 33652 10452 33658 10464
rect 33778 10452 33784 10464
rect 33652 10424 33784 10452
rect 33652 10412 33658 10424
rect 33778 10412 33784 10424
rect 33836 10412 33842 10464
rect 33962 10412 33968 10464
rect 34020 10452 34026 10464
rect 34609 10455 34667 10461
rect 34609 10452 34621 10455
rect 34020 10424 34621 10452
rect 34020 10412 34026 10424
rect 34609 10421 34621 10424
rect 34655 10421 34667 10455
rect 34609 10415 34667 10421
rect 1104 10362 36800 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 36800 10362
rect 1104 10288 36800 10310
rect 4798 10208 4804 10260
rect 4856 10248 4862 10260
rect 6917 10251 6975 10257
rect 4856 10220 6868 10248
rect 4856 10208 4862 10220
rect 5626 10140 5632 10192
rect 5684 10180 5690 10192
rect 6457 10183 6515 10189
rect 6457 10180 6469 10183
rect 5684 10152 6469 10180
rect 5684 10140 5690 10152
rect 6457 10149 6469 10152
rect 6503 10149 6515 10183
rect 6840 10180 6868 10220
rect 6917 10217 6929 10251
rect 6963 10248 6975 10251
rect 7282 10248 7288 10260
rect 6963 10220 7288 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7432 10220 7941 10248
rect 7432 10208 7438 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 9398 10208 9404 10260
rect 9456 10248 9462 10260
rect 12342 10248 12348 10260
rect 9456 10220 12348 10248
rect 9456 10208 9462 10220
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 12526 10208 12532 10260
rect 12584 10208 12590 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 13964 10220 14105 10248
rect 13964 10208 13970 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 14918 10208 14924 10260
rect 14976 10248 14982 10260
rect 15105 10251 15163 10257
rect 15105 10248 15117 10251
rect 14976 10220 15117 10248
rect 14976 10208 14982 10220
rect 15105 10217 15117 10220
rect 15151 10217 15163 10251
rect 15105 10211 15163 10217
rect 16758 10208 16764 10260
rect 16816 10208 16822 10260
rect 17770 10208 17776 10260
rect 17828 10248 17834 10260
rect 17865 10251 17923 10257
rect 17865 10248 17877 10251
rect 17828 10220 17877 10248
rect 17828 10208 17834 10220
rect 17865 10217 17877 10220
rect 17911 10217 17923 10251
rect 22370 10248 22376 10260
rect 17865 10211 17923 10217
rect 20916 10220 22376 10248
rect 7653 10183 7711 10189
rect 6840 10152 7604 10180
rect 6457 10143 6515 10149
rect 4614 10112 4620 10124
rect 3804 10084 4620 10112
rect 3804 10053 3832 10084
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10044 4031 10047
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 4019 10016 4077 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 4065 10013 4077 10016
rect 4111 10044 4123 10047
rect 4154 10044 4160 10056
rect 4111 10016 4160 10044
rect 4111 10013 4123 10016
rect 4065 10007 4123 10013
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4264 10053 4292 10084
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 5905 10115 5963 10121
rect 5905 10112 5917 10115
rect 5132 10084 5917 10112
rect 5132 10072 5138 10084
rect 5905 10081 5917 10084
rect 5951 10112 5963 10115
rect 5951 10084 7052 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10044 4491 10047
rect 4709 10047 4767 10053
rect 4709 10044 4721 10047
rect 4479 10016 4721 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 4709 10013 4721 10016
rect 4755 10044 4767 10047
rect 4798 10044 4804 10056
rect 4755 10016 4804 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 4798 10004 4804 10016
rect 4856 10044 4862 10056
rect 4982 10044 4988 10056
rect 4856 10016 4988 10044
rect 4856 10004 4862 10016
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10013 6147 10047
rect 6089 10007 6147 10013
rect 1486 9936 1492 9988
rect 1544 9936 1550 9988
rect 3881 9979 3939 9985
rect 3881 9945 3893 9979
rect 3927 9976 3939 9979
rect 4525 9979 4583 9985
rect 4525 9976 4537 9979
rect 3927 9948 4537 9976
rect 3927 9945 3939 9948
rect 3881 9939 3939 9945
rect 4525 9945 4537 9948
rect 4571 9945 4583 9979
rect 4525 9939 4583 9945
rect 4893 9979 4951 9985
rect 4893 9945 4905 9979
rect 4939 9976 4951 9979
rect 5077 9979 5135 9985
rect 5077 9976 5089 9979
rect 4939 9948 5089 9976
rect 4939 9945 4951 9948
rect 4893 9939 4951 9945
rect 5077 9945 5089 9948
rect 5123 9945 5135 9979
rect 5077 9939 5135 9945
rect 5261 9979 5319 9985
rect 5261 9945 5273 9979
rect 5307 9976 5319 9979
rect 5718 9976 5724 9988
rect 5307 9948 5724 9976
rect 5307 9945 5319 9948
rect 5261 9939 5319 9945
rect 5718 9936 5724 9948
rect 5776 9976 5782 9988
rect 6104 9976 6132 10007
rect 6362 10004 6368 10056
rect 6420 10044 6426 10056
rect 6733 10047 6791 10053
rect 6733 10044 6745 10047
rect 6420 10016 6745 10044
rect 6420 10004 6426 10016
rect 6733 10013 6745 10016
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 6914 10044 6920 10056
rect 6871 10016 6920 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 7024 10044 7052 10084
rect 7098 10072 7104 10124
rect 7156 10072 7162 10124
rect 7576 10112 7604 10152
rect 7653 10149 7665 10183
rect 7699 10180 7711 10183
rect 7699 10152 13584 10180
rect 7699 10149 7711 10152
rect 7653 10143 7711 10149
rect 7576 10084 8340 10112
rect 7193 10047 7251 10053
rect 7193 10044 7205 10047
rect 7024 10016 7205 10044
rect 7193 10013 7205 10016
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7374 10004 7380 10056
rect 7432 10004 7438 10056
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 6454 9976 6460 9988
rect 5776 9948 6460 9976
rect 5776 9936 5782 9948
rect 6454 9936 6460 9948
rect 6512 9936 6518 9988
rect 7760 9976 7788 10007
rect 7834 10004 7840 10056
rect 7892 10004 7898 10056
rect 8312 10044 8340 10084
rect 8938 10072 8944 10124
rect 8996 10072 9002 10124
rect 11701 10115 11759 10121
rect 11701 10112 11713 10115
rect 9048 10084 11713 10112
rect 9048 10044 9076 10084
rect 11701 10081 11713 10084
rect 11747 10081 11759 10115
rect 13354 10112 13360 10124
rect 11701 10075 11759 10081
rect 12360 10084 13360 10112
rect 12360 10053 12388 10084
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 13446 10072 13452 10124
rect 13504 10072 13510 10124
rect 13556 10112 13584 10152
rect 13630 10140 13636 10192
rect 13688 10180 13694 10192
rect 13688 10152 16620 10180
rect 13688 10140 13694 10152
rect 14737 10115 14795 10121
rect 13556 10084 13768 10112
rect 8312 10016 9076 10044
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 12434 10004 12440 10056
rect 12492 10004 12498 10056
rect 13464 10044 13492 10072
rect 13541 10047 13599 10053
rect 13541 10044 13553 10047
rect 13464 10016 13553 10044
rect 13541 10013 13553 10016
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 13630 10004 13636 10056
rect 13688 10004 13694 10056
rect 9490 9976 9496 9988
rect 7760 9948 9496 9976
rect 9490 9936 9496 9948
rect 9548 9936 9554 9988
rect 11606 9936 11612 9988
rect 11664 9976 11670 9988
rect 11882 9976 11888 9988
rect 11664 9948 11888 9976
rect 11664 9936 11670 9948
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 12253 9979 12311 9985
rect 11992 9948 12204 9976
rect 1578 9868 1584 9920
rect 1636 9868 1642 9920
rect 6273 9911 6331 9917
rect 6273 9877 6285 9911
rect 6319 9908 6331 9911
rect 6546 9908 6552 9920
rect 6319 9880 6552 9908
rect 6319 9877 6331 9880
rect 6273 9871 6331 9877
rect 6546 9868 6552 9880
rect 6604 9908 6610 9920
rect 6641 9911 6699 9917
rect 6641 9908 6653 9911
rect 6604 9880 6653 9908
rect 6604 9868 6610 9880
rect 6641 9877 6653 9880
rect 6687 9908 6699 9911
rect 7101 9911 7159 9917
rect 7101 9908 7113 9911
rect 6687 9880 7113 9908
rect 6687 9877 6699 9880
rect 6641 9871 6699 9877
rect 7101 9877 7113 9880
rect 7147 9877 7159 9911
rect 7101 9871 7159 9877
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 8570 9908 8576 9920
rect 8343 9880 8576 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 8938 9868 8944 9920
rect 8996 9908 9002 9920
rect 11992 9917 12020 9948
rect 9171 9911 9229 9917
rect 9171 9908 9183 9911
rect 8996 9880 9183 9908
rect 8996 9868 9002 9880
rect 9171 9877 9183 9880
rect 9217 9877 9229 9911
rect 9171 9871 9229 9877
rect 11977 9911 12035 9917
rect 11977 9877 11989 9911
rect 12023 9877 12035 9911
rect 11977 9871 12035 9877
rect 12066 9868 12072 9920
rect 12124 9868 12130 9920
rect 12176 9908 12204 9948
rect 12253 9945 12265 9979
rect 12299 9976 12311 9979
rect 13740 9976 13768 10084
rect 14737 10081 14749 10115
rect 14783 10112 14795 10115
rect 15010 10112 15016 10124
rect 14783 10084 15016 10112
rect 14783 10081 14795 10084
rect 14737 10075 14795 10081
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 16592 10112 16620 10152
rect 16592 10084 17264 10112
rect 14274 10004 14280 10056
rect 14332 10004 14338 10056
rect 14918 10004 14924 10056
rect 14976 10004 14982 10056
rect 17126 10004 17132 10056
rect 17184 10004 17190 10056
rect 17236 10044 17264 10084
rect 17310 10072 17316 10124
rect 17368 10112 17374 10124
rect 17586 10112 17592 10124
rect 17368 10084 17592 10112
rect 17368 10072 17374 10084
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 17880 10112 17908 10211
rect 17880 10084 18184 10112
rect 18156 10053 18184 10084
rect 19242 10072 19248 10124
rect 19300 10072 19306 10124
rect 18141 10047 18199 10053
rect 17236 10016 17908 10044
rect 17402 9976 17408 9988
rect 12299 9948 13676 9976
rect 13740 9948 17408 9976
rect 12299 9945 12311 9948
rect 12253 9939 12311 9945
rect 12713 9911 12771 9917
rect 12713 9908 12725 9911
rect 12176 9880 12725 9908
rect 12713 9877 12725 9880
rect 12759 9877 12771 9911
rect 12713 9871 12771 9877
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 13541 9911 13599 9917
rect 13541 9908 13553 9911
rect 12860 9880 13553 9908
rect 12860 9868 12866 9880
rect 13541 9877 13553 9880
rect 13587 9877 13599 9911
rect 13648 9908 13676 9948
rect 17402 9936 17408 9948
rect 17460 9936 17466 9988
rect 17770 9936 17776 9988
rect 17828 9936 17834 9988
rect 17880 9976 17908 10016
rect 18141 10013 18153 10047
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 20806 10004 20812 10056
rect 20864 10044 20870 10056
rect 20916 10053 20944 10220
rect 22370 10208 22376 10220
rect 22428 10248 22434 10260
rect 22428 10220 22784 10248
rect 22428 10208 22434 10220
rect 22094 10180 22100 10192
rect 21560 10152 22100 10180
rect 21560 10121 21588 10152
rect 22094 10140 22100 10152
rect 22152 10180 22158 10192
rect 22554 10180 22560 10192
rect 22152 10152 22560 10180
rect 22152 10140 22158 10152
rect 22554 10140 22560 10152
rect 22612 10140 22618 10192
rect 22756 10189 22784 10220
rect 23198 10208 23204 10260
rect 23256 10248 23262 10260
rect 23256 10220 26280 10248
rect 23256 10208 23262 10220
rect 22741 10183 22799 10189
rect 22741 10149 22753 10183
rect 22787 10149 22799 10183
rect 22741 10143 22799 10149
rect 26145 10183 26203 10189
rect 26145 10149 26157 10183
rect 26191 10149 26203 10183
rect 26252 10180 26280 10220
rect 27706 10208 27712 10260
rect 27764 10248 27770 10260
rect 27801 10251 27859 10257
rect 27801 10248 27813 10251
rect 27764 10220 27813 10248
rect 27764 10208 27770 10220
rect 27801 10217 27813 10220
rect 27847 10217 27859 10251
rect 27801 10211 27859 10217
rect 28626 10208 28632 10260
rect 28684 10248 28690 10260
rect 28721 10251 28779 10257
rect 28721 10248 28733 10251
rect 28684 10220 28733 10248
rect 28684 10208 28690 10220
rect 28721 10217 28733 10220
rect 28767 10217 28779 10251
rect 28721 10211 28779 10217
rect 28810 10208 28816 10260
rect 28868 10248 28874 10260
rect 30650 10248 30656 10260
rect 28868 10220 30656 10248
rect 28868 10208 28874 10220
rect 30650 10208 30656 10220
rect 30708 10208 30714 10260
rect 33229 10251 33287 10257
rect 33229 10217 33241 10251
rect 33275 10248 33287 10251
rect 34790 10248 34796 10260
rect 33275 10220 34796 10248
rect 33275 10217 33287 10220
rect 33229 10211 33287 10217
rect 34790 10208 34796 10220
rect 34848 10208 34854 10260
rect 29362 10180 29368 10192
rect 26252 10152 29368 10180
rect 26145 10143 26203 10149
rect 21545 10115 21603 10121
rect 21545 10112 21557 10115
rect 21100 10084 21557 10112
rect 21100 10053 21128 10084
rect 21545 10081 21557 10084
rect 21591 10081 21603 10115
rect 21545 10075 21603 10081
rect 21818 10072 21824 10124
rect 21876 10072 21882 10124
rect 21913 10115 21971 10121
rect 21913 10081 21925 10115
rect 21959 10112 21971 10115
rect 22002 10112 22008 10124
rect 21959 10084 22008 10112
rect 21959 10081 21971 10084
rect 21913 10075 21971 10081
rect 22002 10072 22008 10084
rect 22060 10112 22066 10124
rect 22060 10084 22784 10112
rect 22060 10072 22066 10084
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 20864 10016 20913 10044
rect 20864 10004 20870 10016
rect 20901 10013 20913 10016
rect 20947 10013 20959 10047
rect 20901 10007 20959 10013
rect 21085 10047 21143 10053
rect 21085 10013 21097 10047
rect 21131 10013 21143 10047
rect 21085 10007 21143 10013
rect 21358 10004 21364 10056
rect 21416 10004 21422 10056
rect 22756 10053 22784 10084
rect 24762 10072 24768 10124
rect 24820 10072 24826 10124
rect 25958 10072 25964 10124
rect 26016 10112 26022 10124
rect 26160 10112 26188 10143
rect 29362 10140 29368 10152
rect 29420 10140 29426 10192
rect 29825 10183 29883 10189
rect 29825 10149 29837 10183
rect 29871 10180 29883 10183
rect 30190 10180 30196 10192
rect 29871 10152 30196 10180
rect 29871 10149 29883 10152
rect 29825 10143 29883 10149
rect 30190 10140 30196 10152
rect 30248 10140 30254 10192
rect 32030 10180 32036 10192
rect 30484 10152 32036 10180
rect 26016 10084 28764 10112
rect 26016 10072 26022 10084
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10013 22615 10047
rect 22557 10007 22615 10013
rect 22741 10047 22799 10053
rect 22741 10013 22753 10047
rect 22787 10013 22799 10047
rect 22741 10007 22799 10013
rect 22925 10047 22983 10053
rect 22925 10013 22937 10047
rect 22971 10038 22983 10047
rect 22971 10013 23060 10038
rect 22925 10010 23060 10013
rect 22925 10007 22983 10010
rect 19512 9979 19570 9985
rect 17880 9948 18368 9976
rect 15654 9908 15660 9920
rect 13648 9880 15660 9908
rect 13541 9871 13599 9877
rect 15654 9868 15660 9880
rect 15712 9868 15718 9920
rect 17221 9911 17279 9917
rect 17221 9877 17233 9911
rect 17267 9908 17279 9911
rect 17494 9908 17500 9920
rect 17267 9880 17500 9908
rect 17267 9877 17279 9880
rect 17221 9871 17279 9877
rect 17494 9868 17500 9880
rect 17552 9868 17558 9920
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 18233 9911 18291 9917
rect 18233 9908 18245 9911
rect 18012 9880 18245 9908
rect 18012 9868 18018 9880
rect 18233 9877 18245 9880
rect 18279 9877 18291 9911
rect 18340 9908 18368 9948
rect 19512 9945 19524 9979
rect 19558 9976 19570 9979
rect 20717 9979 20775 9985
rect 20717 9976 20729 9979
rect 19558 9948 20729 9976
rect 19558 9945 19570 9948
rect 19512 9939 19570 9945
rect 20717 9945 20729 9948
rect 20763 9945 20775 9979
rect 20717 9939 20775 9945
rect 20993 9979 21051 9985
rect 20993 9945 21005 9979
rect 21039 9945 21051 9979
rect 20993 9939 21051 9945
rect 21223 9979 21281 9985
rect 21223 9945 21235 9979
rect 21269 9976 21281 9979
rect 21542 9976 21548 9988
rect 21269 9948 21548 9976
rect 21269 9945 21281 9948
rect 21223 9939 21281 9945
rect 20622 9908 20628 9920
rect 18340 9880 20628 9908
rect 18233 9871 18291 9877
rect 20622 9868 20628 9880
rect 20680 9868 20686 9920
rect 21008 9908 21036 9939
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 21726 9936 21732 9988
rect 21784 9976 21790 9988
rect 22030 9979 22088 9985
rect 22030 9976 22042 9979
rect 21784 9948 22042 9976
rect 21784 9936 21790 9948
rect 22030 9945 22042 9948
rect 22076 9945 22088 9979
rect 22030 9939 22088 9945
rect 21818 9908 21824 9920
rect 21008 9880 21824 9908
rect 21818 9868 21824 9880
rect 21876 9868 21882 9920
rect 22189 9911 22247 9917
rect 22189 9877 22201 9911
rect 22235 9908 22247 9911
rect 22462 9908 22468 9920
rect 22235 9880 22468 9908
rect 22235 9877 22247 9880
rect 22189 9871 22247 9877
rect 22462 9868 22468 9880
rect 22520 9868 22526 9920
rect 22572 9908 22600 10007
rect 23032 9976 23060 10010
rect 23106 10004 23112 10056
rect 23164 10004 23170 10056
rect 23198 10004 23204 10056
rect 23256 10004 23262 10056
rect 23477 10047 23535 10053
rect 23477 10013 23489 10047
rect 23523 10044 23535 10047
rect 23658 10044 23664 10056
rect 23523 10016 23664 10044
rect 23523 10013 23535 10016
rect 23477 10007 23535 10013
rect 23658 10004 23664 10016
rect 23716 10004 23722 10056
rect 24394 10004 24400 10056
rect 24452 10004 24458 10056
rect 26988 10053 27016 10084
rect 26973 10047 27031 10053
rect 26973 10013 26985 10047
rect 27019 10013 27031 10047
rect 26973 10007 27031 10013
rect 27154 10004 27160 10056
rect 27212 10004 27218 10056
rect 27246 10004 27252 10056
rect 27304 10044 27310 10056
rect 27341 10047 27399 10053
rect 27341 10044 27353 10047
rect 27304 10016 27353 10044
rect 27304 10004 27310 10016
rect 27341 10013 27353 10016
rect 27387 10013 27399 10047
rect 27341 10007 27399 10013
rect 27525 10047 27583 10053
rect 27525 10013 27537 10047
rect 27571 10044 27583 10047
rect 27571 10016 28488 10044
rect 27571 10013 27583 10016
rect 27525 10007 27583 10013
rect 23290 9976 23296 9988
rect 23032 9948 23296 9976
rect 23290 9936 23296 9948
rect 23348 9936 23354 9988
rect 25032 9979 25090 9985
rect 25032 9945 25044 9979
rect 25078 9976 25090 9979
rect 26050 9976 26056 9988
rect 25078 9948 26056 9976
rect 25078 9945 25090 9948
rect 25032 9939 25090 9945
rect 26050 9936 26056 9948
rect 26108 9936 26114 9988
rect 27172 9976 27200 10004
rect 27709 9979 27767 9985
rect 27709 9976 27721 9979
rect 27172 9948 27721 9976
rect 27709 9945 27721 9948
rect 27755 9945 27767 9979
rect 27709 9939 27767 9945
rect 22646 9908 22652 9920
rect 22572 9880 22652 9908
rect 22646 9868 22652 9880
rect 22704 9868 22710 9920
rect 23014 9868 23020 9920
rect 23072 9868 23078 9920
rect 23106 9868 23112 9920
rect 23164 9908 23170 9920
rect 23934 9908 23940 9920
rect 23164 9880 23940 9908
rect 23164 9868 23170 9880
rect 23934 9868 23940 9880
rect 23992 9868 23998 9920
rect 24581 9911 24639 9917
rect 24581 9877 24593 9911
rect 24627 9908 24639 9911
rect 24946 9908 24952 9920
rect 24627 9880 24952 9908
rect 24627 9877 24639 9880
rect 24581 9871 24639 9877
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 28460 9908 28488 10016
rect 28534 10004 28540 10056
rect 28592 10044 28598 10056
rect 28629 10047 28687 10053
rect 28629 10044 28641 10047
rect 28592 10016 28641 10044
rect 28592 10004 28598 10016
rect 28629 10013 28641 10016
rect 28675 10013 28687 10047
rect 28736 10044 28764 10084
rect 28902 10072 28908 10124
rect 28960 10072 28966 10124
rect 29086 10072 29092 10124
rect 29144 10112 29150 10124
rect 30484 10121 30512 10152
rect 32030 10140 32036 10152
rect 32088 10140 32094 10192
rect 34425 10183 34483 10189
rect 34425 10180 34437 10183
rect 33428 10152 34437 10180
rect 30469 10115 30527 10121
rect 30469 10112 30481 10115
rect 29144 10084 30481 10112
rect 29144 10072 29150 10084
rect 30469 10081 30481 10084
rect 30515 10081 30527 10115
rect 30469 10075 30527 10081
rect 31481 10115 31539 10121
rect 31481 10081 31493 10115
rect 31527 10112 31539 10115
rect 31662 10112 31668 10124
rect 31527 10084 31668 10112
rect 31527 10081 31539 10084
rect 31481 10075 31539 10081
rect 31662 10072 31668 10084
rect 31720 10072 31726 10124
rect 33134 10112 33140 10124
rect 32600 10084 33140 10112
rect 28736 10016 29960 10044
rect 28629 10007 28687 10013
rect 28905 9979 28963 9985
rect 28905 9945 28917 9979
rect 28951 9976 28963 9979
rect 29822 9976 29828 9988
rect 28951 9948 29828 9976
rect 28951 9945 28963 9948
rect 28905 9939 28963 9945
rect 29822 9936 29828 9948
rect 29880 9936 29886 9988
rect 29932 9976 29960 10016
rect 30098 10004 30104 10056
rect 30156 10004 30162 10056
rect 30193 10047 30251 10053
rect 30193 10013 30205 10047
rect 30239 10044 30251 10047
rect 30282 10044 30288 10056
rect 30239 10016 30288 10044
rect 30239 10013 30251 10016
rect 30193 10007 30251 10013
rect 30282 10004 30288 10016
rect 30340 10004 30346 10056
rect 31018 10004 31024 10056
rect 31076 10044 31082 10056
rect 31113 10047 31171 10053
rect 31113 10044 31125 10047
rect 31076 10016 31125 10044
rect 31076 10004 31082 10016
rect 31113 10013 31125 10016
rect 31159 10044 31171 10047
rect 31202 10044 31208 10056
rect 31159 10016 31208 10044
rect 31159 10013 31171 10016
rect 31113 10007 31171 10013
rect 31202 10004 31208 10016
rect 31260 10004 31266 10056
rect 31941 10047 31999 10053
rect 31941 10013 31953 10047
rect 31987 10044 31999 10047
rect 32214 10044 32220 10056
rect 31987 10016 32220 10044
rect 31987 10013 31999 10016
rect 31941 10007 31999 10013
rect 32214 10004 32220 10016
rect 32272 10044 32278 10056
rect 32600 10053 32628 10084
rect 33134 10072 33140 10084
rect 33192 10072 33198 10124
rect 33428 10121 33456 10152
rect 34425 10149 34437 10152
rect 34471 10149 34483 10183
rect 34425 10143 34483 10149
rect 33413 10115 33471 10121
rect 33413 10081 33425 10115
rect 33459 10081 33471 10115
rect 33413 10075 33471 10081
rect 33505 10115 33563 10121
rect 33505 10081 33517 10115
rect 33551 10112 33563 10115
rect 33778 10112 33784 10124
rect 33551 10084 33784 10112
rect 33551 10081 33563 10084
rect 33505 10075 33563 10081
rect 33778 10072 33784 10084
rect 33836 10072 33842 10124
rect 33962 10072 33968 10124
rect 34020 10072 34026 10124
rect 32401 10047 32459 10053
rect 32401 10044 32413 10047
rect 32272 10016 32413 10044
rect 32272 10004 32278 10016
rect 32401 10013 32413 10016
rect 32447 10013 32459 10047
rect 32401 10007 32459 10013
rect 32585 10047 32643 10053
rect 32585 10013 32597 10047
rect 32631 10013 32643 10047
rect 32585 10007 32643 10013
rect 32674 10004 32680 10056
rect 32732 10004 32738 10056
rect 32769 10047 32827 10053
rect 32769 10013 32781 10047
rect 32815 10044 32827 10047
rect 32858 10044 32864 10056
rect 32815 10016 32864 10044
rect 32815 10013 32827 10016
rect 32769 10007 32827 10013
rect 32858 10004 32864 10016
rect 32916 10004 32922 10056
rect 32950 10004 32956 10056
rect 33008 10004 33014 10056
rect 33597 10047 33655 10053
rect 33597 10013 33609 10047
rect 33643 10013 33655 10047
rect 33597 10007 33655 10013
rect 30742 9976 30748 9988
rect 29932 9948 30748 9976
rect 30742 9936 30748 9948
rect 30800 9976 30806 9988
rect 33612 9976 33640 10007
rect 33686 10004 33692 10056
rect 33744 10004 33750 10056
rect 34057 10047 34115 10053
rect 34057 10013 34069 10047
rect 34103 10044 34115 10047
rect 34330 10044 34336 10056
rect 34103 10016 34336 10044
rect 34103 10013 34115 10016
rect 34057 10007 34115 10013
rect 34330 10004 34336 10016
rect 34388 10004 34394 10056
rect 34793 10047 34851 10053
rect 34793 10013 34805 10047
rect 34839 10044 34851 10047
rect 35894 10044 35900 10056
rect 34839 10016 35900 10044
rect 34839 10013 34851 10016
rect 34793 10007 34851 10013
rect 35894 10004 35900 10016
rect 35952 10004 35958 10056
rect 30800 9948 33640 9976
rect 30800 9936 30806 9948
rect 29914 9908 29920 9920
rect 28460 9880 29920 9908
rect 29914 9868 29920 9880
rect 29972 9868 29978 9920
rect 30006 9868 30012 9920
rect 30064 9868 30070 9920
rect 30282 9868 30288 9920
rect 30340 9908 30346 9920
rect 31297 9911 31355 9917
rect 31297 9908 31309 9911
rect 30340 9880 31309 9908
rect 30340 9868 30346 9880
rect 31297 9877 31309 9880
rect 31343 9908 31355 9911
rect 31386 9908 31392 9920
rect 31343 9880 31392 9908
rect 31343 9877 31355 9880
rect 31297 9871 31355 9877
rect 31386 9868 31392 9880
rect 31444 9868 31450 9920
rect 31754 9868 31760 9920
rect 31812 9868 31818 9920
rect 31849 9911 31907 9917
rect 31849 9877 31861 9911
rect 31895 9908 31907 9911
rect 31938 9908 31944 9920
rect 31895 9880 31944 9908
rect 31895 9877 31907 9880
rect 31849 9871 31907 9877
rect 31938 9868 31944 9880
rect 31996 9868 32002 9920
rect 33134 9868 33140 9920
rect 33192 9868 33198 9920
rect 34882 9868 34888 9920
rect 34940 9868 34946 9920
rect 1104 9818 36800 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 36800 9818
rect 1104 9744 36800 9766
rect 6457 9707 6515 9713
rect 6457 9673 6469 9707
rect 6503 9704 6515 9707
rect 6546 9704 6552 9716
rect 6503 9676 6552 9704
rect 6503 9673 6515 9676
rect 6457 9667 6515 9673
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 8938 9664 8944 9716
rect 8996 9704 9002 9716
rect 11977 9707 12035 9713
rect 8996 9676 9628 9704
rect 8996 9664 9002 9676
rect 5353 9639 5411 9645
rect 5353 9605 5365 9639
rect 5399 9636 5411 9639
rect 5534 9636 5540 9648
rect 5399 9608 5540 9636
rect 5399 9605 5411 9608
rect 5353 9599 5411 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 7926 9636 7932 9648
rect 6748 9608 7932 9636
rect 4798 9528 4804 9580
rect 4856 9568 4862 9580
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 4856 9540 5089 9568
rect 4856 9528 4862 9540
rect 5077 9537 5089 9540
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5626 9568 5632 9580
rect 5215 9540 5632 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 6362 9528 6368 9580
rect 6420 9528 6426 9580
rect 6748 9577 6776 9608
rect 7926 9596 7932 9608
rect 7984 9636 7990 9648
rect 9600 9636 9628 9676
rect 11977 9673 11989 9707
rect 12023 9704 12035 9707
rect 12066 9704 12072 9716
rect 12023 9676 12072 9704
rect 12023 9673 12035 9676
rect 11977 9667 12035 9673
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 14918 9664 14924 9716
rect 14976 9704 14982 9716
rect 15105 9707 15163 9713
rect 15105 9704 15117 9707
rect 14976 9676 15117 9704
rect 14976 9664 14982 9676
rect 15105 9673 15117 9676
rect 15151 9673 15163 9707
rect 17770 9704 17776 9716
rect 15105 9667 15163 9673
rect 15212 9676 17776 9704
rect 10045 9639 10103 9645
rect 7984 9608 9444 9636
rect 9600 9608 9720 9636
rect 7984 9596 7990 9608
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8938 9568 8944 9580
rect 8343 9540 8944 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 9416 9577 9444 9608
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 9582 9528 9588 9580
rect 9640 9528 9646 9580
rect 9692 9577 9720 9608
rect 10045 9605 10057 9639
rect 10091 9636 10103 9639
rect 10091 9608 11836 9636
rect 10091 9605 10103 9608
rect 10045 9599 10103 9605
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9568 9735 9571
rect 9769 9571 9827 9577
rect 9769 9568 9781 9571
rect 9723 9540 9781 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 9769 9537 9781 9540
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 5442 9500 5448 9512
rect 5399 9472 5448 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 5442 9460 5448 9472
rect 5500 9500 5506 9512
rect 5902 9500 5908 9512
rect 5500 9472 5908 9500
rect 5500 9460 5506 9472
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 6549 9503 6607 9509
rect 6549 9500 6561 9503
rect 6512 9472 6561 9500
rect 6512 9460 6518 9472
rect 6549 9469 6561 9472
rect 6595 9469 6607 9503
rect 6549 9463 6607 9469
rect 8570 9460 8576 9512
rect 8628 9460 8634 9512
rect 9030 9460 9036 9512
rect 9088 9460 9094 9512
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9416 9472 10057 9500
rect 6733 9435 6791 9441
rect 6733 9401 6745 9435
rect 6779 9432 6791 9435
rect 7374 9432 7380 9444
rect 6779 9404 7380 9432
rect 6779 9401 6791 9404
rect 6733 9395 6791 9401
rect 7374 9392 7380 9404
rect 7432 9392 7438 9444
rect 8389 9435 8447 9441
rect 8389 9401 8401 9435
rect 8435 9432 8447 9435
rect 9048 9432 9076 9460
rect 9416 9441 9444 9472
rect 10045 9469 10057 9472
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 8435 9404 9076 9432
rect 9401 9435 9459 9441
rect 8435 9401 8447 9404
rect 8389 9395 8447 9401
rect 9401 9401 9413 9435
rect 9447 9401 9459 9435
rect 9401 9395 9459 9401
rect 9582 9392 9588 9444
rect 9640 9432 9646 9444
rect 9861 9435 9919 9441
rect 9861 9432 9873 9435
rect 9640 9404 9873 9432
rect 9640 9392 9646 9404
rect 9861 9401 9873 9404
rect 9907 9401 9919 9435
rect 10704 9432 10732 9531
rect 10778 9528 10784 9580
rect 10836 9528 10842 9580
rect 10870 9528 10876 9580
rect 10928 9528 10934 9580
rect 11514 9528 11520 9580
rect 11572 9528 11578 9580
rect 11808 9577 11836 9608
rect 12526 9596 12532 9648
rect 12584 9636 12590 9648
rect 12897 9639 12955 9645
rect 12897 9636 12909 9639
rect 12584 9608 12909 9636
rect 12584 9596 12590 9608
rect 12897 9605 12909 9608
rect 12943 9605 12955 9639
rect 12897 9599 12955 9605
rect 14550 9596 14556 9648
rect 14608 9636 14614 9648
rect 15212 9636 15240 9676
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 19337 9707 19395 9713
rect 19337 9673 19349 9707
rect 19383 9673 19395 9707
rect 19337 9667 19395 9673
rect 14608 9608 15240 9636
rect 14608 9596 14614 9608
rect 18874 9596 18880 9648
rect 18932 9636 18938 9648
rect 19352 9636 19380 9667
rect 21542 9664 21548 9716
rect 21600 9664 21606 9716
rect 22646 9664 22652 9716
rect 22704 9704 22710 9716
rect 23658 9704 23664 9716
rect 22704 9676 23664 9704
rect 22704 9664 22710 9676
rect 23658 9664 23664 9676
rect 23716 9664 23722 9716
rect 26050 9664 26056 9716
rect 26108 9704 26114 9716
rect 26145 9707 26203 9713
rect 26145 9704 26157 9707
rect 26108 9676 26157 9704
rect 26108 9664 26114 9676
rect 26145 9673 26157 9676
rect 26191 9673 26203 9707
rect 26145 9667 26203 9673
rect 30006 9664 30012 9716
rect 30064 9704 30070 9716
rect 31570 9704 31576 9716
rect 30064 9676 31576 9704
rect 30064 9664 30070 9676
rect 23014 9636 23020 9648
rect 18932 9608 19380 9636
rect 20916 9608 23020 9636
rect 18932 9596 18938 9608
rect 20916 9580 20944 9608
rect 23014 9596 23020 9608
rect 23072 9596 23078 9648
rect 24946 9596 24952 9648
rect 25004 9636 25010 9648
rect 25004 9608 25912 9636
rect 25004 9596 25010 9608
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 12618 9528 12624 9580
rect 12676 9528 12682 9580
rect 12802 9528 12808 9580
rect 12860 9528 12866 9580
rect 12986 9528 12992 9580
rect 13044 9577 13050 9580
rect 13044 9531 13052 9577
rect 13044 9528 13050 9531
rect 14826 9528 14832 9580
rect 14884 9568 14890 9580
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 14884 9540 15301 9568
rect 14884 9528 14890 9540
rect 15289 9537 15301 9540
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 16666 9528 16672 9580
rect 16724 9568 16730 9580
rect 17310 9568 17316 9580
rect 16724 9540 17316 9568
rect 16724 9528 16730 9540
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 18224 9571 18282 9577
rect 18224 9537 18236 9571
rect 18270 9568 18282 9571
rect 18270 9540 20668 9568
rect 18270 9537 18282 9540
rect 18224 9531 18282 9537
rect 11882 9460 11888 9512
rect 11940 9460 11946 9512
rect 12820 9432 12848 9528
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 15562 9500 15568 9512
rect 12943 9472 15568 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 17954 9500 17960 9512
rect 17328 9472 17960 9500
rect 17328 9444 17356 9472
rect 17954 9460 17960 9472
rect 18012 9460 18018 9512
rect 20640 9500 20668 9540
rect 20898 9528 20904 9580
rect 20956 9528 20962 9580
rect 21361 9571 21419 9577
rect 21361 9537 21373 9571
rect 21407 9568 21419 9571
rect 21726 9568 21732 9580
rect 21407 9540 21732 9568
rect 21407 9537 21419 9540
rect 21361 9531 21419 9537
rect 21726 9528 21732 9540
rect 21784 9528 21790 9580
rect 22066 9540 22508 9568
rect 20806 9500 20812 9512
rect 20640 9472 20812 9500
rect 20806 9460 20812 9472
rect 20864 9500 20870 9512
rect 21177 9503 21235 9509
rect 21177 9500 21189 9503
rect 20864 9472 21189 9500
rect 20864 9460 20870 9472
rect 21177 9469 21189 9472
rect 21223 9469 21235 9503
rect 22066 9500 22094 9540
rect 21177 9463 21235 9469
rect 21284 9472 22094 9500
rect 22373 9503 22431 9509
rect 10704 9404 12848 9432
rect 9861 9395 9919 9401
rect 16850 9392 16856 9444
rect 16908 9392 16914 9444
rect 17310 9392 17316 9444
rect 17368 9392 17374 9444
rect 21284 9432 21312 9472
rect 22373 9469 22385 9503
rect 22419 9469 22431 9503
rect 22373 9463 22431 9469
rect 19260 9404 21312 9432
rect 8478 9324 8484 9376
rect 8536 9324 8542 9376
rect 9306 9324 9312 9376
rect 9364 9324 9370 9376
rect 9490 9324 9496 9376
rect 9548 9364 9554 9376
rect 11057 9367 11115 9373
rect 11057 9364 11069 9367
rect 9548 9336 11069 9364
rect 9548 9324 9554 9336
rect 11057 9333 11069 9336
rect 11103 9333 11115 9367
rect 11057 9327 11115 9333
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 11388 9336 11621 9364
rect 11388 9324 11394 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 11609 9327 11667 9333
rect 17218 9324 17224 9376
rect 17276 9364 17282 9376
rect 19260 9364 19288 9404
rect 22002 9392 22008 9444
rect 22060 9432 22066 9444
rect 22388 9432 22416 9463
rect 22060 9404 22416 9432
rect 22060 9392 22066 9404
rect 17276 9336 19288 9364
rect 17276 9324 17282 9336
rect 21082 9324 21088 9376
rect 21140 9324 21146 9376
rect 22480 9364 22508 9540
rect 23566 9528 23572 9580
rect 23624 9528 23630 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 23676 9540 23949 9568
rect 22554 9460 22560 9512
rect 22612 9500 22618 9512
rect 22649 9503 22707 9509
rect 22649 9500 22661 9503
rect 22612 9472 22661 9500
rect 22612 9460 22618 9472
rect 22649 9469 22661 9472
rect 22695 9500 22707 9503
rect 23198 9500 23204 9512
rect 22695 9472 23204 9500
rect 22695 9469 22707 9472
rect 22649 9463 22707 9469
rect 23198 9460 23204 9472
rect 23256 9460 23262 9512
rect 22922 9392 22928 9444
rect 22980 9432 22986 9444
rect 23676 9432 23704 9540
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 24210 9528 24216 9580
rect 24268 9528 24274 9580
rect 24670 9528 24676 9580
rect 24728 9528 24734 9580
rect 25130 9528 25136 9580
rect 25188 9528 25194 9580
rect 25884 9577 25912 9608
rect 30098 9596 30104 9648
rect 30156 9596 30162 9648
rect 30208 9645 30236 9676
rect 31570 9664 31576 9676
rect 31628 9704 31634 9716
rect 31938 9704 31944 9716
rect 31628 9676 31944 9704
rect 31628 9664 31634 9676
rect 31938 9664 31944 9676
rect 31996 9704 32002 9716
rect 32677 9707 32735 9713
rect 32677 9704 32689 9707
rect 31996 9676 32689 9704
rect 31996 9664 32002 9676
rect 32677 9673 32689 9676
rect 32723 9673 32735 9707
rect 32677 9667 32735 9673
rect 33686 9664 33692 9716
rect 33744 9704 33750 9716
rect 33781 9707 33839 9713
rect 33781 9704 33793 9707
rect 33744 9676 33793 9704
rect 33744 9664 33750 9676
rect 33781 9673 33793 9676
rect 33827 9673 33839 9707
rect 34882 9704 34888 9716
rect 33781 9667 33839 9673
rect 33888 9676 34888 9704
rect 30193 9639 30251 9645
rect 30193 9605 30205 9639
rect 30239 9605 30251 9639
rect 33134 9636 33140 9648
rect 30193 9599 30251 9605
rect 30392 9608 30604 9636
rect 25869 9571 25927 9577
rect 25869 9537 25881 9571
rect 25915 9537 25927 9571
rect 25869 9531 25927 9537
rect 25958 9528 25964 9580
rect 26016 9528 26022 9580
rect 29822 9528 29828 9580
rect 29880 9568 29886 9580
rect 30392 9577 30420 9608
rect 30576 9577 30604 9608
rect 32600 9608 33140 9636
rect 30009 9571 30067 9577
rect 30009 9568 30021 9571
rect 29880 9540 30021 9568
rect 29880 9528 29886 9540
rect 30009 9537 30021 9540
rect 30055 9537 30067 9571
rect 30009 9531 30067 9537
rect 30377 9571 30435 9577
rect 30377 9537 30389 9571
rect 30423 9537 30435 9571
rect 30377 9531 30435 9537
rect 30469 9571 30527 9577
rect 30469 9537 30481 9571
rect 30515 9537 30527 9571
rect 30469 9531 30527 9537
rect 30561 9571 30619 9577
rect 30561 9537 30573 9571
rect 30607 9537 30619 9571
rect 30561 9531 30619 9537
rect 24026 9460 24032 9512
rect 24084 9500 24090 9512
rect 25501 9503 25559 9509
rect 25501 9500 25513 9503
rect 24084 9472 25513 9500
rect 24084 9460 24090 9472
rect 25501 9469 25513 9472
rect 25547 9469 25559 9503
rect 25501 9463 25559 9469
rect 29270 9460 29276 9512
rect 29328 9500 29334 9512
rect 30392 9500 30420 9531
rect 29328 9472 30420 9500
rect 29328 9460 29334 9472
rect 22980 9404 23704 9432
rect 23753 9435 23811 9441
rect 22980 9392 22986 9404
rect 23753 9401 23765 9435
rect 23799 9432 23811 9435
rect 24854 9432 24860 9444
rect 23799 9404 24860 9432
rect 23799 9401 23811 9404
rect 23753 9395 23811 9401
rect 24854 9392 24860 9404
rect 24912 9392 24918 9444
rect 27706 9392 27712 9444
rect 27764 9432 27770 9444
rect 28902 9432 28908 9444
rect 27764 9404 28908 9432
rect 27764 9392 27770 9404
rect 28902 9392 28908 9404
rect 28960 9432 28966 9444
rect 30484 9432 30512 9531
rect 30742 9528 30748 9580
rect 30800 9528 30806 9580
rect 31754 9528 31760 9580
rect 31812 9568 31818 9580
rect 32600 9577 32628 9608
rect 33134 9596 33140 9608
rect 33192 9596 33198 9648
rect 33229 9639 33287 9645
rect 33229 9605 33241 9639
rect 33275 9636 33287 9639
rect 33594 9636 33600 9648
rect 33275 9608 33600 9636
rect 33275 9605 33287 9608
rect 33229 9599 33287 9605
rect 33594 9596 33600 9608
rect 33652 9596 33658 9648
rect 32309 9571 32367 9577
rect 32309 9568 32321 9571
rect 31812 9540 32321 9568
rect 31812 9528 31818 9540
rect 32309 9537 32321 9540
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 32585 9571 32643 9577
rect 32585 9537 32597 9571
rect 32631 9537 32643 9571
rect 32585 9531 32643 9537
rect 33042 9528 33048 9580
rect 33100 9568 33106 9580
rect 33505 9571 33563 9577
rect 33505 9568 33517 9571
rect 33100 9540 33517 9568
rect 33100 9528 33106 9540
rect 33505 9537 33517 9540
rect 33551 9568 33563 9571
rect 33888 9568 33916 9676
rect 34882 9664 34888 9676
rect 34940 9664 34946 9716
rect 33551 9540 33916 9568
rect 34149 9571 34207 9577
rect 33551 9537 33563 9540
rect 33505 9531 33563 9537
rect 34149 9537 34161 9571
rect 34195 9537 34207 9571
rect 34149 9531 34207 9537
rect 33226 9460 33232 9512
rect 33284 9500 33290 9512
rect 33321 9503 33379 9509
rect 33321 9500 33333 9503
rect 33284 9472 33333 9500
rect 33284 9460 33290 9472
rect 33321 9469 33333 9472
rect 33367 9469 33379 9503
rect 33321 9463 33379 9469
rect 32401 9435 32459 9441
rect 32401 9432 32413 9435
rect 28960 9404 32413 9432
rect 28960 9392 28966 9404
rect 26418 9364 26424 9376
rect 22480 9336 26424 9364
rect 26418 9324 26424 9336
rect 26476 9324 26482 9376
rect 29825 9367 29883 9373
rect 29825 9333 29837 9367
rect 29871 9364 29883 9367
rect 30466 9364 30472 9376
rect 29871 9336 30472 9364
rect 29871 9333 29883 9336
rect 29825 9327 29883 9333
rect 30466 9324 30472 9336
rect 30524 9324 30530 9376
rect 30576 9373 30604 9404
rect 32401 9401 32413 9404
rect 32447 9401 32459 9435
rect 34164 9432 34192 9531
rect 34238 9460 34244 9512
rect 34296 9460 34302 9512
rect 34330 9460 34336 9512
rect 34388 9460 34394 9512
rect 32401 9395 32459 9401
rect 33152 9404 34192 9432
rect 33152 9376 33180 9404
rect 30561 9367 30619 9373
rect 30561 9333 30573 9367
rect 30607 9333 30619 9367
rect 30561 9327 30619 9333
rect 30926 9324 30932 9376
rect 30984 9324 30990 9376
rect 32125 9367 32183 9373
rect 32125 9333 32137 9367
rect 32171 9364 32183 9367
rect 32306 9364 32312 9376
rect 32171 9336 32312 9364
rect 32171 9333 32183 9336
rect 32125 9327 32183 9333
rect 32306 9324 32312 9336
rect 32364 9324 32370 9376
rect 32493 9367 32551 9373
rect 32493 9333 32505 9367
rect 32539 9364 32551 9367
rect 33134 9364 33140 9376
rect 32539 9336 33140 9364
rect 32539 9333 32551 9336
rect 32493 9327 32551 9333
rect 33134 9324 33140 9336
rect 33192 9324 33198 9376
rect 33410 9324 33416 9376
rect 33468 9324 33474 9376
rect 33689 9367 33747 9373
rect 33689 9333 33701 9367
rect 33735 9364 33747 9367
rect 33870 9364 33876 9376
rect 33735 9336 33876 9364
rect 33735 9333 33747 9336
rect 33689 9327 33747 9333
rect 33870 9324 33876 9336
rect 33928 9324 33934 9376
rect 1104 9274 36800 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 36800 9274
rect 1104 9200 36800 9222
rect 4614 9120 4620 9172
rect 4672 9120 4678 9172
rect 10962 9120 10968 9172
rect 11020 9120 11026 9172
rect 11330 9120 11336 9172
rect 11388 9160 11394 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 11388 9132 13001 9160
rect 11388 9120 11394 9132
rect 12989 9129 13001 9132
rect 13035 9160 13047 9163
rect 13170 9160 13176 9172
rect 13035 9132 13176 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 13357 9163 13415 9169
rect 13357 9129 13369 9163
rect 13403 9160 13415 9163
rect 14274 9160 14280 9172
rect 13403 9132 14280 9160
rect 13403 9129 13415 9132
rect 13357 9123 13415 9129
rect 14274 9120 14280 9132
rect 14332 9120 14338 9172
rect 14458 9120 14464 9172
rect 14516 9120 14522 9172
rect 14826 9120 14832 9172
rect 14884 9120 14890 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 23109 9163 23167 9169
rect 23109 9160 23121 9163
rect 22152 9132 23121 9160
rect 22152 9120 22158 9132
rect 23109 9129 23121 9132
rect 23155 9129 23167 9163
rect 23109 9123 23167 9129
rect 10505 9095 10563 9101
rect 10505 9061 10517 9095
rect 10551 9092 10563 9095
rect 11882 9092 11888 9104
rect 10551 9064 11888 9092
rect 10551 9061 10563 9064
rect 10505 9055 10563 9061
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 11974 9052 11980 9104
rect 12032 9092 12038 9104
rect 12158 9092 12164 9104
rect 12032 9064 12164 9092
rect 12032 9052 12038 9064
rect 12158 9052 12164 9064
rect 12216 9092 12222 9104
rect 16485 9095 16543 9101
rect 16485 9092 16497 9095
rect 12216 9064 16497 9092
rect 12216 9052 12222 9064
rect 16485 9061 16497 9064
rect 16531 9061 16543 9095
rect 16485 9055 16543 9061
rect 16850 9052 16856 9104
rect 16908 9052 16914 9104
rect 20990 9052 20996 9104
rect 21048 9092 21054 9104
rect 22002 9092 22008 9104
rect 21048 9064 22008 9092
rect 21048 9052 21054 9064
rect 22002 9052 22008 9064
rect 22060 9092 22066 9104
rect 22060 9064 23060 9092
rect 22060 9052 22066 9064
rect 7926 8984 7932 9036
rect 7984 9024 7990 9036
rect 11241 9027 11299 9033
rect 7984 8996 10640 9024
rect 7984 8984 7990 8996
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4433 8959 4491 8965
rect 4433 8956 4445 8959
rect 4212 8928 4445 8956
rect 4212 8916 4218 8928
rect 4433 8925 4445 8928
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 4448 8888 4476 8919
rect 10410 8916 10416 8968
rect 10468 8916 10474 8968
rect 10612 8965 10640 8996
rect 11241 8993 11253 9027
rect 11287 9024 11299 9027
rect 11514 9024 11520 9036
rect 11287 8996 11520 9024
rect 11287 8993 11299 8996
rect 11241 8987 11299 8993
rect 11514 8984 11520 8996
rect 11572 9024 11578 9036
rect 16117 9027 16175 9033
rect 11572 8996 12434 9024
rect 11572 8984 11578 8996
rect 10597 8959 10655 8965
rect 10597 8925 10609 8959
rect 10643 8925 10655 8959
rect 10597 8919 10655 8925
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 10502 8888 10508 8900
rect 4448 8860 10508 8888
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 4893 8823 4951 8829
rect 4893 8789 4905 8823
rect 4939 8820 4951 8823
rect 5258 8820 5264 8832
rect 4939 8792 5264 8820
rect 4939 8789 4951 8792
rect 4893 8783 4951 8789
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 10612 8820 10640 8919
rect 11164 8888 11192 8919
rect 11330 8916 11336 8968
rect 11388 8916 11394 8968
rect 11422 8916 11428 8968
rect 11480 8916 11486 8968
rect 11606 8916 11612 8968
rect 11664 8916 11670 8968
rect 12406 8956 12434 8996
rect 16117 8993 16129 9027
rect 16163 9024 16175 9027
rect 16868 9024 16896 9052
rect 16163 8996 16896 9024
rect 21361 9027 21419 9033
rect 16163 8993 16175 8996
rect 16117 8987 16175 8993
rect 21361 8993 21373 9027
rect 21407 9024 21419 9027
rect 21407 8996 21772 9024
rect 21407 8993 21419 8996
rect 21361 8987 21419 8993
rect 12710 8956 12716 8968
rect 12406 8928 12716 8956
rect 12710 8916 12716 8928
rect 12768 8956 12774 8968
rect 12897 8959 12955 8965
rect 12897 8956 12909 8959
rect 12768 8928 12909 8956
rect 12768 8916 12774 8928
rect 12897 8925 12909 8928
rect 12943 8956 12955 8959
rect 14369 8959 14427 8965
rect 14369 8956 14381 8959
rect 12943 8928 14381 8956
rect 12943 8925 12955 8928
rect 12897 8919 12955 8925
rect 14369 8925 14381 8928
rect 14415 8956 14427 8959
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 14415 8928 15853 8956
rect 14415 8925 14427 8928
rect 14369 8919 14427 8925
rect 15841 8925 15853 8928
rect 15887 8925 15899 8959
rect 16577 8959 16635 8965
rect 16577 8956 16589 8959
rect 15841 8919 15899 8925
rect 15948 8928 16589 8956
rect 11974 8888 11980 8900
rect 11164 8860 11980 8888
rect 11974 8848 11980 8860
rect 12032 8848 12038 8900
rect 12434 8888 12440 8900
rect 12268 8860 12440 8888
rect 12268 8820 12296 8860
rect 12434 8848 12440 8860
rect 12492 8848 12498 8900
rect 12618 8848 12624 8900
rect 12676 8888 12682 8900
rect 15948 8888 15976 8928
rect 16577 8925 16589 8928
rect 16623 8956 16635 8959
rect 16853 8959 16911 8965
rect 16623 8928 16804 8956
rect 16623 8925 16635 8928
rect 16577 8919 16635 8925
rect 12676 8860 15976 8888
rect 12676 8848 12682 8860
rect 16206 8848 16212 8900
rect 16264 8888 16270 8900
rect 16301 8891 16359 8897
rect 16301 8888 16313 8891
rect 16264 8860 16313 8888
rect 16264 8848 16270 8860
rect 16301 8857 16313 8860
rect 16347 8857 16359 8891
rect 16301 8851 16359 8857
rect 16482 8848 16488 8900
rect 16540 8888 16546 8900
rect 16669 8891 16727 8897
rect 16669 8888 16681 8891
rect 16540 8860 16681 8888
rect 16540 8848 16546 8860
rect 16669 8857 16681 8860
rect 16715 8857 16727 8891
rect 16776 8888 16804 8928
rect 16853 8925 16865 8959
rect 16899 8956 16911 8959
rect 17218 8956 17224 8968
rect 16899 8928 17224 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 17310 8916 17316 8968
rect 17368 8916 17374 8968
rect 17580 8959 17638 8965
rect 17580 8925 17592 8959
rect 17626 8956 17638 8959
rect 20898 8956 20904 8968
rect 17626 8928 20904 8956
rect 17626 8925 17638 8928
rect 17580 8919 17638 8925
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 21266 8916 21272 8968
rect 21324 8956 21330 8968
rect 21637 8959 21695 8965
rect 21637 8956 21649 8959
rect 21324 8928 21649 8956
rect 21324 8916 21330 8928
rect 21637 8925 21649 8928
rect 21683 8925 21695 8959
rect 21744 8956 21772 8996
rect 21910 8984 21916 9036
rect 21968 9024 21974 9036
rect 22741 9027 22799 9033
rect 22741 9024 22753 9027
rect 21968 8996 22753 9024
rect 21968 8984 21974 8996
rect 22741 8993 22753 8996
rect 22787 8993 22799 9027
rect 22741 8987 22799 8993
rect 22922 8984 22928 9036
rect 22980 8984 22986 9036
rect 22373 8959 22431 8965
rect 22373 8956 22385 8959
rect 21744 8928 22385 8956
rect 21637 8919 21695 8925
rect 22373 8925 22385 8928
rect 22419 8925 22431 8959
rect 22373 8919 22431 8925
rect 17037 8891 17095 8897
rect 17037 8888 17049 8891
rect 16776 8860 17049 8888
rect 16669 8851 16727 8857
rect 17037 8857 17049 8860
rect 17083 8857 17095 8891
rect 22388 8888 22416 8919
rect 22554 8916 22560 8968
rect 22612 8916 22618 8968
rect 23032 8965 23060 9064
rect 23124 9024 23152 9123
rect 23566 9120 23572 9172
rect 23624 9120 23630 9172
rect 23661 9163 23719 9169
rect 23661 9129 23673 9163
rect 23707 9129 23719 9163
rect 23661 9123 23719 9129
rect 23198 9052 23204 9104
rect 23256 9092 23262 9104
rect 23676 9092 23704 9123
rect 24026 9120 24032 9172
rect 24084 9120 24090 9172
rect 26418 9120 26424 9172
rect 26476 9160 26482 9172
rect 26476 9132 28212 9160
rect 26476 9120 26482 9132
rect 23256 9064 23704 9092
rect 23256 9052 23262 9064
rect 27338 9052 27344 9104
rect 27396 9092 27402 9104
rect 27525 9095 27583 9101
rect 27525 9092 27537 9095
rect 27396 9064 27537 9092
rect 27396 9052 27402 9064
rect 27525 9061 27537 9064
rect 27571 9061 27583 9095
rect 28184 9092 28212 9132
rect 29914 9120 29920 9172
rect 29972 9160 29978 9172
rect 34238 9160 34244 9172
rect 29972 9132 34244 9160
rect 29972 9120 29978 9132
rect 34238 9120 34244 9132
rect 34296 9120 34302 9172
rect 27525 9055 27583 9061
rect 27632 9064 28120 9092
rect 28184 9064 31754 9092
rect 23124 8996 23704 9024
rect 23017 8959 23075 8965
rect 23017 8925 23029 8959
rect 23063 8925 23075 8959
rect 23017 8919 23075 8925
rect 23385 8959 23443 8965
rect 23385 8925 23397 8959
rect 23431 8956 23443 8959
rect 23566 8956 23572 8968
rect 23431 8928 23572 8956
rect 23431 8925 23443 8928
rect 23385 8919 23443 8925
rect 23400 8888 23428 8919
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 23676 8965 23704 8996
rect 26786 8984 26792 9036
rect 26844 9024 26850 9036
rect 27632 9024 27660 9064
rect 26844 8996 27660 9024
rect 27816 8996 28028 9024
rect 26844 8984 26850 8996
rect 27816 8968 27844 8996
rect 23661 8959 23719 8965
rect 23661 8925 23673 8959
rect 23707 8925 23719 8959
rect 23661 8919 23719 8925
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 23934 8956 23940 8968
rect 23891 8928 23940 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 23934 8916 23940 8928
rect 23992 8956 23998 8968
rect 25130 8956 25136 8968
rect 23992 8928 25136 8956
rect 23992 8916 23998 8928
rect 25130 8916 25136 8928
rect 25188 8916 25194 8968
rect 27798 8916 27804 8968
rect 27856 8916 27862 8968
rect 27890 8916 27896 8968
rect 27948 8916 27954 8968
rect 28000 8965 28028 8996
rect 27986 8959 28044 8965
rect 27986 8925 27998 8959
rect 28032 8925 28044 8959
rect 28092 8956 28120 9064
rect 31726 9024 31754 9064
rect 36170 9024 36176 9036
rect 31726 8996 36176 9024
rect 36170 8984 36176 8996
rect 36228 8984 36234 9036
rect 28358 8959 28416 8965
rect 28358 8956 28370 8959
rect 28092 8928 28370 8956
rect 27986 8919 28044 8925
rect 28358 8925 28370 8928
rect 28404 8925 28416 8959
rect 28358 8919 28416 8925
rect 30377 8959 30435 8965
rect 30377 8925 30389 8959
rect 30423 8956 30435 8959
rect 30926 8956 30932 8968
rect 30423 8928 30932 8956
rect 30423 8925 30435 8928
rect 30377 8919 30435 8925
rect 30926 8916 30932 8928
rect 30984 8916 30990 8968
rect 22388 8860 23428 8888
rect 27525 8891 27583 8897
rect 17037 8851 17095 8857
rect 27525 8857 27537 8891
rect 27571 8857 27583 8891
rect 27525 8851 27583 8857
rect 27709 8891 27767 8897
rect 27709 8857 27721 8891
rect 27755 8888 27767 8891
rect 28169 8891 28227 8897
rect 28169 8888 28181 8891
rect 27755 8860 28181 8888
rect 27755 8857 27767 8860
rect 27709 8851 27767 8857
rect 28169 8857 28181 8860
rect 28215 8857 28227 8891
rect 28169 8851 28227 8857
rect 10612 8792 12296 8820
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 15194 8820 15200 8832
rect 12400 8792 15200 8820
rect 12400 8780 12406 8792
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 15286 8780 15292 8832
rect 15344 8820 15350 8832
rect 15473 8823 15531 8829
rect 15473 8820 15485 8823
rect 15344 8792 15485 8820
rect 15344 8780 15350 8792
rect 15473 8789 15485 8792
rect 15519 8789 15531 8823
rect 15473 8783 15531 8789
rect 15933 8823 15991 8829
rect 15933 8789 15945 8823
rect 15979 8820 15991 8823
rect 16022 8820 16028 8832
rect 15979 8792 16028 8820
rect 15979 8789 15991 8792
rect 15933 8783 15991 8789
rect 16022 8780 16028 8792
rect 16080 8780 16086 8832
rect 16390 8780 16396 8832
rect 16448 8780 16454 8832
rect 18690 8780 18696 8832
rect 18748 8780 18754 8832
rect 27540 8820 27568 8851
rect 27890 8820 27896 8832
rect 27540 8792 27896 8820
rect 27890 8780 27896 8792
rect 27948 8780 27954 8832
rect 28184 8820 28212 8851
rect 28258 8848 28264 8900
rect 28316 8848 28322 8900
rect 31846 8888 31852 8900
rect 28368 8860 31852 8888
rect 28368 8820 28396 8860
rect 31846 8848 31852 8860
rect 31904 8848 31910 8900
rect 28184 8792 28396 8820
rect 28537 8823 28595 8829
rect 28537 8789 28549 8823
rect 28583 8820 28595 8823
rect 29178 8820 29184 8832
rect 28583 8792 29184 8820
rect 28583 8789 28595 8792
rect 28537 8783 28595 8789
rect 29178 8780 29184 8792
rect 29236 8780 29242 8832
rect 30469 8823 30527 8829
rect 30469 8789 30481 8823
rect 30515 8820 30527 8823
rect 30558 8820 30564 8832
rect 30515 8792 30564 8820
rect 30515 8789 30527 8792
rect 30469 8783 30527 8789
rect 30558 8780 30564 8792
rect 30616 8780 30622 8832
rect 32122 8780 32128 8832
rect 32180 8820 32186 8832
rect 33042 8820 33048 8832
rect 32180 8792 33048 8820
rect 32180 8780 32186 8792
rect 33042 8780 33048 8792
rect 33100 8780 33106 8832
rect 1104 8730 36800 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 36800 8730
rect 1104 8656 36800 8678
rect 10410 8576 10416 8628
rect 10468 8576 10474 8628
rect 12618 8616 12624 8628
rect 10520 8588 12624 8616
rect 8570 8508 8576 8560
rect 8628 8548 8634 8560
rect 10520 8548 10548 8588
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 13817 8619 13875 8625
rect 12952 8588 13037 8616
rect 12952 8576 12958 8588
rect 8628 8520 10548 8548
rect 8628 8508 8634 8520
rect 13009 8511 13037 8588
rect 13817 8585 13829 8619
rect 13863 8616 13875 8619
rect 13998 8616 14004 8628
rect 13863 8588 14004 8616
rect 13863 8585 13875 8588
rect 13817 8579 13875 8585
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8585 15991 8619
rect 15933 8579 15991 8585
rect 15948 8548 15976 8579
rect 16022 8576 16028 8628
rect 16080 8616 16086 8628
rect 16574 8616 16580 8628
rect 16080 8588 16580 8616
rect 16080 8576 16086 8588
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 22554 8616 22560 8628
rect 21836 8588 22560 8616
rect 14016 8520 15976 8548
rect 12993 8505 13051 8511
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8480 7159 8483
rect 7190 8480 7196 8492
rect 7147 8452 7196 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9364 8452 9781 8480
rect 9364 8440 9370 8452
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 9769 8443 9827 8449
rect 9876 8452 12541 8480
rect 5810 8372 5816 8424
rect 5868 8412 5874 8424
rect 9876 8412 9904 8452
rect 12529 8449 12541 8452
rect 12575 8480 12587 8483
rect 12618 8480 12624 8492
rect 12575 8452 12624 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 12618 8440 12624 8452
rect 12676 8440 12682 8492
rect 12802 8440 12808 8492
rect 12860 8440 12866 8492
rect 12993 8471 13005 8505
rect 13039 8471 13051 8505
rect 12993 8465 13051 8471
rect 13357 8483 13415 8489
rect 13357 8449 13369 8483
rect 13403 8480 13415 8483
rect 13722 8480 13728 8492
rect 13403 8452 13728 8480
rect 13403 8449 13415 8452
rect 13357 8443 13415 8449
rect 13722 8440 13728 8452
rect 13780 8480 13786 8492
rect 14016 8489 14044 8520
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 17129 8551 17187 8557
rect 17129 8548 17141 8551
rect 16448 8520 17141 8548
rect 16448 8508 16454 8520
rect 17129 8517 17141 8520
rect 17175 8517 17187 8551
rect 17129 8511 17187 8517
rect 20070 8508 20076 8560
rect 20128 8548 20134 8560
rect 20128 8520 21312 8548
rect 20128 8508 20134 8520
rect 21284 8492 21312 8520
rect 14001 8483 14059 8489
rect 14001 8480 14013 8483
rect 13780 8452 14013 8480
rect 13780 8440 13786 8452
rect 14001 8449 14013 8452
rect 14047 8449 14059 8483
rect 14642 8480 14648 8492
rect 14001 8443 14059 8449
rect 14108 8452 14648 8480
rect 5868 8384 9904 8412
rect 5868 8372 5874 8384
rect 9950 8372 9956 8424
rect 10008 8372 10014 8424
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 14108 8412 14136 8452
rect 12492 8384 14136 8412
rect 12492 8372 12498 8384
rect 14182 8372 14188 8424
rect 14240 8412 14246 8424
rect 14384 8421 14412 8452
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 14820 8483 14878 8489
rect 14820 8449 14832 8483
rect 14866 8480 14878 8483
rect 15102 8480 15108 8492
rect 14866 8452 15108 8480
rect 14866 8449 14878 8452
rect 14820 8443 14878 8449
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 15194 8440 15200 8492
rect 15252 8480 15258 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 15252 8452 16957 8480
rect 15252 8440 15258 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17218 8440 17224 8492
rect 17276 8440 17282 8492
rect 20990 8440 20996 8492
rect 21048 8480 21054 8492
rect 21085 8483 21143 8489
rect 21085 8480 21097 8483
rect 21048 8452 21097 8480
rect 21048 8440 21054 8452
rect 21085 8449 21097 8452
rect 21131 8449 21143 8483
rect 21085 8443 21143 8449
rect 21266 8440 21272 8492
rect 21324 8440 21330 8492
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 21836 8489 21864 8588
rect 22554 8576 22560 8588
rect 22612 8576 22618 8628
rect 23934 8576 23940 8628
rect 23992 8576 23998 8628
rect 26786 8576 26792 8628
rect 26844 8576 26850 8628
rect 28442 8576 28448 8628
rect 28500 8616 28506 8628
rect 29381 8619 29439 8625
rect 29381 8616 29393 8619
rect 28500 8588 29393 8616
rect 28500 8576 28506 8588
rect 29381 8585 29393 8588
rect 29427 8585 29439 8619
rect 29381 8579 29439 8585
rect 32030 8576 32036 8628
rect 32088 8616 32094 8628
rect 32325 8619 32383 8625
rect 32325 8616 32337 8619
rect 32088 8588 32337 8616
rect 32088 8576 32094 8588
rect 32325 8585 32337 8588
rect 32371 8616 32383 8619
rect 32950 8616 32956 8628
rect 32371 8588 32628 8616
rect 32371 8585 32383 8588
rect 32325 8579 32383 8585
rect 27614 8548 27620 8560
rect 26804 8520 27620 8548
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21784 8452 21833 8480
rect 21784 8440 21790 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 22094 8440 22100 8492
rect 22152 8480 22158 8492
rect 22189 8483 22247 8489
rect 22189 8480 22201 8483
rect 22152 8452 22201 8480
rect 22152 8440 22158 8452
rect 22189 8449 22201 8452
rect 22235 8449 22247 8483
rect 22189 8443 22247 8449
rect 22557 8483 22615 8489
rect 22557 8449 22569 8483
rect 22603 8449 22615 8483
rect 22557 8443 22615 8449
rect 14277 8415 14335 8421
rect 14277 8412 14289 8415
rect 14240 8384 14289 8412
rect 14240 8372 14246 8384
rect 14277 8381 14289 8384
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 14369 8415 14427 8421
rect 14369 8381 14381 8415
rect 14415 8381 14427 8415
rect 14369 8375 14427 8381
rect 14550 8372 14556 8424
rect 14608 8372 14614 8424
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 22572 8412 22600 8443
rect 22830 8440 22836 8492
rect 22888 8480 22894 8492
rect 23845 8483 23903 8489
rect 23845 8480 23857 8483
rect 22888 8452 23857 8480
rect 22888 8440 22894 8452
rect 23845 8449 23857 8452
rect 23891 8480 23903 8483
rect 24397 8483 24455 8489
rect 24397 8480 24409 8483
rect 23891 8452 24409 8480
rect 23891 8449 23903 8452
rect 23845 8443 23903 8449
rect 24397 8449 24409 8452
rect 24443 8449 24455 8483
rect 24397 8443 24455 8449
rect 26510 8440 26516 8492
rect 26568 8440 26574 8492
rect 17828 8384 19840 8412
rect 17828 8372 17834 8384
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 12621 8347 12679 8353
rect 12621 8344 12633 8347
rect 12584 8316 12633 8344
rect 12584 8304 12590 8316
rect 12621 8313 12633 8316
rect 12667 8313 12679 8347
rect 12621 8307 12679 8313
rect 12713 8347 12771 8353
rect 12713 8313 12725 8347
rect 12759 8344 12771 8347
rect 13630 8344 13636 8356
rect 12759 8316 13636 8344
rect 12759 8313 12771 8316
rect 12713 8307 12771 8313
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 17221 8347 17279 8353
rect 17221 8313 17233 8347
rect 17267 8344 17279 8347
rect 19058 8344 19064 8356
rect 17267 8316 19064 8344
rect 17267 8313 17279 8316
rect 17221 8307 17279 8313
rect 19058 8304 19064 8316
rect 19116 8304 19122 8356
rect 19812 8344 19840 8384
rect 21100 8384 22600 8412
rect 21100 8356 21128 8384
rect 23566 8372 23572 8424
rect 23624 8412 23630 8424
rect 26804 8421 26832 8520
rect 27614 8508 27620 8520
rect 27672 8548 27678 8560
rect 27672 8520 28856 8548
rect 27672 8508 27678 8520
rect 27338 8440 27344 8492
rect 27396 8440 27402 8492
rect 27706 8440 27712 8492
rect 27764 8440 27770 8492
rect 27893 8483 27951 8489
rect 27893 8449 27905 8483
rect 27939 8449 27951 8483
rect 27893 8443 27951 8449
rect 24121 8415 24179 8421
rect 24121 8412 24133 8415
rect 23624 8384 24133 8412
rect 23624 8372 23630 8384
rect 24121 8381 24133 8384
rect 24167 8381 24179 8415
rect 24121 8375 24179 8381
rect 26789 8415 26847 8421
rect 26789 8381 26801 8415
rect 26835 8381 26847 8415
rect 27522 8412 27528 8424
rect 26789 8375 26847 8381
rect 27172 8384 27528 8412
rect 19812 8316 21036 8344
rect 1486 8236 1492 8288
rect 1544 8276 1550 8288
rect 7006 8276 7012 8288
rect 1544 8248 7012 8276
rect 1544 8236 1550 8248
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 7101 8279 7159 8285
rect 7101 8245 7113 8279
rect 7147 8276 7159 8279
rect 7650 8276 7656 8288
rect 7147 8248 7656 8276
rect 7147 8245 7159 8248
rect 7101 8239 7159 8245
rect 7650 8236 7656 8248
rect 7708 8236 7714 8288
rect 11882 8236 11888 8288
rect 11940 8276 11946 8288
rect 12345 8279 12403 8285
rect 12345 8276 12357 8279
rect 11940 8248 12357 8276
rect 11940 8236 11946 8248
rect 12345 8245 12357 8248
rect 12391 8245 12403 8279
rect 12345 8239 12403 8245
rect 13538 8236 13544 8288
rect 13596 8276 13602 8288
rect 20714 8276 20720 8288
rect 13596 8248 20720 8276
rect 13596 8236 13602 8248
rect 20714 8236 20720 8248
rect 20772 8236 20778 8288
rect 21008 8276 21036 8316
rect 21082 8304 21088 8356
rect 21140 8304 21146 8356
rect 21913 8347 21971 8353
rect 21913 8344 21925 8347
rect 21192 8316 21925 8344
rect 21192 8276 21220 8316
rect 21913 8313 21925 8316
rect 21959 8344 21971 8347
rect 24210 8344 24216 8356
rect 21959 8316 24216 8344
rect 21959 8313 21971 8316
rect 21913 8307 21971 8313
rect 24210 8304 24216 8316
rect 24268 8304 24274 8356
rect 26605 8347 26663 8353
rect 26605 8313 26617 8347
rect 26651 8344 26663 8347
rect 27172 8344 27200 8384
rect 27522 8372 27528 8384
rect 27580 8412 27586 8424
rect 27908 8412 27936 8443
rect 28350 8440 28356 8492
rect 28408 8440 28414 8492
rect 28828 8489 28856 8520
rect 29178 8508 29184 8560
rect 29236 8508 29242 8560
rect 32122 8508 32128 8560
rect 32180 8508 32186 8560
rect 32600 8557 32628 8588
rect 32784 8588 32956 8616
rect 32585 8551 32643 8557
rect 32585 8517 32597 8551
rect 32631 8517 32643 8551
rect 32585 8511 32643 8517
rect 28813 8483 28871 8489
rect 28813 8449 28825 8483
rect 28859 8449 28871 8483
rect 28813 8443 28871 8449
rect 31846 8440 31852 8492
rect 31904 8480 31910 8492
rect 32784 8489 32812 8588
rect 32950 8576 32956 8588
rect 33008 8616 33014 8628
rect 34149 8619 34207 8625
rect 34149 8616 34161 8619
rect 33008 8588 34161 8616
rect 33008 8576 33014 8588
rect 34149 8585 34161 8588
rect 34195 8616 34207 8619
rect 34330 8616 34336 8628
rect 34195 8588 34336 8616
rect 34195 8585 34207 8588
rect 34149 8579 34207 8585
rect 34330 8576 34336 8588
rect 34388 8576 34394 8628
rect 33042 8508 33048 8560
rect 33100 8548 33106 8560
rect 34057 8551 34115 8557
rect 34057 8548 34069 8551
rect 33100 8520 34069 8548
rect 33100 8508 33106 8520
rect 34057 8517 34069 8520
rect 34103 8517 34115 8551
rect 34057 8511 34115 8517
rect 34238 8508 34244 8560
rect 34296 8548 34302 8560
rect 34425 8551 34483 8557
rect 34425 8548 34437 8551
rect 34296 8520 34437 8548
rect 34296 8508 34302 8520
rect 34425 8517 34437 8520
rect 34471 8517 34483 8551
rect 34425 8511 34483 8517
rect 32769 8483 32827 8489
rect 32769 8480 32781 8483
rect 31904 8452 32781 8480
rect 31904 8440 31910 8452
rect 32769 8449 32781 8452
rect 32815 8449 32827 8483
rect 32769 8443 32827 8449
rect 32858 8440 32864 8492
rect 32916 8440 32922 8492
rect 27580 8384 27936 8412
rect 27580 8372 27586 8384
rect 32398 8372 32404 8424
rect 32456 8412 32462 8424
rect 32876 8412 32904 8440
rect 32456 8384 32904 8412
rect 32456 8372 32462 8384
rect 26651 8316 27200 8344
rect 26651 8313 26663 8316
rect 26605 8307 26663 8313
rect 27430 8304 27436 8356
rect 27488 8304 27494 8356
rect 31662 8304 31668 8356
rect 31720 8344 31726 8356
rect 32585 8347 32643 8353
rect 32585 8344 32597 8347
rect 31720 8316 32597 8344
rect 31720 8304 31726 8316
rect 32585 8313 32597 8316
rect 32631 8313 32643 8347
rect 32585 8307 32643 8313
rect 34606 8304 34612 8356
rect 34664 8304 34670 8356
rect 21008 8248 21220 8276
rect 26326 8236 26332 8288
rect 26384 8276 26390 8288
rect 27246 8276 27252 8288
rect 26384 8248 27252 8276
rect 26384 8236 26390 8248
rect 27246 8236 27252 8248
rect 27304 8276 27310 8288
rect 29178 8276 29184 8288
rect 27304 8248 29184 8276
rect 27304 8236 27310 8248
rect 29178 8236 29184 8248
rect 29236 8236 29242 8288
rect 29362 8236 29368 8288
rect 29420 8236 29426 8288
rect 29549 8279 29607 8285
rect 29549 8245 29561 8279
rect 29595 8276 29607 8279
rect 30006 8276 30012 8288
rect 29595 8248 30012 8276
rect 29595 8245 29607 8248
rect 29549 8239 29607 8245
rect 30006 8236 30012 8248
rect 30064 8236 30070 8288
rect 31938 8236 31944 8288
rect 31996 8276 32002 8288
rect 32309 8279 32367 8285
rect 32309 8276 32321 8279
rect 31996 8248 32321 8276
rect 31996 8236 32002 8248
rect 32309 8245 32321 8248
rect 32355 8276 32367 8279
rect 32398 8276 32404 8288
rect 32355 8248 32404 8276
rect 32355 8245 32367 8248
rect 32309 8239 32367 8245
rect 32398 8236 32404 8248
rect 32456 8236 32462 8288
rect 32490 8236 32496 8288
rect 32548 8236 32554 8288
rect 1104 8186 36800 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 36800 8186
rect 1104 8112 36800 8134
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 6181 8075 6239 8081
rect 5408 8044 5948 8072
rect 5408 8032 5414 8044
rect 5442 8004 5448 8016
rect 4908 7976 5448 8004
rect 4709 7939 4767 7945
rect 4709 7936 4721 7939
rect 4448 7908 4721 7936
rect 4448 7877 4476 7908
rect 4709 7905 4721 7908
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 4908 7877 4936 7976
rect 5442 7964 5448 7976
rect 5500 7964 5506 8016
rect 5092 7908 5396 7936
rect 5092 7877 5120 7908
rect 5368 7880 5396 7908
rect 5920 7880 5948 8044
rect 6181 8041 6193 8075
rect 6227 8072 6239 8075
rect 6362 8072 6368 8084
rect 6227 8044 6368 8072
rect 6227 8041 6239 8044
rect 6181 8035 6239 8041
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 7006 8032 7012 8084
rect 7064 8072 7070 8084
rect 10505 8075 10563 8081
rect 7064 8044 8156 8072
rect 7064 8032 7070 8044
rect 8021 8007 8079 8013
rect 7392 7976 7880 8004
rect 7101 7939 7159 7945
rect 7101 7936 7113 7939
rect 6380 7908 7113 7936
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5258 7868 5264 7880
rect 5215 7840 5264 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 4632 7800 4660 7831
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5408 7840 5549 7868
rect 5408 7828 5414 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 5902 7828 5908 7880
rect 5960 7828 5966 7880
rect 6380 7877 6408 7908
rect 7101 7905 7113 7908
rect 7147 7936 7159 7939
rect 7282 7936 7288 7948
rect 7147 7908 7288 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 6365 7871 6423 7877
rect 6365 7868 6377 7871
rect 6135 7840 6377 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 6365 7837 6377 7840
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7868 6699 7871
rect 6730 7868 6736 7880
rect 6687 7840 6736 7868
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 4632 7772 5396 7800
rect 4614 7692 4620 7744
rect 4672 7692 4678 7744
rect 5368 7741 5396 7772
rect 5442 7760 5448 7812
rect 5500 7760 5506 7812
rect 6840 7800 6868 7831
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 7190 7868 7196 7880
rect 6972 7840 7196 7868
rect 6972 7828 6978 7840
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7392 7800 7420 7976
rect 7852 7948 7880 7976
rect 8021 7973 8033 8007
rect 8067 7973 8079 8007
rect 8128 8004 8156 8044
rect 10505 8041 10517 8075
rect 10551 8072 10563 8075
rect 10965 8075 11023 8081
rect 10965 8072 10977 8075
rect 10551 8044 10977 8072
rect 10551 8041 10563 8044
rect 10505 8035 10563 8041
rect 10965 8041 10977 8044
rect 11011 8041 11023 8075
rect 10965 8035 11023 8041
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 11422 8072 11428 8084
rect 11379 8044 11428 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 12158 8032 12164 8084
rect 12216 8072 12222 8084
rect 13814 8072 13820 8084
rect 12216 8044 13820 8072
rect 12216 8032 12222 8044
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 15102 8032 15108 8084
rect 15160 8032 15166 8084
rect 17218 8032 17224 8084
rect 17276 8072 17282 8084
rect 17865 8075 17923 8081
rect 17865 8072 17877 8075
rect 17276 8044 17877 8072
rect 17276 8032 17282 8044
rect 17865 8041 17877 8044
rect 17911 8041 17923 8075
rect 17865 8035 17923 8041
rect 18874 8032 18880 8084
rect 18932 8032 18938 8084
rect 19061 8075 19119 8081
rect 19061 8041 19073 8075
rect 19107 8072 19119 8075
rect 25869 8075 25927 8081
rect 19107 8044 21128 8072
rect 19107 8041 19119 8044
rect 19061 8035 19119 8041
rect 17126 8004 17132 8016
rect 8128 7976 17132 8004
rect 8021 7967 8079 7973
rect 7466 7896 7472 7948
rect 7524 7936 7530 7948
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 7524 7908 7573 7936
rect 7524 7896 7530 7908
rect 7561 7905 7573 7908
rect 7607 7936 7619 7939
rect 7607 7908 7788 7936
rect 7607 7905 7619 7908
rect 7561 7899 7619 7905
rect 7650 7828 7656 7880
rect 7708 7828 7714 7880
rect 7760 7877 7788 7908
rect 7834 7896 7840 7948
rect 7892 7896 7898 7948
rect 8036 7936 8064 7967
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 8205 7939 8263 7945
rect 8036 7908 8156 7936
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 8128 7877 8156 7908
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 8251 7908 12112 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7984 7840 8033 7868
rect 7984 7828 7990 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 7469 7803 7527 7809
rect 7469 7800 7481 7803
rect 6840 7772 7481 7800
rect 7469 7769 7481 7772
rect 7515 7769 7527 7803
rect 8312 7800 8340 7831
rect 8386 7828 8392 7880
rect 8444 7828 8450 7880
rect 8570 7828 8576 7880
rect 8628 7828 8634 7880
rect 9858 7828 9864 7880
rect 9916 7828 9922 7880
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7868 10103 7871
rect 10318 7868 10324 7880
rect 10091 7840 10324 7868
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10778 7828 10784 7880
rect 10836 7868 10842 7880
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 10836 7840 10885 7868
rect 10836 7828 10842 7840
rect 10873 7837 10885 7840
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 7469 7763 7527 7769
rect 7668 7772 8340 7800
rect 5353 7735 5411 7741
rect 5353 7701 5365 7735
rect 5399 7701 5411 7735
rect 5353 7695 5411 7701
rect 6917 7735 6975 7741
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7668 7732 7696 7772
rect 6963 7704 7696 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7834 7692 7840 7744
rect 7892 7732 7898 7744
rect 8481 7735 8539 7741
rect 8481 7732 8493 7735
rect 7892 7704 8493 7732
rect 7892 7692 7898 7704
rect 8481 7701 8493 7704
rect 8527 7701 8539 7735
rect 10888 7732 10916 7831
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 12084 7877 12112 7908
rect 12158 7896 12164 7948
rect 12216 7896 12222 7948
rect 13538 7936 13544 7948
rect 12268 7908 13544 7936
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 11977 7803 12035 7809
rect 11977 7769 11989 7803
rect 12023 7800 12035 7803
rect 12268 7800 12296 7908
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 13630 7896 13636 7948
rect 13688 7936 13694 7948
rect 17497 7939 17555 7945
rect 13688 7908 14136 7936
rect 13688 7896 13694 7908
rect 13722 7828 13728 7880
rect 13780 7828 13786 7880
rect 14108 7877 14136 7908
rect 17497 7905 17509 7939
rect 17543 7936 17555 7939
rect 18230 7936 18236 7948
rect 17543 7908 18236 7936
rect 17543 7905 17555 7908
rect 17497 7899 17555 7905
rect 18230 7896 18236 7908
rect 18288 7936 18294 7948
rect 18892 7936 18920 8032
rect 18288 7908 18920 7936
rect 18288 7896 18294 7908
rect 19058 7896 19064 7948
rect 19116 7936 19122 7948
rect 21100 7945 21128 8044
rect 25869 8041 25881 8075
rect 25915 8072 25927 8075
rect 26326 8072 26332 8084
rect 25915 8044 26332 8072
rect 25915 8041 25927 8044
rect 25869 8035 25927 8041
rect 26326 8032 26332 8044
rect 26384 8032 26390 8084
rect 26510 8032 26516 8084
rect 26568 8072 26574 8084
rect 26605 8075 26663 8081
rect 26605 8072 26617 8075
rect 26568 8044 26617 8072
rect 26568 8032 26574 8044
rect 26605 8041 26617 8044
rect 26651 8072 26663 8075
rect 27617 8075 27675 8081
rect 27617 8072 27629 8075
rect 26651 8044 27629 8072
rect 26651 8041 26663 8044
rect 26605 8035 26663 8041
rect 27617 8041 27629 8044
rect 27663 8072 27675 8075
rect 28350 8072 28356 8084
rect 27663 8044 28356 8072
rect 27663 8041 27675 8044
rect 27617 8035 27675 8041
rect 28350 8032 28356 8044
rect 28408 8032 28414 8084
rect 30193 8075 30251 8081
rect 30193 8041 30205 8075
rect 30239 8072 30251 8075
rect 30558 8072 30564 8084
rect 30239 8044 30564 8072
rect 30239 8041 30251 8044
rect 30193 8035 30251 8041
rect 30558 8032 30564 8044
rect 30616 8072 30622 8084
rect 31754 8072 31760 8084
rect 30616 8044 31760 8072
rect 30616 8032 30622 8044
rect 31754 8032 31760 8044
rect 31812 8072 31818 8084
rect 33505 8075 33563 8081
rect 33505 8072 33517 8075
rect 31812 8044 33517 8072
rect 31812 8032 31818 8044
rect 33505 8041 33517 8044
rect 33551 8041 33563 8075
rect 33505 8035 33563 8041
rect 21453 8007 21511 8013
rect 21453 7973 21465 8007
rect 21499 8004 21511 8007
rect 21910 8004 21916 8016
rect 21499 7976 21916 8004
rect 21499 7973 21511 7976
rect 21453 7967 21511 7973
rect 21910 7964 21916 7976
rect 21968 7964 21974 8016
rect 26421 8007 26479 8013
rect 26421 7973 26433 8007
rect 26467 8004 26479 8007
rect 27341 8007 27399 8013
rect 26467 7976 26648 8004
rect 26467 7973 26479 7976
rect 26421 7967 26479 7973
rect 26620 7948 26648 7976
rect 27341 7973 27353 8007
rect 27387 8004 27399 8007
rect 27706 8004 27712 8016
rect 27387 7976 27712 8004
rect 27387 7973 27399 7976
rect 27341 7967 27399 7973
rect 27706 7964 27712 7976
rect 27764 8004 27770 8016
rect 28077 8007 28135 8013
rect 28077 8004 28089 8007
rect 27764 7976 28089 8004
rect 27764 7964 27770 7976
rect 28077 7973 28089 7976
rect 28123 7973 28135 8007
rect 30837 8007 30895 8013
rect 30837 8004 30849 8007
rect 28077 7967 28135 7973
rect 29932 7976 30849 8004
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 19116 7908 19380 7936
rect 19116 7896 19122 7908
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7868 14151 7871
rect 14274 7868 14280 7880
rect 14139 7840 14280 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7868 14427 7871
rect 14458 7868 14464 7880
rect 14415 7840 14464 7868
rect 14415 7837 14427 7840
rect 14369 7831 14427 7837
rect 12023 7772 12296 7800
rect 12023 7769 12035 7772
rect 11977 7763 12035 7769
rect 13170 7760 13176 7812
rect 13228 7800 13234 7812
rect 14384 7800 14412 7831
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 15286 7828 15292 7880
rect 15344 7828 15350 7880
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7868 17279 7871
rect 18414 7868 18420 7880
rect 17267 7840 18420 7868
rect 17267 7837 17279 7840
rect 17221 7831 17279 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7837 18567 7871
rect 18509 7831 18567 7837
rect 13228 7772 14412 7800
rect 17706 7803 17764 7809
rect 13228 7760 13234 7772
rect 17706 7769 17718 7803
rect 17752 7800 17764 7803
rect 18524 7800 18552 7831
rect 18598 7828 18604 7880
rect 18656 7868 18662 7880
rect 18877 7871 18935 7877
rect 18877 7868 18889 7871
rect 18656 7840 18889 7868
rect 18656 7828 18662 7840
rect 18877 7837 18889 7840
rect 18923 7837 18935 7871
rect 18877 7831 18935 7837
rect 19242 7828 19248 7880
rect 19300 7828 19306 7880
rect 19352 7868 19380 7908
rect 20732 7908 20913 7936
rect 20732 7868 20760 7908
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 20901 7899 20959 7905
rect 21085 7939 21143 7945
rect 21085 7905 21097 7939
rect 21131 7936 21143 7939
rect 21266 7936 21272 7948
rect 21131 7908 21272 7936
rect 21131 7905 21143 7908
rect 21085 7899 21143 7905
rect 19352 7840 20760 7868
rect 20806 7828 20812 7880
rect 20864 7828 20870 7880
rect 20916 7868 20944 7899
rect 21266 7896 21272 7908
rect 21324 7896 21330 7948
rect 26602 7896 26608 7948
rect 26660 7896 26666 7948
rect 27614 7896 27620 7948
rect 27672 7896 27678 7948
rect 27890 7896 27896 7948
rect 27948 7936 27954 7948
rect 27948 7908 28580 7936
rect 27948 7896 27954 7908
rect 20916 7840 21312 7868
rect 18690 7800 18696 7812
rect 17752 7772 18696 7800
rect 17752 7769 17764 7772
rect 17706 7763 17764 7769
rect 18690 7760 18696 7772
rect 18748 7760 18754 7812
rect 19512 7803 19570 7809
rect 19512 7769 19524 7803
rect 19558 7800 19570 7803
rect 21082 7800 21088 7812
rect 19558 7772 21088 7800
rect 19558 7769 19570 7772
rect 19512 7763 19570 7769
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 21284 7800 21312 7840
rect 21358 7828 21364 7880
rect 21416 7868 21422 7880
rect 21453 7871 21511 7877
rect 21453 7868 21465 7871
rect 21416 7840 21465 7868
rect 21416 7828 21422 7840
rect 21453 7837 21465 7840
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 21634 7828 21640 7880
rect 21692 7828 21698 7880
rect 21818 7828 21824 7880
rect 21876 7828 21882 7880
rect 22738 7828 22744 7880
rect 22796 7828 22802 7880
rect 22830 7828 22836 7880
rect 22888 7828 22894 7880
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7837 23167 7871
rect 23109 7831 23167 7837
rect 22370 7800 22376 7812
rect 21284 7772 22376 7800
rect 12391 7735 12449 7741
rect 12391 7732 12403 7735
rect 10888 7704 12403 7732
rect 8481 7695 8539 7701
rect 12391 7701 12403 7704
rect 12437 7732 12449 7735
rect 12526 7732 12532 7744
rect 12437 7704 12532 7732
rect 12437 7701 12449 7704
rect 12391 7695 12449 7701
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 17586 7692 17592 7744
rect 17644 7692 17650 7744
rect 18414 7692 18420 7744
rect 18472 7732 18478 7744
rect 20625 7735 20683 7741
rect 20625 7732 20637 7735
rect 18472 7704 20637 7732
rect 18472 7692 18478 7704
rect 20625 7701 20637 7704
rect 20671 7701 20683 7735
rect 21284 7732 21312 7772
rect 22370 7760 22376 7772
rect 22428 7760 22434 7812
rect 23124 7800 23152 7831
rect 23474 7828 23480 7880
rect 23532 7868 23538 7880
rect 23937 7871 23995 7877
rect 23937 7868 23949 7871
rect 23532 7840 23949 7868
rect 23532 7828 23538 7840
rect 23937 7837 23949 7840
rect 23983 7837 23995 7871
rect 23937 7831 23995 7837
rect 24489 7871 24547 7877
rect 24489 7837 24501 7871
rect 24535 7868 24547 7871
rect 25038 7868 25044 7880
rect 24535 7840 25044 7868
rect 24535 7837 24547 7840
rect 24489 7831 24547 7837
rect 25038 7828 25044 7840
rect 25096 7828 25102 7880
rect 26786 7828 26792 7880
rect 26844 7868 26850 7880
rect 27249 7871 27307 7877
rect 27249 7868 27261 7871
rect 26844 7840 27261 7868
rect 26844 7828 26850 7840
rect 27249 7837 27261 7840
rect 27295 7837 27307 7871
rect 27249 7831 27307 7837
rect 27433 7871 27491 7877
rect 27433 7837 27445 7871
rect 27479 7837 27491 7871
rect 27433 7831 27491 7837
rect 22572 7772 23152 7800
rect 21450 7732 21456 7744
rect 21284 7704 21456 7732
rect 20625 7695 20683 7701
rect 21450 7692 21456 7704
rect 21508 7692 21514 7744
rect 21729 7735 21787 7741
rect 21729 7701 21741 7735
rect 21775 7732 21787 7735
rect 22186 7732 22192 7744
rect 21775 7704 22192 7732
rect 21775 7701 21787 7704
rect 21729 7695 21787 7701
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 22572 7741 22600 7772
rect 24118 7760 24124 7812
rect 24176 7800 24182 7812
rect 24734 7803 24792 7809
rect 24734 7800 24746 7803
rect 24176 7772 24746 7800
rect 24176 7760 24182 7772
rect 24734 7769 24746 7772
rect 24780 7769 24792 7803
rect 24734 7763 24792 7769
rect 25958 7760 25964 7812
rect 26016 7800 26022 7812
rect 26145 7803 26203 7809
rect 26145 7800 26157 7803
rect 26016 7772 26157 7800
rect 26016 7760 26022 7772
rect 26145 7769 26157 7772
rect 26191 7769 26203 7803
rect 27448 7800 27476 7831
rect 27522 7828 27528 7880
rect 27580 7828 27586 7880
rect 28552 7877 28580 7908
rect 29932 7877 29960 7976
rect 30837 7973 30849 7976
rect 30883 7973 30895 8007
rect 32769 8007 32827 8013
rect 32769 8004 32781 8007
rect 30837 7967 30895 7973
rect 30944 7976 32781 8004
rect 30190 7896 30196 7948
rect 30248 7936 30254 7948
rect 30377 7939 30435 7945
rect 30377 7936 30389 7939
rect 30248 7908 30389 7936
rect 30248 7896 30254 7908
rect 30377 7905 30389 7908
rect 30423 7905 30435 7939
rect 30377 7899 30435 7905
rect 30466 7896 30472 7948
rect 30524 7936 30530 7948
rect 30561 7939 30619 7945
rect 30561 7936 30573 7939
rect 30524 7908 30573 7936
rect 30524 7896 30530 7908
rect 30561 7905 30573 7908
rect 30607 7905 30619 7939
rect 30561 7899 30619 7905
rect 30653 7939 30711 7945
rect 30653 7905 30665 7939
rect 30699 7936 30711 7939
rect 30944 7936 30972 7976
rect 32769 7973 32781 7976
rect 32815 7973 32827 8007
rect 32769 7967 32827 7973
rect 32950 7964 32956 8016
rect 33008 8004 33014 8016
rect 33594 8004 33600 8016
rect 33008 7976 33600 8004
rect 33008 7964 33014 7976
rect 33594 7964 33600 7976
rect 33652 8004 33658 8016
rect 34054 8004 34060 8016
rect 33652 7976 34060 8004
rect 33652 7964 33658 7976
rect 34054 7964 34060 7976
rect 34112 7964 34118 8016
rect 30699 7908 30972 7936
rect 31021 7939 31079 7945
rect 30699 7905 30711 7908
rect 30653 7899 30711 7905
rect 28353 7871 28411 7877
rect 28353 7837 28365 7871
rect 28399 7837 28411 7871
rect 28353 7831 28411 7837
rect 28537 7871 28595 7877
rect 28537 7837 28549 7871
rect 28583 7837 28595 7871
rect 29917 7871 29975 7877
rect 28537 7831 28595 7837
rect 28644 7840 29592 7868
rect 28368 7800 28396 7831
rect 28644 7800 28672 7840
rect 27448 7772 27936 7800
rect 28368 7772 28672 7800
rect 26145 7763 26203 7769
rect 27908 7741 27936 7772
rect 29178 7760 29184 7812
rect 29236 7760 29242 7812
rect 29564 7800 29592 7840
rect 29917 7837 29929 7871
rect 29963 7837 29975 7871
rect 29917 7831 29975 7837
rect 30006 7828 30012 7880
rect 30064 7828 30070 7880
rect 30208 7800 30236 7896
rect 30852 7880 30880 7908
rect 31021 7905 31033 7939
rect 31067 7936 31079 7939
rect 31481 7939 31539 7945
rect 31481 7936 31493 7939
rect 31067 7908 31493 7936
rect 31067 7905 31079 7908
rect 31021 7899 31079 7905
rect 31481 7905 31493 7908
rect 31527 7905 31539 7939
rect 33137 7939 33195 7945
rect 31481 7899 31539 7905
rect 31588 7908 33088 7936
rect 31588 7880 31616 7908
rect 30285 7871 30343 7877
rect 30285 7837 30297 7871
rect 30331 7868 30343 7871
rect 30331 7840 30696 7868
rect 30331 7837 30343 7840
rect 30285 7831 30343 7837
rect 30466 7809 30472 7812
rect 29564 7772 30236 7800
rect 30447 7803 30472 7809
rect 30447 7769 30459 7803
rect 30447 7763 30472 7769
rect 30466 7760 30472 7763
rect 30524 7760 30530 7812
rect 30668 7800 30696 7840
rect 30742 7828 30748 7880
rect 30800 7828 30806 7880
rect 30834 7828 30840 7880
rect 30892 7828 30898 7880
rect 31110 7828 31116 7880
rect 31168 7828 31174 7880
rect 31202 7828 31208 7880
rect 31260 7828 31266 7880
rect 31297 7871 31355 7877
rect 31297 7837 31309 7871
rect 31343 7868 31355 7871
rect 31570 7868 31576 7880
rect 31343 7840 31576 7868
rect 31343 7837 31355 7840
rect 31297 7831 31355 7837
rect 31570 7828 31576 7840
rect 31628 7828 31634 7880
rect 31665 7871 31723 7877
rect 31665 7837 31677 7871
rect 31711 7837 31723 7871
rect 31665 7831 31723 7837
rect 31757 7871 31815 7877
rect 31757 7837 31769 7871
rect 31803 7868 31815 7871
rect 31846 7868 31852 7880
rect 31803 7840 31852 7868
rect 31803 7837 31815 7840
rect 31757 7831 31815 7837
rect 31386 7800 31392 7812
rect 30668 7772 31392 7800
rect 31386 7760 31392 7772
rect 31444 7800 31450 7812
rect 31680 7800 31708 7831
rect 31846 7828 31852 7840
rect 31904 7828 31910 7880
rect 32030 7828 32036 7880
rect 32088 7828 32094 7880
rect 32125 7871 32183 7877
rect 32125 7837 32137 7871
rect 32171 7868 32183 7871
rect 32585 7871 32643 7877
rect 32585 7868 32597 7871
rect 32171 7840 32597 7868
rect 32171 7837 32183 7840
rect 32125 7831 32183 7837
rect 32585 7837 32597 7840
rect 32631 7837 32643 7871
rect 32585 7831 32643 7837
rect 32140 7800 32168 7831
rect 31444 7772 31708 7800
rect 31864 7772 32168 7800
rect 31444 7760 31450 7772
rect 22557 7735 22615 7741
rect 22557 7701 22569 7735
rect 22603 7701 22615 7735
rect 22557 7695 22615 7701
rect 27893 7735 27951 7741
rect 27893 7701 27905 7735
rect 27939 7732 27951 7735
rect 28166 7732 28172 7744
rect 27939 7704 28172 7732
rect 27939 7701 27951 7704
rect 27893 7695 27951 7701
rect 28166 7692 28172 7704
rect 28224 7692 28230 7744
rect 28261 7735 28319 7741
rect 28261 7701 28273 7735
rect 28307 7732 28319 7735
rect 28442 7732 28448 7744
rect 28307 7704 28448 7732
rect 28307 7701 28319 7704
rect 28261 7695 28319 7701
rect 28442 7692 28448 7704
rect 28500 7692 28506 7744
rect 29086 7692 29092 7744
rect 29144 7732 29150 7744
rect 29273 7735 29331 7741
rect 29273 7732 29285 7735
rect 29144 7704 29285 7732
rect 29144 7692 29150 7704
rect 29273 7701 29285 7704
rect 29319 7701 29331 7735
rect 29273 7695 29331 7701
rect 29730 7692 29736 7744
rect 29788 7692 29794 7744
rect 31478 7692 31484 7744
rect 31536 7732 31542 7744
rect 31864 7732 31892 7772
rect 32214 7760 32220 7812
rect 32272 7760 32278 7812
rect 32493 7803 32551 7809
rect 32493 7800 32505 7803
rect 32324 7772 32505 7800
rect 31536 7704 31892 7732
rect 31536 7692 31542 7704
rect 31938 7692 31944 7744
rect 31996 7692 32002 7744
rect 32030 7692 32036 7744
rect 32088 7732 32094 7744
rect 32324 7732 32352 7772
rect 32493 7769 32505 7772
rect 32539 7800 32551 7803
rect 32674 7800 32680 7812
rect 32539 7772 32680 7800
rect 32539 7769 32551 7772
rect 32493 7763 32551 7769
rect 32674 7760 32680 7772
rect 32732 7760 32738 7812
rect 32950 7800 32956 7812
rect 32784 7772 32956 7800
rect 32088 7704 32352 7732
rect 32401 7735 32459 7741
rect 32088 7692 32094 7704
rect 32401 7701 32413 7735
rect 32447 7732 32459 7735
rect 32784 7732 32812 7772
rect 32950 7760 32956 7772
rect 33008 7760 33014 7812
rect 33060 7800 33088 7908
rect 33137 7905 33149 7939
rect 33183 7936 33195 7939
rect 33183 7908 34836 7936
rect 33183 7905 33195 7908
rect 33137 7899 33195 7905
rect 33318 7828 33324 7880
rect 33376 7828 33382 7880
rect 33597 7871 33655 7877
rect 33597 7837 33609 7871
rect 33643 7868 33655 7871
rect 34514 7868 34520 7880
rect 33643 7840 34520 7868
rect 33643 7837 33655 7840
rect 33597 7831 33655 7837
rect 34514 7828 34520 7840
rect 34572 7828 34578 7880
rect 34698 7828 34704 7880
rect 34756 7828 34762 7880
rect 34808 7868 34836 7908
rect 34957 7871 35015 7877
rect 34957 7868 34969 7871
rect 34808 7840 34969 7868
rect 34957 7837 34969 7840
rect 35003 7837 35015 7871
rect 34957 7831 35015 7837
rect 36446 7828 36452 7880
rect 36504 7828 36510 7880
rect 33686 7800 33692 7812
rect 33060 7772 33692 7800
rect 33686 7760 33692 7772
rect 33744 7760 33750 7812
rect 33781 7803 33839 7809
rect 33781 7769 33793 7803
rect 33827 7800 33839 7803
rect 34054 7800 34060 7812
rect 33827 7772 34060 7800
rect 33827 7769 33839 7772
rect 33781 7763 33839 7769
rect 34054 7760 34060 7772
rect 34112 7800 34118 7812
rect 34112 7772 36124 7800
rect 34112 7760 34118 7772
rect 32447 7704 32812 7732
rect 32447 7701 32459 7704
rect 32401 7695 32459 7701
rect 32858 7692 32864 7744
rect 32916 7732 32922 7744
rect 33873 7735 33931 7741
rect 33873 7732 33885 7735
rect 32916 7704 33885 7732
rect 32916 7692 32922 7704
rect 33873 7701 33885 7704
rect 33919 7732 33931 7735
rect 34514 7732 34520 7744
rect 33919 7704 34520 7732
rect 33919 7701 33931 7704
rect 33873 7695 33931 7701
rect 34514 7692 34520 7704
rect 34572 7692 34578 7744
rect 36096 7741 36124 7772
rect 36081 7735 36139 7741
rect 36081 7701 36093 7735
rect 36127 7701 36139 7735
rect 36081 7695 36139 7701
rect 36262 7692 36268 7744
rect 36320 7692 36326 7744
rect 1104 7642 36800 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 36800 7642
rect 1104 7568 36800 7590
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 7193 7531 7251 7537
rect 7193 7528 7205 7531
rect 7156 7500 7205 7528
rect 7156 7488 7162 7500
rect 7193 7497 7205 7500
rect 7239 7497 7251 7531
rect 7193 7491 7251 7497
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7616 7500 7849 7528
rect 7616 7488 7622 7500
rect 7837 7497 7849 7500
rect 7883 7497 7895 7531
rect 7837 7491 7895 7497
rect 9950 7488 9956 7540
rect 10008 7528 10014 7540
rect 10045 7531 10103 7537
rect 10045 7528 10057 7531
rect 10008 7500 10057 7528
rect 10008 7488 10014 7500
rect 10045 7497 10057 7500
rect 10091 7497 10103 7531
rect 10045 7491 10103 7497
rect 10318 7488 10324 7540
rect 10376 7488 10382 7540
rect 11790 7488 11796 7540
rect 11848 7488 11854 7540
rect 12802 7488 12808 7540
rect 12860 7528 12866 7540
rect 13725 7531 13783 7537
rect 13725 7528 13737 7531
rect 12860 7500 13737 7528
rect 12860 7488 12866 7500
rect 13725 7497 13737 7500
rect 13771 7497 13783 7531
rect 13725 7491 13783 7497
rect 19978 7488 19984 7540
rect 20036 7488 20042 7540
rect 20990 7488 20996 7540
rect 21048 7488 21054 7540
rect 21266 7488 21272 7540
rect 21324 7528 21330 7540
rect 21324 7500 22324 7528
rect 21324 7488 21330 7500
rect 5997 7463 6055 7469
rect 5997 7429 6009 7463
rect 6043 7460 6055 7463
rect 7469 7463 7527 7469
rect 6043 7432 7144 7460
rect 6043 7429 6055 7432
rect 5997 7423 6055 7429
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 5902 7392 5908 7404
rect 5500 7364 5908 7392
rect 5500 7352 5506 7364
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 7116 7401 7144 7432
rect 7469 7429 7481 7463
rect 7515 7460 7527 7463
rect 7515 7432 7972 7460
rect 7515 7429 7527 7432
rect 7469 7423 7527 7429
rect 6089 7395 6147 7401
rect 6089 7361 6101 7395
rect 6135 7361 6147 7395
rect 6089 7355 6147 7361
rect 7101 7395 7159 7401
rect 7101 7361 7113 7395
rect 7147 7392 7159 7395
rect 7190 7392 7196 7404
rect 7147 7364 7196 7392
rect 7147 7361 7159 7364
rect 7101 7355 7159 7361
rect 5810 7284 5816 7336
rect 5868 7324 5874 7336
rect 6104 7324 6132 7355
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7558 7392 7564 7404
rect 7423 7364 7564 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 7558 7352 7564 7364
rect 7616 7392 7622 7404
rect 7944 7401 7972 7432
rect 16574 7420 16580 7472
rect 16632 7460 16638 7472
rect 16936 7463 16994 7469
rect 16936 7460 16948 7463
rect 16632 7432 16948 7460
rect 16632 7420 16638 7432
rect 16936 7429 16948 7432
rect 16982 7460 16994 7463
rect 19996 7460 20024 7488
rect 16982 7432 20024 7460
rect 16982 7429 16994 7432
rect 16936 7423 16994 7429
rect 20438 7420 20444 7472
rect 20496 7460 20502 7472
rect 21913 7463 21971 7469
rect 20496 7432 21588 7460
rect 20496 7420 20502 7432
rect 7745 7395 7803 7401
rect 7745 7392 7757 7395
rect 7616 7364 7757 7392
rect 7616 7352 7622 7364
rect 7745 7361 7757 7364
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 8110 7392 8116 7404
rect 7975 7364 8116 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 10226 7352 10232 7404
rect 10284 7352 10290 7404
rect 10502 7352 10508 7404
rect 10560 7352 10566 7404
rect 11974 7352 11980 7404
rect 12032 7352 12038 7404
rect 12345 7395 12403 7401
rect 12345 7361 12357 7395
rect 12391 7392 12403 7395
rect 12526 7392 12532 7404
rect 12391 7364 12532 7392
rect 12391 7361 12403 7364
rect 12345 7355 12403 7361
rect 12526 7352 12532 7364
rect 12584 7352 12590 7404
rect 12621 7395 12679 7401
rect 12621 7361 12633 7395
rect 12667 7392 12679 7395
rect 12710 7392 12716 7404
rect 12667 7364 12716 7392
rect 12667 7361 12679 7364
rect 12621 7355 12679 7361
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7392 13323 7395
rect 13814 7392 13820 7404
rect 13311 7364 13820 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 14369 7395 14427 7401
rect 14369 7392 14381 7395
rect 14332 7364 14381 7392
rect 14332 7352 14338 7364
rect 14369 7361 14381 7364
rect 14415 7361 14427 7395
rect 17310 7392 17316 7404
rect 14369 7355 14427 7361
rect 16684 7364 17316 7392
rect 5868 7296 6132 7324
rect 5868 7284 5874 7296
rect 7282 7284 7288 7336
rect 7340 7284 7346 7336
rect 14093 7327 14151 7333
rect 14093 7293 14105 7327
rect 14139 7324 14151 7327
rect 14182 7324 14188 7336
rect 14139 7296 14188 7324
rect 14139 7293 14151 7296
rect 14093 7287 14151 7293
rect 14182 7284 14188 7296
rect 14240 7284 14246 7336
rect 16574 7284 16580 7336
rect 16632 7324 16638 7336
rect 16684 7333 16712 7364
rect 17310 7352 17316 7364
rect 17368 7352 17374 7404
rect 19886 7352 19892 7404
rect 19944 7352 19950 7404
rect 20070 7352 20076 7404
rect 20128 7392 20134 7404
rect 20530 7392 20536 7404
rect 20128 7364 20536 7392
rect 20128 7352 20134 7364
rect 20530 7352 20536 7364
rect 20588 7352 20594 7404
rect 21177 7395 21235 7401
rect 21177 7361 21189 7395
rect 21223 7361 21235 7395
rect 21177 7355 21235 7361
rect 16669 7327 16727 7333
rect 16669 7324 16681 7327
rect 16632 7296 16681 7324
rect 16632 7284 16638 7296
rect 16669 7293 16681 7296
rect 16715 7293 16727 7327
rect 21192 7324 21220 7355
rect 21266 7352 21272 7404
rect 21324 7392 21330 7404
rect 21361 7395 21419 7401
rect 21361 7392 21373 7395
rect 21324 7364 21373 7392
rect 21324 7352 21330 7364
rect 21361 7361 21373 7364
rect 21407 7361 21419 7395
rect 21361 7355 21419 7361
rect 21450 7352 21456 7404
rect 21508 7352 21514 7404
rect 21560 7392 21588 7432
rect 21913 7429 21925 7463
rect 21959 7460 21971 7463
rect 22002 7460 22008 7472
rect 21959 7432 22008 7460
rect 21959 7429 21971 7432
rect 21913 7423 21971 7429
rect 22002 7420 22008 7432
rect 22060 7420 22066 7472
rect 21637 7395 21695 7401
rect 21637 7392 21649 7395
rect 21560 7364 21649 7392
rect 21637 7361 21649 7364
rect 21683 7361 21695 7395
rect 21637 7355 21695 7361
rect 22094 7352 22100 7404
rect 22152 7352 22158 7404
rect 22186 7352 22192 7404
rect 22244 7352 22250 7404
rect 22296 7401 22324 7500
rect 22738 7488 22744 7540
rect 22796 7528 22802 7540
rect 23109 7531 23167 7537
rect 23109 7528 23121 7531
rect 22796 7500 23121 7528
rect 22796 7488 22802 7500
rect 23109 7497 23121 7500
rect 23155 7497 23167 7531
rect 23109 7491 23167 7497
rect 23474 7488 23480 7540
rect 23532 7488 23538 7540
rect 24118 7488 24124 7540
rect 24176 7488 24182 7540
rect 27433 7531 27491 7537
rect 27433 7497 27445 7531
rect 27479 7528 27491 7531
rect 27522 7528 27528 7540
rect 27479 7500 27528 7528
rect 27479 7497 27491 7500
rect 27433 7491 27491 7497
rect 27522 7488 27528 7500
rect 27580 7488 27586 7540
rect 29917 7531 29975 7537
rect 29917 7497 29929 7531
rect 29963 7528 29975 7531
rect 30466 7528 30472 7540
rect 29963 7500 30472 7528
rect 29963 7497 29975 7500
rect 29917 7491 29975 7497
rect 30466 7488 30472 7500
rect 30524 7488 30530 7540
rect 30742 7488 30748 7540
rect 30800 7488 30806 7540
rect 33318 7488 33324 7540
rect 33376 7528 33382 7540
rect 33505 7531 33563 7537
rect 33505 7528 33517 7531
rect 33376 7500 33517 7528
rect 33376 7488 33382 7500
rect 33505 7497 33517 7500
rect 33551 7497 33563 7531
rect 33505 7491 33563 7497
rect 33686 7488 33692 7540
rect 33744 7528 33750 7540
rect 34606 7528 34612 7540
rect 33744 7500 34612 7528
rect 33744 7488 33750 7500
rect 23569 7463 23627 7469
rect 23569 7429 23581 7463
rect 23615 7460 23627 7463
rect 23842 7460 23848 7472
rect 23615 7432 23848 7460
rect 23615 7429 23627 7432
rect 23569 7423 23627 7429
rect 23842 7420 23848 7432
rect 23900 7420 23906 7472
rect 25216 7463 25274 7469
rect 25216 7429 25228 7463
rect 25262 7460 25274 7463
rect 29730 7460 29736 7472
rect 25262 7432 29736 7460
rect 25262 7429 25274 7432
rect 25216 7423 25274 7429
rect 29730 7420 29736 7432
rect 29788 7420 29794 7472
rect 30009 7463 30067 7469
rect 30009 7429 30021 7463
rect 30055 7460 30067 7463
rect 31849 7463 31907 7469
rect 30055 7432 30420 7460
rect 30055 7429 30067 7432
rect 30009 7423 30067 7429
rect 30392 7404 30420 7432
rect 31128 7432 31524 7460
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7361 22339 7395
rect 22281 7355 22339 7361
rect 22370 7352 22376 7404
rect 22428 7352 22434 7404
rect 24121 7395 24179 7401
rect 24121 7392 24133 7395
rect 23768 7364 24133 7392
rect 21192 7296 21680 7324
rect 16669 7287 16727 7293
rect 4614 7216 4620 7268
rect 4672 7256 4678 7268
rect 9858 7256 9864 7268
rect 4672 7228 9864 7256
rect 4672 7216 4678 7228
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 21269 7259 21327 7265
rect 21269 7225 21281 7259
rect 21315 7225 21327 7259
rect 21652 7256 21680 7296
rect 23566 7284 23572 7336
rect 23624 7324 23630 7336
rect 23768 7333 23796 7364
rect 24121 7361 24133 7364
rect 24167 7392 24179 7395
rect 24302 7392 24308 7404
rect 24167 7364 24308 7392
rect 24167 7361 24179 7364
rect 24121 7355 24179 7361
rect 24302 7352 24308 7364
rect 24360 7352 24366 7404
rect 24397 7395 24455 7401
rect 24397 7361 24409 7395
rect 24443 7361 24455 7395
rect 24397 7355 24455 7361
rect 24581 7395 24639 7401
rect 24581 7361 24593 7395
rect 24627 7392 24639 7395
rect 24627 7364 28396 7392
rect 24627 7361 24639 7364
rect 24581 7355 24639 7361
rect 23753 7327 23811 7333
rect 23753 7324 23765 7327
rect 23624 7296 23765 7324
rect 23624 7284 23630 7296
rect 23753 7293 23765 7296
rect 23799 7293 23811 7327
rect 23753 7287 23811 7293
rect 24210 7284 24216 7336
rect 24268 7284 24274 7336
rect 22370 7256 22376 7268
rect 21652 7228 22376 7256
rect 21269 7219 21327 7225
rect 12802 7148 12808 7200
rect 12860 7188 12866 7200
rect 13357 7191 13415 7197
rect 13357 7188 13369 7191
rect 12860 7160 13369 7188
rect 12860 7148 12866 7160
rect 13357 7157 13369 7160
rect 13403 7157 13415 7191
rect 13357 7151 13415 7157
rect 17586 7148 17592 7200
rect 17644 7188 17650 7200
rect 18049 7191 18107 7197
rect 18049 7188 18061 7191
rect 17644 7160 18061 7188
rect 17644 7148 17650 7160
rect 18049 7157 18061 7160
rect 18095 7188 18107 7191
rect 18506 7188 18512 7200
rect 18095 7160 18512 7188
rect 18095 7157 18107 7160
rect 18049 7151 18107 7157
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 21284 7188 21312 7219
rect 22370 7216 22376 7228
rect 22428 7216 22434 7268
rect 24412 7256 24440 7355
rect 24946 7284 24952 7336
rect 25004 7284 25010 7336
rect 26602 7284 26608 7336
rect 26660 7324 26666 7336
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26660 7296 26985 7324
rect 26660 7284 26666 7296
rect 26973 7293 26985 7296
rect 27019 7293 27031 7327
rect 28368 7324 28396 7364
rect 29086 7352 29092 7404
rect 29144 7392 29150 7404
rect 29144 7364 30236 7392
rect 29144 7352 29150 7364
rect 28368 7296 28994 7324
rect 26973 7287 27031 7293
rect 23216 7228 24440 7256
rect 21634 7188 21640 7200
rect 21284 7160 21640 7188
rect 21634 7148 21640 7160
rect 21692 7188 21698 7200
rect 21910 7188 21916 7200
rect 21692 7160 21916 7188
rect 21692 7148 21698 7160
rect 21910 7148 21916 7160
rect 21968 7148 21974 7200
rect 22002 7148 22008 7200
rect 22060 7188 22066 7200
rect 23216 7188 23244 7228
rect 26694 7216 26700 7268
rect 26752 7256 26758 7268
rect 27249 7259 27307 7265
rect 27249 7256 27261 7259
rect 26752 7228 27261 7256
rect 26752 7216 26758 7228
rect 27249 7225 27261 7228
rect 27295 7225 27307 7259
rect 28966 7256 28994 7296
rect 29914 7284 29920 7336
rect 29972 7324 29978 7336
rect 30101 7327 30159 7333
rect 30101 7324 30113 7327
rect 29972 7296 30113 7324
rect 29972 7284 29978 7296
rect 30101 7293 30113 7296
rect 30147 7293 30159 7327
rect 30208 7324 30236 7364
rect 30374 7352 30380 7404
rect 30432 7392 30438 7404
rect 30469 7395 30527 7401
rect 30469 7392 30481 7395
rect 30432 7364 30481 7392
rect 30432 7352 30438 7364
rect 30469 7361 30481 7364
rect 30515 7361 30527 7395
rect 30469 7355 30527 7361
rect 30558 7352 30564 7404
rect 30616 7392 30622 7404
rect 30834 7392 30840 7404
rect 30616 7364 30840 7392
rect 30616 7352 30622 7364
rect 30834 7352 30840 7364
rect 30892 7392 30898 7404
rect 31021 7395 31079 7401
rect 31021 7392 31033 7395
rect 30892 7364 31033 7392
rect 30892 7352 30898 7364
rect 31021 7361 31033 7364
rect 31067 7361 31079 7395
rect 31021 7355 31079 7361
rect 30742 7324 30748 7336
rect 30208 7296 30748 7324
rect 30101 7287 30159 7293
rect 30742 7284 30748 7296
rect 30800 7284 30806 7336
rect 29181 7259 29239 7265
rect 29181 7256 29193 7259
rect 28966 7228 29193 7256
rect 27249 7219 27307 7225
rect 29181 7225 29193 7228
rect 29227 7256 29239 7259
rect 31128 7256 31156 7432
rect 31202 7352 31208 7404
rect 31260 7390 31266 7404
rect 31386 7392 31392 7404
rect 31312 7390 31392 7392
rect 31260 7364 31392 7390
rect 31260 7362 31340 7364
rect 31260 7352 31266 7362
rect 31386 7352 31392 7364
rect 31444 7352 31450 7404
rect 31496 7401 31524 7432
rect 31849 7429 31861 7463
rect 31895 7460 31907 7463
rect 31895 7432 32352 7460
rect 31895 7429 31907 7432
rect 31849 7423 31907 7429
rect 31481 7395 31539 7401
rect 31481 7361 31493 7395
rect 31527 7361 31539 7395
rect 31481 7355 31539 7361
rect 31938 7352 31944 7404
rect 31996 7352 32002 7404
rect 32324 7401 32352 7432
rect 33870 7420 33876 7472
rect 33928 7420 33934 7472
rect 32309 7395 32367 7401
rect 32309 7361 32321 7395
rect 32355 7361 32367 7395
rect 32309 7355 32367 7361
rect 32398 7352 32404 7404
rect 32456 7352 32462 7404
rect 32674 7352 32680 7404
rect 32732 7352 32738 7404
rect 33689 7395 33747 7401
rect 33689 7361 33701 7395
rect 33735 7361 33747 7395
rect 33689 7355 33747 7361
rect 31662 7333 31668 7336
rect 31619 7327 31668 7333
rect 31619 7293 31631 7327
rect 31665 7293 31668 7327
rect 31619 7287 31668 7293
rect 31662 7284 31668 7287
rect 31720 7284 31726 7336
rect 31956 7324 31984 7352
rect 32585 7327 32643 7333
rect 32585 7324 32597 7327
rect 31956 7296 32597 7324
rect 32585 7293 32597 7296
rect 32631 7293 32643 7327
rect 33704 7324 33732 7355
rect 33778 7352 33784 7404
rect 33836 7352 33842 7404
rect 34164 7401 34192 7500
rect 34606 7488 34612 7500
rect 34664 7488 34670 7540
rect 34790 7488 34796 7540
rect 34848 7528 34854 7540
rect 34848 7500 35020 7528
rect 34848 7488 34854 7500
rect 34241 7463 34299 7469
rect 34241 7429 34253 7463
rect 34287 7460 34299 7463
rect 34885 7463 34943 7469
rect 34885 7460 34897 7463
rect 34287 7432 34897 7460
rect 34287 7429 34299 7432
rect 34241 7423 34299 7429
rect 34885 7429 34897 7432
rect 34931 7429 34943 7463
rect 34885 7423 34943 7429
rect 34057 7395 34115 7401
rect 34057 7361 34069 7395
rect 34103 7361 34115 7395
rect 34057 7355 34115 7361
rect 34149 7395 34207 7401
rect 34149 7361 34161 7395
rect 34195 7361 34207 7395
rect 34149 7355 34207 7361
rect 33962 7324 33968 7336
rect 33704 7296 33968 7324
rect 32585 7287 32643 7293
rect 33962 7284 33968 7296
rect 34020 7284 34026 7336
rect 34072 7324 34100 7355
rect 34330 7352 34336 7404
rect 34388 7392 34394 7404
rect 34425 7395 34483 7401
rect 34425 7392 34437 7395
rect 34388 7364 34437 7392
rect 34388 7352 34394 7364
rect 34425 7361 34437 7364
rect 34471 7361 34483 7395
rect 34425 7355 34483 7361
rect 34514 7352 34520 7404
rect 34572 7352 34578 7404
rect 34609 7395 34667 7401
rect 34609 7361 34621 7395
rect 34655 7392 34667 7395
rect 34992 7392 35020 7500
rect 34655 7364 35020 7392
rect 34655 7361 34667 7364
rect 34609 7355 34667 7361
rect 34532 7324 34560 7352
rect 34701 7327 34759 7333
rect 34701 7324 34713 7327
rect 34072 7296 34284 7324
rect 34532 7296 34713 7324
rect 29227 7228 31156 7256
rect 29227 7225 29239 7228
rect 29181 7219 29239 7225
rect 31754 7216 31760 7268
rect 31812 7256 31818 7268
rect 32490 7256 32496 7268
rect 31812 7228 32496 7256
rect 31812 7216 31818 7228
rect 32490 7216 32496 7228
rect 32548 7216 32554 7268
rect 34256 7265 34284 7296
rect 34701 7293 34713 7296
rect 34747 7293 34759 7327
rect 34701 7287 34759 7293
rect 34790 7284 34796 7336
rect 34848 7324 34854 7336
rect 34885 7327 34943 7333
rect 34885 7324 34897 7327
rect 34848 7296 34897 7324
rect 34848 7284 34854 7296
rect 34885 7293 34897 7296
rect 34931 7293 34943 7327
rect 34885 7287 34943 7293
rect 34241 7259 34299 7265
rect 34241 7225 34253 7259
rect 34287 7225 34299 7259
rect 34241 7219 34299 7225
rect 22060 7160 23244 7188
rect 22060 7148 22066 7160
rect 23934 7148 23940 7200
rect 23992 7188 23998 7200
rect 24305 7191 24363 7197
rect 24305 7188 24317 7191
rect 23992 7160 24317 7188
rect 23992 7148 23998 7160
rect 24305 7157 24317 7160
rect 24351 7157 24363 7191
rect 24305 7151 24363 7157
rect 25958 7148 25964 7200
rect 26016 7188 26022 7200
rect 26329 7191 26387 7197
rect 26329 7188 26341 7191
rect 26016 7160 26341 7188
rect 26016 7148 26022 7160
rect 26329 7157 26341 7160
rect 26375 7157 26387 7191
rect 26329 7151 26387 7157
rect 29454 7148 29460 7200
rect 29512 7188 29518 7200
rect 29549 7191 29607 7197
rect 29549 7188 29561 7191
rect 29512 7160 29561 7188
rect 29512 7148 29518 7160
rect 29549 7157 29561 7160
rect 29595 7157 29607 7191
rect 29549 7151 29607 7157
rect 30558 7148 30564 7200
rect 30616 7148 30622 7200
rect 31113 7191 31171 7197
rect 31113 7157 31125 7191
rect 31159 7188 31171 7191
rect 31294 7188 31300 7200
rect 31159 7160 31300 7188
rect 31159 7157 31171 7160
rect 31113 7151 31171 7157
rect 31294 7148 31300 7160
rect 31352 7148 31358 7200
rect 32125 7191 32183 7197
rect 32125 7157 32137 7191
rect 32171 7188 32183 7191
rect 32306 7188 32312 7200
rect 32171 7160 32312 7188
rect 32171 7157 32183 7160
rect 32125 7151 32183 7157
rect 32306 7148 32312 7160
rect 32364 7148 32370 7200
rect 1104 7098 36800 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 36800 7098
rect 1104 7024 36800 7046
rect 10137 6987 10195 6993
rect 10137 6953 10149 6987
rect 10183 6953 10195 6987
rect 10137 6947 10195 6953
rect 5721 6919 5779 6925
rect 5721 6885 5733 6919
rect 5767 6916 5779 6919
rect 5810 6916 5816 6928
rect 5767 6888 5816 6916
rect 5767 6885 5779 6888
rect 5721 6879 5779 6885
rect 5810 6876 5816 6888
rect 5868 6876 5874 6928
rect 10152 6916 10180 6947
rect 10226 6944 10232 6996
rect 10284 6984 10290 6996
rect 10413 6987 10471 6993
rect 10413 6984 10425 6987
rect 10284 6956 10425 6984
rect 10284 6944 10290 6956
rect 10413 6953 10425 6956
rect 10459 6953 10471 6987
rect 10413 6947 10471 6953
rect 11241 6987 11299 6993
rect 11241 6953 11253 6987
rect 11287 6953 11299 6987
rect 11241 6947 11299 6953
rect 11425 6987 11483 6993
rect 11425 6953 11437 6987
rect 11471 6984 11483 6987
rect 11974 6984 11980 6996
rect 11471 6956 11980 6984
rect 11471 6953 11483 6956
rect 11425 6947 11483 6953
rect 11256 6916 11284 6947
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 19242 6984 19248 6996
rect 15028 6956 19248 6984
rect 11790 6916 11796 6928
rect 10152 6888 11796 6916
rect 11790 6876 11796 6888
rect 11848 6876 11854 6928
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5442 6848 5448 6860
rect 5399 6820 5448 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 11517 6851 11575 6857
rect 11517 6817 11529 6851
rect 11563 6848 11575 6851
rect 12710 6848 12716 6860
rect 11563 6820 12716 6848
rect 11563 6817 11575 6820
rect 11517 6811 11575 6817
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 14458 6808 14464 6860
rect 14516 6848 14522 6860
rect 15028 6857 15056 6956
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 20898 6944 20904 6996
rect 20956 6984 20962 6996
rect 22002 6984 22008 6996
rect 20956 6956 22008 6984
rect 20956 6944 20962 6956
rect 22002 6944 22008 6956
rect 22060 6944 22066 6996
rect 23566 6944 23572 6996
rect 23624 6944 23630 6996
rect 31018 6944 31024 6996
rect 31076 6984 31082 6996
rect 33594 6984 33600 6996
rect 31076 6956 33600 6984
rect 31076 6944 31082 6956
rect 33594 6944 33600 6956
rect 33652 6944 33658 6996
rect 17126 6876 17132 6928
rect 17184 6916 17190 6928
rect 25958 6916 25964 6928
rect 17184 6888 25964 6916
rect 17184 6876 17190 6888
rect 25958 6876 25964 6888
rect 26016 6876 26022 6928
rect 29362 6876 29368 6928
rect 29420 6916 29426 6928
rect 33778 6916 33784 6928
rect 29420 6888 33784 6916
rect 29420 6876 29426 6888
rect 33778 6876 33784 6888
rect 33836 6876 33842 6928
rect 15013 6851 15071 6857
rect 14516 6820 14964 6848
rect 14516 6808 14522 6820
rect 9953 6783 10011 6789
rect 2746 6752 5488 6780
rect 1946 6672 1952 6724
rect 2004 6712 2010 6724
rect 2746 6712 2774 6752
rect 2004 6684 2774 6712
rect 5460 6712 5488 6752
rect 9953 6749 9965 6783
rect 9999 6780 10011 6783
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 9999 6752 10977 6780
rect 9999 6749 10011 6752
rect 9953 6743 10011 6749
rect 10965 6749 10977 6752
rect 11011 6780 11023 6783
rect 11054 6780 11060 6792
rect 11011 6752 11060 6780
rect 11011 6749 11023 6752
rect 10965 6743 11023 6749
rect 11054 6740 11060 6752
rect 11112 6780 11118 6792
rect 14936 6789 14964 6820
rect 15013 6817 15025 6851
rect 15059 6817 15071 6851
rect 15013 6811 15071 6817
rect 15197 6851 15255 6857
rect 15197 6817 15209 6851
rect 15243 6848 15255 6851
rect 16666 6848 16672 6860
rect 15243 6820 16672 6848
rect 15243 6817 15255 6820
rect 15197 6811 15255 6817
rect 16666 6808 16672 6820
rect 16724 6808 16730 6860
rect 18230 6808 18236 6860
rect 18288 6848 18294 6860
rect 18417 6851 18475 6857
rect 18417 6848 18429 6851
rect 18288 6820 18429 6848
rect 18288 6808 18294 6820
rect 18417 6817 18429 6820
rect 18463 6817 18475 6851
rect 18417 6811 18475 6817
rect 18765 6851 18823 6857
rect 18765 6817 18777 6851
rect 18811 6848 18823 6851
rect 20438 6848 20444 6860
rect 18811 6820 20444 6848
rect 18811 6817 18823 6820
rect 18765 6811 18823 6817
rect 20438 6808 20444 6820
rect 20496 6808 20502 6860
rect 21453 6851 21511 6857
rect 21453 6817 21465 6851
rect 21499 6848 21511 6851
rect 22094 6848 22100 6860
rect 21499 6820 22100 6848
rect 21499 6817 21511 6820
rect 21453 6811 21511 6817
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 22370 6808 22376 6860
rect 22428 6808 22434 6860
rect 11793 6783 11851 6789
rect 11793 6780 11805 6783
rect 11112 6752 11805 6780
rect 11112 6740 11118 6752
rect 11793 6749 11805 6752
rect 11839 6749 11851 6783
rect 11793 6743 11851 6749
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6780 14335 6783
rect 14921 6783 14979 6789
rect 14323 6752 14596 6780
rect 14323 6749 14335 6752
rect 14277 6743 14335 6749
rect 14458 6712 14464 6724
rect 5460 6684 14464 6712
rect 2004 6672 2010 6684
rect 14458 6672 14464 6684
rect 14516 6672 14522 6724
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5813 6647 5871 6653
rect 5813 6644 5825 6647
rect 5316 6616 5825 6644
rect 5316 6604 5322 6616
rect 5813 6613 5825 6616
rect 5859 6644 5871 6647
rect 6362 6644 6368 6656
rect 5859 6616 6368 6644
rect 5859 6613 5871 6616
rect 5813 6607 5871 6613
rect 6362 6604 6368 6616
rect 6420 6604 6426 6656
rect 7282 6604 7288 6656
rect 7340 6644 7346 6656
rect 7834 6644 7840 6656
rect 7340 6616 7840 6644
rect 7340 6604 7346 6616
rect 7834 6604 7840 6616
rect 7892 6644 7898 6656
rect 8570 6644 8576 6656
rect 7892 6616 8576 6644
rect 7892 6604 7898 6616
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 14568 6653 14596 6752
rect 14921 6749 14933 6783
rect 14967 6749 14979 6783
rect 14921 6743 14979 6749
rect 18322 6740 18328 6792
rect 18380 6740 18386 6792
rect 18506 6740 18512 6792
rect 18564 6740 18570 6792
rect 18966 6780 18972 6792
rect 18616 6752 18972 6780
rect 18141 6715 18199 6721
rect 18141 6681 18153 6715
rect 18187 6712 18199 6715
rect 18616 6712 18644 6752
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 20806 6740 20812 6792
rect 20864 6780 20870 6792
rect 21637 6783 21695 6789
rect 21637 6780 21649 6783
rect 20864 6752 21649 6780
rect 20864 6740 20870 6752
rect 21637 6749 21649 6752
rect 21683 6749 21695 6783
rect 21637 6743 21695 6749
rect 18187 6684 18644 6712
rect 18187 6681 18199 6684
rect 18141 6675 18199 6681
rect 18690 6672 18696 6724
rect 18748 6672 18754 6724
rect 21652 6712 21680 6743
rect 21910 6740 21916 6792
rect 21968 6740 21974 6792
rect 22462 6740 22468 6792
rect 22520 6780 22526 6792
rect 25976 6789 26004 6876
rect 30558 6808 30564 6860
rect 30616 6848 30622 6860
rect 31297 6851 31355 6857
rect 31297 6848 31309 6851
rect 30616 6820 31309 6848
rect 30616 6808 30622 6820
rect 31297 6817 31309 6820
rect 31343 6848 31355 6851
rect 31754 6848 31760 6860
rect 31343 6820 31760 6848
rect 31343 6817 31355 6820
rect 31297 6811 31355 6817
rect 31754 6808 31760 6820
rect 31812 6808 31818 6860
rect 23385 6783 23443 6789
rect 23385 6780 23397 6783
rect 22520 6752 23397 6780
rect 22520 6740 22526 6752
rect 23385 6749 23397 6752
rect 23431 6749 23443 6783
rect 23385 6743 23443 6749
rect 25961 6783 26019 6789
rect 25961 6749 25973 6783
rect 26007 6749 26019 6783
rect 25961 6743 26019 6749
rect 28902 6740 28908 6792
rect 28960 6740 28966 6792
rect 29086 6740 29092 6792
rect 29144 6740 29150 6792
rect 31202 6740 31208 6792
rect 31260 6780 31266 6792
rect 31389 6783 31447 6789
rect 31389 6780 31401 6783
rect 31260 6752 31401 6780
rect 31260 6740 31266 6752
rect 31389 6749 31401 6752
rect 31435 6749 31447 6783
rect 31389 6743 31447 6749
rect 31478 6740 31484 6792
rect 31536 6740 31542 6792
rect 31573 6783 31631 6789
rect 31573 6749 31585 6783
rect 31619 6780 31631 6783
rect 31662 6780 31668 6792
rect 31619 6752 31668 6780
rect 31619 6749 31631 6752
rect 31573 6743 31631 6749
rect 31662 6740 31668 6752
rect 31720 6740 31726 6792
rect 33870 6740 33876 6792
rect 33928 6780 33934 6792
rect 34790 6780 34796 6792
rect 33928 6752 34796 6780
rect 33928 6740 33934 6752
rect 34790 6740 34796 6752
rect 34848 6740 34854 6792
rect 22002 6712 22008 6724
rect 21652 6684 22008 6712
rect 22002 6672 22008 6684
rect 22060 6672 22066 6724
rect 22189 6715 22247 6721
rect 22189 6681 22201 6715
rect 22235 6712 22247 6715
rect 22554 6712 22560 6724
rect 22235 6684 22560 6712
rect 22235 6681 22247 6684
rect 22189 6675 22247 6681
rect 22554 6672 22560 6684
rect 22612 6672 22618 6724
rect 26145 6715 26203 6721
rect 26145 6681 26157 6715
rect 26191 6712 26203 6715
rect 26694 6712 26700 6724
rect 26191 6684 26700 6712
rect 26191 6681 26203 6684
rect 26145 6675 26203 6681
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 30374 6672 30380 6724
rect 30432 6712 30438 6724
rect 31496 6712 31524 6740
rect 30432 6684 31524 6712
rect 30432 6672 30438 6684
rect 14553 6647 14611 6653
rect 14553 6613 14565 6647
rect 14599 6613 14611 6647
rect 14553 6607 14611 6613
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 18877 6647 18935 6653
rect 18877 6644 18889 6647
rect 18380 6616 18889 6644
rect 18380 6604 18386 6616
rect 18877 6613 18889 6616
rect 18923 6613 18935 6647
rect 18877 6607 18935 6613
rect 21818 6604 21824 6656
rect 21876 6644 21882 6656
rect 22094 6644 22100 6656
rect 21876 6616 22100 6644
rect 21876 6604 21882 6616
rect 22094 6604 22100 6616
rect 22152 6604 22158 6656
rect 28994 6604 29000 6656
rect 29052 6644 29058 6656
rect 29089 6647 29147 6653
rect 29089 6644 29101 6647
rect 29052 6616 29101 6644
rect 29052 6604 29058 6616
rect 29089 6613 29101 6616
rect 29135 6644 29147 6647
rect 29362 6644 29368 6656
rect 29135 6616 29368 6644
rect 29135 6613 29147 6616
rect 29089 6607 29147 6613
rect 29362 6604 29368 6616
rect 29420 6604 29426 6656
rect 31113 6647 31171 6653
rect 31113 6613 31125 6647
rect 31159 6644 31171 6647
rect 31386 6644 31392 6656
rect 31159 6616 31392 6644
rect 31159 6613 31171 6616
rect 31113 6607 31171 6613
rect 31386 6604 31392 6616
rect 31444 6604 31450 6656
rect 33962 6604 33968 6656
rect 34020 6604 34026 6656
rect 1104 6554 36800 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 36800 6554
rect 1104 6480 36800 6502
rect 5350 6400 5356 6452
rect 5408 6440 5414 6452
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 5408 6412 5457 6440
rect 5408 6400 5414 6412
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 5644 6412 6592 6440
rect 1670 6381 1676 6384
rect 1664 6372 1676 6381
rect 1631 6344 1676 6372
rect 1664 6335 1676 6344
rect 1670 6332 1676 6335
rect 1728 6332 1734 6384
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6304 1455 6307
rect 4062 6304 4068 6316
rect 1443 6276 4068 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5184 6236 5212 6267
rect 5258 6264 5264 6316
rect 5316 6264 5322 6316
rect 5644 6304 5672 6412
rect 5368 6276 5672 6304
rect 5368 6236 5396 6276
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 6564 6313 6592 6412
rect 7558 6400 7564 6452
rect 7616 6400 7622 6452
rect 10413 6443 10471 6449
rect 7668 6412 9674 6440
rect 7668 6372 7696 6412
rect 9646 6372 9674 6412
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 10502 6440 10508 6452
rect 10459 6412 10508 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 14182 6400 14188 6452
rect 14240 6440 14246 6452
rect 14553 6443 14611 6449
rect 14553 6440 14565 6443
rect 14240 6412 14565 6440
rect 14240 6400 14246 6412
rect 14553 6409 14565 6412
rect 14599 6409 14611 6443
rect 14553 6403 14611 6409
rect 15381 6443 15439 6449
rect 15381 6409 15393 6443
rect 15427 6409 15439 6443
rect 15381 6403 15439 6409
rect 15473 6443 15531 6449
rect 15473 6409 15485 6443
rect 15519 6440 15531 6443
rect 15654 6440 15660 6452
rect 15519 6412 15660 6440
rect 15519 6409 15531 6412
rect 15473 6403 15531 6409
rect 13440 6375 13498 6381
rect 7576 6344 7696 6372
rect 8128 6344 8708 6372
rect 9646 6344 11652 6372
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6304 6607 6307
rect 7374 6304 7380 6316
rect 6595 6276 7380 6304
rect 6595 6273 6607 6276
rect 6549 6267 6607 6273
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 7466 6264 7472 6316
rect 7524 6264 7530 6316
rect 5184 6208 5396 6236
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6236 5503 6239
rect 5736 6236 5764 6264
rect 5491 6208 5764 6236
rect 5813 6239 5871 6245
rect 5491 6205 5503 6208
rect 5445 6199 5503 6205
rect 5813 6205 5825 6239
rect 5859 6236 5871 6239
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 5859 6208 6469 6236
rect 5859 6205 5871 6208
rect 5813 6199 5871 6205
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 7576 6236 7604 6344
rect 8128 6316 8156 6344
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 7834 6304 7840 6316
rect 7699 6276 7840 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 7834 6264 7840 6276
rect 7892 6264 7898 6316
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6304 7987 6307
rect 8018 6304 8024 6316
rect 7975 6276 8024 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8110 6264 8116 6316
rect 8168 6264 8174 6316
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8478 6304 8484 6316
rect 8251 6276 8484 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 8680 6313 8708 6344
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 9953 6307 10011 6313
rect 9953 6273 9965 6307
rect 9999 6304 10011 6307
rect 11054 6304 11060 6316
rect 9999 6276 11060 6304
rect 9999 6273 10011 6276
rect 9953 6267 10011 6273
rect 11054 6264 11060 6276
rect 11112 6264 11118 6316
rect 11330 6264 11336 6316
rect 11388 6304 11394 6316
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 11388 6276 11529 6304
rect 11388 6264 11394 6276
rect 11517 6273 11529 6276
rect 11563 6273 11575 6307
rect 11624 6304 11652 6344
rect 13440 6341 13452 6375
rect 13486 6372 13498 6375
rect 14090 6372 14096 6384
rect 13486 6344 14096 6372
rect 13486 6341 13498 6344
rect 13440 6335 13498 6341
rect 14090 6332 14096 6344
rect 14148 6332 14154 6384
rect 14458 6332 14464 6384
rect 14516 6372 14522 6384
rect 15105 6375 15163 6381
rect 15105 6372 15117 6375
rect 14516 6344 15117 6372
rect 14516 6332 14522 6344
rect 15105 6341 15117 6344
rect 15151 6341 15163 6375
rect 15396 6372 15424 6403
rect 15654 6400 15660 6412
rect 15712 6440 15718 6452
rect 16298 6440 16304 6452
rect 15712 6412 16304 6440
rect 15712 6400 15718 6412
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 17313 6443 17371 6449
rect 17313 6409 17325 6443
rect 17359 6440 17371 6443
rect 19978 6440 19984 6452
rect 17359 6412 19984 6440
rect 17359 6409 17371 6412
rect 17313 6403 17371 6409
rect 19978 6400 19984 6412
rect 20036 6400 20042 6452
rect 22002 6400 22008 6452
rect 22060 6400 22066 6452
rect 22094 6400 22100 6452
rect 22152 6440 22158 6452
rect 22649 6443 22707 6449
rect 22649 6440 22661 6443
rect 22152 6412 22661 6440
rect 22152 6400 22158 6412
rect 22649 6409 22661 6412
rect 22695 6409 22707 6443
rect 22649 6403 22707 6409
rect 23569 6443 23627 6449
rect 23569 6409 23581 6443
rect 23615 6440 23627 6443
rect 24210 6440 24216 6452
rect 23615 6412 24216 6440
rect 23615 6409 23627 6412
rect 23569 6403 23627 6409
rect 24210 6400 24216 6412
rect 24268 6400 24274 6452
rect 27801 6443 27859 6449
rect 27801 6409 27813 6443
rect 27847 6440 27859 6443
rect 28166 6440 28172 6452
rect 27847 6412 28172 6440
rect 27847 6409 27859 6412
rect 27801 6403 27859 6409
rect 28166 6400 28172 6412
rect 28224 6440 28230 6452
rect 33134 6440 33140 6452
rect 28224 6412 28396 6440
rect 28224 6400 28230 6412
rect 15562 6372 15568 6384
rect 15396 6344 15568 6372
rect 15105 6335 15163 6341
rect 15562 6332 15568 6344
rect 15620 6372 15626 6384
rect 16758 6372 16764 6384
rect 15620 6344 16764 6372
rect 15620 6332 15626 6344
rect 16758 6332 16764 6344
rect 16816 6332 16822 6384
rect 18509 6375 18567 6381
rect 18509 6341 18521 6375
rect 18555 6372 18567 6375
rect 18690 6372 18696 6384
rect 18555 6344 18696 6372
rect 18555 6341 18567 6344
rect 18509 6335 18567 6341
rect 18690 6332 18696 6344
rect 18748 6372 18754 6384
rect 19245 6375 19303 6381
rect 19245 6372 19257 6375
rect 18748 6344 19257 6372
rect 18748 6332 18754 6344
rect 19245 6341 19257 6344
rect 19291 6341 19303 6375
rect 22020 6372 22048 6400
rect 28368 6381 28396 6412
rect 31312 6412 33140 6440
rect 28353 6375 28411 6381
rect 22020 6344 22324 6372
rect 19245 6335 19303 6341
rect 14550 6304 14556 6316
rect 11624 6276 14556 6304
rect 11517 6267 11575 6273
rect 14550 6264 14556 6276
rect 14608 6264 14614 6316
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6304 15347 6307
rect 15378 6304 15384 6316
rect 15335 6276 15384 6304
rect 15335 6273 15347 6276
rect 15289 6267 15347 6273
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6304 15715 6307
rect 16206 6304 16212 6316
rect 15703 6276 16212 6304
rect 15703 6273 15715 6276
rect 15657 6267 15715 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 17221 6307 17279 6313
rect 17221 6273 17233 6307
rect 17267 6304 17279 6307
rect 17310 6304 17316 6316
rect 17267 6276 17316 6304
rect 17267 6273 17279 6276
rect 17221 6267 17279 6273
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17405 6307 17463 6313
rect 17405 6273 17417 6307
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 17589 6307 17647 6313
rect 17589 6273 17601 6307
rect 17635 6304 17647 6307
rect 18230 6304 18236 6316
rect 17635 6276 18236 6304
rect 17635 6273 17647 6276
rect 17589 6267 17647 6273
rect 6457 6199 6515 6205
rect 6564 6208 7604 6236
rect 8128 6236 8156 6264
rect 8297 6239 8355 6245
rect 8297 6236 8309 6239
rect 8128 6208 8309 6236
rect 6086 6128 6092 6180
rect 6144 6128 6150 6180
rect 2777 6103 2835 6109
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 6564 6100 6592 6208
rect 8297 6205 8309 6208
rect 8343 6205 8355 6239
rect 8496 6236 8524 6264
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8496 6208 8953 6236
rect 8297 6199 8355 6205
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 11790 6196 11796 6248
rect 11848 6196 11854 6248
rect 13173 6239 13231 6245
rect 13173 6205 13185 6239
rect 13219 6205 13231 6239
rect 16574 6236 16580 6248
rect 13173 6199 13231 6205
rect 14200 6208 16580 6236
rect 8570 6128 8576 6180
rect 8628 6128 8634 6180
rect 8662 6128 8668 6180
rect 8720 6168 8726 6180
rect 8849 6171 8907 6177
rect 8849 6168 8861 6171
rect 8720 6140 8861 6168
rect 8720 6128 8726 6140
rect 8849 6137 8861 6140
rect 8895 6137 8907 6171
rect 8849 6131 8907 6137
rect 2823 6072 6592 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 8205 6103 8263 6109
rect 8205 6100 8217 6103
rect 7616 6072 8217 6100
rect 7616 6060 7622 6072
rect 8205 6069 8217 6072
rect 8251 6100 8263 6103
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 8251 6072 8769 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 8757 6063 8815 6069
rect 10226 6060 10232 6112
rect 10284 6060 10290 6112
rect 13188 6100 13216 6199
rect 14200 6100 14228 6208
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 17126 6196 17132 6248
rect 17184 6236 17190 6248
rect 17420 6236 17448 6267
rect 18230 6264 18236 6276
rect 18288 6264 18294 6316
rect 18874 6264 18880 6316
rect 18932 6264 18938 6316
rect 18969 6310 19027 6313
rect 19058 6310 19064 6316
rect 18969 6307 19064 6310
rect 18969 6273 18981 6307
rect 19015 6282 19064 6307
rect 19015 6273 19027 6282
rect 18969 6267 19027 6273
rect 19058 6264 19064 6282
rect 19116 6264 19122 6316
rect 20625 6307 20683 6313
rect 20625 6273 20637 6307
rect 20671 6304 20683 6307
rect 20714 6304 20720 6316
rect 20671 6276 20720 6304
rect 20671 6273 20683 6276
rect 20625 6267 20683 6273
rect 20714 6264 20720 6276
rect 20772 6264 20778 6316
rect 20809 6307 20867 6313
rect 20809 6273 20821 6307
rect 20855 6304 20867 6307
rect 21818 6304 21824 6316
rect 20855 6276 21824 6304
rect 20855 6273 20867 6276
rect 20809 6267 20867 6273
rect 17865 6239 17923 6245
rect 17865 6236 17877 6239
rect 17184 6208 17877 6236
rect 17184 6196 17190 6208
rect 17865 6205 17877 6208
rect 17911 6205 17923 6239
rect 18248 6236 18276 6264
rect 18693 6239 18751 6245
rect 18693 6236 18705 6239
rect 18248 6208 18705 6236
rect 17865 6199 17923 6205
rect 18693 6205 18705 6208
rect 18739 6205 18751 6239
rect 18693 6199 18751 6205
rect 18782 6196 18788 6248
rect 18840 6196 18846 6248
rect 19242 6196 19248 6248
rect 19300 6236 19306 6248
rect 20824 6236 20852 6267
rect 21818 6264 21824 6276
rect 21876 6264 21882 6316
rect 21910 6264 21916 6316
rect 21968 6304 21974 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21968 6276 22017 6304
rect 21968 6264 21974 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22094 6264 22100 6316
rect 22152 6264 22158 6316
rect 22296 6313 22324 6344
rect 27632 6344 28212 6372
rect 22281 6307 22339 6313
rect 22281 6273 22293 6307
rect 22327 6273 22339 6307
rect 22281 6267 22339 6273
rect 22373 6307 22431 6313
rect 22373 6273 22385 6307
rect 22419 6273 22431 6307
rect 22373 6267 22431 6273
rect 19300 6208 20852 6236
rect 22388 6236 22416 6267
rect 22554 6264 22560 6316
rect 22612 6264 22618 6316
rect 22646 6264 22652 6316
rect 22704 6304 22710 6316
rect 23385 6307 23443 6313
rect 23385 6304 23397 6307
rect 22704 6276 23397 6304
rect 22704 6264 22710 6276
rect 23385 6273 23397 6276
rect 23431 6273 23443 6307
rect 23385 6267 23443 6273
rect 23934 6264 23940 6316
rect 23992 6264 23998 6316
rect 25038 6264 25044 6316
rect 25096 6304 25102 6316
rect 25317 6307 25375 6313
rect 25317 6304 25329 6307
rect 25096 6276 25329 6304
rect 25096 6264 25102 6276
rect 25317 6273 25329 6276
rect 25363 6273 25375 6307
rect 25317 6267 25375 6273
rect 25501 6307 25559 6313
rect 25501 6273 25513 6307
rect 25547 6304 25559 6307
rect 25682 6304 25688 6316
rect 25547 6276 25688 6304
rect 25547 6273 25559 6276
rect 25501 6267 25559 6273
rect 25682 6264 25688 6276
rect 25740 6264 25746 6316
rect 27522 6264 27528 6316
rect 27580 6304 27586 6316
rect 27632 6313 27660 6344
rect 28184 6313 28212 6344
rect 28353 6341 28365 6375
rect 28399 6341 28411 6375
rect 29086 6372 29092 6384
rect 28353 6335 28411 6341
rect 28552 6344 29092 6372
rect 27617 6307 27675 6313
rect 27617 6304 27629 6307
rect 27580 6276 27629 6304
rect 27580 6264 27586 6276
rect 27617 6273 27629 6276
rect 27663 6273 27675 6307
rect 27617 6267 27675 6273
rect 27893 6307 27951 6313
rect 27893 6273 27905 6307
rect 27939 6273 27951 6307
rect 27893 6267 27951 6273
rect 28169 6307 28227 6313
rect 28169 6273 28181 6307
rect 28215 6273 28227 6307
rect 28169 6267 28227 6273
rect 28261 6307 28319 6313
rect 28261 6273 28273 6307
rect 28307 6304 28319 6307
rect 28442 6304 28448 6316
rect 28307 6276 28448 6304
rect 28307 6273 28319 6276
rect 28261 6267 28319 6273
rect 24210 6236 24216 6248
rect 22388 6208 24216 6236
rect 19300 6196 19306 6208
rect 24210 6196 24216 6208
rect 24268 6196 24274 6248
rect 27908 6236 27936 6267
rect 28276 6236 28304 6267
rect 28442 6264 28448 6276
rect 28500 6264 28506 6316
rect 28552 6313 28580 6344
rect 29086 6332 29092 6344
rect 29144 6332 29150 6384
rect 31312 6316 31340 6412
rect 33134 6400 33140 6412
rect 33192 6440 33198 6452
rect 33962 6440 33968 6452
rect 33192 6412 33968 6440
rect 33192 6400 33198 6412
rect 33962 6400 33968 6412
rect 34020 6400 34026 6452
rect 28537 6307 28595 6313
rect 28537 6273 28549 6307
rect 28583 6273 28595 6307
rect 28537 6267 28595 6273
rect 28629 6307 28687 6313
rect 28629 6273 28641 6307
rect 28675 6304 28687 6307
rect 28902 6304 28908 6316
rect 28675 6276 28908 6304
rect 28675 6273 28687 6276
rect 28629 6267 28687 6273
rect 28902 6264 28908 6276
rect 28960 6264 28966 6316
rect 29454 6264 29460 6316
rect 29512 6264 29518 6316
rect 31110 6264 31116 6316
rect 31168 6304 31174 6316
rect 31294 6304 31300 6316
rect 31168 6276 31300 6304
rect 31168 6264 31174 6276
rect 31294 6264 31300 6276
rect 31352 6264 31358 6316
rect 31386 6264 31392 6316
rect 31444 6264 31450 6316
rect 31481 6307 31539 6313
rect 31481 6273 31493 6307
rect 31527 6304 31539 6307
rect 31570 6304 31576 6316
rect 31527 6276 31576 6304
rect 31527 6273 31539 6276
rect 31481 6267 31539 6273
rect 31570 6264 31576 6276
rect 31628 6264 31634 6316
rect 27908 6208 28304 6236
rect 31205 6239 31263 6245
rect 31205 6205 31217 6239
rect 31251 6205 31263 6239
rect 31205 6199 31263 6205
rect 14550 6128 14556 6180
rect 14608 6168 14614 6180
rect 24854 6168 24860 6180
rect 14608 6140 24860 6168
rect 14608 6128 14614 6140
rect 24854 6128 24860 6140
rect 24912 6128 24918 6180
rect 26694 6128 26700 6180
rect 26752 6168 26758 6180
rect 30834 6168 30840 6180
rect 26752 6140 30840 6168
rect 26752 6128 26758 6140
rect 30834 6128 30840 6140
rect 30892 6128 30898 6180
rect 31220 6168 31248 6199
rect 31846 6168 31852 6180
rect 31220 6140 31852 6168
rect 31846 6128 31852 6140
rect 31904 6128 31910 6180
rect 13188 6072 14228 6100
rect 16298 6060 16304 6112
rect 16356 6100 16362 6112
rect 18322 6100 18328 6112
rect 16356 6072 18328 6100
rect 16356 6060 16362 6072
rect 18322 6060 18328 6072
rect 18380 6060 18386 6112
rect 19334 6060 19340 6112
rect 19392 6060 19398 6112
rect 20622 6060 20628 6112
rect 20680 6060 20686 6112
rect 21174 6060 21180 6112
rect 21232 6100 21238 6112
rect 21821 6103 21879 6109
rect 21821 6100 21833 6103
rect 21232 6072 21833 6100
rect 21232 6060 21238 6072
rect 21821 6069 21833 6072
rect 21867 6069 21879 6103
rect 21821 6063 21879 6069
rect 23658 6060 23664 6112
rect 23716 6100 23722 6112
rect 23753 6103 23811 6109
rect 23753 6100 23765 6103
rect 23716 6072 23765 6100
rect 23716 6060 23722 6072
rect 23753 6069 23765 6072
rect 23799 6069 23811 6103
rect 23753 6063 23811 6069
rect 25317 6103 25375 6109
rect 25317 6069 25329 6103
rect 25363 6100 25375 6103
rect 25866 6100 25872 6112
rect 25363 6072 25872 6100
rect 25363 6069 25375 6072
rect 25317 6063 25375 6069
rect 25866 6060 25872 6072
rect 25924 6060 25930 6112
rect 27614 6060 27620 6112
rect 27672 6060 27678 6112
rect 27706 6060 27712 6112
rect 27764 6100 27770 6112
rect 27985 6103 28043 6109
rect 27985 6100 27997 6103
rect 27764 6072 27997 6100
rect 27764 6060 27770 6072
rect 27985 6069 27997 6072
rect 28031 6069 28043 6103
rect 27985 6063 28043 6069
rect 29273 6103 29331 6109
rect 29273 6069 29285 6103
rect 29319 6100 29331 6103
rect 29638 6100 29644 6112
rect 29319 6072 29644 6100
rect 29319 6069 29331 6072
rect 29273 6063 29331 6069
rect 29638 6060 29644 6072
rect 29696 6060 29702 6112
rect 31018 6060 31024 6112
rect 31076 6060 31082 6112
rect 31294 6060 31300 6112
rect 31352 6100 31358 6112
rect 31938 6100 31944 6112
rect 31352 6072 31944 6100
rect 31352 6060 31358 6072
rect 31938 6060 31944 6072
rect 31996 6060 32002 6112
rect 1104 6010 36800 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 36800 6010
rect 1104 5936 36800 5958
rect 1302 5856 1308 5908
rect 1360 5896 1366 5908
rect 1581 5899 1639 5905
rect 1581 5896 1593 5899
rect 1360 5868 1593 5896
rect 1360 5856 1366 5868
rect 1581 5865 1593 5868
rect 1627 5865 1639 5899
rect 1581 5859 1639 5865
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 7561 5899 7619 5905
rect 7561 5896 7573 5899
rect 7524 5868 7573 5896
rect 7524 5856 7530 5868
rect 7561 5865 7573 5868
rect 7607 5896 7619 5899
rect 8018 5896 8024 5908
rect 7607 5868 8024 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 8481 5899 8539 5905
rect 8481 5896 8493 5899
rect 8128 5868 8493 5896
rect 1854 5788 1860 5840
rect 1912 5828 1918 5840
rect 8128 5837 8156 5868
rect 8481 5865 8493 5868
rect 8527 5865 8539 5899
rect 8481 5859 8539 5865
rect 10689 5899 10747 5905
rect 10689 5865 10701 5899
rect 10735 5896 10747 5899
rect 10870 5896 10876 5908
rect 10735 5868 10876 5896
rect 10735 5865 10747 5868
rect 10689 5859 10747 5865
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11241 5899 11299 5905
rect 11241 5865 11253 5899
rect 11287 5896 11299 5899
rect 11790 5896 11796 5908
rect 11287 5868 11796 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 12161 5899 12219 5905
rect 12161 5865 12173 5899
rect 12207 5896 12219 5899
rect 12802 5896 12808 5908
rect 12207 5868 12808 5896
rect 12207 5865 12219 5868
rect 12161 5859 12219 5865
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 12897 5899 12955 5905
rect 12897 5865 12909 5899
rect 12943 5896 12955 5899
rect 12986 5896 12992 5908
rect 12943 5868 12992 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 15841 5899 15899 5905
rect 15841 5896 15853 5899
rect 14292 5868 15853 5896
rect 8113 5831 8171 5837
rect 1912 5800 2774 5828
rect 1912 5788 1918 5800
rect 2746 5760 2774 5800
rect 8113 5797 8125 5831
rect 8159 5797 8171 5831
rect 14292 5828 14320 5868
rect 15841 5865 15853 5868
rect 15887 5865 15899 5899
rect 18506 5896 18512 5908
rect 15841 5859 15899 5865
rect 17144 5868 18512 5896
rect 17144 5837 17172 5868
rect 18506 5856 18512 5868
rect 18564 5896 18570 5908
rect 18782 5896 18788 5908
rect 18564 5868 18788 5896
rect 18564 5856 18570 5868
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 20993 5899 21051 5905
rect 20993 5865 21005 5899
rect 21039 5896 21051 5899
rect 21358 5896 21364 5908
rect 21039 5868 21364 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 21358 5856 21364 5868
rect 21416 5856 21422 5908
rect 22462 5896 22468 5908
rect 21468 5868 22468 5896
rect 8113 5791 8171 5797
rect 8220 5800 14320 5828
rect 14737 5831 14795 5837
rect 8220 5760 8248 5800
rect 14737 5797 14749 5831
rect 14783 5797 14795 5831
rect 17129 5831 17187 5837
rect 17129 5828 17141 5831
rect 14737 5791 14795 5797
rect 16776 5800 17141 5828
rect 2746 5732 8248 5760
rect 8570 5720 8576 5772
rect 8628 5760 8634 5772
rect 8628 5732 9168 5760
rect 8628 5720 8634 5732
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 5810 5692 5816 5704
rect 1443 5664 5816 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 7282 5652 7288 5704
rect 7340 5652 7346 5704
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 7432 5664 7849 5692
rect 7432 5652 7438 5664
rect 7837 5661 7849 5664
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 7926 5652 7932 5704
rect 7984 5692 7990 5704
rect 7984 5664 8616 5692
rect 7984 5652 7990 5664
rect 8588 5633 8616 5664
rect 8662 5652 8668 5704
rect 8720 5692 8726 5704
rect 9140 5701 9168 5732
rect 9214 5720 9220 5772
rect 9272 5760 9278 5772
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 9272 5732 10057 5760
rect 9272 5720 9278 5732
rect 10045 5729 10057 5732
rect 10091 5729 10103 5763
rect 10045 5723 10103 5729
rect 11425 5763 11483 5769
rect 11425 5729 11437 5763
rect 11471 5760 11483 5763
rect 12526 5760 12532 5772
rect 11471 5732 12532 5760
rect 11471 5729 11483 5732
rect 11425 5723 11483 5729
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 14752 5760 14780 5791
rect 14752 5732 15884 5760
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8720 5664 8953 5692
rect 8720 5652 8726 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9950 5652 9956 5704
rect 10008 5652 10014 5704
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 10229 5655 10287 5661
rect 10965 5695 11023 5701
rect 10965 5661 10977 5695
rect 11011 5692 11023 5695
rect 11054 5692 11060 5704
rect 11011 5664 11060 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 8389 5627 8447 5633
rect 8389 5624 8401 5627
rect 7944 5596 8401 5624
rect 7742 5516 7748 5568
rect 7800 5556 7806 5568
rect 7944 5556 7972 5596
rect 8389 5593 8401 5596
rect 8435 5593 8447 5627
rect 8389 5587 8447 5593
rect 8573 5627 8631 5633
rect 8573 5593 8585 5627
rect 8619 5593 8631 5627
rect 10244 5624 10272 5655
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 8573 5587 8631 5593
rect 9784 5596 10272 5624
rect 7800 5528 7972 5556
rect 7800 5516 7806 5528
rect 8294 5516 8300 5568
rect 8352 5516 8358 5568
rect 9309 5559 9367 5565
rect 9309 5525 9321 5559
rect 9355 5556 9367 5559
rect 9674 5556 9680 5568
rect 9355 5528 9680 5556
rect 9355 5525 9367 5528
rect 9309 5519 9367 5525
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 9784 5565 9812 5596
rect 9769 5559 9827 5565
rect 9769 5525 9781 5559
rect 9815 5525 9827 5559
rect 9769 5519 9827 5525
rect 9858 5516 9864 5568
rect 9916 5556 9922 5568
rect 11532 5556 11560 5655
rect 11716 5624 11744 5655
rect 12250 5652 12256 5704
rect 12308 5652 12314 5704
rect 12434 5652 12440 5704
rect 12492 5652 12498 5704
rect 14918 5652 14924 5704
rect 14976 5652 14982 5704
rect 15013 5695 15071 5701
rect 15013 5661 15025 5695
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 15105 5695 15163 5701
rect 15105 5661 15117 5695
rect 15151 5692 15163 5695
rect 15470 5692 15476 5704
rect 15151 5664 15476 5692
rect 15151 5661 15163 5664
rect 15105 5655 15163 5661
rect 12618 5624 12624 5636
rect 11716 5596 12624 5624
rect 12618 5584 12624 5596
rect 12676 5584 12682 5636
rect 14737 5627 14795 5633
rect 14737 5593 14749 5627
rect 14783 5624 14795 5627
rect 15028 5624 15056 5655
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 15562 5652 15568 5704
rect 15620 5701 15626 5704
rect 15856 5701 15884 5732
rect 16776 5701 16804 5800
rect 17129 5797 17141 5800
rect 17175 5797 17187 5831
rect 17129 5791 17187 5797
rect 17865 5831 17923 5837
rect 17865 5797 17877 5831
rect 17911 5828 17923 5831
rect 20162 5828 20168 5840
rect 17911 5800 20168 5828
rect 17911 5797 17923 5800
rect 17865 5791 17923 5797
rect 20162 5788 20168 5800
rect 20220 5788 20226 5840
rect 17218 5720 17224 5772
rect 17276 5760 17282 5772
rect 17681 5763 17739 5769
rect 17681 5760 17693 5763
rect 17276 5732 17693 5760
rect 17276 5720 17282 5732
rect 17681 5729 17693 5732
rect 17727 5760 17739 5763
rect 18874 5760 18880 5772
rect 17727 5732 18880 5760
rect 17727 5729 17739 5732
rect 17681 5723 17739 5729
rect 18064 5701 18092 5732
rect 18874 5720 18880 5732
rect 18932 5720 18938 5772
rect 18966 5720 18972 5772
rect 19024 5760 19030 5772
rect 19429 5763 19487 5769
rect 19429 5760 19441 5763
rect 19024 5732 19441 5760
rect 19024 5720 19030 5732
rect 19429 5729 19441 5732
rect 19475 5729 19487 5763
rect 20180 5760 20208 5788
rect 20180 5732 21312 5760
rect 19429 5723 19487 5729
rect 15620 5695 15648 5701
rect 15636 5661 15648 5695
rect 15620 5655 15648 5661
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5661 16083 5695
rect 16025 5655 16083 5661
rect 16761 5695 16819 5701
rect 16761 5661 16773 5695
rect 16807 5661 16819 5695
rect 16761 5655 16819 5661
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5692 18107 5695
rect 18233 5695 18291 5701
rect 18095 5664 18129 5692
rect 18095 5661 18107 5664
rect 18049 5655 18107 5661
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 18322 5692 18328 5704
rect 18279 5664 18328 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 15620 5652 15626 5655
rect 15580 5624 15608 5652
rect 16040 5624 16068 5655
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5692 19303 5695
rect 19334 5692 19340 5704
rect 19291 5664 19340 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 19702 5652 19708 5704
rect 19760 5652 19766 5704
rect 19978 5652 19984 5704
rect 20036 5652 20042 5704
rect 20070 5652 20076 5704
rect 20128 5692 20134 5704
rect 20165 5695 20223 5701
rect 20165 5692 20177 5695
rect 20128 5664 20177 5692
rect 20128 5652 20134 5664
rect 20165 5661 20177 5664
rect 20211 5661 20223 5695
rect 20165 5655 20223 5661
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 20548 5701 20576 5732
rect 20533 5695 20591 5701
rect 20312 5664 20357 5692
rect 20312 5652 20318 5664
rect 20533 5661 20545 5695
rect 20579 5661 20591 5695
rect 20533 5655 20591 5661
rect 20622 5652 20628 5704
rect 20680 5701 20686 5704
rect 20680 5692 20688 5701
rect 20680 5664 20725 5692
rect 20680 5655 20688 5664
rect 20680 5652 20686 5655
rect 21174 5652 21180 5704
rect 21232 5652 21238 5704
rect 21284 5701 21312 5732
rect 21468 5701 21496 5868
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 22554 5856 22560 5908
rect 22612 5896 22618 5908
rect 22925 5899 22983 5905
rect 22925 5896 22937 5899
rect 22612 5868 22937 5896
rect 22612 5856 22618 5868
rect 22925 5865 22937 5868
rect 22971 5865 22983 5899
rect 22925 5859 22983 5865
rect 24210 5856 24216 5908
rect 24268 5856 24274 5908
rect 25685 5899 25743 5905
rect 25685 5865 25697 5899
rect 25731 5896 25743 5899
rect 27617 5899 27675 5905
rect 25731 5868 26740 5896
rect 25731 5865 25743 5868
rect 25685 5859 25743 5865
rect 24857 5831 24915 5837
rect 24857 5797 24869 5831
rect 24903 5828 24915 5831
rect 25038 5828 25044 5840
rect 24903 5800 25044 5828
rect 24903 5797 24915 5800
rect 24857 5791 24915 5797
rect 25038 5788 25044 5800
rect 25096 5788 25102 5840
rect 25866 5788 25872 5840
rect 25924 5828 25930 5840
rect 26513 5831 26571 5837
rect 26513 5828 26525 5831
rect 25924 5800 26525 5828
rect 25924 5788 25930 5800
rect 26513 5797 26525 5800
rect 26559 5797 26571 5831
rect 26513 5791 26571 5797
rect 26145 5763 26203 5769
rect 26145 5760 26157 5763
rect 23860 5732 26157 5760
rect 23860 5704 23888 5732
rect 26145 5729 26157 5732
rect 26191 5760 26203 5763
rect 26602 5760 26608 5772
rect 26191 5732 26608 5760
rect 26191 5729 26203 5732
rect 26145 5723 26203 5729
rect 26602 5720 26608 5732
rect 26660 5720 26666 5772
rect 26712 5760 26740 5868
rect 27617 5865 27629 5899
rect 27663 5896 27675 5899
rect 27663 5868 30512 5896
rect 27663 5865 27675 5868
rect 27617 5859 27675 5865
rect 30484 5828 30512 5868
rect 31294 5856 31300 5908
rect 31352 5896 31358 5908
rect 31573 5899 31631 5905
rect 31573 5896 31585 5899
rect 31352 5868 31585 5896
rect 31352 5856 31358 5868
rect 31573 5865 31585 5868
rect 31619 5865 31631 5899
rect 31573 5859 31631 5865
rect 31846 5856 31852 5908
rect 31904 5856 31910 5908
rect 33594 5856 33600 5908
rect 33652 5856 33658 5908
rect 30484 5800 31432 5828
rect 27157 5763 27215 5769
rect 26712 5732 26832 5760
rect 21269 5695 21327 5701
rect 21269 5661 21281 5695
rect 21315 5661 21327 5695
rect 21269 5655 21327 5661
rect 21453 5695 21511 5701
rect 21453 5661 21465 5695
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 21542 5652 21548 5704
rect 21600 5652 21606 5704
rect 21818 5652 21824 5704
rect 21876 5652 21882 5704
rect 21913 5695 21971 5701
rect 21913 5661 21925 5695
rect 21959 5661 21971 5695
rect 21913 5655 21971 5661
rect 14783 5596 14964 5624
rect 15028 5596 15608 5624
rect 15764 5596 16068 5624
rect 14783 5593 14795 5596
rect 14737 5587 14795 5593
rect 9916 5528 11560 5556
rect 14936 5556 14964 5596
rect 15378 5556 15384 5568
rect 14936 5528 15384 5556
rect 9916 5516 9922 5528
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 15473 5559 15531 5565
rect 15473 5525 15485 5559
rect 15519 5556 15531 5559
rect 15654 5556 15660 5568
rect 15519 5528 15660 5556
rect 15519 5525 15531 5528
rect 15473 5519 15531 5525
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 15764 5565 15792 5596
rect 16206 5584 16212 5636
rect 16264 5624 16270 5636
rect 17126 5624 17132 5636
rect 16264 5596 17132 5624
rect 16264 5584 16270 5596
rect 17126 5584 17132 5596
rect 17184 5584 17190 5636
rect 17402 5584 17408 5636
rect 17460 5624 17466 5636
rect 17589 5627 17647 5633
rect 17589 5624 17601 5627
rect 17460 5596 17601 5624
rect 17460 5584 17466 5596
rect 17589 5593 17601 5596
rect 17635 5624 17647 5627
rect 18414 5624 18420 5636
rect 17635 5596 18420 5624
rect 17635 5593 17647 5596
rect 17589 5587 17647 5593
rect 18414 5584 18420 5596
rect 18472 5624 18478 5636
rect 19058 5624 19064 5636
rect 18472 5596 19064 5624
rect 18472 5584 18478 5596
rect 19058 5584 19064 5596
rect 19116 5584 19122 5636
rect 19996 5624 20024 5652
rect 20441 5627 20499 5633
rect 20441 5624 20453 5627
rect 19996 5596 20453 5624
rect 20441 5593 20453 5596
rect 20487 5593 20499 5627
rect 20898 5624 20904 5636
rect 20441 5587 20499 5593
rect 20640 5596 20904 5624
rect 15749 5559 15807 5565
rect 15749 5525 15761 5559
rect 15795 5525 15807 5559
rect 15749 5519 15807 5525
rect 16758 5516 16764 5568
rect 16816 5556 16822 5568
rect 16853 5559 16911 5565
rect 16853 5556 16865 5559
rect 16816 5528 16865 5556
rect 16816 5516 16822 5528
rect 16853 5525 16865 5528
rect 16899 5525 16911 5559
rect 16853 5519 16911 5525
rect 19521 5559 19579 5565
rect 19521 5525 19533 5559
rect 19567 5556 19579 5559
rect 20640 5556 20668 5596
rect 20898 5584 20904 5596
rect 20956 5584 20962 5636
rect 21726 5624 21732 5636
rect 21560 5596 21732 5624
rect 19567 5528 20668 5556
rect 20809 5559 20867 5565
rect 19567 5525 19579 5528
rect 19521 5519 19579 5525
rect 20809 5525 20821 5559
rect 20855 5556 20867 5559
rect 21560 5556 21588 5596
rect 21726 5584 21732 5596
rect 21784 5584 21790 5636
rect 21928 5624 21956 5655
rect 22186 5652 22192 5704
rect 22244 5692 22250 5704
rect 23201 5695 23259 5701
rect 22244 5664 22287 5692
rect 22244 5652 22250 5664
rect 23201 5661 23213 5695
rect 23247 5661 23259 5695
rect 23201 5655 23259 5661
rect 23477 5695 23535 5701
rect 23477 5661 23489 5695
rect 23523 5692 23535 5695
rect 23658 5692 23664 5704
rect 23523 5664 23664 5692
rect 23523 5661 23535 5664
rect 23477 5655 23535 5661
rect 22002 5624 22008 5636
rect 21928 5596 22008 5624
rect 22002 5584 22008 5596
rect 22060 5584 22066 5636
rect 22278 5584 22284 5636
rect 22336 5624 22342 5636
rect 22830 5624 22836 5636
rect 22336 5596 22836 5624
rect 22336 5584 22342 5596
rect 22830 5584 22836 5596
rect 22888 5624 22894 5636
rect 23216 5624 23244 5655
rect 23658 5652 23664 5664
rect 23716 5652 23722 5704
rect 23842 5652 23848 5704
rect 23900 5652 23906 5704
rect 24673 5695 24731 5701
rect 24673 5661 24685 5695
rect 24719 5692 24731 5695
rect 24854 5692 24860 5704
rect 24719 5664 24860 5692
rect 24719 5661 24731 5664
rect 24673 5655 24731 5661
rect 24854 5652 24860 5664
rect 24912 5652 24918 5704
rect 25866 5652 25872 5704
rect 25924 5652 25930 5704
rect 25958 5652 25964 5704
rect 26016 5652 26022 5704
rect 26804 5701 26832 5732
rect 27157 5729 27169 5763
rect 27203 5760 27215 5763
rect 27522 5760 27528 5772
rect 27203 5732 27528 5760
rect 27203 5729 27215 5732
rect 27157 5723 27215 5729
rect 27522 5720 27528 5732
rect 27580 5760 27586 5772
rect 27580 5732 28028 5760
rect 27580 5720 27586 5732
rect 26237 5695 26295 5701
rect 26237 5661 26249 5695
rect 26283 5692 26295 5695
rect 26789 5695 26847 5701
rect 26283 5664 26740 5692
rect 26283 5661 26295 5664
rect 26237 5655 26295 5661
rect 22888 5596 23244 5624
rect 25976 5624 26004 5652
rect 26712 5636 26740 5664
rect 26789 5661 26801 5695
rect 26835 5692 26847 5695
rect 27246 5692 27252 5704
rect 26835 5664 27252 5692
rect 26835 5661 26847 5664
rect 26789 5655 26847 5661
rect 27246 5652 27252 5664
rect 27304 5652 27310 5704
rect 27617 5695 27675 5701
rect 27617 5661 27629 5695
rect 27663 5692 27675 5695
rect 27706 5692 27712 5704
rect 27663 5664 27712 5692
rect 27663 5661 27675 5664
rect 27617 5655 27675 5661
rect 27706 5652 27712 5664
rect 27764 5652 27770 5704
rect 28000 5701 28028 5732
rect 31018 5720 31024 5772
rect 31076 5726 31082 5772
rect 31404 5760 31432 5800
rect 31662 5788 31668 5840
rect 31720 5788 31726 5840
rect 31754 5788 31760 5840
rect 31812 5788 31818 5840
rect 31404 5732 31524 5760
rect 31076 5720 31340 5726
rect 27893 5695 27951 5701
rect 27893 5661 27905 5695
rect 27939 5661 27951 5695
rect 27893 5655 27951 5661
rect 27985 5695 28043 5701
rect 27985 5661 27997 5695
rect 28031 5661 28043 5695
rect 27985 5655 28043 5661
rect 26329 5627 26387 5633
rect 26329 5624 26341 5627
rect 25976 5596 26341 5624
rect 22888 5584 22894 5596
rect 26329 5593 26341 5596
rect 26375 5593 26387 5627
rect 26329 5587 26387 5593
rect 26694 5584 26700 5636
rect 26752 5584 26758 5636
rect 26973 5627 27031 5633
rect 26973 5593 26985 5627
rect 27019 5593 27031 5627
rect 26973 5587 27031 5593
rect 20855 5528 21588 5556
rect 21637 5559 21695 5565
rect 20855 5525 20867 5528
rect 20809 5519 20867 5525
rect 21637 5525 21649 5559
rect 21683 5556 21695 5559
rect 22186 5556 22192 5568
rect 21683 5528 22192 5556
rect 21683 5525 21695 5528
rect 21637 5519 21695 5525
rect 22186 5516 22192 5528
rect 22244 5516 22250 5568
rect 26421 5559 26479 5565
rect 26421 5525 26433 5559
rect 26467 5556 26479 5559
rect 26988 5556 27016 5587
rect 27430 5584 27436 5636
rect 27488 5624 27494 5636
rect 27908 5624 27936 5655
rect 28534 5652 28540 5704
rect 28592 5692 28598 5704
rect 29454 5692 29460 5704
rect 28592 5664 29460 5692
rect 28592 5652 28598 5664
rect 29454 5652 29460 5664
rect 29512 5692 29518 5704
rect 29549 5695 29607 5701
rect 29549 5692 29561 5695
rect 29512 5664 29561 5692
rect 29512 5652 29518 5664
rect 29549 5661 29561 5664
rect 29595 5661 29607 5695
rect 29549 5655 29607 5661
rect 29638 5652 29644 5704
rect 29696 5692 29702 5704
rect 31036 5701 31340 5720
rect 29805 5695 29863 5701
rect 31036 5698 31355 5701
rect 29805 5692 29817 5695
rect 29696 5664 29817 5692
rect 29696 5652 29702 5664
rect 29805 5661 29817 5664
rect 29851 5661 29863 5695
rect 29805 5655 29863 5661
rect 31297 5695 31355 5698
rect 31297 5661 31309 5695
rect 31343 5661 31355 5695
rect 31297 5655 31355 5661
rect 31389 5695 31447 5701
rect 31389 5661 31401 5695
rect 31435 5686 31447 5695
rect 31496 5686 31524 5732
rect 31680 5701 31708 5788
rect 31772 5701 31800 5788
rect 33689 5763 33747 5769
rect 33689 5729 33701 5763
rect 33735 5760 33747 5763
rect 34698 5760 34704 5772
rect 33735 5732 34704 5760
rect 33735 5729 33747 5732
rect 33689 5723 33747 5729
rect 34698 5720 34704 5732
rect 34756 5720 34762 5772
rect 31435 5661 31524 5686
rect 31389 5658 31524 5661
rect 31665 5695 31723 5701
rect 31665 5661 31677 5695
rect 31711 5661 31723 5695
rect 31389 5655 31447 5658
rect 31665 5655 31723 5661
rect 31757 5695 31815 5701
rect 31757 5661 31769 5695
rect 31803 5661 31815 5695
rect 31757 5655 31815 5661
rect 31938 5652 31944 5704
rect 31996 5692 32002 5704
rect 32125 5695 32183 5701
rect 32125 5692 32137 5695
rect 31996 5664 32137 5692
rect 31996 5652 32002 5664
rect 32125 5661 32137 5664
rect 32171 5661 32183 5695
rect 32125 5655 32183 5661
rect 32214 5652 32220 5704
rect 32272 5652 32278 5704
rect 32306 5652 32312 5704
rect 32364 5692 32370 5704
rect 32473 5695 32531 5701
rect 32473 5692 32485 5695
rect 32364 5664 32485 5692
rect 32364 5652 32370 5664
rect 32473 5661 32485 5664
rect 32519 5661 32531 5695
rect 32473 5655 32531 5661
rect 33965 5695 34023 5701
rect 33965 5661 33977 5695
rect 34011 5661 34023 5695
rect 33965 5655 34023 5661
rect 27488 5596 27936 5624
rect 27488 5584 27494 5596
rect 31846 5584 31852 5636
rect 31904 5584 31910 5636
rect 32232 5624 32260 5652
rect 33980 5624 34008 5655
rect 32232 5596 34008 5624
rect 26467 5528 27016 5556
rect 26467 5525 26479 5528
rect 26421 5519 26479 5525
rect 27798 5516 27804 5568
rect 27856 5556 27862 5568
rect 28077 5559 28135 5565
rect 28077 5556 28089 5559
rect 27856 5528 28089 5556
rect 27856 5516 27862 5528
rect 28077 5525 28089 5528
rect 28123 5525 28135 5559
rect 28077 5519 28135 5525
rect 30650 5516 30656 5568
rect 30708 5556 30714 5568
rect 30929 5559 30987 5565
rect 30929 5556 30941 5559
rect 30708 5528 30941 5556
rect 30708 5516 30714 5528
rect 30929 5525 30941 5528
rect 30975 5525 30987 5559
rect 30929 5519 30987 5525
rect 31110 5516 31116 5568
rect 31168 5516 31174 5568
rect 31202 5516 31208 5568
rect 31260 5556 31266 5568
rect 31941 5559 31999 5565
rect 31941 5556 31953 5559
rect 31260 5528 31953 5556
rect 31260 5516 31266 5528
rect 31941 5525 31953 5528
rect 31987 5525 31999 5559
rect 31941 5519 31999 5525
rect 1104 5466 36800 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 36800 5466
rect 1104 5392 36800 5414
rect 7653 5355 7711 5361
rect 7653 5321 7665 5355
rect 7699 5352 7711 5355
rect 8662 5352 8668 5364
rect 7699 5324 8668 5352
rect 7699 5321 7711 5324
rect 7653 5315 7711 5321
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 9217 5355 9275 5361
rect 9217 5321 9229 5355
rect 9263 5352 9275 5355
rect 9858 5352 9864 5364
rect 9263 5324 9864 5352
rect 9263 5321 9275 5324
rect 9217 5315 9275 5321
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 10505 5355 10563 5361
rect 10505 5352 10517 5355
rect 10008 5324 10517 5352
rect 10008 5312 10014 5324
rect 10505 5321 10517 5324
rect 10551 5321 10563 5355
rect 10505 5315 10563 5321
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12434 5352 12440 5364
rect 12299 5324 12440 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 12434 5312 12440 5324
rect 12492 5312 12498 5364
rect 12529 5355 12587 5361
rect 12529 5321 12541 5355
rect 12575 5352 12587 5355
rect 12618 5352 12624 5364
rect 12575 5324 12624 5352
rect 12575 5321 12587 5324
rect 12529 5315 12587 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 15378 5312 15384 5364
rect 15436 5352 15442 5364
rect 17310 5352 17316 5364
rect 15436 5324 17316 5352
rect 15436 5312 15442 5324
rect 14918 5244 14924 5296
rect 14976 5284 14982 5296
rect 15105 5287 15163 5293
rect 15105 5284 15117 5287
rect 14976 5256 15117 5284
rect 14976 5244 14982 5256
rect 15105 5253 15117 5256
rect 15151 5284 15163 5287
rect 15654 5284 15660 5296
rect 15151 5256 15660 5284
rect 15151 5253 15163 5256
rect 15105 5247 15163 5253
rect 15654 5244 15660 5256
rect 15712 5244 15718 5296
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5216 7527 5219
rect 7650 5216 7656 5228
rect 7515 5188 7656 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 7742 5176 7748 5228
rect 7800 5176 7806 5228
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 8352 5188 9413 5216
rect 8352 5176 8358 5188
rect 9401 5185 9413 5188
rect 9447 5185 9459 5219
rect 9401 5179 9459 5185
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 9732 5188 9873 5216
rect 9732 5176 9738 5188
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 11054 5216 11060 5228
rect 10091 5188 11060 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 11054 5176 11060 5188
rect 11112 5216 11118 5228
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 11112 5188 11529 5216
rect 11112 5176 11118 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5216 12495 5219
rect 12526 5216 12532 5228
rect 12483 5188 12532 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 16132 5225 16160 5324
rect 17310 5312 17316 5324
rect 17368 5352 17374 5364
rect 17497 5355 17555 5361
rect 17497 5352 17509 5355
rect 17368 5324 17509 5352
rect 17368 5312 17374 5324
rect 17497 5321 17509 5324
rect 17543 5321 17555 5355
rect 17497 5315 17555 5321
rect 19886 5312 19892 5364
rect 19944 5352 19950 5364
rect 19981 5355 20039 5361
rect 19981 5352 19993 5355
rect 19944 5324 19993 5352
rect 19944 5312 19950 5324
rect 19981 5321 19993 5324
rect 20027 5321 20039 5355
rect 20254 5352 20260 5364
rect 19981 5315 20039 5321
rect 20088 5324 20260 5352
rect 19702 5284 19708 5296
rect 16960 5256 19708 5284
rect 16960 5228 16988 5256
rect 19702 5244 19708 5256
rect 19760 5284 19766 5296
rect 20088 5284 20116 5324
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 21818 5312 21824 5364
rect 21876 5352 21882 5364
rect 22005 5355 22063 5361
rect 22005 5352 22017 5355
rect 21876 5324 22017 5352
rect 21876 5312 21882 5324
rect 22005 5321 22017 5324
rect 22051 5321 22063 5355
rect 22005 5315 22063 5321
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 22373 5355 22431 5361
rect 22373 5352 22385 5355
rect 22152 5324 22385 5352
rect 22152 5312 22158 5324
rect 22373 5321 22385 5324
rect 22419 5321 22431 5355
rect 22373 5315 22431 5321
rect 23477 5355 23535 5361
rect 23477 5321 23489 5355
rect 23523 5352 23535 5355
rect 23934 5352 23940 5364
rect 23523 5324 23940 5352
rect 23523 5321 23535 5324
rect 23477 5315 23535 5321
rect 23934 5312 23940 5324
rect 23992 5312 23998 5364
rect 25409 5355 25467 5361
rect 25409 5321 25421 5355
rect 25455 5352 25467 5355
rect 25958 5352 25964 5364
rect 25455 5324 25964 5352
rect 25455 5321 25467 5324
rect 25409 5315 25467 5321
rect 25958 5312 25964 5324
rect 26016 5312 26022 5364
rect 27430 5312 27436 5364
rect 27488 5312 27494 5364
rect 30837 5355 30895 5361
rect 30837 5321 30849 5355
rect 30883 5352 30895 5355
rect 31478 5352 31484 5364
rect 30883 5324 31484 5352
rect 30883 5321 30895 5324
rect 30837 5315 30895 5321
rect 31478 5312 31484 5324
rect 31536 5352 31542 5364
rect 31938 5352 31944 5364
rect 31536 5324 31944 5352
rect 31536 5312 31542 5324
rect 31938 5312 31944 5324
rect 31996 5312 32002 5364
rect 34149 5355 34207 5361
rect 34149 5352 34161 5355
rect 32324 5324 34161 5352
rect 19760 5256 20116 5284
rect 19760 5244 19766 5256
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5185 12771 5219
rect 12713 5179 12771 5185
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5216 14887 5219
rect 15749 5219 15807 5225
rect 15749 5216 15761 5219
rect 14875 5188 15761 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 15749 5185 15761 5188
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5148 12035 5151
rect 12728 5148 12756 5179
rect 12023 5120 12756 5148
rect 12023 5117 12035 5120
rect 11977 5111 12035 5117
rect 13078 5108 13084 5160
rect 13136 5148 13142 5160
rect 15010 5148 15016 5160
rect 13136 5120 15016 5148
rect 13136 5108 13142 5120
rect 15010 5108 15016 5120
rect 15068 5108 15074 5160
rect 15470 5108 15476 5160
rect 15528 5108 15534 5160
rect 15565 5151 15623 5157
rect 15565 5117 15577 5151
rect 15611 5148 15623 5151
rect 16132 5148 16160 5179
rect 16206 5176 16212 5228
rect 16264 5176 16270 5228
rect 16298 5176 16304 5228
rect 16356 5176 16362 5228
rect 16393 5219 16451 5225
rect 16393 5185 16405 5219
rect 16439 5216 16451 5219
rect 16758 5216 16764 5228
rect 16439 5188 16764 5216
rect 16439 5185 16451 5188
rect 16393 5179 16451 5185
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 16942 5176 16948 5228
rect 17000 5176 17006 5228
rect 17218 5176 17224 5228
rect 17276 5176 17282 5228
rect 17402 5176 17408 5228
rect 17460 5176 17466 5228
rect 17494 5176 17500 5228
rect 17552 5216 17558 5228
rect 18598 5216 18604 5228
rect 17552 5188 18604 5216
rect 17552 5176 17558 5188
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 19904 5225 19932 5256
rect 20162 5244 20168 5296
rect 20220 5244 20226 5296
rect 20622 5284 20628 5296
rect 20272 5256 20628 5284
rect 19797 5219 19855 5225
rect 19797 5185 19809 5219
rect 19843 5185 19855 5219
rect 19797 5179 19855 5185
rect 19889 5219 19947 5225
rect 19889 5185 19901 5219
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 15611 5120 16160 5148
rect 15611 5117 15623 5120
rect 15565 5111 15623 5117
rect 7374 5040 7380 5092
rect 7432 5080 7438 5092
rect 7469 5083 7527 5089
rect 7469 5080 7481 5083
rect 7432 5052 7481 5080
rect 7432 5040 7438 5052
rect 7469 5049 7481 5052
rect 7515 5049 7527 5083
rect 7469 5043 7527 5049
rect 9677 5083 9735 5089
rect 9677 5049 9689 5083
rect 9723 5080 9735 5083
rect 12250 5080 12256 5092
rect 9723 5052 12256 5080
rect 9723 5049 9735 5052
rect 9677 5043 9735 5049
rect 12250 5040 12256 5052
rect 12308 5040 12314 5092
rect 15488 5080 15516 5108
rect 16224 5080 16252 5176
rect 19812 5148 19840 5179
rect 19978 5176 19984 5228
rect 20036 5216 20042 5228
rect 20272 5225 20300 5256
rect 20622 5244 20628 5256
rect 20680 5244 20686 5296
rect 23845 5287 23903 5293
rect 23845 5253 23857 5287
rect 23891 5284 23903 5287
rect 24210 5284 24216 5296
rect 23891 5256 24216 5284
rect 23891 5253 23903 5256
rect 23845 5247 23903 5253
rect 24210 5244 24216 5256
rect 24268 5244 24274 5296
rect 27246 5244 27252 5296
rect 27304 5244 27310 5296
rect 30190 5244 30196 5296
rect 30248 5284 30254 5296
rect 31294 5284 31300 5296
rect 30248 5256 31300 5284
rect 30248 5244 30254 5256
rect 31294 5244 31300 5256
rect 31352 5244 31358 5296
rect 31757 5287 31815 5293
rect 31757 5253 31769 5287
rect 31803 5284 31815 5287
rect 32324 5284 32352 5324
rect 34149 5321 34161 5324
rect 34195 5352 34207 5355
rect 36538 5352 36544 5364
rect 34195 5324 36544 5352
rect 34195 5321 34207 5324
rect 34149 5315 34207 5321
rect 36538 5312 36544 5324
rect 36596 5312 36602 5364
rect 31803 5256 32352 5284
rect 31803 5253 31815 5256
rect 31757 5247 31815 5253
rect 20073 5219 20131 5225
rect 20073 5216 20085 5219
rect 20036 5188 20085 5216
rect 20036 5176 20042 5188
rect 20073 5185 20085 5188
rect 20119 5185 20131 5219
rect 20073 5179 20131 5185
rect 20257 5219 20315 5225
rect 20257 5185 20269 5219
rect 20303 5185 20315 5219
rect 20257 5179 20315 5185
rect 20438 5176 20444 5228
rect 20496 5216 20502 5228
rect 20533 5219 20591 5225
rect 20533 5216 20545 5219
rect 20496 5188 20545 5216
rect 20496 5176 20502 5188
rect 20533 5185 20545 5188
rect 20579 5216 20591 5219
rect 21542 5216 21548 5228
rect 20579 5188 21548 5216
rect 20579 5185 20591 5188
rect 20533 5179 20591 5185
rect 21542 5176 21548 5188
rect 21600 5176 21606 5228
rect 24854 5176 24860 5228
rect 24912 5216 24918 5228
rect 25225 5219 25283 5225
rect 25225 5216 25237 5219
rect 24912 5188 25237 5216
rect 24912 5176 24918 5188
rect 25225 5185 25237 5188
rect 25271 5185 25283 5219
rect 25225 5179 25283 5185
rect 27525 5219 27583 5225
rect 27525 5185 27537 5219
rect 27571 5216 27583 5219
rect 27798 5216 27804 5228
rect 27571 5188 27804 5216
rect 27571 5185 27583 5188
rect 27525 5179 27583 5185
rect 27798 5176 27804 5188
rect 27856 5176 27862 5228
rect 30650 5176 30656 5228
rect 30708 5216 30714 5228
rect 30745 5219 30803 5225
rect 30745 5216 30757 5219
rect 30708 5188 30757 5216
rect 30708 5176 30714 5188
rect 30745 5185 30757 5188
rect 30791 5185 30803 5219
rect 30745 5179 30803 5185
rect 32214 5176 32220 5228
rect 32272 5216 32278 5228
rect 32766 5216 32772 5228
rect 32272 5188 32772 5216
rect 32272 5176 32278 5188
rect 32766 5176 32772 5188
rect 32824 5176 32830 5228
rect 33025 5219 33083 5225
rect 33025 5216 33037 5219
rect 32876 5188 33037 5216
rect 19812 5120 20760 5148
rect 20088 5092 20116 5120
rect 15488 5052 16252 5080
rect 20070 5040 20076 5092
rect 20128 5040 20134 5092
rect 20732 5089 20760 5120
rect 22002 5108 22008 5160
rect 22060 5148 22066 5160
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 22060 5120 22477 5148
rect 22060 5108 22066 5120
rect 22465 5117 22477 5120
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 22646 5108 22652 5160
rect 22704 5108 22710 5160
rect 23934 5108 23940 5160
rect 23992 5108 23998 5160
rect 24118 5108 24124 5160
rect 24176 5108 24182 5160
rect 25041 5151 25099 5157
rect 25041 5117 25053 5151
rect 25087 5117 25099 5151
rect 25041 5111 25099 5117
rect 20717 5083 20775 5089
rect 20717 5049 20729 5083
rect 20763 5080 20775 5083
rect 21082 5080 21088 5092
rect 20763 5052 21088 5080
rect 20763 5049 20775 5052
rect 20717 5043 20775 5049
rect 21082 5040 21088 5052
rect 21140 5080 21146 5092
rect 22664 5080 22692 5108
rect 21140 5052 22692 5080
rect 25056 5080 25084 5111
rect 31110 5108 31116 5160
rect 31168 5148 31174 5160
rect 32876 5148 32904 5188
rect 33025 5185 33037 5188
rect 33071 5185 33083 5219
rect 33025 5179 33083 5185
rect 36170 5176 36176 5228
rect 36228 5176 36234 5228
rect 31168 5120 32904 5148
rect 31168 5108 31174 5120
rect 25682 5080 25688 5092
rect 25056 5052 25688 5080
rect 21140 5040 21146 5052
rect 25682 5040 25688 5052
rect 25740 5080 25746 5092
rect 25740 5052 31340 5080
rect 25740 5040 25746 5052
rect 31312 5024 31340 5052
rect 10226 4972 10232 5024
rect 10284 5012 10290 5024
rect 10321 5015 10379 5021
rect 10321 5012 10333 5015
rect 10284 4984 10333 5012
rect 10284 4972 10290 4984
rect 10321 4981 10333 4984
rect 10367 5012 10379 5015
rect 11790 5012 11796 5024
rect 10367 4984 11796 5012
rect 10367 4981 10379 4984
rect 10321 4975 10379 4981
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 15933 5015 15991 5021
rect 15933 4981 15945 5015
rect 15979 5012 15991 5015
rect 20438 5012 20444 5024
rect 15979 4984 20444 5012
rect 15979 4981 15991 4984
rect 15933 4975 15991 4981
rect 20438 4972 20444 4984
rect 20496 4972 20502 5024
rect 26234 4972 26240 5024
rect 26292 5012 26298 5024
rect 27249 5015 27307 5021
rect 27249 5012 27261 5015
rect 26292 4984 27261 5012
rect 26292 4972 26298 4984
rect 27249 4981 27261 4984
rect 27295 4981 27307 5015
rect 27249 4975 27307 4981
rect 31294 4972 31300 5024
rect 31352 5012 31358 5024
rect 31849 5015 31907 5021
rect 31849 5012 31861 5015
rect 31352 4984 31861 5012
rect 31352 4972 31358 4984
rect 31849 4981 31861 4984
rect 31895 4981 31907 5015
rect 31849 4975 31907 4981
rect 36354 4972 36360 5024
rect 36412 4972 36418 5024
rect 1104 4922 36800 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 36800 4922
rect 1104 4848 36800 4870
rect 10134 4768 10140 4820
rect 10192 4808 10198 4820
rect 18322 4808 18328 4820
rect 10192 4780 18328 4808
rect 10192 4768 10198 4780
rect 18322 4768 18328 4780
rect 18380 4768 18386 4820
rect 25038 4768 25044 4820
rect 25096 4808 25102 4820
rect 25501 4811 25559 4817
rect 25501 4808 25513 4811
rect 25096 4780 25513 4808
rect 25096 4768 25102 4780
rect 25501 4777 25513 4780
rect 25547 4777 25559 4811
rect 25501 4771 25559 4777
rect 27614 4768 27620 4820
rect 27672 4808 27678 4820
rect 28353 4811 28411 4817
rect 28353 4808 28365 4811
rect 27672 4780 28365 4808
rect 27672 4768 27678 4780
rect 28353 4777 28365 4780
rect 28399 4777 28411 4811
rect 28353 4771 28411 4777
rect 16758 4632 16764 4684
rect 16816 4672 16822 4684
rect 25056 4672 25084 4768
rect 25682 4740 25688 4752
rect 25148 4712 25688 4740
rect 25148 4681 25176 4712
rect 25682 4700 25688 4712
rect 25740 4700 25746 4752
rect 28258 4740 28264 4752
rect 27540 4712 28264 4740
rect 16816 4644 17264 4672
rect 16816 4632 16822 4644
rect 16942 4564 16948 4616
rect 17000 4564 17006 4616
rect 17236 4613 17264 4644
rect 22066 4644 25084 4672
rect 22066 4616 22094 4644
rect 17221 4607 17279 4613
rect 17221 4573 17233 4607
rect 17267 4573 17279 4607
rect 17221 4567 17279 4573
rect 21358 4564 21364 4616
rect 21416 4604 21422 4616
rect 22002 4604 22008 4616
rect 21416 4576 22008 4604
rect 21416 4564 21422 4576
rect 22002 4564 22008 4576
rect 22060 4576 22094 4616
rect 25056 4613 25084 4644
rect 25133 4675 25191 4681
rect 25133 4641 25145 4675
rect 25179 4641 25191 4675
rect 25133 4635 25191 4641
rect 25317 4675 25375 4681
rect 25317 4641 25329 4675
rect 25363 4672 25375 4675
rect 26694 4672 26700 4684
rect 25363 4644 26700 4672
rect 25363 4641 25375 4644
rect 25317 4635 25375 4641
rect 26694 4632 26700 4644
rect 26752 4632 26758 4684
rect 25041 4607 25099 4613
rect 22060 4564 22066 4576
rect 25041 4573 25053 4607
rect 25087 4604 25099 4607
rect 25222 4604 25228 4616
rect 25087 4576 25228 4604
rect 25087 4573 25099 4576
rect 25041 4567 25099 4573
rect 25222 4564 25228 4576
rect 25280 4564 25286 4616
rect 25501 4607 25559 4613
rect 25501 4604 25513 4607
rect 25424 4576 25513 4604
rect 16761 4539 16819 4545
rect 16761 4505 16773 4539
rect 16807 4536 16819 4539
rect 23842 4536 23848 4548
rect 16807 4508 23848 4536
rect 16807 4505 16819 4508
rect 16761 4499 16819 4505
rect 23842 4496 23848 4508
rect 23900 4496 23906 4548
rect 25424 4545 25452 4576
rect 25501 4573 25513 4576
rect 25547 4573 25559 4607
rect 25501 4567 25559 4573
rect 25682 4564 25688 4616
rect 25740 4564 25746 4616
rect 27246 4564 27252 4616
rect 27304 4604 27310 4616
rect 27540 4613 27568 4712
rect 28258 4700 28264 4712
rect 28316 4700 28322 4752
rect 28721 4743 28779 4749
rect 28721 4709 28733 4743
rect 28767 4709 28779 4743
rect 28721 4703 28779 4709
rect 27798 4632 27804 4684
rect 27856 4632 27862 4684
rect 28350 4632 28356 4684
rect 28408 4672 28414 4684
rect 28629 4675 28687 4681
rect 28629 4672 28641 4675
rect 28408 4644 28641 4672
rect 28408 4632 28414 4644
rect 28629 4641 28641 4644
rect 28675 4641 28687 4675
rect 28629 4635 28687 4641
rect 27525 4607 27583 4613
rect 27525 4604 27537 4607
rect 27304 4576 27537 4604
rect 27304 4564 27310 4576
rect 27525 4573 27537 4576
rect 27571 4573 27583 4607
rect 27525 4567 27583 4573
rect 27673 4607 27731 4613
rect 27673 4573 27685 4607
rect 27719 4604 27731 4607
rect 27816 4604 27844 4632
rect 27719 4576 27844 4604
rect 27990 4607 28048 4613
rect 27719 4573 27731 4576
rect 27673 4567 27731 4573
rect 27990 4573 28002 4607
rect 28036 4604 28048 4607
rect 28166 4604 28172 4616
rect 28036 4576 28172 4604
rect 28036 4573 28048 4576
rect 27990 4567 28048 4573
rect 25409 4539 25467 4545
rect 25409 4505 25421 4539
rect 25455 4505 25467 4539
rect 25409 4499 25467 4505
rect 15010 4428 15016 4480
rect 15068 4468 15074 4480
rect 17129 4471 17187 4477
rect 17129 4468 17141 4471
rect 15068 4440 17141 4468
rect 15068 4428 15074 4440
rect 17129 4437 17141 4440
rect 17175 4437 17187 4471
rect 17129 4431 17187 4437
rect 25038 4428 25044 4480
rect 25096 4468 25102 4480
rect 25424 4468 25452 4499
rect 27430 4496 27436 4548
rect 27488 4536 27494 4548
rect 27801 4539 27859 4545
rect 27801 4536 27813 4539
rect 27488 4508 27813 4536
rect 27488 4496 27494 4508
rect 27801 4505 27813 4508
rect 27847 4505 27859 4539
rect 27801 4499 27859 4505
rect 27890 4496 27896 4548
rect 27948 4496 27954 4548
rect 25096 4440 25452 4468
rect 25869 4471 25927 4477
rect 25096 4428 25102 4440
rect 25869 4437 25881 4471
rect 25915 4468 25927 4471
rect 26510 4468 26516 4480
rect 25915 4440 26516 4468
rect 25915 4437 25927 4440
rect 25869 4431 25927 4437
rect 26510 4428 26516 4440
rect 26568 4468 26574 4480
rect 28005 4468 28033 4567
rect 28166 4564 28172 4576
rect 28224 4564 28230 4616
rect 28258 4564 28264 4616
rect 28316 4564 28322 4616
rect 28442 4564 28448 4616
rect 28500 4604 28506 4616
rect 28537 4607 28595 4613
rect 28537 4604 28549 4607
rect 28500 4576 28549 4604
rect 28500 4564 28506 4576
rect 28537 4573 28549 4576
rect 28583 4573 28595 4607
rect 28736 4604 28764 4703
rect 31110 4700 31116 4752
rect 31168 4740 31174 4752
rect 31389 4743 31447 4749
rect 31389 4740 31401 4743
rect 31168 4712 31401 4740
rect 31168 4700 31174 4712
rect 31389 4709 31401 4712
rect 31435 4740 31447 4743
rect 31662 4740 31668 4752
rect 31435 4712 31668 4740
rect 31435 4709 31447 4712
rect 31389 4703 31447 4709
rect 31662 4700 31668 4712
rect 31720 4700 31726 4752
rect 29089 4607 29147 4613
rect 29089 4604 29101 4607
rect 28736 4576 29101 4604
rect 28537 4567 28595 4573
rect 29089 4573 29101 4576
rect 29135 4573 29147 4607
rect 29089 4567 29147 4573
rect 31205 4607 31263 4613
rect 31205 4573 31217 4607
rect 31251 4604 31263 4607
rect 31294 4604 31300 4616
rect 31251 4576 31300 4604
rect 31251 4573 31263 4576
rect 31205 4567 31263 4573
rect 31294 4564 31300 4576
rect 31352 4564 31358 4616
rect 28813 4539 28871 4545
rect 28813 4536 28825 4539
rect 28184 4508 28825 4536
rect 28184 4477 28212 4508
rect 28813 4505 28825 4508
rect 28859 4505 28871 4539
rect 28813 4499 28871 4505
rect 28994 4496 29000 4548
rect 29052 4496 29058 4548
rect 26568 4440 28033 4468
rect 28169 4471 28227 4477
rect 26568 4428 26574 4440
rect 28169 4437 28181 4471
rect 28215 4437 28227 4471
rect 28169 4431 28227 4437
rect 29089 4471 29147 4477
rect 29089 4437 29101 4471
rect 29135 4468 29147 4471
rect 29730 4468 29736 4480
rect 29135 4440 29736 4468
rect 29135 4437 29147 4440
rect 29089 4431 29147 4437
rect 29730 4428 29736 4440
rect 29788 4428 29794 4480
rect 1104 4378 36800 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 36800 4378
rect 1104 4304 36800 4326
rect 19426 4224 19432 4276
rect 19484 4264 19490 4276
rect 19978 4264 19984 4276
rect 19484 4236 19984 4264
rect 19484 4224 19490 4236
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 20073 4267 20131 4273
rect 20073 4233 20085 4267
rect 20119 4264 20131 4267
rect 21358 4264 21364 4276
rect 20119 4236 21364 4264
rect 20119 4233 20131 4236
rect 20073 4227 20131 4233
rect 21358 4224 21364 4236
rect 21416 4224 21422 4276
rect 22833 4267 22891 4273
rect 22833 4233 22845 4267
rect 22879 4264 22891 4267
rect 22922 4264 22928 4276
rect 22879 4236 22928 4264
rect 22879 4233 22891 4236
rect 22833 4227 22891 4233
rect 22922 4224 22928 4236
rect 22980 4224 22986 4276
rect 22741 4199 22799 4205
rect 18524 4168 18736 4196
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 6621 4131 6679 4137
rect 6621 4128 6633 4131
rect 5960 4100 6633 4128
rect 5960 4088 5966 4100
rect 6621 4097 6633 4100
rect 6667 4097 6679 4131
rect 6621 4091 6679 4097
rect 9122 4088 9128 4140
rect 9180 4128 9186 4140
rect 9565 4131 9623 4137
rect 9565 4128 9577 4131
rect 9180 4100 9577 4128
rect 9180 4088 9186 4100
rect 9565 4097 9577 4100
rect 9611 4097 9623 4131
rect 9565 4091 9623 4097
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 4120 4032 6377 4060
rect 4120 4020 4126 4032
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 6380 3924 6408 4023
rect 9306 4020 9312 4072
rect 9364 4020 9370 4072
rect 18524 4060 18552 4168
rect 18598 4088 18604 4140
rect 18656 4088 18662 4140
rect 18708 4128 18736 4168
rect 19904 4168 20116 4196
rect 19904 4128 19932 4168
rect 18708 4100 19932 4128
rect 20088 4128 20116 4168
rect 21744 4168 22140 4196
rect 21744 4128 21772 4168
rect 20088 4100 21772 4128
rect 21818 4088 21824 4140
rect 21876 4128 21882 4140
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 21876 4100 22017 4128
rect 21876 4088 21882 4100
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 22112 4128 22140 4168
rect 22741 4165 22753 4199
rect 22787 4196 22799 4199
rect 23474 4196 23480 4208
rect 22787 4168 23480 4196
rect 22787 4165 22799 4168
rect 22741 4159 22799 4165
rect 23474 4156 23480 4168
rect 23532 4156 23538 4208
rect 27890 4196 27896 4208
rect 26712 4168 27896 4196
rect 26712 4140 26740 4168
rect 27890 4156 27896 4168
rect 27948 4196 27954 4208
rect 28442 4196 28448 4208
rect 27948 4168 28448 4196
rect 27948 4156 27954 4168
rect 28442 4156 28448 4168
rect 28500 4156 28506 4208
rect 30558 4196 30564 4208
rect 30392 4168 30564 4196
rect 23934 4128 23940 4140
rect 22112 4100 23940 4128
rect 22005 4091 22063 4097
rect 23934 4088 23940 4100
rect 23992 4088 23998 4140
rect 25038 4088 25044 4140
rect 25096 4088 25102 4140
rect 25222 4088 25228 4140
rect 25280 4088 25286 4140
rect 25317 4131 25375 4137
rect 25317 4097 25329 4131
rect 25363 4128 25375 4131
rect 25682 4128 25688 4140
rect 25363 4100 25688 4128
rect 25363 4097 25375 4100
rect 25317 4091 25375 4097
rect 25682 4088 25688 4100
rect 25740 4088 25746 4140
rect 26234 4088 26240 4140
rect 26292 4088 26298 4140
rect 26421 4131 26479 4137
rect 26421 4097 26433 4131
rect 26467 4097 26479 4131
rect 26421 4091 26479 4097
rect 10704 4032 18552 4060
rect 9324 3992 9352 4020
rect 10704 4001 10732 4032
rect 18690 4020 18696 4072
rect 18748 4020 18754 4072
rect 18877 4063 18935 4069
rect 18877 4029 18889 4063
rect 18923 4060 18935 4063
rect 19334 4060 19340 4072
rect 18923 4032 19340 4060
rect 18923 4029 18935 4032
rect 18877 4023 18935 4029
rect 19334 4020 19340 4032
rect 19392 4060 19398 4072
rect 20257 4063 20315 4069
rect 20257 4060 20269 4063
rect 19392 4032 20269 4060
rect 19392 4020 19398 4032
rect 20257 4029 20269 4032
rect 20303 4060 20315 4063
rect 22462 4060 22468 4072
rect 20303 4032 22468 4060
rect 20303 4029 20315 4032
rect 20257 4023 20315 4029
rect 22462 4020 22468 4032
rect 22520 4060 22526 4072
rect 22925 4063 22983 4069
rect 22925 4060 22937 4063
rect 22520 4032 22937 4060
rect 22520 4020 22526 4032
rect 22925 4029 22937 4032
rect 22971 4029 22983 4063
rect 26436 4060 26464 4091
rect 26510 4088 26516 4140
rect 26568 4088 26574 4140
rect 26694 4088 26700 4140
rect 26752 4088 26758 4140
rect 30282 4088 30288 4140
rect 30340 4088 30346 4140
rect 30392 4137 30420 4168
rect 30558 4156 30564 4168
rect 30616 4196 30622 4208
rect 31110 4196 31116 4208
rect 30616 4168 31116 4196
rect 30616 4156 30622 4168
rect 31110 4156 31116 4168
rect 31168 4156 31174 4208
rect 30377 4131 30435 4137
rect 30377 4097 30389 4131
rect 30423 4097 30435 4131
rect 30377 4091 30435 4097
rect 30469 4131 30527 4137
rect 30469 4097 30481 4131
rect 30515 4128 30527 4131
rect 30837 4131 30895 4137
rect 30515 4100 30788 4128
rect 30515 4097 30527 4100
rect 30469 4091 30527 4097
rect 26602 4060 26608 4072
rect 22925 4023 22983 4029
rect 24780 4032 26372 4060
rect 26436 4032 26608 4060
rect 7300 3964 9352 3992
rect 10689 3995 10747 4001
rect 7300 3924 7328 3964
rect 10689 3961 10701 3995
rect 10735 3961 10747 3995
rect 24780 3992 24808 4032
rect 10689 3955 10747 3961
rect 12406 3964 24808 3992
rect 24857 3995 24915 4001
rect 6380 3896 7328 3924
rect 7745 3927 7803 3933
rect 7745 3893 7757 3927
rect 7791 3924 7803 3927
rect 12406 3924 12434 3964
rect 24857 3961 24869 3995
rect 24903 3992 24915 3995
rect 25961 3995 26019 4001
rect 25961 3992 25973 3995
rect 24903 3964 25973 3992
rect 24903 3961 24915 3964
rect 24857 3955 24915 3961
rect 25961 3961 25973 3964
rect 26007 3961 26019 3995
rect 26344 3992 26372 4032
rect 26602 4020 26608 4032
rect 26660 4020 26666 4072
rect 30561 4063 30619 4069
rect 30561 4029 30573 4063
rect 30607 4029 30619 4063
rect 30760 4060 30788 4100
rect 30837 4097 30849 4131
rect 30883 4128 30895 4131
rect 30926 4128 30932 4140
rect 30883 4100 30932 4128
rect 30883 4097 30895 4100
rect 30837 4091 30895 4097
rect 30926 4088 30932 4100
rect 30984 4088 30990 4140
rect 31021 4063 31079 4069
rect 31021 4060 31033 4063
rect 30760 4032 31033 4060
rect 30561 4023 30619 4029
rect 31021 4029 31033 4032
rect 31067 4060 31079 4063
rect 31202 4060 31208 4072
rect 31067 4032 31208 4060
rect 31067 4029 31079 4032
rect 31021 4023 31079 4029
rect 27982 3992 27988 4004
rect 26344 3964 27988 3992
rect 25961 3955 26019 3961
rect 27982 3952 27988 3964
rect 28040 3952 28046 4004
rect 30374 3952 30380 4004
rect 30432 3992 30438 4004
rect 30576 3992 30604 4023
rect 31202 4020 31208 4032
rect 31260 4020 31266 4072
rect 30432 3964 30604 3992
rect 30432 3952 30438 3964
rect 7791 3896 12434 3924
rect 7791 3893 7803 3896
rect 7745 3887 7803 3893
rect 18230 3884 18236 3936
rect 18288 3884 18294 3936
rect 19610 3884 19616 3936
rect 19668 3884 19674 3936
rect 21542 3884 21548 3936
rect 21600 3924 21606 3936
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 21600 3896 21833 3924
rect 21600 3884 21606 3896
rect 21821 3893 21833 3896
rect 21867 3893 21879 3927
rect 21821 3887 21879 3893
rect 22373 3927 22431 3933
rect 22373 3893 22385 3927
rect 22419 3924 22431 3927
rect 22830 3924 22836 3936
rect 22419 3896 22836 3924
rect 22419 3893 22431 3896
rect 22373 3887 22431 3893
rect 22830 3884 22836 3896
rect 22888 3884 22894 3936
rect 26142 3884 26148 3936
rect 26200 3924 26206 3936
rect 26237 3927 26295 3933
rect 26237 3924 26249 3927
rect 26200 3896 26249 3924
rect 26200 3884 26206 3896
rect 26237 3893 26249 3896
rect 26283 3893 26295 3927
rect 26237 3887 26295 3893
rect 30101 3927 30159 3933
rect 30101 3893 30113 3927
rect 30147 3924 30159 3927
rect 30742 3924 30748 3936
rect 30147 3896 30748 3924
rect 30147 3893 30159 3896
rect 30101 3887 30159 3893
rect 30742 3884 30748 3896
rect 30800 3884 30806 3936
rect 1104 3834 36800 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 36800 3834
rect 1104 3760 36800 3782
rect 18690 3680 18696 3732
rect 18748 3720 18754 3732
rect 18748 3692 20208 3720
rect 18748 3680 18754 3692
rect 19242 3584 19248 3596
rect 18432 3556 19248 3584
rect 15749 3519 15807 3525
rect 15749 3485 15761 3519
rect 15795 3516 15807 3519
rect 16574 3516 16580 3528
rect 15795 3488 16580 3516
rect 15795 3485 15807 3488
rect 15749 3479 15807 3485
rect 16574 3476 16580 3488
rect 16632 3516 16638 3528
rect 17586 3516 17592 3528
rect 16632 3488 17592 3516
rect 16632 3476 16638 3488
rect 17586 3476 17592 3488
rect 17644 3476 17650 3528
rect 17681 3519 17739 3525
rect 17681 3485 17693 3519
rect 17727 3485 17739 3519
rect 17681 3479 17739 3485
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3516 17831 3519
rect 17819 3488 18000 3516
rect 17819 3485 17831 3488
rect 17773 3479 17831 3485
rect 16016 3451 16074 3457
rect 16016 3417 16028 3451
rect 16062 3448 16074 3451
rect 16206 3448 16212 3460
rect 16062 3420 16212 3448
rect 16062 3417 16074 3420
rect 16016 3411 16074 3417
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 17126 3340 17132 3392
rect 17184 3340 17190 3392
rect 17494 3340 17500 3392
rect 17552 3340 17558 3392
rect 17688 3380 17716 3479
rect 17972 3448 18000 3488
rect 18046 3476 18052 3528
rect 18104 3476 18110 3528
rect 18432 3516 18460 3556
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 20180 3584 20208 3692
rect 22002 3680 22008 3732
rect 22060 3720 22066 3732
rect 22281 3723 22339 3729
rect 22281 3720 22293 3723
rect 22060 3692 22293 3720
rect 22060 3680 22066 3692
rect 22281 3689 22293 3692
rect 22327 3689 22339 3723
rect 22281 3683 22339 3689
rect 23474 3680 23480 3732
rect 23532 3720 23538 3732
rect 24486 3720 24492 3732
rect 23532 3692 24492 3720
rect 23532 3680 23538 3692
rect 24486 3680 24492 3692
rect 24544 3680 24550 3732
rect 30282 3720 30288 3732
rect 26068 3692 30288 3720
rect 20898 3584 20904 3596
rect 20180 3556 20904 3584
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 21082 3544 21088 3596
rect 21140 3544 21146 3596
rect 22094 3544 22100 3596
rect 22152 3584 22158 3596
rect 22465 3587 22523 3593
rect 22465 3584 22477 3587
rect 22152 3556 22477 3584
rect 22152 3544 22158 3556
rect 22465 3553 22477 3556
rect 22511 3553 22523 3587
rect 22465 3547 22523 3553
rect 18248 3488 18460 3516
rect 18248 3448 18276 3488
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 19484 3488 19533 3516
rect 19484 3476 19490 3488
rect 19521 3485 19533 3488
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 19978 3476 19984 3528
rect 20036 3516 20042 3528
rect 20349 3519 20407 3525
rect 20349 3516 20361 3519
rect 20036 3488 20361 3516
rect 20036 3476 20042 3488
rect 20349 3485 20361 3488
rect 20395 3485 20407 3519
rect 20349 3479 20407 3485
rect 20530 3476 20536 3528
rect 20588 3516 20594 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 20588 3488 21281 3516
rect 20588 3476 20594 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 21542 3476 21548 3528
rect 21600 3476 21606 3528
rect 22646 3476 22652 3528
rect 22704 3516 22710 3528
rect 22741 3519 22799 3525
rect 22741 3516 22753 3519
rect 22704 3488 22753 3516
rect 22704 3476 22710 3488
rect 22741 3485 22753 3488
rect 22787 3485 22799 3519
rect 22741 3479 22799 3485
rect 25682 3476 25688 3528
rect 25740 3516 25746 3528
rect 25869 3519 25927 3525
rect 25869 3516 25881 3519
rect 25740 3488 25881 3516
rect 25740 3476 25746 3488
rect 25869 3485 25881 3488
rect 25915 3485 25927 3519
rect 25869 3479 25927 3485
rect 25958 3476 25964 3528
rect 26016 3476 26022 3528
rect 17972 3420 18276 3448
rect 18322 3408 18328 3460
rect 18380 3448 18386 3460
rect 26068 3448 26096 3692
rect 30282 3680 30288 3692
rect 30340 3680 30346 3732
rect 30374 3680 30380 3732
rect 30432 3720 30438 3732
rect 31294 3720 31300 3732
rect 30432 3692 31300 3720
rect 30432 3680 30438 3692
rect 31294 3680 31300 3692
rect 31352 3680 31358 3732
rect 31846 3680 31852 3732
rect 31904 3720 31910 3732
rect 34149 3723 34207 3729
rect 34149 3720 34161 3723
rect 31904 3692 34161 3720
rect 31904 3680 31910 3692
rect 34149 3689 34161 3692
rect 34195 3720 34207 3723
rect 36078 3720 36084 3732
rect 34195 3692 36084 3720
rect 34195 3689 34207 3692
rect 34149 3683 34207 3689
rect 36078 3680 36084 3692
rect 36136 3680 36142 3732
rect 26881 3655 26939 3661
rect 26881 3621 26893 3655
rect 26927 3652 26939 3655
rect 28445 3655 28503 3661
rect 26927 3624 28212 3652
rect 26927 3621 26939 3624
rect 26881 3615 26939 3621
rect 26142 3544 26148 3596
rect 26200 3544 26206 3596
rect 26234 3544 26240 3596
rect 26292 3584 26298 3596
rect 26973 3587 27031 3593
rect 26292 3556 26832 3584
rect 26292 3544 26298 3556
rect 26510 3476 26516 3528
rect 26568 3476 26574 3528
rect 26602 3476 26608 3528
rect 26660 3516 26666 3528
rect 26804 3525 26832 3556
rect 26973 3553 26985 3587
rect 27019 3584 27031 3587
rect 27522 3584 27528 3596
rect 27019 3556 27528 3584
rect 27019 3553 27031 3556
rect 26973 3547 27031 3553
rect 27522 3544 27528 3556
rect 27580 3544 27586 3596
rect 26697 3519 26755 3525
rect 26697 3516 26709 3519
rect 26660 3488 26709 3516
rect 26660 3476 26666 3488
rect 26697 3485 26709 3488
rect 26743 3485 26755 3519
rect 26697 3479 26755 3485
rect 26789 3519 26847 3525
rect 26789 3485 26801 3519
rect 26835 3485 26847 3519
rect 26789 3479 26847 3485
rect 27062 3476 27068 3528
rect 27120 3476 27126 3528
rect 28184 3525 28212 3624
rect 28445 3621 28457 3655
rect 28491 3652 28503 3655
rect 32214 3652 32220 3664
rect 28491 3624 32220 3652
rect 28491 3621 28503 3624
rect 28445 3615 28503 3621
rect 32214 3612 32220 3624
rect 32272 3612 32278 3664
rect 30101 3587 30159 3593
rect 30101 3553 30113 3587
rect 30147 3584 30159 3587
rect 30466 3584 30472 3596
rect 30147 3556 30472 3584
rect 30147 3553 30159 3556
rect 30101 3547 30159 3553
rect 30466 3544 30472 3556
rect 30524 3544 30530 3596
rect 30742 3544 30748 3596
rect 30800 3584 30806 3596
rect 31573 3587 31631 3593
rect 31573 3584 31585 3587
rect 30800 3556 31585 3584
rect 30800 3544 30806 3556
rect 31573 3553 31585 3556
rect 31619 3553 31631 3587
rect 31573 3547 31631 3553
rect 31662 3544 31668 3596
rect 31720 3584 31726 3596
rect 32309 3587 32367 3593
rect 31720 3556 31800 3584
rect 31720 3544 31726 3556
rect 28169 3519 28227 3525
rect 28169 3485 28181 3519
rect 28215 3485 28227 3519
rect 28445 3519 28503 3525
rect 28445 3516 28457 3519
rect 28169 3479 28227 3485
rect 28276 3488 28457 3516
rect 18380 3420 26096 3448
rect 26145 3451 26203 3457
rect 18380 3408 18386 3420
rect 26145 3417 26157 3451
rect 26191 3448 26203 3451
rect 28276 3448 28304 3488
rect 28445 3485 28457 3488
rect 28491 3485 28503 3519
rect 28445 3479 28503 3485
rect 29730 3519 29788 3525
rect 29730 3485 29742 3519
rect 29776 3516 29788 3519
rect 29822 3516 29828 3528
rect 29776 3488 29828 3516
rect 29776 3485 29788 3488
rect 29730 3479 29788 3485
rect 29822 3476 29828 3488
rect 29880 3476 29886 3528
rect 30190 3476 30196 3528
rect 30248 3476 30254 3528
rect 30834 3476 30840 3528
rect 30892 3476 30898 3528
rect 30926 3476 30932 3528
rect 30984 3476 30990 3528
rect 31294 3476 31300 3528
rect 31352 3476 31358 3528
rect 31386 3476 31392 3528
rect 31444 3476 31450 3528
rect 31478 3476 31484 3528
rect 31536 3476 31542 3528
rect 31772 3525 31800 3556
rect 32309 3553 32321 3587
rect 32355 3584 32367 3587
rect 32355 3556 32904 3584
rect 32355 3553 32367 3556
rect 32309 3547 32367 3553
rect 31757 3519 31815 3525
rect 31757 3485 31769 3519
rect 31803 3485 31815 3519
rect 31757 3479 31815 3485
rect 31846 3476 31852 3528
rect 31904 3476 31910 3528
rect 31941 3519 31999 3525
rect 31941 3485 31953 3519
rect 31987 3516 31999 3519
rect 32140 3516 32352 3518
rect 32398 3516 32404 3528
rect 31987 3490 32404 3516
rect 31987 3488 32168 3490
rect 32324 3488 32404 3490
rect 31987 3485 31999 3488
rect 31941 3479 31999 3485
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 32498 3497 32556 3503
rect 26191 3420 28304 3448
rect 28353 3451 28411 3457
rect 26191 3417 26203 3420
rect 26145 3411 26203 3417
rect 28353 3417 28365 3451
rect 28399 3448 28411 3451
rect 28994 3448 29000 3460
rect 28399 3420 29000 3448
rect 28399 3417 28411 3420
rect 28353 3411 28411 3417
rect 28994 3408 29000 3420
rect 29052 3408 29058 3460
rect 30852 3448 30880 3476
rect 32498 3463 32510 3497
rect 32544 3463 32556 3497
rect 32766 3476 32772 3528
rect 32824 3476 32830 3528
rect 32876 3516 32904 3556
rect 33025 3519 33083 3525
rect 33025 3516 33037 3519
rect 32876 3488 33037 3516
rect 33025 3485 33037 3488
rect 33071 3485 33083 3519
rect 33025 3479 33083 3485
rect 29472 3420 29868 3448
rect 18230 3380 18236 3392
rect 17688 3352 18236 3380
rect 18230 3340 18236 3352
rect 18288 3340 18294 3392
rect 18598 3340 18604 3392
rect 18656 3380 18662 3392
rect 18785 3383 18843 3389
rect 18785 3380 18797 3383
rect 18656 3352 18797 3380
rect 18656 3340 18662 3352
rect 18785 3349 18797 3352
rect 18831 3349 18843 3383
rect 18785 3343 18843 3349
rect 20070 3340 20076 3392
rect 20128 3380 20134 3392
rect 20441 3383 20499 3389
rect 20441 3380 20453 3383
rect 20128 3352 20453 3380
rect 20128 3340 20134 3352
rect 20441 3349 20453 3352
rect 20487 3349 20499 3383
rect 20441 3343 20499 3349
rect 20806 3340 20812 3392
rect 20864 3340 20870 3392
rect 20898 3340 20904 3392
rect 20956 3380 20962 3392
rect 23382 3380 23388 3392
rect 20956 3352 23388 3380
rect 20956 3340 20962 3352
rect 23382 3340 23388 3352
rect 23440 3340 23446 3392
rect 25130 3340 25136 3392
rect 25188 3380 25194 3392
rect 29472 3380 29500 3420
rect 25188 3352 29500 3380
rect 25188 3340 25194 3352
rect 29546 3340 29552 3392
rect 29604 3340 29610 3392
rect 29730 3340 29736 3392
rect 29788 3340 29794 3392
rect 29840 3380 29868 3420
rect 30576 3420 30880 3448
rect 30576 3380 30604 3420
rect 31570 3408 31576 3460
rect 31628 3448 31634 3460
rect 32125 3451 32183 3457
rect 32125 3448 32137 3451
rect 31628 3420 32137 3448
rect 31628 3408 31634 3420
rect 32125 3417 32137 3420
rect 32171 3417 32183 3451
rect 32125 3411 32183 3417
rect 32214 3408 32220 3460
rect 32272 3448 32278 3460
rect 32498 3457 32556 3463
rect 32309 3451 32367 3457
rect 32309 3448 32321 3451
rect 32272 3420 32321 3448
rect 32272 3408 32278 3420
rect 32309 3417 32321 3420
rect 32355 3417 32367 3451
rect 32309 3411 32367 3417
rect 29840 3352 30604 3380
rect 30650 3340 30656 3392
rect 30708 3340 30714 3392
rect 31110 3340 31116 3392
rect 31168 3340 31174 3392
rect 31202 3340 31208 3392
rect 31260 3340 31266 3392
rect 31294 3340 31300 3392
rect 31352 3380 31358 3392
rect 31665 3383 31723 3389
rect 31665 3380 31677 3383
rect 31352 3352 31677 3380
rect 31352 3340 31358 3352
rect 31665 3349 31677 3352
rect 31711 3349 31723 3383
rect 31665 3343 31723 3349
rect 31754 3340 31760 3392
rect 31812 3380 31818 3392
rect 32508 3380 32536 3457
rect 31812 3352 32536 3380
rect 31812 3340 31818 3352
rect 1104 3290 36800 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 36800 3290
rect 1104 3216 36800 3238
rect 1397 3179 1455 3185
rect 1397 3145 1409 3179
rect 1443 3145 1455 3179
rect 1397 3139 1455 3145
rect 1412 3108 1440 3139
rect 16206 3136 16212 3188
rect 16264 3136 16270 3188
rect 17037 3179 17095 3185
rect 17037 3145 17049 3179
rect 17083 3176 17095 3179
rect 18598 3176 18604 3188
rect 17083 3148 18604 3176
rect 17083 3145 17095 3148
rect 17037 3139 17095 3145
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 18690 3136 18696 3188
rect 18748 3176 18754 3188
rect 18969 3179 19027 3185
rect 18969 3176 18981 3179
rect 18748 3148 18981 3176
rect 18748 3136 18754 3148
rect 18969 3145 18981 3148
rect 19015 3145 19027 3179
rect 18969 3139 19027 3145
rect 19426 3136 19432 3188
rect 19484 3136 19490 3188
rect 19889 3179 19947 3185
rect 19889 3145 19901 3179
rect 19935 3145 19947 3179
rect 19889 3139 19947 3145
rect 3114 3111 3172 3117
rect 3114 3108 3126 3111
rect 1412 3080 3126 3108
rect 3114 3077 3126 3080
rect 3160 3077 3172 3111
rect 3114 3071 3172 3077
rect 16022 3068 16028 3120
rect 16080 3108 16086 3120
rect 17126 3108 17132 3120
rect 16080 3080 17132 3108
rect 16080 3068 16086 3080
rect 17126 3068 17132 3080
rect 17184 3068 17190 3120
rect 17770 3108 17776 3120
rect 17328 3080 17776 3108
rect 934 3000 940 3052
rect 992 3040 998 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 992 3012 1593 3040
rect 992 3000 998 3012
rect 1581 3009 1593 3012
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 4062 3040 4068 3052
rect 2915 3012 4068 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 16393 3043 16451 3049
rect 16393 3009 16405 3043
rect 16439 3040 16451 3043
rect 16439 3012 16712 3040
rect 16439 3009 16451 3012
rect 16393 3003 16451 3009
rect 4246 2864 4252 2916
rect 4304 2864 4310 2916
rect 16684 2913 16712 3012
rect 17328 2981 17356 3080
rect 17770 3068 17776 3080
rect 17828 3068 17834 3120
rect 19904 3108 19932 3139
rect 20806 3136 20812 3188
rect 20864 3176 20870 3188
rect 21177 3179 21235 3185
rect 21177 3176 21189 3179
rect 20864 3148 21189 3176
rect 20864 3136 20870 3148
rect 21177 3145 21189 3148
rect 21223 3145 21235 3179
rect 21177 3139 21235 3145
rect 21818 3136 21824 3188
rect 21876 3136 21882 3188
rect 22002 3136 22008 3188
rect 22060 3176 22066 3188
rect 22189 3179 22247 3185
rect 22189 3176 22201 3179
rect 22060 3148 22201 3176
rect 22060 3136 22066 3148
rect 22189 3145 22201 3148
rect 22235 3145 22247 3179
rect 22189 3139 22247 3145
rect 22646 3136 22652 3188
rect 22704 3136 22710 3188
rect 24765 3179 24823 3185
rect 24765 3145 24777 3179
rect 24811 3176 24823 3179
rect 25038 3176 25044 3188
rect 24811 3148 25044 3176
rect 24811 3145 24823 3148
rect 24765 3139 24823 3145
rect 25038 3136 25044 3148
rect 25096 3136 25102 3188
rect 25409 3179 25467 3185
rect 25409 3145 25421 3179
rect 25455 3145 25467 3179
rect 25409 3139 25467 3145
rect 19904 3080 20484 3108
rect 17586 3000 17592 3052
rect 17644 3000 17650 3052
rect 17856 3043 17914 3049
rect 17856 3009 17868 3043
rect 17902 3040 17914 3043
rect 18138 3040 18144 3052
rect 17902 3012 18144 3040
rect 17902 3009 17914 3012
rect 17856 3003 17914 3009
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 19610 3000 19616 3052
rect 19668 3000 19674 3052
rect 20070 3000 20076 3052
rect 20128 3000 20134 3052
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3040 20223 3043
rect 20346 3040 20352 3052
rect 20211 3012 20352 3040
rect 20211 3009 20223 3012
rect 20165 3003 20223 3009
rect 17313 2975 17371 2981
rect 17313 2941 17325 2975
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 20180 2972 20208 3003
rect 20346 3000 20352 3012
rect 20404 3000 20410 3052
rect 20456 3049 20484 3080
rect 23382 3068 23388 3120
rect 23440 3108 23446 3120
rect 25424 3108 25452 3139
rect 25682 3136 25688 3188
rect 25740 3136 25746 3188
rect 26142 3136 26148 3188
rect 26200 3136 26206 3188
rect 26973 3179 27031 3185
rect 26973 3145 26985 3179
rect 27019 3176 27031 3179
rect 27062 3176 27068 3188
rect 27019 3148 27068 3176
rect 27019 3145 27031 3148
rect 26973 3139 27031 3145
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 27522 3136 27528 3188
rect 27580 3136 27586 3188
rect 30466 3176 30472 3188
rect 28460 3148 30472 3176
rect 26160 3108 26188 3136
rect 23440 3080 25084 3108
rect 25424 3080 27200 3108
rect 23440 3068 23446 3080
rect 20441 3043 20499 3049
rect 20441 3009 20453 3043
rect 20487 3009 20499 3043
rect 20441 3003 20499 3009
rect 22066 3012 22416 3040
rect 19392 2944 20208 2972
rect 19392 2932 19398 2944
rect 21082 2932 21088 2984
rect 21140 2972 21146 2984
rect 22066 2972 22094 3012
rect 22388 2981 22416 3012
rect 22830 3000 22836 3052
rect 22888 3000 22894 3052
rect 23934 3000 23940 3052
rect 23992 3040 23998 3052
rect 25056 3049 25084 3080
rect 25884 3049 25912 3080
rect 24397 3043 24455 3049
rect 24397 3040 24409 3043
rect 23992 3012 24409 3040
rect 23992 3000 23998 3012
rect 24397 3009 24409 3012
rect 24443 3009 24455 3043
rect 24397 3003 24455 3009
rect 25041 3043 25099 3049
rect 25041 3009 25053 3043
rect 25087 3009 25099 3043
rect 25041 3003 25099 3009
rect 25869 3043 25927 3049
rect 25869 3009 25881 3043
rect 25915 3009 25927 3043
rect 25869 3003 25927 3009
rect 26050 3000 26056 3052
rect 26108 3040 26114 3052
rect 26145 3043 26203 3049
rect 26145 3040 26157 3043
rect 26108 3012 26157 3040
rect 26108 3000 26114 3012
rect 26145 3009 26157 3012
rect 26191 3009 26203 3043
rect 26145 3003 26203 3009
rect 21140 2944 22094 2972
rect 22281 2975 22339 2981
rect 21140 2932 21146 2944
rect 22281 2941 22293 2975
rect 22327 2941 22339 2975
rect 22281 2935 22339 2941
rect 22373 2975 22431 2981
rect 22373 2941 22385 2975
rect 22419 2941 22431 2975
rect 22373 2935 22431 2941
rect 16669 2907 16727 2913
rect 16669 2873 16681 2907
rect 16715 2873 16727 2907
rect 22296 2904 22324 2935
rect 24302 2932 24308 2984
rect 24360 2932 24366 2984
rect 25130 2932 25136 2984
rect 25188 2932 25194 2984
rect 22922 2904 22928 2916
rect 22296 2876 22928 2904
rect 16669 2867 16727 2873
rect 22922 2864 22928 2876
rect 22980 2904 22986 2916
rect 24121 2907 24179 2913
rect 24121 2904 24133 2907
rect 22980 2876 24133 2904
rect 22980 2864 22986 2876
rect 24121 2873 24133 2876
rect 24167 2904 24179 2907
rect 25314 2904 25320 2916
rect 24167 2876 25320 2904
rect 24167 2873 24179 2876
rect 24121 2867 24179 2873
rect 25314 2864 25320 2876
rect 25372 2864 25378 2916
rect 26160 2904 26188 3003
rect 26234 3000 26240 3052
rect 26292 3040 26298 3052
rect 27172 3049 27200 3080
rect 26329 3043 26387 3049
rect 26329 3040 26341 3043
rect 26292 3012 26341 3040
rect 26292 3000 26298 3012
rect 26329 3009 26341 3012
rect 26375 3009 26387 3043
rect 26329 3003 26387 3009
rect 27157 3043 27215 3049
rect 27157 3009 27169 3043
rect 27203 3040 27215 3043
rect 27525 3043 27583 3049
rect 27525 3040 27537 3043
rect 27203 3012 27537 3040
rect 27203 3009 27215 3012
rect 27157 3003 27215 3009
rect 27525 3009 27537 3012
rect 27571 3009 27583 3043
rect 27525 3003 27583 3009
rect 26344 2972 26372 3003
rect 27433 2975 27491 2981
rect 27433 2972 27445 2975
rect 26344 2944 27445 2972
rect 27433 2941 27445 2944
rect 27479 2972 27491 2975
rect 27801 2975 27859 2981
rect 27801 2972 27813 2975
rect 27479 2944 27813 2972
rect 27479 2941 27491 2944
rect 27433 2935 27491 2941
rect 27801 2941 27813 2944
rect 27847 2941 27859 2975
rect 27801 2935 27859 2941
rect 27617 2907 27675 2913
rect 27617 2904 27629 2907
rect 26160 2876 27629 2904
rect 27617 2873 27629 2876
rect 27663 2904 27675 2907
rect 28460 2904 28488 3148
rect 30466 3136 30472 3148
rect 30524 3136 30530 3188
rect 30558 3136 30564 3188
rect 30616 3136 30622 3188
rect 30650 3136 30656 3188
rect 30708 3176 30714 3188
rect 31389 3179 31447 3185
rect 31389 3176 31401 3179
rect 30708 3148 31401 3176
rect 30708 3136 30714 3148
rect 31389 3145 31401 3148
rect 31435 3145 31447 3179
rect 31389 3139 31447 3145
rect 31570 3136 31576 3188
rect 31628 3136 31634 3188
rect 34146 3136 34152 3188
rect 34204 3136 34210 3188
rect 28804 3111 28862 3117
rect 28804 3077 28816 3111
rect 28850 3108 28862 3111
rect 29546 3108 29552 3120
rect 28850 3080 29552 3108
rect 28850 3077 28862 3080
rect 28804 3071 28862 3077
rect 29546 3068 29552 3080
rect 29604 3068 29610 3120
rect 31478 3108 31484 3120
rect 30668 3080 31484 3108
rect 28534 3000 28540 3052
rect 28592 3000 28598 3052
rect 30374 3000 30380 3052
rect 30432 3000 30438 3052
rect 30469 3043 30527 3049
rect 30469 3009 30481 3043
rect 30515 3009 30527 3043
rect 30469 3003 30527 3009
rect 30484 2972 30512 3003
rect 27663 2876 28488 2904
rect 30208 2944 30512 2972
rect 27663 2873 27675 2876
rect 27617 2867 27675 2873
rect 30208 2848 30236 2944
rect 30668 2913 30696 3080
rect 31478 3068 31484 3080
rect 31536 3108 31542 3120
rect 32125 3111 32183 3117
rect 32125 3108 32137 3111
rect 31536 3080 32137 3108
rect 31536 3068 31542 3080
rect 32125 3077 32137 3080
rect 32171 3077 32183 3111
rect 32125 3071 32183 3077
rect 32309 3111 32367 3117
rect 32309 3077 32321 3111
rect 32355 3108 32367 3111
rect 32398 3108 32404 3120
rect 32355 3080 32404 3108
rect 32355 3077 32367 3080
rect 32309 3071 32367 3077
rect 32398 3068 32404 3080
rect 32456 3068 32462 3120
rect 30745 3043 30803 3049
rect 30745 3009 30757 3043
rect 30791 3040 30803 3043
rect 30926 3040 30932 3052
rect 30791 3012 30932 3040
rect 30791 3009 30803 3012
rect 30745 3003 30803 3009
rect 30926 3000 30932 3012
rect 30984 3000 30990 3052
rect 31297 3043 31355 3049
rect 31297 3009 31309 3043
rect 31343 3040 31355 3043
rect 31386 3040 31392 3052
rect 31343 3012 31392 3040
rect 31343 3009 31355 3012
rect 31297 3003 31355 3009
rect 31386 3000 31392 3012
rect 31444 3000 31450 3052
rect 31662 3000 31668 3052
rect 31720 3000 31726 3052
rect 32766 3000 32772 3052
rect 32824 3000 32830 3052
rect 33042 3049 33048 3052
rect 33036 3003 33048 3049
rect 33042 3000 33048 3003
rect 33100 3000 33106 3052
rect 36081 3043 36139 3049
rect 36081 3040 36093 3043
rect 35636 3012 36093 3040
rect 35636 2981 35664 3012
rect 36081 3009 36093 3012
rect 36127 3009 36139 3043
rect 36081 3003 36139 3009
rect 31481 2975 31539 2981
rect 31481 2941 31493 2975
rect 31527 2972 31539 2975
rect 32493 2975 32551 2981
rect 32493 2972 32505 2975
rect 31527 2944 32505 2972
rect 31527 2941 31539 2944
rect 31481 2935 31539 2941
rect 32493 2941 32505 2944
rect 32539 2941 32551 2975
rect 35621 2975 35679 2981
rect 35621 2972 35633 2975
rect 32493 2935 32551 2941
rect 34072 2944 35633 2972
rect 30653 2907 30711 2913
rect 30653 2873 30665 2907
rect 30699 2873 30711 2907
rect 30653 2867 30711 2873
rect 24302 2796 24308 2848
rect 24360 2836 24366 2848
rect 27341 2839 27399 2845
rect 27341 2836 27353 2839
rect 24360 2808 27353 2836
rect 24360 2796 24366 2808
rect 27341 2805 27353 2808
rect 27387 2836 27399 2839
rect 29917 2839 29975 2845
rect 29917 2836 29929 2839
rect 27387 2808 29929 2836
rect 27387 2805 27399 2808
rect 27341 2799 27399 2805
rect 29917 2805 29929 2808
rect 29963 2836 29975 2839
rect 30190 2836 30196 2848
rect 29963 2808 30196 2836
rect 29963 2805 29975 2808
rect 29917 2799 29975 2805
rect 30190 2796 30196 2808
rect 30248 2796 30254 2848
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 34072 2836 34100 2944
rect 35621 2941 35633 2944
rect 35667 2941 35679 2975
rect 35621 2935 35679 2941
rect 35434 2864 35440 2916
rect 35492 2904 35498 2916
rect 36265 2907 36323 2913
rect 36265 2904 36277 2907
rect 35492 2876 36277 2904
rect 35492 2864 35498 2876
rect 36265 2873 36277 2876
rect 36311 2873 36323 2907
rect 36265 2867 36323 2873
rect 30340 2808 34100 2836
rect 30340 2796 30346 2808
rect 1104 2746 36800 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 36800 2746
rect 1104 2672 36800 2694
rect 5902 2592 5908 2644
rect 5960 2592 5966 2644
rect 9122 2592 9128 2644
rect 9180 2592 9186 2644
rect 18138 2592 18144 2644
rect 18196 2592 18202 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 21361 2635 21419 2641
rect 21361 2632 21373 2635
rect 19576 2604 21373 2632
rect 19576 2592 19582 2604
rect 21361 2601 21373 2604
rect 21407 2601 21419 2635
rect 21361 2595 21419 2601
rect 25777 2635 25835 2641
rect 25777 2601 25789 2635
rect 25823 2632 25835 2635
rect 25958 2632 25964 2644
rect 25823 2604 25964 2632
rect 25823 2601 25835 2604
rect 25777 2595 25835 2601
rect 25958 2592 25964 2604
rect 26016 2592 26022 2644
rect 32953 2635 33011 2641
rect 32953 2601 32965 2635
rect 32999 2632 33011 2635
rect 33042 2632 33048 2644
rect 32999 2604 33048 2632
rect 32999 2601 33011 2604
rect 32953 2595 33011 2601
rect 33042 2592 33048 2604
rect 33100 2592 33106 2644
rect 3329 2567 3387 2573
rect 3329 2533 3341 2567
rect 3375 2564 3387 2567
rect 29914 2564 29920 2576
rect 3375 2536 29920 2564
rect 3375 2533 3387 2536
rect 3329 2527 3387 2533
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 3344 2428 3372 2527
rect 29914 2524 29920 2536
rect 29972 2524 29978 2576
rect 30377 2567 30435 2573
rect 30377 2533 30389 2567
rect 30423 2564 30435 2567
rect 30466 2564 30472 2576
rect 30423 2536 30472 2564
rect 30423 2533 30435 2536
rect 30377 2527 30435 2533
rect 30466 2524 30472 2536
rect 30524 2564 30530 2576
rect 31202 2564 31208 2576
rect 30524 2536 31208 2564
rect 30524 2524 30530 2536
rect 31202 2524 31208 2536
rect 31260 2524 31266 2576
rect 24302 2496 24308 2508
rect 11716 2468 24308 2496
rect 2915 2400 3372 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6089 2431 6147 2437
rect 6089 2428 6101 2431
rect 5868 2400 6101 2428
rect 5868 2388 5874 2400
rect 6089 2397 6101 2400
rect 6135 2397 6147 2431
rect 6089 2391 6147 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 11716 2437 11744 2468
rect 24302 2456 24308 2468
rect 24360 2456 24366 2508
rect 25958 2456 25964 2508
rect 26016 2456 26022 2508
rect 26142 2456 26148 2508
rect 26200 2456 26206 2508
rect 35621 2499 35679 2505
rect 35621 2465 35633 2499
rect 35667 2496 35679 2499
rect 36078 2496 36084 2508
rect 35667 2468 36084 2496
rect 35667 2465 35679 2468
rect 35621 2459 35679 2465
rect 36078 2456 36084 2468
rect 36136 2456 36142 2508
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9088 2400 9321 2428
rect 9088 2388 9094 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 16022 2428 16028 2440
rect 14967 2400 16028 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 18104 2400 18337 2428
rect 18104 2388 18110 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 21545 2431 21603 2437
rect 21545 2428 21557 2431
rect 21324 2400 21557 2428
rect 21324 2388 21330 2400
rect 21545 2397 21557 2400
rect 21591 2397 21603 2431
rect 21545 2391 21603 2397
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 23937 2431 23995 2437
rect 23937 2428 23949 2431
rect 23900 2400 23949 2428
rect 23900 2388 23906 2400
rect 23937 2397 23949 2400
rect 23983 2397 23995 2431
rect 23937 2391 23995 2397
rect 25314 2388 25320 2440
rect 25372 2428 25378 2440
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 25372 2400 26065 2428
rect 25372 2388 25378 2400
rect 26053 2397 26065 2400
rect 26099 2428 26111 2431
rect 26234 2428 26240 2440
rect 26099 2400 26240 2428
rect 26099 2397 26111 2400
rect 26053 2391 26111 2397
rect 26234 2388 26240 2400
rect 26292 2388 26298 2440
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27120 2400 27353 2428
rect 27120 2388 27126 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 30561 2431 30619 2437
rect 30561 2428 30573 2431
rect 29696 2400 30573 2428
rect 29696 2388 29702 2400
rect 30561 2397 30573 2400
rect 30607 2397 30619 2431
rect 30561 2391 30619 2397
rect 32858 2388 32864 2440
rect 32916 2428 32922 2440
rect 33137 2431 33195 2437
rect 33137 2428 33149 2431
rect 32916 2400 33149 2428
rect 32916 2388 32922 2400
rect 33137 2397 33149 2400
rect 33183 2397 33195 2431
rect 33137 2391 33195 2397
rect 35894 2388 35900 2440
rect 35952 2388 35958 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 72 2332 1409 2360
rect 72 2320 78 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 1765 2363 1823 2369
rect 1765 2329 1777 2363
rect 1811 2360 1823 2363
rect 1811 2332 2268 2360
rect 1811 2329 1823 2332
rect 1765 2323 1823 2329
rect 2240 2304 2268 2332
rect 19150 2320 19156 2372
rect 19208 2360 19214 2372
rect 19208 2332 26234 2360
rect 19208 2320 19214 2332
rect 2222 2252 2228 2304
rect 2280 2252 2286 2304
rect 2590 2252 2596 2304
rect 2648 2252 2654 2304
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11885 2295 11943 2301
rect 11885 2292 11897 2295
rect 11664 2264 11897 2292
rect 11664 2252 11670 2264
rect 11885 2261 11897 2264
rect 11931 2261 11943 2295
rect 11885 2255 11943 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14884 2264 15117 2292
rect 14884 2252 14890 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24121 2295 24179 2301
rect 24121 2292 24133 2295
rect 23900 2264 24133 2292
rect 23900 2252 23906 2264
rect 24121 2261 24133 2264
rect 24167 2261 24179 2295
rect 26206 2292 26234 2332
rect 30190 2320 30196 2372
rect 30248 2320 30254 2372
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26206 2264 27169 2292
rect 24121 2255 24179 2261
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 30374 2252 30380 2304
rect 30432 2292 30438 2304
rect 30653 2295 30711 2301
rect 30653 2292 30665 2295
rect 30432 2264 30665 2292
rect 30432 2252 30438 2264
rect 30653 2261 30665 2264
rect 30699 2261 30711 2295
rect 30653 2255 30711 2261
rect 1104 2202 36800 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 36800 2202
rect 1104 2128 36800 2150
rect 2222 1980 2228 2032
rect 2280 2020 2286 2032
rect 30742 2020 30748 2032
rect 2280 1992 30748 2020
rect 2280 1980 2286 1992
rect 30742 1980 30748 1992
rect 30800 1980 30806 2032
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 940 37408 992 37460
rect 21272 37408 21324 37460
rect 4620 37315 4672 37324
rect 4620 37281 4629 37315
rect 4629 37281 4663 37315
rect 4663 37281 4672 37315
rect 4620 37272 4672 37281
rect 17040 37272 17092 37324
rect 1308 37136 1360 37188
rect 5448 37204 5500 37256
rect 6828 37204 6880 37256
rect 10416 37247 10468 37256
rect 10416 37213 10425 37247
rect 10425 37213 10459 37247
rect 10459 37213 10468 37247
rect 10416 37204 10468 37213
rect 12808 37204 12860 37256
rect 17224 37136 17276 37188
rect 17868 37204 17920 37256
rect 29920 37340 29972 37392
rect 31760 37383 31812 37392
rect 31760 37349 31769 37383
rect 31769 37349 31803 37383
rect 31803 37349 31812 37383
rect 31760 37340 31812 37349
rect 28448 37315 28500 37324
rect 28448 37281 28457 37315
rect 28457 37281 28491 37315
rect 28491 37281 28500 37315
rect 28448 37272 28500 37281
rect 19340 37204 19392 37256
rect 19616 37204 19668 37256
rect 22284 37204 22336 37256
rect 25872 37247 25924 37256
rect 25872 37213 25881 37247
rect 25881 37213 25915 37247
rect 25915 37213 25924 37247
rect 25872 37204 25924 37213
rect 28632 37204 28684 37256
rect 34796 37204 34848 37256
rect 36176 37247 36228 37256
rect 36176 37213 36185 37247
rect 36185 37213 36219 37247
rect 36219 37213 36228 37247
rect 36176 37204 36228 37213
rect 20628 37136 20680 37188
rect 25136 37136 25188 37188
rect 31484 37136 31536 37188
rect 37372 37136 37424 37188
rect 2320 37111 2372 37120
rect 2320 37077 2329 37111
rect 2329 37077 2363 37111
rect 2363 37077 2372 37111
rect 2320 37068 2372 37077
rect 7380 37111 7432 37120
rect 7380 37077 7389 37111
rect 7389 37077 7423 37111
rect 7423 37077 7432 37111
rect 7380 37068 7432 37077
rect 10600 37111 10652 37120
rect 10600 37077 10609 37111
rect 10609 37077 10643 37111
rect 10643 37077 10652 37111
rect 10600 37068 10652 37077
rect 13544 37068 13596 37120
rect 16396 37111 16448 37120
rect 16396 37077 16405 37111
rect 16405 37077 16439 37111
rect 16439 37077 16448 37111
rect 16396 37068 16448 37077
rect 20168 37111 20220 37120
rect 20168 37077 20177 37111
rect 20177 37077 20211 37111
rect 20211 37077 20220 37111
rect 20168 37068 20220 37077
rect 22928 37111 22980 37120
rect 22928 37077 22937 37111
rect 22937 37077 22971 37111
rect 22971 37077 22980 37111
rect 22928 37068 22980 37077
rect 26056 37111 26108 37120
rect 26056 37077 26065 37111
rect 26065 37077 26099 37111
rect 26099 37077 26108 37111
rect 26056 37068 26108 37077
rect 30104 37068 30156 37120
rect 36360 37111 36412 37120
rect 36360 37077 36369 37111
rect 36369 37077 36403 37111
rect 36403 37077 36412 37111
rect 36360 37068 36412 37077
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 6828 36907 6880 36916
rect 6828 36873 6837 36907
rect 6837 36873 6871 36907
rect 6871 36873 6880 36907
rect 6828 36864 6880 36873
rect 6920 36728 6972 36780
rect 17040 36796 17092 36848
rect 20628 36907 20680 36916
rect 20628 36873 20637 36907
rect 20637 36873 20671 36907
rect 20671 36873 20680 36907
rect 20628 36864 20680 36873
rect 22284 36907 22336 36916
rect 22284 36873 22293 36907
rect 22293 36873 22327 36907
rect 22327 36873 22336 36907
rect 22284 36864 22336 36873
rect 20168 36796 20220 36848
rect 30104 36839 30156 36848
rect 30104 36805 30113 36839
rect 30113 36805 30147 36839
rect 30147 36805 30156 36839
rect 30104 36796 30156 36805
rect 16672 36728 16724 36780
rect 17960 36728 18012 36780
rect 19156 36771 19208 36780
rect 19156 36737 19165 36771
rect 19165 36737 19199 36771
rect 19199 36737 19208 36771
rect 19156 36728 19208 36737
rect 17408 36703 17460 36712
rect 17408 36669 17417 36703
rect 17417 36669 17451 36703
rect 17451 36669 17460 36703
rect 17408 36660 17460 36669
rect 19248 36703 19300 36712
rect 19248 36669 19257 36703
rect 19257 36669 19291 36703
rect 19291 36669 19300 36703
rect 19248 36660 19300 36669
rect 10416 36592 10468 36644
rect 22560 36728 22612 36780
rect 22836 36728 22888 36780
rect 16120 36524 16172 36576
rect 22744 36592 22796 36644
rect 30840 36592 30892 36644
rect 18328 36524 18380 36576
rect 21548 36524 21600 36576
rect 24124 36567 24176 36576
rect 24124 36533 24133 36567
rect 24133 36533 24167 36567
rect 24167 36533 24176 36567
rect 24124 36524 24176 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 17224 36363 17276 36372
rect 17224 36329 17233 36363
rect 17233 36329 17267 36363
rect 17267 36329 17276 36363
rect 17224 36320 17276 36329
rect 17960 36363 18012 36372
rect 17960 36329 17969 36363
rect 17969 36329 18003 36363
rect 18003 36329 18012 36363
rect 17960 36320 18012 36329
rect 19156 36320 19208 36372
rect 19064 36184 19116 36236
rect 20628 36252 20680 36304
rect 22284 36320 22336 36372
rect 22744 36320 22796 36372
rect 30288 36320 30340 36372
rect 3792 36116 3844 36168
rect 8484 36116 8536 36168
rect 16120 36159 16172 36168
rect 16120 36125 16154 36159
rect 16154 36125 16172 36159
rect 6368 36048 6420 36100
rect 16120 36116 16172 36125
rect 17316 36116 17368 36168
rect 17868 36116 17920 36168
rect 18420 36116 18472 36168
rect 21272 36227 21324 36236
rect 21272 36193 21281 36227
rect 21281 36193 21315 36227
rect 21315 36193 21324 36227
rect 21272 36184 21324 36193
rect 29276 36184 29328 36236
rect 21548 36159 21600 36168
rect 21548 36125 21582 36159
rect 21582 36125 21600 36159
rect 21548 36116 21600 36125
rect 29920 36159 29972 36168
rect 29920 36125 29929 36159
rect 29929 36125 29963 36159
rect 29963 36125 29972 36159
rect 32772 36184 32824 36236
rect 29920 36116 29972 36125
rect 30840 36159 30892 36168
rect 30840 36125 30849 36159
rect 30849 36125 30883 36159
rect 30883 36125 30892 36159
rect 30840 36116 30892 36125
rect 7196 36023 7248 36032
rect 7196 35989 7205 36023
rect 7205 35989 7239 36023
rect 7239 35989 7248 36023
rect 7196 35980 7248 35989
rect 17408 35980 17460 36032
rect 18328 35980 18380 36032
rect 19524 35980 19576 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 6368 35819 6420 35828
rect 6368 35785 6377 35819
rect 6377 35785 6411 35819
rect 6411 35785 6420 35819
rect 6368 35776 6420 35785
rect 16672 35819 16724 35828
rect 16672 35785 16681 35819
rect 16681 35785 16715 35819
rect 16715 35785 16724 35819
rect 16672 35776 16724 35785
rect 17224 35776 17276 35828
rect 19248 35708 19300 35760
rect 6184 35640 6236 35692
rect 16948 35640 17000 35692
rect 21272 35708 21324 35760
rect 30196 35776 30248 35828
rect 36176 35776 36228 35828
rect 19708 35683 19760 35692
rect 19708 35649 19742 35683
rect 19742 35649 19760 35683
rect 19708 35640 19760 35649
rect 29276 35683 29328 35692
rect 29276 35649 29285 35683
rect 29285 35649 29319 35683
rect 29319 35649 29328 35683
rect 29276 35640 29328 35649
rect 29736 35640 29788 35692
rect 19064 35572 19116 35624
rect 20996 35436 21048 35488
rect 30564 35436 30616 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 6184 35275 6236 35284
rect 6184 35241 6193 35275
rect 6193 35241 6227 35275
rect 6227 35241 6236 35275
rect 6184 35232 6236 35241
rect 10324 35232 10376 35284
rect 19708 35275 19760 35284
rect 19708 35241 19717 35275
rect 19717 35241 19751 35275
rect 19751 35241 19760 35275
rect 19708 35232 19760 35241
rect 6736 35139 6788 35148
rect 6736 35105 6745 35139
rect 6745 35105 6779 35139
rect 6779 35105 6788 35139
rect 6736 35096 6788 35105
rect 2136 35028 2188 35080
rect 7196 35028 7248 35080
rect 11704 35096 11756 35148
rect 7288 34960 7340 35012
rect 11060 35028 11112 35080
rect 17132 35028 17184 35080
rect 19800 35096 19852 35148
rect 24492 35232 24544 35284
rect 29736 35275 29788 35284
rect 29736 35241 29745 35275
rect 29745 35241 29779 35275
rect 29779 35241 29788 35275
rect 29736 35232 29788 35241
rect 18788 35028 18840 35080
rect 9864 34960 9916 35012
rect 12900 34960 12952 35012
rect 17040 34960 17092 35012
rect 940 34892 992 34944
rect 9220 34935 9272 34944
rect 9220 34901 9229 34935
rect 9229 34901 9263 34935
rect 9263 34901 9272 34935
rect 9220 34892 9272 34901
rect 13820 34892 13872 34944
rect 14556 34935 14608 34944
rect 14556 34901 14565 34935
rect 14565 34901 14599 34935
rect 14599 34901 14608 34935
rect 14556 34892 14608 34901
rect 15568 34892 15620 34944
rect 17316 34892 17368 34944
rect 18696 34892 18748 34944
rect 20996 35028 21048 35080
rect 21088 35071 21140 35080
rect 21088 35037 21097 35071
rect 21097 35037 21131 35071
rect 21131 35037 21140 35071
rect 21088 35028 21140 35037
rect 21272 35028 21324 35080
rect 22836 35071 22888 35080
rect 22836 35037 22845 35071
rect 22845 35037 22879 35071
rect 22879 35037 22888 35071
rect 22836 35028 22888 35037
rect 23940 35028 23992 35080
rect 24952 35071 25004 35080
rect 24952 35037 24961 35071
rect 24961 35037 24995 35071
rect 24995 35037 25004 35071
rect 24952 35028 25004 35037
rect 30196 35139 30248 35148
rect 30196 35105 30205 35139
rect 30205 35105 30239 35139
rect 30239 35105 30248 35139
rect 30196 35096 30248 35105
rect 30288 35139 30340 35148
rect 30288 35105 30297 35139
rect 30297 35105 30331 35139
rect 30331 35105 30340 35139
rect 30288 35096 30340 35105
rect 20352 34935 20404 34944
rect 20352 34901 20361 34935
rect 20361 34901 20395 34935
rect 20395 34901 20404 34935
rect 20352 34892 20404 34901
rect 22100 34892 22152 34944
rect 24308 34892 24360 34944
rect 25504 34960 25556 35012
rect 24860 34892 24912 34944
rect 25596 34892 25648 34944
rect 26516 34892 26568 34944
rect 30104 34935 30156 34944
rect 30104 34901 30113 34935
rect 30113 34901 30147 34935
rect 30147 34901 30156 34935
rect 30104 34892 30156 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 6368 34688 6420 34740
rect 9864 34731 9916 34740
rect 9864 34697 9873 34731
rect 9873 34697 9907 34731
rect 9907 34697 9916 34731
rect 9864 34688 9916 34697
rect 10048 34688 10100 34740
rect 9220 34620 9272 34672
rect 4620 34552 4672 34604
rect 5632 34595 5684 34604
rect 5632 34561 5641 34595
rect 5641 34561 5675 34595
rect 5675 34561 5684 34595
rect 5632 34552 5684 34561
rect 7012 34552 7064 34604
rect 8484 34595 8536 34604
rect 8484 34561 8493 34595
rect 8493 34561 8527 34595
rect 8527 34561 8536 34595
rect 8484 34552 8536 34561
rect 10232 34595 10284 34604
rect 10232 34561 10266 34595
rect 10266 34561 10284 34595
rect 10232 34552 10284 34561
rect 3792 34527 3844 34536
rect 3792 34493 3801 34527
rect 3801 34493 3835 34527
rect 3835 34493 3844 34527
rect 3792 34484 3844 34493
rect 6736 34484 6788 34536
rect 6920 34527 6972 34536
rect 6920 34493 6929 34527
rect 6929 34493 6963 34527
rect 6963 34493 6972 34527
rect 6920 34484 6972 34493
rect 14004 34688 14056 34740
rect 14556 34688 14608 34740
rect 11704 34595 11756 34604
rect 11704 34561 11713 34595
rect 11713 34561 11747 34595
rect 11747 34561 11756 34595
rect 11704 34552 11756 34561
rect 12164 34595 12216 34604
rect 12164 34561 12198 34595
rect 12198 34561 12216 34595
rect 12164 34552 12216 34561
rect 14096 34620 14148 34672
rect 17040 34731 17092 34740
rect 17040 34697 17049 34731
rect 17049 34697 17083 34731
rect 17083 34697 17092 34731
rect 17040 34688 17092 34697
rect 13728 34595 13780 34604
rect 13728 34561 13762 34595
rect 13762 34561 13780 34595
rect 13728 34552 13780 34561
rect 16856 34595 16908 34604
rect 16856 34561 16865 34595
rect 16865 34561 16899 34595
rect 16899 34561 16908 34595
rect 16856 34552 16908 34561
rect 18328 34688 18380 34740
rect 21088 34688 21140 34740
rect 23940 34688 23992 34740
rect 24308 34731 24360 34740
rect 24308 34697 24317 34731
rect 24317 34697 24351 34731
rect 24351 34697 24360 34731
rect 24308 34688 24360 34697
rect 24952 34688 25004 34740
rect 18696 34663 18748 34672
rect 18696 34629 18705 34663
rect 18705 34629 18739 34663
rect 18739 34629 18748 34663
rect 18696 34620 18748 34629
rect 20352 34620 20404 34672
rect 25412 34620 25464 34672
rect 17132 34484 17184 34536
rect 4712 34348 4764 34400
rect 17316 34527 17368 34536
rect 17316 34493 17325 34527
rect 17325 34493 17359 34527
rect 17359 34493 17368 34527
rect 17316 34484 17368 34493
rect 17684 34484 17736 34536
rect 18788 34527 18840 34536
rect 18788 34493 18797 34527
rect 18797 34493 18831 34527
rect 18831 34493 18840 34527
rect 18788 34484 18840 34493
rect 19800 34595 19852 34604
rect 19800 34561 19809 34595
rect 19809 34561 19843 34595
rect 19843 34561 19852 34595
rect 19800 34552 19852 34561
rect 23848 34552 23900 34604
rect 24768 34552 24820 34604
rect 29276 34620 29328 34672
rect 22100 34484 22152 34536
rect 24492 34527 24544 34536
rect 24492 34493 24501 34527
rect 24501 34493 24535 34527
rect 24535 34493 24544 34527
rect 24492 34484 24544 34493
rect 25044 34484 25096 34536
rect 25596 34552 25648 34604
rect 25504 34484 25556 34536
rect 26332 34484 26384 34536
rect 26516 34527 26568 34536
rect 26516 34493 26525 34527
rect 26525 34493 26559 34527
rect 26559 34493 26568 34527
rect 26516 34484 26568 34493
rect 7104 34348 7156 34400
rect 7564 34348 7616 34400
rect 11612 34391 11664 34400
rect 11612 34357 11621 34391
rect 11621 34357 11655 34391
rect 11655 34357 11664 34391
rect 11612 34348 11664 34357
rect 12992 34348 13044 34400
rect 16672 34348 16724 34400
rect 26608 34416 26660 34468
rect 28632 34416 28684 34468
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 4620 34144 4672 34196
rect 7012 34144 7064 34196
rect 8484 34144 8536 34196
rect 10232 34144 10284 34196
rect 12164 34144 12216 34196
rect 10324 34119 10376 34128
rect 10324 34085 10333 34119
rect 10333 34085 10367 34119
rect 10367 34085 10376 34119
rect 10324 34076 10376 34085
rect 11060 34076 11112 34128
rect 3792 34008 3844 34060
rect 4712 33940 4764 33992
rect 5632 33940 5684 33992
rect 7012 34008 7064 34060
rect 7564 34051 7616 34060
rect 7564 34017 7573 34051
rect 7573 34017 7607 34051
rect 7607 34017 7616 34051
rect 7564 34008 7616 34017
rect 11612 34008 11664 34060
rect 12992 34051 13044 34060
rect 12992 34017 13001 34051
rect 13001 34017 13035 34051
rect 13035 34017 13044 34051
rect 12992 34008 13044 34017
rect 13728 34144 13780 34196
rect 16856 34144 16908 34196
rect 26608 34144 26660 34196
rect 30288 34144 30340 34196
rect 17868 34076 17920 34128
rect 5264 33872 5316 33924
rect 5356 33804 5408 33856
rect 7104 33872 7156 33924
rect 9772 33872 9824 33924
rect 12900 33983 12952 33992
rect 12900 33949 12909 33983
rect 12909 33949 12943 33983
rect 12943 33949 12952 33983
rect 12900 33940 12952 33949
rect 13084 33940 13136 33992
rect 13820 33983 13872 33992
rect 13820 33949 13829 33983
rect 13829 33949 13863 33983
rect 13863 33949 13872 33983
rect 13820 33940 13872 33949
rect 14096 33983 14148 33992
rect 14096 33949 14105 33983
rect 14105 33949 14139 33983
rect 14139 33949 14148 33983
rect 14096 33940 14148 33949
rect 16672 34051 16724 34060
rect 16672 34017 16681 34051
rect 16681 34017 16715 34051
rect 16715 34017 16724 34051
rect 16672 34008 16724 34017
rect 18328 34008 18380 34060
rect 11704 33872 11756 33924
rect 14372 33915 14424 33924
rect 14372 33881 14406 33915
rect 14406 33881 14424 33915
rect 14372 33872 14424 33881
rect 17684 33872 17736 33924
rect 6276 33847 6328 33856
rect 6276 33813 6285 33847
rect 6285 33813 6319 33847
rect 6319 33813 6328 33847
rect 6276 33804 6328 33813
rect 7288 33804 7340 33856
rect 15200 33804 15252 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 5264 33600 5316 33652
rect 14372 33600 14424 33652
rect 6276 33464 6328 33516
rect 14464 33507 14516 33516
rect 14464 33473 14473 33507
rect 14473 33473 14507 33507
rect 14507 33473 14516 33507
rect 14464 33464 14516 33473
rect 17316 33507 17368 33516
rect 17316 33473 17325 33507
rect 17325 33473 17359 33507
rect 17359 33473 17368 33507
rect 17316 33464 17368 33473
rect 17408 33507 17460 33516
rect 17408 33473 17417 33507
rect 17417 33473 17451 33507
rect 17451 33473 17460 33507
rect 17408 33464 17460 33473
rect 18880 33464 18932 33516
rect 21272 33464 21324 33516
rect 22744 33464 22796 33516
rect 24400 33464 24452 33516
rect 26700 33507 26752 33516
rect 26700 33473 26709 33507
rect 26709 33473 26743 33507
rect 26743 33473 26752 33507
rect 26700 33464 26752 33473
rect 35992 33464 36044 33516
rect 19156 33439 19208 33448
rect 19156 33405 19165 33439
rect 19165 33405 19199 33439
rect 19199 33405 19208 33439
rect 19156 33396 19208 33405
rect 24308 33439 24360 33448
rect 24308 33405 24317 33439
rect 24317 33405 24351 33439
rect 24351 33405 24360 33439
rect 24308 33396 24360 33405
rect 26332 33396 26384 33448
rect 26424 33328 26476 33380
rect 26884 33328 26936 33380
rect 36360 33371 36412 33380
rect 36360 33337 36369 33371
rect 36369 33337 36403 33371
rect 36403 33337 36412 33371
rect 36360 33328 36412 33337
rect 18788 33303 18840 33312
rect 18788 33269 18797 33303
rect 18797 33269 18831 33303
rect 18831 33269 18840 33303
rect 18788 33260 18840 33269
rect 20260 33260 20312 33312
rect 22284 33260 22336 33312
rect 24216 33260 24268 33312
rect 28356 33303 28408 33312
rect 28356 33269 28365 33303
rect 28365 33269 28399 33303
rect 28399 33269 28408 33303
rect 28356 33260 28408 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2688 33056 2740 33108
rect 3792 32963 3844 32972
rect 3792 32929 3801 32963
rect 3801 32929 3835 32963
rect 3835 32929 3844 32963
rect 3792 32920 3844 32929
rect 3608 32895 3660 32904
rect 3608 32861 3617 32895
rect 3617 32861 3651 32895
rect 3651 32861 3660 32895
rect 3608 32852 3660 32861
rect 6828 32988 6880 33040
rect 7380 33056 7432 33108
rect 9496 33056 9548 33108
rect 9680 33056 9732 33108
rect 7196 32988 7248 33040
rect 9864 32988 9916 33040
rect 8024 32920 8076 32972
rect 10692 32963 10744 32972
rect 10692 32929 10701 32963
rect 10701 32929 10735 32963
rect 10735 32929 10744 32963
rect 10692 32920 10744 32929
rect 11428 32920 11480 32972
rect 11796 33056 11848 33108
rect 14188 33056 14240 33108
rect 14464 33056 14516 33108
rect 17316 33056 17368 33108
rect 18880 33099 18932 33108
rect 18880 33065 18889 33099
rect 18889 33065 18923 33099
rect 18923 33065 18932 33099
rect 18880 33056 18932 33065
rect 17040 32988 17092 33040
rect 18696 32988 18748 33040
rect 18052 32963 18104 32972
rect 18052 32929 18061 32963
rect 18061 32929 18095 32963
rect 18095 32929 18104 32963
rect 18052 32920 18104 32929
rect 6828 32895 6880 32904
rect 6828 32861 6837 32895
rect 6837 32861 6871 32895
rect 6871 32861 6880 32895
rect 6828 32852 6880 32861
rect 7656 32895 7708 32904
rect 7656 32861 7690 32895
rect 7690 32861 7708 32895
rect 7656 32852 7708 32861
rect 10048 32895 10100 32904
rect 10048 32861 10057 32895
rect 10057 32861 10091 32895
rect 10091 32861 10100 32895
rect 10048 32852 10100 32861
rect 10232 32895 10284 32904
rect 10232 32861 10241 32895
rect 10241 32861 10275 32895
rect 10275 32861 10284 32895
rect 10232 32852 10284 32861
rect 10968 32895 11020 32904
rect 10968 32861 10977 32895
rect 10977 32861 11011 32895
rect 11011 32861 11020 32895
rect 10968 32852 11020 32861
rect 11060 32895 11112 32904
rect 11060 32861 11094 32895
rect 11094 32861 11112 32895
rect 11060 32852 11112 32861
rect 12440 32895 12492 32904
rect 12440 32861 12449 32895
rect 12449 32861 12483 32895
rect 12483 32861 12492 32895
rect 12440 32852 12492 32861
rect 15200 32852 15252 32904
rect 15476 32895 15528 32904
rect 15476 32861 15485 32895
rect 15485 32861 15519 32895
rect 15519 32861 15528 32895
rect 15476 32852 15528 32861
rect 1952 32827 2004 32836
rect 1952 32793 1986 32827
rect 1986 32793 2004 32827
rect 1952 32784 2004 32793
rect 12900 32784 12952 32836
rect 4252 32716 4304 32768
rect 7656 32716 7708 32768
rect 9588 32716 9640 32768
rect 11520 32716 11572 32768
rect 12256 32759 12308 32768
rect 12256 32725 12265 32759
rect 12265 32725 12299 32759
rect 12299 32725 12308 32759
rect 12256 32716 12308 32725
rect 13176 32716 13228 32768
rect 16028 32784 16080 32836
rect 16212 32784 16264 32836
rect 17960 32852 18012 32904
rect 18788 32852 18840 32904
rect 19984 32963 20036 32972
rect 19984 32929 19993 32963
rect 19993 32929 20027 32963
rect 20027 32929 20036 32963
rect 19984 32920 20036 32929
rect 22100 33056 22152 33108
rect 22192 33056 22244 33108
rect 20260 32988 20312 33040
rect 20812 32963 20864 32972
rect 20812 32929 20821 32963
rect 20821 32929 20855 32963
rect 20855 32929 20864 32963
rect 20812 32920 20864 32929
rect 22100 32963 22152 32972
rect 22100 32929 22109 32963
rect 22109 32929 22143 32963
rect 22143 32929 22152 32963
rect 22100 32920 22152 32929
rect 22284 32963 22336 32972
rect 22284 32929 22293 32963
rect 22293 32929 22327 32963
rect 22327 32929 22336 32963
rect 22284 32920 22336 32929
rect 22652 32920 22704 32972
rect 23480 32920 23532 32972
rect 25688 33056 25740 33108
rect 26148 33056 26200 33108
rect 26700 33056 26752 33108
rect 24768 32920 24820 32972
rect 20260 32852 20312 32904
rect 16856 32759 16908 32768
rect 16856 32725 16865 32759
rect 16865 32725 16899 32759
rect 16899 32725 16908 32759
rect 16856 32716 16908 32725
rect 19156 32784 19208 32836
rect 18328 32716 18380 32768
rect 18880 32716 18932 32768
rect 19892 32716 19944 32768
rect 21088 32895 21140 32904
rect 21088 32861 21097 32895
rect 21097 32861 21131 32895
rect 21131 32861 21140 32895
rect 21088 32852 21140 32861
rect 21364 32895 21416 32904
rect 21364 32861 21373 32895
rect 21373 32861 21407 32895
rect 21407 32861 21416 32895
rect 21364 32852 21416 32861
rect 23020 32895 23072 32904
rect 23020 32861 23029 32895
rect 23029 32861 23063 32895
rect 23063 32861 23072 32895
rect 23020 32852 23072 32861
rect 24216 32895 24268 32904
rect 24216 32861 24225 32895
rect 24225 32861 24259 32895
rect 24259 32861 24268 32895
rect 24216 32852 24268 32861
rect 24492 32895 24544 32904
rect 24492 32861 24501 32895
rect 24501 32861 24535 32895
rect 24535 32861 24544 32895
rect 24492 32852 24544 32861
rect 22284 32784 22336 32836
rect 23940 32784 23992 32836
rect 25412 32895 25464 32904
rect 25412 32861 25421 32895
rect 25421 32861 25455 32895
rect 25455 32861 25464 32895
rect 25412 32852 25464 32861
rect 25504 32895 25556 32904
rect 25504 32861 25538 32895
rect 25538 32861 25556 32895
rect 25504 32852 25556 32861
rect 25688 32895 25740 32904
rect 25688 32861 25697 32895
rect 25697 32861 25731 32895
rect 25731 32861 25740 32895
rect 25688 32852 25740 32861
rect 26884 32963 26936 32972
rect 26884 32929 26893 32963
rect 26893 32929 26927 32963
rect 26927 32929 26936 32963
rect 26884 32920 26936 32929
rect 27620 32920 27672 32972
rect 28172 32920 28224 32972
rect 28356 32852 28408 32904
rect 22008 32759 22060 32768
rect 22008 32725 22017 32759
rect 22017 32725 22051 32759
rect 22051 32725 22060 32759
rect 22008 32716 22060 32725
rect 22100 32716 22152 32768
rect 23020 32716 23072 32768
rect 24032 32759 24084 32768
rect 24032 32725 24041 32759
rect 24041 32725 24075 32759
rect 24075 32725 24084 32759
rect 24032 32716 24084 32725
rect 24400 32716 24452 32768
rect 25504 32716 25556 32768
rect 25688 32716 25740 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 1952 32555 2004 32564
rect 1952 32521 1961 32555
rect 1961 32521 1995 32555
rect 1995 32521 2004 32555
rect 1952 32512 2004 32521
rect 2688 32555 2740 32564
rect 2688 32521 2697 32555
rect 2697 32521 2731 32555
rect 2731 32521 2740 32555
rect 2688 32512 2740 32521
rect 3608 32512 3660 32564
rect 4252 32555 4304 32564
rect 4252 32521 4261 32555
rect 4261 32521 4295 32555
rect 4295 32521 4304 32555
rect 4252 32512 4304 32521
rect 3332 32444 3384 32496
rect 1492 32376 1544 32428
rect 2596 32376 2648 32428
rect 6920 32512 6972 32564
rect 8208 32512 8260 32564
rect 8944 32512 8996 32564
rect 9496 32512 9548 32564
rect 13820 32512 13872 32564
rect 6828 32376 6880 32428
rect 7564 32376 7616 32428
rect 940 32172 992 32224
rect 7196 32308 7248 32360
rect 7840 32308 7892 32360
rect 11244 32444 11296 32496
rect 12256 32444 12308 32496
rect 8484 32376 8536 32428
rect 8944 32376 8996 32428
rect 8392 32351 8444 32360
rect 8392 32317 8401 32351
rect 8401 32317 8435 32351
rect 8435 32317 8444 32351
rect 8392 32308 8444 32317
rect 6920 32240 6972 32292
rect 7104 32283 7156 32292
rect 7104 32249 7113 32283
rect 7113 32249 7147 32283
rect 7147 32249 7156 32283
rect 7104 32240 7156 32249
rect 9772 32376 9824 32428
rect 11980 32376 12032 32428
rect 14280 32512 14332 32564
rect 15200 32512 15252 32564
rect 16856 32512 16908 32564
rect 15476 32444 15528 32496
rect 16212 32487 16264 32496
rect 16212 32453 16221 32487
rect 16221 32453 16255 32487
rect 16255 32453 16264 32487
rect 16212 32444 16264 32453
rect 14740 32419 14792 32428
rect 14740 32385 14774 32419
rect 14774 32385 14792 32419
rect 14740 32376 14792 32385
rect 9496 32308 9548 32360
rect 12992 32308 13044 32360
rect 14004 32308 14056 32360
rect 14648 32351 14700 32360
rect 14648 32317 14657 32351
rect 14657 32317 14691 32351
rect 14691 32317 14700 32351
rect 14648 32308 14700 32317
rect 16304 32308 16356 32360
rect 17960 32512 18012 32564
rect 18052 32512 18104 32564
rect 21088 32512 21140 32564
rect 22100 32512 22152 32564
rect 22284 32512 22336 32564
rect 22744 32512 22796 32564
rect 24492 32512 24544 32564
rect 18880 32487 18932 32496
rect 18880 32453 18889 32487
rect 18889 32453 18923 32487
rect 18923 32453 18932 32487
rect 18880 32444 18932 32453
rect 19892 32444 19944 32496
rect 17040 32419 17092 32428
rect 17040 32385 17049 32419
rect 17049 32385 17083 32419
rect 17083 32385 17092 32419
rect 17040 32376 17092 32385
rect 17224 32419 17276 32428
rect 17224 32385 17233 32419
rect 17233 32385 17267 32419
rect 17267 32385 17276 32419
rect 17224 32376 17276 32385
rect 17960 32419 18012 32428
rect 17960 32385 17969 32419
rect 17969 32385 18003 32419
rect 18003 32385 18012 32419
rect 17960 32376 18012 32385
rect 18052 32351 18104 32360
rect 4620 32172 4672 32224
rect 8208 32172 8260 32224
rect 8760 32172 8812 32224
rect 9128 32172 9180 32224
rect 11060 32172 11112 32224
rect 18052 32317 18086 32351
rect 18086 32317 18104 32351
rect 18052 32308 18104 32317
rect 18604 32308 18656 32360
rect 12992 32172 13044 32224
rect 13268 32215 13320 32224
rect 13268 32181 13277 32215
rect 13277 32181 13311 32215
rect 13311 32181 13320 32215
rect 13268 32172 13320 32181
rect 15568 32215 15620 32224
rect 15568 32181 15577 32215
rect 15577 32181 15611 32215
rect 15611 32181 15620 32215
rect 15568 32172 15620 32181
rect 16212 32172 16264 32224
rect 16672 32172 16724 32224
rect 16856 32240 16908 32292
rect 17500 32240 17552 32292
rect 19984 32376 20036 32428
rect 24032 32444 24084 32496
rect 26516 32512 26568 32564
rect 24768 32419 24820 32428
rect 24768 32385 24777 32419
rect 24777 32385 24811 32419
rect 24811 32385 24820 32419
rect 24768 32376 24820 32385
rect 25596 32419 25648 32428
rect 25596 32385 25630 32419
rect 25630 32385 25648 32419
rect 25596 32376 25648 32385
rect 28540 32376 28592 32428
rect 22836 32308 22888 32360
rect 25504 32351 25556 32360
rect 25504 32317 25513 32351
rect 25513 32317 25547 32351
rect 25547 32317 25556 32351
rect 25504 32308 25556 32317
rect 25780 32351 25832 32360
rect 25780 32317 25789 32351
rect 25789 32317 25823 32351
rect 25823 32317 25832 32351
rect 25780 32308 25832 32317
rect 26884 32308 26936 32360
rect 24400 32240 24452 32292
rect 25228 32283 25280 32292
rect 25228 32249 25237 32283
rect 25237 32249 25271 32283
rect 25271 32249 25280 32283
rect 25228 32240 25280 32249
rect 27620 32240 27672 32292
rect 27252 32172 27304 32224
rect 29276 32172 29328 32224
rect 29368 32215 29420 32224
rect 29368 32181 29377 32215
rect 29377 32181 29411 32215
rect 29411 32181 29420 32215
rect 29368 32172 29420 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 6644 31968 6696 32020
rect 7840 31968 7892 32020
rect 8484 31968 8536 32020
rect 4620 31832 4672 31884
rect 7104 31900 7156 31952
rect 9312 31943 9364 31952
rect 9312 31909 9321 31943
rect 9321 31909 9355 31943
rect 9355 31909 9364 31943
rect 9312 31900 9364 31909
rect 11796 31968 11848 32020
rect 12440 32011 12492 32020
rect 12440 31977 12449 32011
rect 12449 31977 12483 32011
rect 12483 31977 12492 32011
rect 12440 31968 12492 31977
rect 13268 31968 13320 32020
rect 14740 31968 14792 32020
rect 22652 31968 22704 32020
rect 23940 31968 23992 32020
rect 15752 31900 15804 31952
rect 17776 31900 17828 31952
rect 7196 31832 7248 31884
rect 7380 31832 7432 31884
rect 5356 31764 5408 31816
rect 2780 31696 2832 31748
rect 6368 31807 6420 31816
rect 6368 31773 6377 31807
rect 6377 31773 6411 31807
rect 6411 31773 6420 31807
rect 6368 31764 6420 31773
rect 6460 31807 6512 31816
rect 6460 31773 6494 31807
rect 6494 31773 6512 31807
rect 6460 31764 6512 31773
rect 6644 31807 6696 31816
rect 6644 31773 6653 31807
rect 6653 31773 6687 31807
rect 6687 31773 6696 31807
rect 6644 31764 6696 31773
rect 7472 31764 7524 31816
rect 8944 31807 8996 31816
rect 8944 31773 8953 31807
rect 8953 31773 8987 31807
rect 8987 31773 8996 31807
rect 8944 31764 8996 31773
rect 9128 31807 9180 31816
rect 9128 31773 9137 31807
rect 9137 31773 9171 31807
rect 9171 31773 9180 31807
rect 9128 31764 9180 31773
rect 10048 31875 10100 31884
rect 10048 31841 10057 31875
rect 10057 31841 10091 31875
rect 10091 31841 10100 31875
rect 10048 31832 10100 31841
rect 10968 31875 11020 31884
rect 10968 31841 10977 31875
rect 10977 31841 11011 31875
rect 11011 31841 11020 31875
rect 10968 31832 11020 31841
rect 11060 31875 11112 31884
rect 11060 31841 11094 31875
rect 11094 31841 11112 31875
rect 11060 31832 11112 31841
rect 11244 31875 11296 31884
rect 11244 31841 11253 31875
rect 11253 31841 11287 31875
rect 11287 31841 11296 31875
rect 11244 31832 11296 31841
rect 9680 31764 9732 31816
rect 10232 31807 10284 31816
rect 10232 31773 10241 31807
rect 10241 31773 10275 31807
rect 10275 31773 10284 31807
rect 10232 31764 10284 31773
rect 12900 31875 12952 31884
rect 12900 31841 12909 31875
rect 12909 31841 12943 31875
rect 12943 31841 12952 31875
rect 12900 31832 12952 31841
rect 12992 31875 13044 31884
rect 12992 31841 13001 31875
rect 13001 31841 13035 31875
rect 13035 31841 13044 31875
rect 12992 31832 13044 31841
rect 13176 31764 13228 31816
rect 3424 31628 3476 31680
rect 5540 31628 5592 31680
rect 5632 31628 5684 31680
rect 8576 31671 8628 31680
rect 8576 31637 8585 31671
rect 8585 31637 8619 31671
rect 8619 31637 8628 31671
rect 8576 31628 8628 31637
rect 13176 31628 13228 31680
rect 14004 31832 14056 31884
rect 14280 31875 14332 31884
rect 14280 31841 14289 31875
rect 14289 31841 14323 31875
rect 14323 31841 14332 31875
rect 14280 31832 14332 31841
rect 14740 31875 14792 31884
rect 14740 31841 14749 31875
rect 14749 31841 14783 31875
rect 14783 31841 14792 31875
rect 14740 31832 14792 31841
rect 14832 31832 14884 31884
rect 17040 31875 17092 31884
rect 17040 31841 17049 31875
rect 17049 31841 17083 31875
rect 17083 31841 17092 31875
rect 17040 31832 17092 31841
rect 17224 31875 17276 31884
rect 17224 31841 17233 31875
rect 17233 31841 17267 31875
rect 17267 31841 17276 31875
rect 17224 31832 17276 31841
rect 17960 31875 18012 31884
rect 17960 31841 17969 31875
rect 17969 31841 18003 31875
rect 18003 31841 18012 31875
rect 17960 31832 18012 31841
rect 18052 31875 18104 31884
rect 18052 31841 18086 31875
rect 18086 31841 18104 31875
rect 18052 31832 18104 31841
rect 18788 31832 18840 31884
rect 19156 31900 19208 31952
rect 23480 31900 23532 31952
rect 24308 31900 24360 31952
rect 28540 32011 28592 32020
rect 28540 31977 28549 32011
rect 28549 31977 28583 32011
rect 28583 31977 28592 32011
rect 28540 31968 28592 31977
rect 31852 31968 31904 32020
rect 25780 31832 25832 31884
rect 28632 31832 28684 31884
rect 15016 31807 15068 31816
rect 15016 31773 15025 31807
rect 15025 31773 15059 31807
rect 15059 31773 15068 31807
rect 15016 31764 15068 31773
rect 15292 31807 15344 31816
rect 15292 31773 15301 31807
rect 15301 31773 15335 31807
rect 15335 31773 15344 31807
rect 15292 31764 15344 31773
rect 16028 31764 16080 31816
rect 16212 31807 16264 31816
rect 16212 31773 16221 31807
rect 16221 31773 16255 31807
rect 16255 31773 16264 31807
rect 16212 31764 16264 31773
rect 16304 31764 16356 31816
rect 15108 31628 15160 31680
rect 18236 31807 18288 31816
rect 18236 31773 18245 31807
rect 18245 31773 18279 31807
rect 18279 31773 18288 31807
rect 18236 31764 18288 31773
rect 26884 31764 26936 31816
rect 28080 31764 28132 31816
rect 31944 31900 31996 31952
rect 32588 31832 32640 31884
rect 29828 31807 29880 31816
rect 29828 31773 29837 31807
rect 29837 31773 29871 31807
rect 29871 31773 29880 31807
rect 29828 31764 29880 31773
rect 31208 31807 31260 31816
rect 31208 31773 31217 31807
rect 31217 31773 31251 31807
rect 31251 31773 31260 31807
rect 31208 31764 31260 31773
rect 27344 31739 27396 31748
rect 27344 31705 27378 31739
rect 27378 31705 27396 31739
rect 27344 31696 27396 31705
rect 29368 31696 29420 31748
rect 18512 31628 18564 31680
rect 27896 31628 27948 31680
rect 29644 31671 29696 31680
rect 29644 31637 29653 31671
rect 29653 31637 29687 31671
rect 29687 31637 29696 31671
rect 29644 31628 29696 31637
rect 30012 31628 30064 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 1768 31356 1820 31408
rect 10232 31424 10284 31476
rect 23480 31424 23532 31476
rect 1860 31331 1912 31340
rect 1860 31297 1894 31331
rect 1894 31297 1912 31331
rect 1860 31288 1912 31297
rect 7288 31356 7340 31408
rect 3424 31331 3476 31340
rect 3424 31297 3433 31331
rect 3433 31297 3467 31331
rect 3467 31297 3476 31331
rect 3424 31288 3476 31297
rect 7380 31331 7432 31340
rect 7380 31297 7389 31331
rect 7389 31297 7423 31331
rect 7423 31297 7432 31331
rect 7380 31288 7432 31297
rect 9312 31356 9364 31408
rect 7656 31288 7708 31340
rect 3516 31263 3568 31272
rect 3516 31229 3525 31263
rect 3525 31229 3559 31263
rect 3559 31229 3568 31263
rect 3516 31220 3568 31229
rect 7564 31263 7616 31272
rect 7564 31229 7573 31263
rect 7573 31229 7607 31263
rect 7607 31229 7616 31263
rect 7564 31220 7616 31229
rect 8392 31220 8444 31272
rect 9404 31288 9456 31340
rect 19892 31331 19944 31340
rect 19892 31297 19901 31331
rect 19901 31297 19935 31331
rect 19935 31297 19944 31331
rect 19892 31288 19944 31297
rect 23848 31331 23900 31340
rect 23848 31297 23857 31331
rect 23857 31297 23891 31331
rect 23891 31297 23900 31331
rect 23848 31288 23900 31297
rect 24768 31288 24820 31340
rect 27344 31424 27396 31476
rect 27896 31467 27948 31476
rect 27896 31433 27905 31467
rect 27905 31433 27939 31467
rect 27939 31433 27948 31467
rect 27896 31424 27948 31433
rect 28080 31356 28132 31408
rect 29644 31399 29696 31408
rect 29644 31365 29678 31399
rect 29678 31365 29696 31399
rect 29644 31356 29696 31365
rect 25320 31288 25372 31340
rect 26148 31331 26200 31340
rect 26148 31297 26157 31331
rect 26157 31297 26191 31331
rect 26191 31297 26200 31331
rect 26148 31288 26200 31297
rect 24952 31263 25004 31272
rect 24952 31229 24961 31263
rect 24961 31229 24995 31263
rect 24995 31229 25004 31263
rect 24952 31220 25004 31229
rect 5540 31152 5592 31204
rect 6460 31152 6512 31204
rect 23296 31195 23348 31204
rect 23296 31161 23305 31195
rect 23305 31161 23339 31195
rect 23339 31161 23348 31195
rect 23296 31152 23348 31161
rect 23940 31152 23992 31204
rect 2688 31084 2740 31136
rect 5632 31084 5684 31136
rect 8024 31084 8076 31136
rect 19708 31127 19760 31136
rect 19708 31093 19717 31127
rect 19717 31093 19751 31127
rect 19751 31093 19760 31127
rect 19708 31084 19760 31093
rect 26056 31220 26108 31272
rect 26056 31084 26108 31136
rect 26516 31084 26568 31136
rect 29276 31288 29328 31340
rect 30196 31288 30248 31340
rect 31944 31331 31996 31340
rect 31944 31297 31953 31331
rect 31953 31297 31987 31331
rect 31987 31297 31996 31331
rect 31944 31288 31996 31297
rect 28172 31263 28224 31272
rect 28172 31229 28181 31263
rect 28181 31229 28215 31263
rect 28215 31229 28224 31263
rect 28172 31220 28224 31229
rect 28540 31220 28592 31272
rect 30564 31220 30616 31272
rect 29368 31084 29420 31136
rect 30748 31127 30800 31136
rect 30748 31093 30757 31127
rect 30757 31093 30791 31127
rect 30791 31093 30800 31127
rect 30748 31084 30800 31093
rect 31760 31127 31812 31136
rect 31760 31093 31769 31127
rect 31769 31093 31803 31127
rect 31803 31093 31812 31127
rect 31760 31084 31812 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1860 30880 1912 30932
rect 7380 30880 7432 30932
rect 26056 30880 26108 30932
rect 25228 30812 25280 30864
rect 29828 30880 29880 30932
rect 2596 30744 2648 30796
rect 5356 30744 5408 30796
rect 5632 30744 5684 30796
rect 5816 30744 5868 30796
rect 6184 30787 6236 30796
rect 6184 30753 6193 30787
rect 6193 30753 6227 30787
rect 6227 30753 6236 30787
rect 6184 30744 6236 30753
rect 6368 30744 6420 30796
rect 6644 30744 6696 30796
rect 2688 30719 2740 30728
rect 2688 30685 2697 30719
rect 2697 30685 2731 30719
rect 2731 30685 2740 30719
rect 2688 30676 2740 30685
rect 2780 30719 2832 30728
rect 2780 30685 2789 30719
rect 2789 30685 2823 30719
rect 2823 30685 2832 30719
rect 2780 30676 2832 30685
rect 7196 30719 7248 30728
rect 7196 30685 7205 30719
rect 7205 30685 7239 30719
rect 7239 30685 7248 30719
rect 7196 30676 7248 30685
rect 11336 30676 11388 30728
rect 12072 30676 12124 30728
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 15476 30676 15528 30728
rect 19432 30719 19484 30728
rect 19432 30685 19441 30719
rect 19441 30685 19475 30719
rect 19475 30685 19484 30719
rect 19432 30676 19484 30685
rect 19708 30719 19760 30728
rect 19708 30685 19742 30719
rect 19742 30685 19760 30719
rect 19708 30676 19760 30685
rect 5264 30608 5316 30660
rect 7840 30608 7892 30660
rect 12348 30608 12400 30660
rect 21180 30719 21232 30728
rect 21180 30685 21189 30719
rect 21189 30685 21223 30719
rect 21223 30685 21232 30719
rect 21180 30676 21232 30685
rect 25320 30787 25372 30796
rect 25320 30753 25329 30787
rect 25329 30753 25363 30787
rect 25363 30753 25372 30787
rect 25320 30744 25372 30753
rect 25780 30787 25832 30796
rect 25780 30753 25789 30787
rect 25789 30753 25823 30787
rect 25823 30753 25832 30787
rect 25780 30744 25832 30753
rect 25872 30744 25924 30796
rect 30748 30812 30800 30864
rect 30288 30787 30340 30796
rect 30288 30753 30297 30787
rect 30297 30753 30331 30787
rect 30331 30753 30340 30787
rect 30288 30744 30340 30753
rect 22652 30676 22704 30728
rect 24584 30719 24636 30728
rect 24584 30685 24593 30719
rect 24593 30685 24627 30719
rect 24627 30685 24636 30719
rect 24584 30676 24636 30685
rect 24952 30676 25004 30728
rect 25136 30719 25188 30728
rect 25136 30685 25145 30719
rect 25145 30685 25179 30719
rect 25179 30685 25188 30719
rect 25136 30676 25188 30685
rect 26056 30719 26108 30728
rect 26056 30685 26065 30719
rect 26065 30685 26099 30719
rect 26099 30685 26108 30719
rect 26056 30676 26108 30685
rect 26148 30719 26200 30728
rect 26148 30685 26182 30719
rect 26182 30685 26200 30719
rect 26148 30676 26200 30685
rect 4804 30540 4856 30592
rect 7104 30583 7156 30592
rect 7104 30549 7113 30583
rect 7113 30549 7147 30583
rect 7147 30549 7156 30583
rect 7104 30540 7156 30549
rect 13360 30583 13412 30592
rect 13360 30549 13369 30583
rect 13369 30549 13403 30583
rect 13403 30549 13412 30583
rect 13360 30540 13412 30549
rect 14096 30583 14148 30592
rect 14096 30549 14105 30583
rect 14105 30549 14139 30583
rect 14139 30549 14148 30583
rect 14096 30540 14148 30549
rect 17224 30540 17276 30592
rect 20720 30540 20772 30592
rect 30380 30676 30432 30728
rect 31760 30676 31812 30728
rect 22192 30540 22244 30592
rect 24216 30583 24268 30592
rect 24216 30549 24225 30583
rect 24225 30549 24259 30583
rect 24259 30549 24268 30583
rect 24216 30540 24268 30549
rect 32404 30608 32456 30660
rect 25780 30540 25832 30592
rect 26240 30540 26292 30592
rect 26608 30540 26660 30592
rect 29828 30540 29880 30592
rect 30012 30540 30064 30592
rect 31208 30540 31260 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 3516 30200 3568 30252
rect 4804 30268 4856 30320
rect 7840 30379 7892 30388
rect 7840 30345 7849 30379
rect 7849 30345 7883 30379
rect 7883 30345 7892 30379
rect 7840 30336 7892 30345
rect 11336 30336 11388 30388
rect 11888 30336 11940 30388
rect 12348 30379 12400 30388
rect 12348 30345 12357 30379
rect 12357 30345 12391 30379
rect 12391 30345 12400 30379
rect 12348 30336 12400 30345
rect 13360 30336 13412 30388
rect 7196 30268 7248 30320
rect 7012 30200 7064 30252
rect 8024 30243 8076 30252
rect 8024 30209 8033 30243
rect 8033 30209 8067 30243
rect 8067 30209 8076 30243
rect 8024 30200 8076 30209
rect 9128 30200 9180 30252
rect 12164 30268 12216 30320
rect 10232 30243 10284 30252
rect 10232 30209 10266 30243
rect 10266 30209 10284 30243
rect 10232 30200 10284 30209
rect 10508 30200 10560 30252
rect 8392 30132 8444 30184
rect 5356 29996 5408 30048
rect 9864 30039 9916 30048
rect 9864 30005 9873 30039
rect 9873 30005 9907 30039
rect 9907 30005 9916 30039
rect 9864 29996 9916 30005
rect 10140 29996 10192 30048
rect 12992 30243 13044 30252
rect 12992 30209 13001 30243
rect 13001 30209 13035 30243
rect 13035 30209 13044 30243
rect 12992 30200 13044 30209
rect 14096 30268 14148 30320
rect 19892 30379 19944 30388
rect 19892 30345 19901 30379
rect 19901 30345 19935 30379
rect 19935 30345 19944 30379
rect 19892 30336 19944 30345
rect 20720 30336 20772 30388
rect 21180 30336 21232 30388
rect 22192 30379 22244 30388
rect 13268 30175 13320 30184
rect 13268 30141 13277 30175
rect 13277 30141 13311 30175
rect 13311 30141 13320 30175
rect 13268 30132 13320 30141
rect 11520 30039 11572 30048
rect 11520 30005 11529 30039
rect 11529 30005 11563 30039
rect 11563 30005 11572 30039
rect 11520 29996 11572 30005
rect 14556 29996 14608 30048
rect 16856 30243 16908 30252
rect 16856 30209 16865 30243
rect 16865 30209 16899 30243
rect 16899 30209 16908 30243
rect 16856 30200 16908 30209
rect 17132 30243 17184 30252
rect 17132 30209 17141 30243
rect 17141 30209 17175 30243
rect 17175 30209 17184 30243
rect 17132 30200 17184 30209
rect 17224 30175 17276 30184
rect 17224 30141 17233 30175
rect 17233 30141 17267 30175
rect 17267 30141 17276 30175
rect 17224 30132 17276 30141
rect 20260 30243 20312 30252
rect 20260 30209 20269 30243
rect 20269 30209 20303 30243
rect 20303 30209 20312 30243
rect 20260 30200 20312 30209
rect 20628 30268 20680 30320
rect 22192 30345 22201 30379
rect 22201 30345 22235 30379
rect 22235 30345 22244 30379
rect 22192 30336 22244 30345
rect 24584 30336 24636 30388
rect 25136 30336 25188 30388
rect 31208 30336 31260 30388
rect 22284 30311 22336 30320
rect 22284 30277 22293 30311
rect 22293 30277 22327 30311
rect 22327 30277 22336 30311
rect 22284 30268 22336 30277
rect 24768 30268 24820 30320
rect 22468 30175 22520 30184
rect 22468 30141 22477 30175
rect 22477 30141 22511 30175
rect 22511 30141 22520 30175
rect 22468 30132 22520 30141
rect 23756 30200 23808 30252
rect 24032 30200 24084 30252
rect 24216 30243 24268 30252
rect 24216 30209 24225 30243
rect 24225 30209 24259 30243
rect 24259 30209 24268 30243
rect 24216 30200 24268 30209
rect 24400 30200 24452 30252
rect 26148 30268 26200 30320
rect 25044 30243 25096 30252
rect 25044 30209 25053 30243
rect 25053 30209 25087 30243
rect 25087 30209 25096 30243
rect 25044 30200 25096 30209
rect 24952 30132 25004 30184
rect 23388 30107 23440 30116
rect 23388 30073 23397 30107
rect 23397 30073 23431 30107
rect 23431 30073 23440 30107
rect 27804 30243 27856 30252
rect 27804 30209 27813 30243
rect 27813 30209 27847 30243
rect 27847 30209 27856 30243
rect 27804 30200 27856 30209
rect 28080 30200 28132 30252
rect 36544 30200 36596 30252
rect 27988 30175 28040 30184
rect 27988 30141 27997 30175
rect 27997 30141 28031 30175
rect 28031 30141 28040 30175
rect 27988 30132 28040 30141
rect 23388 30064 23440 30073
rect 15476 29996 15528 30048
rect 16580 29996 16632 30048
rect 17868 29996 17920 30048
rect 18880 30039 18932 30048
rect 18880 30005 18889 30039
rect 18889 30005 18923 30039
rect 18923 30005 18932 30039
rect 18880 29996 18932 30005
rect 19708 30039 19760 30048
rect 19708 30005 19717 30039
rect 19717 30005 19751 30039
rect 19751 30005 19760 30039
rect 19708 29996 19760 30005
rect 20260 29996 20312 30048
rect 20904 29996 20956 30048
rect 22284 29996 22336 30048
rect 27160 30039 27212 30048
rect 27160 30005 27169 30039
rect 27169 30005 27203 30039
rect 27203 30005 27212 30039
rect 27160 29996 27212 30005
rect 28448 29996 28500 30048
rect 36360 30039 36412 30048
rect 36360 30005 36369 30039
rect 36369 30005 36403 30039
rect 36403 30005 36412 30039
rect 36360 29996 36412 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 5264 29835 5316 29844
rect 5264 29801 5273 29835
rect 5273 29801 5307 29835
rect 5307 29801 5316 29835
rect 5264 29792 5316 29801
rect 9128 29835 9180 29844
rect 9128 29801 9137 29835
rect 9137 29801 9171 29835
rect 9171 29801 9180 29835
rect 9128 29792 9180 29801
rect 10232 29792 10284 29844
rect 14280 29792 14332 29844
rect 16856 29792 16908 29844
rect 17132 29792 17184 29844
rect 27804 29792 27856 29844
rect 28264 29835 28316 29844
rect 28264 29801 28273 29835
rect 28273 29801 28307 29835
rect 28307 29801 28316 29835
rect 28264 29792 28316 29801
rect 5908 29724 5960 29776
rect 3516 29656 3568 29708
rect 5724 29699 5776 29708
rect 5724 29665 5733 29699
rect 5733 29665 5767 29699
rect 5767 29665 5776 29699
rect 5724 29656 5776 29665
rect 7564 29724 7616 29776
rect 6368 29656 6420 29708
rect 3608 29631 3660 29640
rect 3608 29597 3617 29631
rect 3617 29597 3651 29631
rect 3651 29597 3660 29631
rect 3608 29588 3660 29597
rect 5356 29588 5408 29640
rect 7656 29588 7708 29640
rect 8208 29588 8260 29640
rect 9496 29588 9548 29640
rect 13268 29724 13320 29776
rect 11520 29656 11572 29708
rect 7564 29520 7616 29572
rect 10600 29631 10652 29640
rect 10600 29597 10609 29631
rect 10609 29597 10643 29631
rect 10643 29597 10652 29631
rect 10600 29588 10652 29597
rect 6184 29452 6236 29504
rect 7840 29452 7892 29504
rect 9864 29520 9916 29572
rect 10968 29520 11020 29572
rect 10508 29495 10560 29504
rect 10508 29461 10517 29495
rect 10517 29461 10551 29495
rect 10551 29461 10560 29495
rect 14556 29588 14608 29640
rect 16580 29699 16632 29708
rect 16580 29665 16589 29699
rect 16589 29665 16623 29699
rect 16623 29665 16632 29699
rect 16580 29656 16632 29665
rect 19708 29724 19760 29776
rect 18880 29656 18932 29708
rect 22652 29656 22704 29708
rect 24952 29699 25004 29708
rect 24952 29665 24961 29699
rect 24961 29665 24995 29699
rect 24995 29665 25004 29699
rect 24952 29656 25004 29665
rect 26884 29699 26936 29708
rect 26884 29665 26893 29699
rect 26893 29665 26927 29699
rect 26927 29665 26936 29699
rect 26884 29656 26936 29665
rect 21088 29588 21140 29640
rect 23296 29588 23348 29640
rect 24860 29631 24912 29640
rect 24860 29597 24869 29631
rect 24869 29597 24903 29631
rect 24903 29597 24912 29631
rect 24860 29588 24912 29597
rect 27160 29631 27212 29640
rect 27160 29597 27194 29631
rect 27194 29597 27212 29631
rect 27160 29588 27212 29597
rect 29368 29631 29420 29640
rect 29368 29597 29377 29631
rect 29377 29597 29411 29631
rect 29411 29597 29420 29631
rect 29368 29588 29420 29597
rect 30196 29588 30248 29640
rect 31208 29631 31260 29640
rect 31208 29597 31217 29631
rect 31217 29597 31251 29631
rect 31251 29597 31260 29631
rect 31208 29588 31260 29597
rect 16948 29520 17000 29572
rect 17776 29563 17828 29572
rect 17776 29529 17785 29563
rect 17785 29529 17819 29563
rect 17819 29529 17828 29563
rect 17776 29520 17828 29529
rect 10508 29452 10560 29461
rect 12992 29452 13044 29504
rect 17316 29452 17368 29504
rect 17684 29452 17736 29504
rect 20444 29452 20496 29504
rect 20812 29452 20864 29504
rect 25504 29452 25556 29504
rect 29920 29452 29972 29504
rect 31024 29495 31076 29504
rect 31024 29461 31033 29495
rect 31033 29461 31067 29495
rect 31067 29461 31076 29495
rect 31024 29452 31076 29461
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 3608 29248 3660 29300
rect 4712 29248 4764 29300
rect 5724 29248 5776 29300
rect 7840 29291 7892 29300
rect 7840 29257 7849 29291
rect 7849 29257 7883 29291
rect 7883 29257 7892 29291
rect 7840 29248 7892 29257
rect 9496 29248 9548 29300
rect 10324 29248 10376 29300
rect 10600 29248 10652 29300
rect 1584 29155 1636 29164
rect 1584 29121 1593 29155
rect 1593 29121 1627 29155
rect 1627 29121 1636 29155
rect 1584 29112 1636 29121
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 2044 29155 2096 29164
rect 2044 29121 2078 29155
rect 2078 29121 2096 29155
rect 2044 29112 2096 29121
rect 5908 29112 5960 29164
rect 6184 29155 6236 29164
rect 6184 29121 6193 29155
rect 6193 29121 6227 29155
rect 6227 29121 6236 29155
rect 6184 29112 6236 29121
rect 8392 29112 8444 29164
rect 12532 29155 12584 29164
rect 12532 29121 12541 29155
rect 12541 29121 12575 29155
rect 12575 29121 12584 29155
rect 12532 29112 12584 29121
rect 19432 29180 19484 29232
rect 19156 29112 19208 29164
rect 20628 29248 20680 29300
rect 24860 29248 24912 29300
rect 25504 29291 25556 29300
rect 25504 29257 25513 29291
rect 25513 29257 25547 29291
rect 25547 29257 25556 29291
rect 25504 29248 25556 29257
rect 22468 29180 22520 29232
rect 20996 29155 21048 29164
rect 20996 29121 21005 29155
rect 21005 29121 21039 29155
rect 21039 29121 21048 29155
rect 20996 29112 21048 29121
rect 22652 29155 22704 29164
rect 22652 29121 22661 29155
rect 22661 29121 22695 29155
rect 22695 29121 22704 29155
rect 22652 29112 22704 29121
rect 22928 29155 22980 29164
rect 22928 29121 22962 29155
rect 22962 29121 22980 29155
rect 22928 29112 22980 29121
rect 23296 29112 23348 29164
rect 24492 29180 24544 29232
rect 27436 29248 27488 29300
rect 29368 29248 29420 29300
rect 29920 29291 29972 29300
rect 29920 29257 29929 29291
rect 29929 29257 29963 29291
rect 29963 29257 29972 29291
rect 29920 29248 29972 29257
rect 31024 29180 31076 29232
rect 6368 29044 6420 29096
rect 20536 29044 20588 29096
rect 20720 29087 20772 29096
rect 20720 29053 20729 29087
rect 20729 29053 20763 29087
rect 20763 29053 20772 29087
rect 20720 29044 20772 29053
rect 20812 29087 20864 29096
rect 20812 29053 20846 29087
rect 20846 29053 20864 29087
rect 20812 29044 20864 29053
rect 21180 29044 21232 29096
rect 1676 28976 1728 29028
rect 12440 28976 12492 29028
rect 20444 29019 20496 29028
rect 3148 28951 3200 28960
rect 3148 28917 3157 28951
rect 3157 28917 3191 28951
rect 3191 28917 3200 28951
rect 3148 28908 3200 28917
rect 5816 28908 5868 28960
rect 10692 28908 10744 28960
rect 20444 28985 20453 29019
rect 20453 28985 20487 29019
rect 20487 28985 20496 29019
rect 20444 28976 20496 28985
rect 24032 29044 24084 29096
rect 25044 29044 25096 29096
rect 27528 29044 27580 29096
rect 28172 29155 28224 29164
rect 28172 29121 28181 29155
rect 28181 29121 28215 29155
rect 28215 29121 28224 29155
rect 28172 29112 28224 29121
rect 28264 29155 28316 29164
rect 28264 29121 28298 29155
rect 28298 29121 28316 29155
rect 28264 29112 28316 29121
rect 28448 29155 28500 29164
rect 28448 29121 28457 29155
rect 28457 29121 28491 29155
rect 28491 29121 28500 29155
rect 28448 29112 28500 29121
rect 29828 29044 29880 29096
rect 30564 29155 30616 29164
rect 30564 29121 30573 29155
rect 30573 29121 30607 29155
rect 30607 29121 30616 29155
rect 30564 29112 30616 29121
rect 30472 29044 30524 29096
rect 29092 29019 29144 29028
rect 29092 28985 29101 29019
rect 29101 28985 29135 29019
rect 29135 28985 29144 29019
rect 29092 28976 29144 28985
rect 19892 28908 19944 28960
rect 20812 28908 20864 28960
rect 21548 28908 21600 28960
rect 23664 28908 23716 28960
rect 24584 28908 24636 28960
rect 25504 28908 25556 28960
rect 28172 28908 28224 28960
rect 28816 28908 28868 28960
rect 31944 28951 31996 28960
rect 31944 28917 31953 28951
rect 31953 28917 31987 28951
rect 31987 28917 31996 28951
rect 31944 28908 31996 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2044 28747 2096 28756
rect 2044 28713 2053 28747
rect 2053 28713 2087 28747
rect 2087 28713 2096 28747
rect 2044 28704 2096 28713
rect 3516 28568 3568 28620
rect 5356 28636 5408 28688
rect 5816 28679 5868 28688
rect 5816 28645 5825 28679
rect 5825 28645 5859 28679
rect 5859 28645 5868 28679
rect 5816 28636 5868 28645
rect 8944 28679 8996 28688
rect 8944 28645 8953 28679
rect 8953 28645 8987 28679
rect 8987 28645 8996 28679
rect 8944 28636 8996 28645
rect 5908 28568 5960 28620
rect 6552 28568 6604 28620
rect 5356 28543 5408 28552
rect 5356 28509 5365 28543
rect 5365 28509 5399 28543
rect 5399 28509 5408 28543
rect 5356 28500 5408 28509
rect 6184 28543 6236 28552
rect 10876 28611 10928 28620
rect 10876 28577 10885 28611
rect 10885 28577 10919 28611
rect 10919 28577 10928 28611
rect 10876 28568 10928 28577
rect 14372 28636 14424 28688
rect 17500 28704 17552 28756
rect 11244 28611 11296 28620
rect 11244 28577 11278 28611
rect 11278 28577 11296 28611
rect 11244 28568 11296 28577
rect 11612 28568 11664 28620
rect 12164 28611 12216 28620
rect 12164 28577 12173 28611
rect 12173 28577 12207 28611
rect 12207 28577 12216 28611
rect 12164 28568 12216 28577
rect 14096 28611 14148 28620
rect 14096 28577 14105 28611
rect 14105 28577 14139 28611
rect 14139 28577 14148 28611
rect 14096 28568 14148 28577
rect 14464 28568 14516 28620
rect 16580 28636 16632 28688
rect 19156 28704 19208 28756
rect 6184 28509 6218 28543
rect 6218 28509 6236 28543
rect 6184 28500 6236 28509
rect 9312 28543 9364 28552
rect 9312 28509 9321 28543
rect 9321 28509 9355 28543
rect 9355 28509 9364 28543
rect 9312 28500 9364 28509
rect 9772 28500 9824 28552
rect 10048 28500 10100 28552
rect 10416 28543 10468 28552
rect 10416 28509 10425 28543
rect 10425 28509 10459 28543
rect 10459 28509 10468 28543
rect 10416 28500 10468 28509
rect 11152 28543 11204 28552
rect 11152 28509 11161 28543
rect 11161 28509 11195 28543
rect 11195 28509 11204 28543
rect 11152 28500 11204 28509
rect 12440 28543 12492 28552
rect 12440 28509 12474 28543
rect 12474 28509 12492 28543
rect 12440 28500 12492 28509
rect 13912 28500 13964 28552
rect 15016 28543 15068 28552
rect 15016 28509 15025 28543
rect 15025 28509 15059 28543
rect 15059 28509 15068 28543
rect 15016 28500 15068 28509
rect 3148 28432 3200 28484
rect 2872 28407 2924 28416
rect 2872 28373 2881 28407
rect 2881 28373 2915 28407
rect 2915 28373 2924 28407
rect 2872 28364 2924 28373
rect 6092 28364 6144 28416
rect 7104 28364 7156 28416
rect 8576 28364 8628 28416
rect 12072 28407 12124 28416
rect 12072 28373 12081 28407
rect 12081 28373 12115 28407
rect 12115 28373 12124 28407
rect 12072 28364 12124 28373
rect 13360 28364 13412 28416
rect 14280 28364 14332 28416
rect 15016 28364 15068 28416
rect 15292 28364 15344 28416
rect 16948 28611 17000 28620
rect 16948 28577 16957 28611
rect 16957 28577 16991 28611
rect 16991 28577 17000 28611
rect 16948 28568 17000 28577
rect 17592 28611 17644 28620
rect 17592 28577 17601 28611
rect 17601 28577 17635 28611
rect 17635 28577 17644 28611
rect 17592 28568 17644 28577
rect 17684 28568 17736 28620
rect 18696 28568 18748 28620
rect 17132 28543 17184 28552
rect 17132 28509 17141 28543
rect 17141 28509 17175 28543
rect 17175 28509 17184 28543
rect 17132 28500 17184 28509
rect 17960 28543 18012 28552
rect 17960 28509 17994 28543
rect 17994 28509 18012 28543
rect 17960 28500 18012 28509
rect 18144 28543 18196 28552
rect 18144 28509 18153 28543
rect 18153 28509 18187 28543
rect 18187 28509 18196 28543
rect 18144 28500 18196 28509
rect 18052 28364 18104 28416
rect 18604 28364 18656 28416
rect 18880 28364 18932 28416
rect 19984 28611 20036 28620
rect 19984 28577 19993 28611
rect 19993 28577 20027 28611
rect 20027 28577 20036 28611
rect 19984 28568 20036 28577
rect 19892 28543 19944 28552
rect 19892 28509 19901 28543
rect 19901 28509 19935 28543
rect 19935 28509 19944 28543
rect 19892 28500 19944 28509
rect 20720 28636 20772 28688
rect 22928 28704 22980 28756
rect 25872 28704 25924 28756
rect 26148 28704 26200 28756
rect 20168 28611 20220 28620
rect 20168 28577 20177 28611
rect 20177 28577 20211 28611
rect 20211 28577 20220 28611
rect 20168 28568 20220 28577
rect 21088 28568 21140 28620
rect 21548 28611 21600 28620
rect 21548 28577 21582 28611
rect 21582 28577 21600 28611
rect 21548 28568 21600 28577
rect 23388 28568 23440 28620
rect 27988 28636 28040 28688
rect 31208 28704 31260 28756
rect 20628 28500 20680 28552
rect 20720 28543 20772 28552
rect 20720 28509 20729 28543
rect 20729 28509 20763 28543
rect 20763 28509 20772 28543
rect 20720 28500 20772 28509
rect 21732 28543 21784 28552
rect 21732 28509 21741 28543
rect 21741 28509 21775 28543
rect 21775 28509 21784 28543
rect 21732 28500 21784 28509
rect 21732 28364 21784 28416
rect 22376 28407 22428 28416
rect 22376 28373 22385 28407
rect 22385 28373 22419 28407
rect 22419 28373 22428 28407
rect 22376 28364 22428 28373
rect 26424 28568 26476 28620
rect 27436 28611 27488 28620
rect 27436 28577 27445 28611
rect 27445 28577 27479 28611
rect 27479 28577 27488 28611
rect 27436 28568 27488 28577
rect 27528 28568 27580 28620
rect 28172 28568 28224 28620
rect 28448 28611 28500 28620
rect 28448 28577 28482 28611
rect 28482 28577 28500 28611
rect 28448 28568 28500 28577
rect 28816 28568 28868 28620
rect 23664 28475 23716 28484
rect 23664 28441 23673 28475
rect 23673 28441 23707 28475
rect 23707 28441 23716 28475
rect 23664 28432 23716 28441
rect 23388 28364 23440 28416
rect 25780 28500 25832 28552
rect 26056 28432 26108 28484
rect 25412 28364 25464 28416
rect 27620 28543 27672 28552
rect 27620 28509 27629 28543
rect 27629 28509 27663 28543
rect 27663 28509 27672 28543
rect 27620 28500 27672 28509
rect 28632 28543 28684 28552
rect 28632 28509 28641 28543
rect 28641 28509 28675 28543
rect 28675 28509 28684 28543
rect 28632 28500 28684 28509
rect 32036 28568 32088 28620
rect 31944 28500 31996 28552
rect 28632 28364 28684 28416
rect 29276 28407 29328 28416
rect 29276 28373 29285 28407
rect 29285 28373 29319 28407
rect 29319 28373 29328 28407
rect 29276 28364 29328 28373
rect 29828 28364 29880 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 5356 28160 5408 28212
rect 9772 28203 9824 28212
rect 9772 28169 9781 28203
rect 9781 28169 9815 28203
rect 9815 28169 9824 28203
rect 9772 28160 9824 28169
rect 12532 28203 12584 28212
rect 12532 28169 12541 28203
rect 12541 28169 12575 28203
rect 12575 28169 12584 28203
rect 12532 28160 12584 28169
rect 14372 28160 14424 28212
rect 16120 28160 16172 28212
rect 8944 28092 8996 28144
rect 9312 28092 9364 28144
rect 3884 28067 3936 28076
rect 3884 28033 3918 28067
rect 3918 28033 3936 28067
rect 3884 28024 3936 28033
rect 8392 28067 8444 28076
rect 8392 28033 8401 28067
rect 8401 28033 8435 28067
rect 8435 28033 8444 28067
rect 8392 28024 8444 28033
rect 12900 28024 12952 28076
rect 3056 27956 3108 28008
rect 14280 28067 14332 28076
rect 14280 28033 14289 28067
rect 14289 28033 14323 28067
rect 14323 28033 14332 28067
rect 14280 28024 14332 28033
rect 14372 28067 14424 28076
rect 14372 28033 14406 28067
rect 14406 28033 14424 28067
rect 14372 28024 14424 28033
rect 14096 27956 14148 28008
rect 14556 27999 14608 28008
rect 14556 27965 14565 27999
rect 14565 27965 14599 27999
rect 14599 27965 14608 27999
rect 16488 28092 16540 28144
rect 14556 27956 14608 27965
rect 13912 27888 13964 27940
rect 14004 27931 14056 27940
rect 14004 27897 14013 27931
rect 14013 27897 14047 27931
rect 14047 27897 14056 27931
rect 14004 27888 14056 27897
rect 16580 28024 16632 28076
rect 20444 28203 20496 28212
rect 20444 28169 20453 28203
rect 20453 28169 20487 28203
rect 20487 28169 20496 28203
rect 20444 28160 20496 28169
rect 20996 28203 21048 28212
rect 20996 28169 21005 28203
rect 21005 28169 21039 28203
rect 21039 28169 21048 28203
rect 20996 28160 21048 28169
rect 16948 28024 17000 28076
rect 17776 28067 17828 28076
rect 17776 28033 17785 28067
rect 17785 28033 17819 28067
rect 17819 28033 17828 28067
rect 17776 28024 17828 28033
rect 17868 28067 17920 28076
rect 17868 28033 17902 28067
rect 17902 28033 17920 28067
rect 17868 28024 17920 28033
rect 18052 28067 18104 28076
rect 18052 28033 18061 28067
rect 18061 28033 18095 28067
rect 18095 28033 18104 28067
rect 18052 28024 18104 28033
rect 15200 27863 15252 27872
rect 15200 27829 15209 27863
rect 15209 27829 15243 27863
rect 15243 27829 15252 27863
rect 15200 27820 15252 27829
rect 15476 27863 15528 27872
rect 15476 27829 15485 27863
rect 15485 27829 15519 27863
rect 15519 27829 15528 27863
rect 15476 27820 15528 27829
rect 17132 27956 17184 28008
rect 17500 27999 17552 28008
rect 17500 27965 17509 27999
rect 17509 27965 17543 27999
rect 17543 27965 17552 27999
rect 17500 27956 17552 27965
rect 18236 27956 18288 28008
rect 19340 28067 19392 28076
rect 19340 28033 19349 28067
rect 19349 28033 19383 28067
rect 19383 28033 19392 28067
rect 19340 28024 19392 28033
rect 20168 28024 20220 28076
rect 20352 28067 20404 28076
rect 20352 28033 20361 28067
rect 20361 28033 20395 28067
rect 20395 28033 20404 28067
rect 20352 28024 20404 28033
rect 23388 28160 23440 28212
rect 21732 28092 21784 28144
rect 21548 28067 21600 28076
rect 21548 28033 21557 28067
rect 21557 28033 21591 28067
rect 21591 28033 21600 28067
rect 21548 28024 21600 28033
rect 24492 28160 24544 28212
rect 24952 28160 25004 28212
rect 26240 28160 26292 28212
rect 27528 28092 27580 28144
rect 27620 28092 27672 28144
rect 28908 28092 28960 28144
rect 24400 28067 24452 28076
rect 24400 28033 24409 28067
rect 24409 28033 24443 28067
rect 24443 28033 24452 28067
rect 24400 28024 24452 28033
rect 24584 28024 24636 28076
rect 25964 28024 26016 28076
rect 16488 27888 16540 27940
rect 16672 27820 16724 27872
rect 17500 27820 17552 27872
rect 19984 27888 20036 27940
rect 20812 27888 20864 27940
rect 21640 27888 21692 27940
rect 21732 27888 21784 27940
rect 23664 27999 23716 28008
rect 23664 27965 23673 27999
rect 23673 27965 23707 27999
rect 23707 27965 23716 27999
rect 23664 27956 23716 27965
rect 24860 27956 24912 28008
rect 25412 27999 25464 28008
rect 23848 27888 23900 27940
rect 24216 27888 24268 27940
rect 18144 27820 18196 27872
rect 18696 27863 18748 27872
rect 18696 27829 18705 27863
rect 18705 27829 18739 27863
rect 18739 27829 18748 27863
rect 18696 27820 18748 27829
rect 18972 27863 19024 27872
rect 18972 27829 18981 27863
rect 18981 27829 19015 27863
rect 19015 27829 19024 27863
rect 18972 27820 19024 27829
rect 20720 27820 20772 27872
rect 24032 27820 24084 27872
rect 24860 27820 24912 27872
rect 25412 27965 25421 27999
rect 25421 27965 25455 27999
rect 25455 27965 25464 27999
rect 25412 27956 25464 27965
rect 28816 27999 28868 28008
rect 28816 27965 28825 27999
rect 28825 27965 28859 27999
rect 28859 27965 28868 27999
rect 28816 27956 28868 27965
rect 28632 27888 28684 27940
rect 25136 27820 25188 27872
rect 26792 27863 26844 27872
rect 26792 27829 26801 27863
rect 26801 27829 26835 27863
rect 26835 27829 26844 27863
rect 26792 27820 26844 27829
rect 27896 27820 27948 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3884 27659 3936 27668
rect 3884 27625 3893 27659
rect 3893 27625 3927 27659
rect 3927 27625 3936 27659
rect 3884 27616 3936 27625
rect 3516 27523 3568 27532
rect 3516 27489 3525 27523
rect 3525 27489 3559 27523
rect 3559 27489 3568 27523
rect 3516 27480 3568 27489
rect 3056 27412 3108 27464
rect 3240 27412 3292 27464
rect 7288 27548 7340 27600
rect 7380 27548 7432 27600
rect 14004 27616 14056 27668
rect 16672 27616 16724 27668
rect 17132 27616 17184 27668
rect 18604 27616 18656 27668
rect 19340 27616 19392 27668
rect 4804 27523 4856 27532
rect 4804 27489 4813 27523
rect 4813 27489 4847 27523
rect 4847 27489 4856 27523
rect 4804 27480 4856 27489
rect 5356 27480 5408 27532
rect 5908 27523 5960 27532
rect 5908 27489 5917 27523
rect 5917 27489 5951 27523
rect 5951 27489 5960 27523
rect 5908 27480 5960 27489
rect 6092 27480 6144 27532
rect 6920 27523 6972 27532
rect 6920 27489 6929 27523
rect 6929 27489 6963 27523
rect 6963 27489 6972 27523
rect 6920 27480 6972 27489
rect 21548 27616 21600 27668
rect 21732 27616 21784 27668
rect 24032 27616 24084 27668
rect 10048 27523 10100 27532
rect 10048 27489 10057 27523
rect 10057 27489 10091 27523
rect 10091 27489 10100 27523
rect 10048 27480 10100 27489
rect 10416 27480 10468 27532
rect 10692 27523 10744 27532
rect 10692 27489 10701 27523
rect 10701 27489 10735 27523
rect 10735 27489 10744 27523
rect 10692 27480 10744 27489
rect 11060 27523 11112 27532
rect 11060 27489 11094 27523
rect 11094 27489 11112 27523
rect 11060 27480 11112 27489
rect 5080 27412 5132 27464
rect 6184 27455 6236 27464
rect 6184 27421 6193 27455
rect 6193 27421 6227 27455
rect 6227 27421 6236 27455
rect 6184 27412 6236 27421
rect 7012 27412 7064 27464
rect 7840 27455 7892 27464
rect 7840 27421 7849 27455
rect 7849 27421 7883 27455
rect 7883 27421 7892 27455
rect 7840 27412 7892 27421
rect 7932 27455 7984 27464
rect 7932 27421 7966 27455
rect 7966 27421 7984 27455
rect 7932 27412 7984 27421
rect 8116 27455 8168 27464
rect 8116 27421 8125 27455
rect 8125 27421 8159 27455
rect 8159 27421 8168 27455
rect 8116 27412 8168 27421
rect 10968 27455 11020 27464
rect 10968 27421 10977 27455
rect 10977 27421 11011 27455
rect 11011 27421 11020 27455
rect 10968 27412 11020 27421
rect 11244 27455 11296 27464
rect 11244 27421 11253 27455
rect 11253 27421 11287 27455
rect 11287 27421 11296 27455
rect 11244 27412 11296 27421
rect 1768 27344 1820 27396
rect 2872 27319 2924 27328
rect 2872 27285 2881 27319
rect 2881 27285 2915 27319
rect 2915 27285 2924 27319
rect 2872 27276 2924 27285
rect 4252 27276 4304 27328
rect 6828 27319 6880 27328
rect 6828 27285 6837 27319
rect 6837 27285 6871 27319
rect 6871 27285 6880 27319
rect 6828 27276 6880 27285
rect 7656 27276 7708 27328
rect 7932 27276 7984 27328
rect 8116 27276 8168 27328
rect 8760 27319 8812 27328
rect 8760 27285 8769 27319
rect 8769 27285 8803 27319
rect 8803 27285 8812 27319
rect 8760 27276 8812 27285
rect 14556 27480 14608 27532
rect 14280 27455 14332 27464
rect 14280 27421 14289 27455
rect 14289 27421 14323 27455
rect 14323 27421 14332 27455
rect 14280 27412 14332 27421
rect 15476 27455 15528 27464
rect 15476 27421 15510 27455
rect 15510 27421 15528 27455
rect 13636 27344 13688 27396
rect 15476 27412 15528 27421
rect 23572 27480 23624 27532
rect 23664 27480 23716 27532
rect 24952 27480 25004 27532
rect 25504 27480 25556 27532
rect 25780 27480 25832 27532
rect 24492 27412 24544 27464
rect 25320 27455 25372 27464
rect 25320 27421 25329 27455
rect 25329 27421 25363 27455
rect 25363 27421 25372 27455
rect 25320 27412 25372 27421
rect 28908 27616 28960 27668
rect 27988 27548 28040 27600
rect 26884 27523 26936 27532
rect 26884 27489 26893 27523
rect 26893 27489 26927 27523
rect 26927 27489 26936 27523
rect 26884 27480 26936 27489
rect 26792 27412 26844 27464
rect 27896 27455 27948 27464
rect 27896 27421 27905 27455
rect 27905 27421 27939 27455
rect 27939 27421 27948 27455
rect 27896 27412 27948 27421
rect 27988 27455 28040 27464
rect 27988 27421 27997 27455
rect 27997 27421 28031 27455
rect 28031 27421 28040 27455
rect 27988 27412 28040 27421
rect 31852 27591 31904 27600
rect 31852 27557 31861 27591
rect 31861 27557 31895 27591
rect 31895 27557 31904 27591
rect 31852 27548 31904 27557
rect 30932 27480 30984 27532
rect 17408 27344 17460 27396
rect 17592 27387 17644 27396
rect 17592 27353 17626 27387
rect 17626 27353 17644 27387
rect 17592 27344 17644 27353
rect 20720 27344 20772 27396
rect 11980 27276 12032 27328
rect 14096 27319 14148 27328
rect 14096 27285 14105 27319
rect 14105 27285 14139 27319
rect 14139 27285 14148 27319
rect 14096 27276 14148 27285
rect 14740 27276 14792 27328
rect 15568 27276 15620 27328
rect 16580 27319 16632 27328
rect 16580 27285 16589 27319
rect 16589 27285 16623 27319
rect 16623 27285 16632 27319
rect 16580 27276 16632 27285
rect 17868 27276 17920 27328
rect 19432 27319 19484 27328
rect 19432 27285 19441 27319
rect 19441 27285 19475 27319
rect 19475 27285 19484 27319
rect 19432 27276 19484 27285
rect 20628 27276 20680 27328
rect 24400 27276 24452 27328
rect 25228 27276 25280 27328
rect 25872 27276 25924 27328
rect 26332 27319 26384 27328
rect 26332 27285 26341 27319
rect 26341 27285 26375 27319
rect 26375 27285 26384 27319
rect 26332 27276 26384 27285
rect 26792 27319 26844 27328
rect 26792 27285 26801 27319
rect 26801 27285 26835 27319
rect 26835 27285 26844 27319
rect 26792 27276 26844 27285
rect 35440 27412 35492 27464
rect 31116 27344 31168 27396
rect 33324 27344 33376 27396
rect 30656 27319 30708 27328
rect 30656 27285 30665 27319
rect 30665 27285 30699 27319
rect 30699 27285 30708 27319
rect 30656 27276 30708 27285
rect 30748 27319 30800 27328
rect 30748 27285 30757 27319
rect 30757 27285 30791 27319
rect 30791 27285 30800 27319
rect 30748 27276 30800 27285
rect 31576 27276 31628 27328
rect 36360 27319 36412 27328
rect 36360 27285 36369 27319
rect 36369 27285 36403 27319
rect 36403 27285 36412 27319
rect 36360 27276 36412 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 1768 27115 1820 27124
rect 1768 27081 1777 27115
rect 1777 27081 1811 27115
rect 1811 27081 1820 27115
rect 1768 27072 1820 27081
rect 10416 27072 10468 27124
rect 14004 27072 14056 27124
rect 14464 27072 14516 27124
rect 15108 27072 15160 27124
rect 18236 27072 18288 27124
rect 18604 27115 18656 27124
rect 18604 27081 18613 27115
rect 18613 27081 18647 27115
rect 18647 27081 18656 27115
rect 18604 27072 18656 27081
rect 23664 27072 23716 27124
rect 24768 27072 24820 27124
rect 25964 27115 26016 27124
rect 25964 27081 25973 27115
rect 25973 27081 26007 27115
rect 26007 27081 26016 27115
rect 25964 27072 26016 27081
rect 26332 27072 26384 27124
rect 26424 27115 26476 27124
rect 26424 27081 26433 27115
rect 26433 27081 26467 27115
rect 26467 27081 26476 27115
rect 26424 27072 26476 27081
rect 26884 27072 26936 27124
rect 28632 27072 28684 27124
rect 31116 27115 31168 27124
rect 31116 27081 31125 27115
rect 31125 27081 31159 27115
rect 31159 27081 31168 27115
rect 31116 27072 31168 27081
rect 2872 26936 2924 26988
rect 2964 26979 3016 26988
rect 2964 26945 2973 26979
rect 2973 26945 3007 26979
rect 3007 26945 3016 26979
rect 2964 26936 3016 26945
rect 3056 26911 3108 26920
rect 3056 26877 3065 26911
rect 3065 26877 3099 26911
rect 3099 26877 3108 26911
rect 3056 26868 3108 26877
rect 7012 26936 7064 26988
rect 7564 26979 7616 26988
rect 7564 26945 7573 26979
rect 7573 26945 7607 26979
rect 7607 26945 7616 26979
rect 7564 26936 7616 26945
rect 7656 26979 7708 26988
rect 7656 26945 7690 26979
rect 7690 26945 7708 26979
rect 7656 26936 7708 26945
rect 8484 26936 8536 26988
rect 10232 26979 10284 26988
rect 10232 26945 10266 26979
rect 10266 26945 10284 26979
rect 10232 26936 10284 26945
rect 11244 26936 11296 26988
rect 14096 27004 14148 27056
rect 12440 26979 12492 26988
rect 12440 26945 12449 26979
rect 12449 26945 12483 26979
rect 12483 26945 12492 26979
rect 12440 26936 12492 26945
rect 15016 26936 15068 26988
rect 18972 27004 19024 27056
rect 19708 27004 19760 27056
rect 20628 27004 20680 27056
rect 22836 27004 22888 27056
rect 17408 26936 17460 26988
rect 19892 26979 19944 26988
rect 19892 26945 19901 26979
rect 19901 26945 19935 26979
rect 19935 26945 19944 26979
rect 19892 26936 19944 26945
rect 20812 26936 20864 26988
rect 22744 26936 22796 26988
rect 6920 26868 6972 26920
rect 4620 26800 4672 26852
rect 6184 26800 6236 26852
rect 7288 26843 7340 26852
rect 7288 26809 7297 26843
rect 7297 26809 7331 26843
rect 7331 26809 7340 26843
rect 7288 26800 7340 26809
rect 7656 26732 7708 26784
rect 9496 26775 9548 26784
rect 9496 26741 9505 26775
rect 9505 26741 9539 26775
rect 9539 26741 9548 26775
rect 9496 26732 9548 26741
rect 11336 26868 11388 26920
rect 13636 26911 13688 26920
rect 13636 26877 13645 26911
rect 13645 26877 13679 26911
rect 13679 26877 13688 26911
rect 13636 26868 13688 26877
rect 17684 26868 17736 26920
rect 10968 26800 11020 26852
rect 11336 26732 11388 26784
rect 11520 26775 11572 26784
rect 11520 26741 11529 26775
rect 11529 26741 11563 26775
rect 11563 26741 11572 26775
rect 11520 26732 11572 26741
rect 12164 26732 12216 26784
rect 14648 26800 14700 26852
rect 19432 26868 19484 26920
rect 24768 26936 24820 26988
rect 32588 27047 32640 27056
rect 32588 27013 32597 27047
rect 32597 27013 32631 27047
rect 32631 27013 32640 27047
rect 32588 27004 32640 27013
rect 26792 26936 26844 26988
rect 28816 26936 28868 26988
rect 30196 26936 30248 26988
rect 30840 26936 30892 26988
rect 31300 26936 31352 26988
rect 31668 26936 31720 26988
rect 30748 26868 30800 26920
rect 30932 26868 30984 26920
rect 31852 26868 31904 26920
rect 33324 26979 33376 26988
rect 33324 26945 33333 26979
rect 33333 26945 33367 26979
rect 33367 26945 33376 26979
rect 33324 26936 33376 26945
rect 32864 26868 32916 26920
rect 29092 26800 29144 26852
rect 29828 26843 29880 26852
rect 29828 26809 29837 26843
rect 29837 26809 29871 26843
rect 29871 26809 29880 26843
rect 29828 26800 29880 26809
rect 15108 26732 15160 26784
rect 17776 26732 17828 26784
rect 19616 26732 19668 26784
rect 20996 26732 21048 26784
rect 23480 26732 23532 26784
rect 25044 26732 25096 26784
rect 28080 26732 28132 26784
rect 28448 26775 28500 26784
rect 28448 26741 28457 26775
rect 28457 26741 28491 26775
rect 28491 26741 28500 26775
rect 28448 26732 28500 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2964 26528 3016 26580
rect 10232 26528 10284 26580
rect 12900 26528 12952 26580
rect 14280 26528 14332 26580
rect 16120 26528 16172 26580
rect 17592 26571 17644 26580
rect 17592 26537 17601 26571
rect 17601 26537 17635 26571
rect 17635 26537 17644 26571
rect 17592 26528 17644 26537
rect 21272 26528 21324 26580
rect 22376 26528 22428 26580
rect 32404 26571 32456 26580
rect 32404 26537 32413 26571
rect 32413 26537 32447 26571
rect 32447 26537 32456 26571
rect 32404 26528 32456 26537
rect 7288 26460 7340 26512
rect 7932 26460 7984 26512
rect 4620 26392 4672 26444
rect 4804 26435 4856 26444
rect 4804 26401 4813 26435
rect 4813 26401 4847 26435
rect 4847 26401 4856 26435
rect 4804 26392 4856 26401
rect 8576 26392 8628 26444
rect 10968 26460 11020 26512
rect 22744 26503 22796 26512
rect 4620 26299 4672 26308
rect 4620 26265 4629 26299
rect 4629 26265 4663 26299
rect 4663 26265 4672 26299
rect 4620 26256 4672 26265
rect 8484 26256 8536 26308
rect 9220 26367 9272 26376
rect 9220 26333 9229 26367
rect 9229 26333 9263 26367
rect 9263 26333 9272 26367
rect 9220 26324 9272 26333
rect 11520 26392 11572 26444
rect 14648 26435 14700 26444
rect 11244 26324 11296 26376
rect 11336 26324 11388 26376
rect 11888 26367 11940 26376
rect 11888 26333 11897 26367
rect 11897 26333 11931 26367
rect 11931 26333 11940 26367
rect 11888 26324 11940 26333
rect 12164 26367 12216 26376
rect 12164 26333 12198 26367
rect 12198 26333 12216 26367
rect 12164 26324 12216 26333
rect 14648 26401 14657 26435
rect 14657 26401 14691 26435
rect 14691 26401 14700 26435
rect 14648 26392 14700 26401
rect 17316 26392 17368 26444
rect 22744 26469 22753 26503
rect 22753 26469 22787 26503
rect 22787 26469 22796 26503
rect 22744 26460 22796 26469
rect 14464 26367 14516 26376
rect 14464 26333 14473 26367
rect 14473 26333 14507 26367
rect 14507 26333 14516 26367
rect 14464 26324 14516 26333
rect 17776 26367 17828 26376
rect 17776 26333 17785 26367
rect 17785 26333 17819 26367
rect 17819 26333 17828 26367
rect 17776 26324 17828 26333
rect 19340 26367 19392 26376
rect 19340 26333 19349 26367
rect 19349 26333 19383 26367
rect 19383 26333 19392 26367
rect 19340 26324 19392 26333
rect 19616 26367 19668 26376
rect 19616 26333 19650 26367
rect 19650 26333 19668 26367
rect 19616 26324 19668 26333
rect 21824 26435 21876 26444
rect 21824 26401 21833 26435
rect 21833 26401 21867 26435
rect 21867 26401 21876 26435
rect 21824 26392 21876 26401
rect 23204 26392 23256 26444
rect 13360 26256 13412 26308
rect 16856 26256 16908 26308
rect 17684 26256 17736 26308
rect 17868 26256 17920 26308
rect 21364 26367 21416 26376
rect 21364 26333 21373 26367
rect 21373 26333 21407 26367
rect 21407 26333 21416 26367
rect 21364 26324 21416 26333
rect 21916 26367 21968 26376
rect 21916 26333 21925 26367
rect 21925 26333 21959 26367
rect 21959 26333 21968 26367
rect 21916 26324 21968 26333
rect 21180 26256 21232 26308
rect 21548 26256 21600 26308
rect 22468 26256 22520 26308
rect 25596 26392 25648 26444
rect 31944 26460 31996 26512
rect 32864 26460 32916 26512
rect 30656 26392 30708 26444
rect 31208 26392 31260 26444
rect 31668 26392 31720 26444
rect 24584 26367 24636 26376
rect 24584 26333 24593 26367
rect 24593 26333 24627 26367
rect 24627 26333 24636 26367
rect 24584 26324 24636 26333
rect 28540 26324 28592 26376
rect 22928 26256 22980 26308
rect 30840 26299 30892 26308
rect 30840 26265 30849 26299
rect 30849 26265 30883 26299
rect 30883 26265 30892 26299
rect 30840 26256 30892 26265
rect 31300 26256 31352 26308
rect 31576 26324 31628 26376
rect 31852 26367 31904 26376
rect 31852 26333 31861 26367
rect 31861 26333 31895 26367
rect 31895 26333 31904 26367
rect 31852 26324 31904 26333
rect 33324 26392 33376 26444
rect 32864 26324 32916 26376
rect 13176 26188 13228 26240
rect 20720 26231 20772 26240
rect 20720 26197 20729 26231
rect 20729 26197 20763 26231
rect 20763 26197 20772 26231
rect 20720 26188 20772 26197
rect 21272 26231 21324 26240
rect 21272 26197 21281 26231
rect 21281 26197 21315 26231
rect 21315 26197 21324 26231
rect 21272 26188 21324 26197
rect 24400 26231 24452 26240
rect 24400 26197 24409 26231
rect 24409 26197 24443 26231
rect 24443 26197 24452 26231
rect 24400 26188 24452 26197
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 6828 26027 6880 26036
rect 6828 25993 6837 26027
rect 6837 25993 6871 26027
rect 6871 25993 6880 26027
rect 6828 25984 6880 25993
rect 2780 25916 2832 25968
rect 4988 25916 5040 25968
rect 9404 25984 9456 26036
rect 12440 26027 12492 26036
rect 12440 25993 12449 26027
rect 12449 25993 12483 26027
rect 12483 25993 12492 26027
rect 12440 25984 12492 25993
rect 12992 25984 13044 26036
rect 13544 25984 13596 26036
rect 17316 25984 17368 26036
rect 18696 25984 18748 26036
rect 19892 26027 19944 26036
rect 19892 25993 19901 26027
rect 19901 25993 19935 26027
rect 19935 25993 19944 26027
rect 19892 25984 19944 25993
rect 20720 25984 20772 26036
rect 22744 25984 22796 26036
rect 2872 25848 2924 25900
rect 6368 25848 6420 25900
rect 7564 25848 7616 25900
rect 8208 25848 8260 25900
rect 9128 25891 9180 25900
rect 9128 25857 9162 25891
rect 9162 25857 9180 25891
rect 9128 25848 9180 25857
rect 9404 25848 9456 25900
rect 3148 25780 3200 25832
rect 7288 25780 7340 25832
rect 8668 25780 8720 25832
rect 10324 25891 10376 25900
rect 10324 25857 10333 25891
rect 10333 25857 10367 25891
rect 10367 25857 10376 25891
rect 10324 25848 10376 25857
rect 11796 25848 11848 25900
rect 8208 25712 8260 25764
rect 11520 25823 11572 25832
rect 11520 25789 11529 25823
rect 11529 25789 11563 25823
rect 11563 25789 11572 25823
rect 11520 25780 11572 25789
rect 12164 25780 12216 25832
rect 13360 25848 13412 25900
rect 15108 25891 15160 25900
rect 15108 25857 15117 25891
rect 15117 25857 15151 25891
rect 15151 25857 15160 25891
rect 15108 25848 15160 25857
rect 15844 25848 15896 25900
rect 13176 25712 13228 25764
rect 14740 25823 14792 25832
rect 14740 25789 14749 25823
rect 14749 25789 14783 25823
rect 14783 25789 14792 25823
rect 14740 25780 14792 25789
rect 14924 25780 14976 25832
rect 17132 25823 17184 25832
rect 17132 25789 17141 25823
rect 17141 25789 17175 25823
rect 17175 25789 17184 25823
rect 17132 25780 17184 25789
rect 18328 25916 18380 25968
rect 17868 25823 17920 25832
rect 1768 25644 1820 25696
rect 6644 25644 6696 25696
rect 7380 25644 7432 25696
rect 8668 25644 8720 25696
rect 9220 25644 9272 25696
rect 10324 25644 10376 25696
rect 10416 25687 10468 25696
rect 10416 25653 10425 25687
rect 10425 25653 10459 25687
rect 10459 25653 10468 25687
rect 10416 25644 10468 25653
rect 10692 25644 10744 25696
rect 13544 25687 13596 25696
rect 13544 25653 13553 25687
rect 13553 25653 13587 25687
rect 13587 25653 13596 25687
rect 13544 25644 13596 25653
rect 14648 25644 14700 25696
rect 16672 25687 16724 25696
rect 16672 25653 16681 25687
rect 16681 25653 16715 25687
rect 16715 25653 16724 25687
rect 16672 25644 16724 25653
rect 17868 25789 17877 25823
rect 17877 25789 17911 25823
rect 17911 25789 17920 25823
rect 17868 25780 17920 25789
rect 18328 25823 18380 25832
rect 18328 25789 18337 25823
rect 18337 25789 18371 25823
rect 18371 25789 18380 25823
rect 18972 25848 19024 25900
rect 21364 25916 21416 25968
rect 22836 25959 22888 25968
rect 22836 25925 22845 25959
rect 22845 25925 22879 25959
rect 22879 25925 22888 25959
rect 22836 25916 22888 25925
rect 20996 25848 21048 25900
rect 21732 25848 21784 25900
rect 22100 25848 22152 25900
rect 26516 25984 26568 26036
rect 24400 25959 24452 25968
rect 24400 25925 24434 25959
rect 24434 25925 24452 25959
rect 24400 25916 24452 25925
rect 24860 25848 24912 25900
rect 25964 25848 26016 25900
rect 33324 26027 33376 26036
rect 33324 25993 33333 26027
rect 33333 25993 33367 26027
rect 33367 25993 33376 26027
rect 33324 25984 33376 25993
rect 27344 25891 27396 25900
rect 27344 25857 27353 25891
rect 27353 25857 27387 25891
rect 27387 25857 27396 25891
rect 27344 25848 27396 25857
rect 28080 25891 28132 25900
rect 28080 25857 28089 25891
rect 28089 25857 28123 25891
rect 28123 25857 28132 25891
rect 28080 25848 28132 25857
rect 31300 25848 31352 25900
rect 33140 25891 33192 25900
rect 33140 25857 33149 25891
rect 33149 25857 33183 25891
rect 33183 25857 33192 25891
rect 33140 25848 33192 25857
rect 18328 25780 18380 25789
rect 20168 25780 20220 25832
rect 20536 25823 20588 25832
rect 20536 25789 20545 25823
rect 20545 25789 20579 25823
rect 20579 25789 20588 25823
rect 20536 25780 20588 25789
rect 18512 25687 18564 25696
rect 18512 25653 18521 25687
rect 18521 25653 18555 25687
rect 18555 25653 18564 25687
rect 18512 25644 18564 25653
rect 18604 25687 18656 25696
rect 18604 25653 18613 25687
rect 18613 25653 18647 25687
rect 18647 25653 18656 25687
rect 18604 25644 18656 25653
rect 20812 25644 20864 25696
rect 21916 25644 21968 25696
rect 23204 25712 23256 25764
rect 26424 25780 26476 25832
rect 27528 25823 27580 25832
rect 27528 25789 27537 25823
rect 27537 25789 27571 25823
rect 27571 25789 27580 25823
rect 27528 25780 27580 25789
rect 30012 25780 30064 25832
rect 31116 25712 31168 25764
rect 32404 25780 32456 25832
rect 32956 25823 33008 25832
rect 32956 25789 32965 25823
rect 32965 25789 32999 25823
rect 32999 25789 33008 25823
rect 32956 25780 33008 25789
rect 23572 25687 23624 25696
rect 23572 25653 23581 25687
rect 23581 25653 23615 25687
rect 23615 25653 23624 25687
rect 23572 25644 23624 25653
rect 25504 25687 25556 25696
rect 25504 25653 25513 25687
rect 25513 25653 25547 25687
rect 25547 25653 25556 25687
rect 25504 25644 25556 25653
rect 26240 25644 26292 25696
rect 27896 25687 27948 25696
rect 27896 25653 27905 25687
rect 27905 25653 27939 25687
rect 27939 25653 27948 25687
rect 27896 25644 27948 25653
rect 31208 25644 31260 25696
rect 33876 25755 33928 25764
rect 33876 25721 33885 25755
rect 33885 25721 33919 25755
rect 33919 25721 33928 25755
rect 33876 25712 33928 25721
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2872 25483 2924 25492
rect 2872 25449 2881 25483
rect 2881 25449 2915 25483
rect 2915 25449 2924 25483
rect 2872 25440 2924 25449
rect 1768 25279 1820 25288
rect 1768 25245 1802 25279
rect 1802 25245 1820 25279
rect 1768 25236 1820 25245
rect 4988 25304 5040 25356
rect 5448 25304 5500 25356
rect 7196 25440 7248 25492
rect 5816 25347 5868 25356
rect 5816 25313 5825 25347
rect 5825 25313 5859 25347
rect 5859 25313 5868 25347
rect 5816 25304 5868 25313
rect 8024 25440 8076 25492
rect 9128 25440 9180 25492
rect 11520 25440 11572 25492
rect 17684 25440 17736 25492
rect 7472 25347 7524 25356
rect 7472 25313 7481 25347
rect 7481 25313 7515 25347
rect 7515 25313 7524 25347
rect 7472 25304 7524 25313
rect 7564 25347 7616 25356
rect 7564 25313 7573 25347
rect 7573 25313 7607 25347
rect 7607 25313 7616 25347
rect 7564 25304 7616 25313
rect 2872 25168 2924 25220
rect 3792 25143 3844 25152
rect 3792 25109 3801 25143
rect 3801 25109 3835 25143
rect 3835 25109 3844 25143
rect 3792 25100 3844 25109
rect 4804 25236 4856 25288
rect 5264 25236 5316 25288
rect 5908 25279 5960 25288
rect 5908 25245 5942 25279
rect 5942 25245 5960 25279
rect 5908 25236 5960 25245
rect 7288 25236 7340 25288
rect 10416 25372 10468 25424
rect 9312 25304 9364 25356
rect 9496 25236 9548 25288
rect 12164 25372 12216 25424
rect 20812 25440 20864 25492
rect 24584 25440 24636 25492
rect 24676 25440 24728 25492
rect 27344 25483 27396 25492
rect 27344 25449 27353 25483
rect 27353 25449 27387 25483
rect 27387 25449 27396 25483
rect 27344 25440 27396 25449
rect 11244 25304 11296 25356
rect 11520 25304 11572 25356
rect 4712 25168 4764 25220
rect 7012 25168 7064 25220
rect 10692 25279 10744 25288
rect 10692 25245 10701 25279
rect 10701 25245 10735 25279
rect 10735 25245 10744 25279
rect 10692 25236 10744 25245
rect 12072 25168 12124 25220
rect 4528 25143 4580 25152
rect 4528 25109 4537 25143
rect 4537 25109 4571 25143
rect 4571 25109 4580 25143
rect 4528 25100 4580 25109
rect 5816 25100 5868 25152
rect 6920 25100 6972 25152
rect 7196 25100 7248 25152
rect 9956 25100 10008 25152
rect 11152 25143 11204 25152
rect 11152 25109 11161 25143
rect 11161 25109 11195 25143
rect 11195 25109 11204 25143
rect 11152 25100 11204 25109
rect 14464 25100 14516 25152
rect 14924 25236 14976 25288
rect 15292 25168 15344 25220
rect 18972 25304 19024 25356
rect 16672 25236 16724 25288
rect 20536 25304 20588 25356
rect 27988 25440 28040 25492
rect 19248 25279 19300 25288
rect 19248 25245 19257 25279
rect 19257 25245 19291 25279
rect 19291 25245 19300 25279
rect 19248 25236 19300 25245
rect 19340 25236 19392 25288
rect 25504 25236 25556 25288
rect 15844 25168 15896 25220
rect 18972 25100 19024 25152
rect 22100 25168 22152 25220
rect 25964 25279 26016 25288
rect 25964 25245 25973 25279
rect 25973 25245 26007 25279
rect 26007 25245 26016 25279
rect 25964 25236 26016 25245
rect 26240 25279 26292 25288
rect 26240 25245 26274 25279
rect 26274 25245 26292 25279
rect 26240 25236 26292 25245
rect 27896 25279 27948 25288
rect 27896 25245 27930 25279
rect 27930 25245 27948 25279
rect 27896 25236 27948 25245
rect 29368 25279 29420 25288
rect 29368 25245 29377 25279
rect 29377 25245 29411 25279
rect 29411 25245 29420 25279
rect 29368 25236 29420 25245
rect 30472 25440 30524 25492
rect 32312 25483 32364 25492
rect 32312 25449 32321 25483
rect 32321 25449 32355 25483
rect 32355 25449 32364 25483
rect 32312 25440 32364 25449
rect 31116 25304 31168 25356
rect 32404 25372 32456 25424
rect 32772 25347 32824 25356
rect 32772 25313 32781 25347
rect 32781 25313 32815 25347
rect 32815 25313 32824 25347
rect 32772 25304 32824 25313
rect 32956 25304 33008 25356
rect 30380 25236 30432 25288
rect 30748 25236 30800 25288
rect 29092 25168 29144 25220
rect 19984 25100 20036 25152
rect 25044 25100 25096 25152
rect 28264 25100 28316 25152
rect 31392 25168 31444 25220
rect 33048 25279 33100 25288
rect 33048 25245 33057 25279
rect 33057 25245 33091 25279
rect 33091 25245 33100 25279
rect 33048 25236 33100 25245
rect 33876 25236 33928 25288
rect 33140 25168 33192 25220
rect 30932 25143 30984 25152
rect 30932 25109 30941 25143
rect 30941 25109 30975 25143
rect 30975 25109 30984 25143
rect 30932 25100 30984 25109
rect 31576 25100 31628 25152
rect 32036 25143 32088 25152
rect 32036 25109 32045 25143
rect 32045 25109 32079 25143
rect 32079 25109 32088 25143
rect 32036 25100 32088 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 4528 24896 4580 24948
rect 8208 24896 8260 24948
rect 11520 24896 11572 24948
rect 18972 24896 19024 24948
rect 19340 24896 19392 24948
rect 19984 24939 20036 24948
rect 19984 24905 19993 24939
rect 19993 24905 20027 24939
rect 20027 24905 20036 24939
rect 19984 24896 20036 24905
rect 20904 24896 20956 24948
rect 3792 24828 3844 24880
rect 7748 24828 7800 24880
rect 1400 24803 1452 24812
rect 1400 24769 1409 24803
rect 1409 24769 1443 24803
rect 1443 24769 1452 24803
rect 1400 24760 1452 24769
rect 1860 24692 1912 24744
rect 2872 24692 2924 24744
rect 3332 24735 3384 24744
rect 3332 24701 3341 24735
rect 3341 24701 3375 24735
rect 3375 24701 3384 24735
rect 3332 24692 3384 24701
rect 6644 24803 6696 24812
rect 6644 24769 6653 24803
rect 6653 24769 6687 24803
rect 6687 24769 6696 24803
rect 6644 24760 6696 24769
rect 7196 24760 7248 24812
rect 7656 24803 7708 24812
rect 7656 24769 7665 24803
rect 7665 24769 7699 24803
rect 7699 24769 7708 24803
rect 7656 24760 7708 24769
rect 11888 24760 11940 24812
rect 12348 24803 12400 24812
rect 12348 24769 12382 24803
rect 12382 24769 12400 24803
rect 12348 24760 12400 24769
rect 12624 24760 12676 24812
rect 7012 24692 7064 24744
rect 8208 24692 8260 24744
rect 14464 24803 14516 24812
rect 14464 24769 14473 24803
rect 14473 24769 14507 24803
rect 14507 24769 14516 24803
rect 14464 24760 14516 24769
rect 14648 24735 14700 24744
rect 14648 24701 14657 24735
rect 14657 24701 14691 24735
rect 14691 24701 14700 24735
rect 14648 24692 14700 24701
rect 14832 24735 14884 24744
rect 14832 24701 14841 24735
rect 14841 24701 14875 24735
rect 14875 24701 14884 24735
rect 14832 24692 14884 24701
rect 18604 24828 18656 24880
rect 7564 24624 7616 24676
rect 10876 24624 10928 24676
rect 11888 24624 11940 24676
rect 14004 24667 14056 24676
rect 14004 24633 14013 24667
rect 14013 24633 14047 24667
rect 14047 24633 14056 24667
rect 14004 24624 14056 24633
rect 14464 24624 14516 24676
rect 16488 24624 16540 24676
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 18512 24692 18564 24744
rect 6276 24556 6328 24608
rect 7104 24556 7156 24608
rect 12992 24556 13044 24608
rect 14096 24556 14148 24608
rect 16672 24556 16724 24608
rect 18604 24624 18656 24676
rect 20168 24760 20220 24812
rect 21180 24803 21232 24812
rect 21180 24769 21189 24803
rect 21189 24769 21223 24803
rect 21223 24769 21232 24803
rect 21180 24760 21232 24769
rect 21824 24760 21876 24812
rect 25136 24896 25188 24948
rect 28080 24896 28132 24948
rect 28264 24939 28316 24948
rect 28264 24905 28273 24939
rect 28273 24905 28307 24939
rect 28307 24905 28316 24939
rect 28264 24896 28316 24905
rect 29368 24896 29420 24948
rect 29828 24939 29880 24948
rect 29828 24905 29837 24939
rect 29837 24905 29871 24939
rect 29871 24905 29880 24939
rect 29828 24896 29880 24905
rect 31576 24896 31628 24948
rect 32036 24896 32088 24948
rect 33876 24939 33928 24948
rect 33876 24905 33885 24939
rect 33885 24905 33919 24939
rect 33919 24905 33928 24939
rect 33876 24896 33928 24905
rect 25228 24828 25280 24880
rect 22928 24803 22980 24812
rect 22928 24769 22937 24803
rect 22937 24769 22971 24803
rect 22971 24769 22980 24803
rect 22928 24760 22980 24769
rect 23112 24760 23164 24812
rect 21272 24692 21324 24744
rect 21548 24692 21600 24744
rect 23204 24692 23256 24744
rect 23940 24692 23992 24744
rect 27528 24760 27580 24812
rect 20904 24599 20956 24608
rect 20904 24565 20913 24599
rect 20913 24565 20947 24599
rect 20947 24565 20956 24599
rect 20904 24556 20956 24565
rect 20996 24556 21048 24608
rect 21548 24556 21600 24608
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 22836 24599 22888 24608
rect 22836 24565 22845 24599
rect 22845 24565 22879 24599
rect 22879 24565 22888 24599
rect 22836 24556 22888 24565
rect 23756 24624 23808 24676
rect 26056 24692 26108 24744
rect 28172 24692 28224 24744
rect 28356 24735 28408 24744
rect 28356 24701 28365 24735
rect 28365 24701 28399 24735
rect 28399 24701 28408 24735
rect 28356 24692 28408 24701
rect 27528 24624 27580 24676
rect 30932 24760 30984 24812
rect 32220 24760 32272 24812
rect 33048 24828 33100 24880
rect 32588 24760 32640 24812
rect 30012 24735 30064 24744
rect 30012 24701 30021 24735
rect 30021 24701 30055 24735
rect 30055 24701 30064 24735
rect 30012 24692 30064 24701
rect 25412 24556 25464 24608
rect 27804 24556 27856 24608
rect 29092 24556 29144 24608
rect 30656 24735 30708 24744
rect 30656 24701 30665 24735
rect 30665 24701 30699 24735
rect 30699 24701 30708 24735
rect 30656 24692 30708 24701
rect 30748 24735 30800 24744
rect 30748 24701 30757 24735
rect 30757 24701 30791 24735
rect 30791 24701 30800 24735
rect 30748 24692 30800 24701
rect 31300 24692 31352 24744
rect 31392 24735 31444 24744
rect 31392 24701 31401 24735
rect 31401 24701 31435 24735
rect 31435 24701 31444 24735
rect 31392 24692 31444 24701
rect 30380 24556 30432 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3332 24352 3384 24404
rect 2504 24284 2556 24336
rect 5264 24284 5316 24336
rect 5172 24216 5224 24268
rect 5724 24259 5776 24268
rect 5724 24225 5733 24259
rect 5733 24225 5767 24259
rect 5767 24225 5776 24259
rect 5724 24216 5776 24225
rect 7288 24259 7340 24268
rect 7288 24225 7297 24259
rect 7297 24225 7331 24259
rect 7331 24225 7340 24259
rect 7288 24216 7340 24225
rect 11244 24352 11296 24404
rect 12348 24395 12400 24404
rect 12348 24361 12357 24395
rect 12357 24361 12391 24395
rect 12391 24361 12400 24395
rect 12348 24352 12400 24361
rect 11704 24284 11756 24336
rect 14832 24352 14884 24404
rect 17960 24352 18012 24404
rect 18604 24395 18656 24404
rect 18604 24361 18613 24395
rect 18613 24361 18647 24395
rect 18647 24361 18656 24395
rect 18604 24352 18656 24361
rect 21272 24395 21324 24404
rect 21272 24361 21281 24395
rect 21281 24361 21315 24395
rect 21315 24361 21324 24395
rect 21272 24352 21324 24361
rect 21824 24395 21876 24404
rect 21824 24361 21833 24395
rect 21833 24361 21867 24395
rect 21867 24361 21876 24395
rect 21824 24352 21876 24361
rect 22100 24395 22152 24404
rect 22100 24361 22109 24395
rect 22109 24361 22143 24395
rect 22143 24361 22152 24395
rect 22100 24352 22152 24361
rect 23112 24352 23164 24404
rect 23572 24352 23624 24404
rect 23940 24352 23992 24404
rect 32588 24352 32640 24404
rect 2964 24148 3016 24200
rect 4804 24191 4856 24200
rect 4804 24157 4813 24191
rect 4813 24157 4847 24191
rect 4847 24157 4856 24191
rect 4804 24148 4856 24157
rect 5816 24191 5868 24200
rect 5816 24157 5850 24191
rect 5850 24157 5868 24191
rect 5816 24148 5868 24157
rect 6000 24191 6052 24200
rect 6000 24157 6009 24191
rect 6009 24157 6043 24191
rect 6043 24157 6052 24191
rect 6000 24148 6052 24157
rect 7012 24191 7064 24200
rect 7012 24157 7021 24191
rect 7021 24157 7055 24191
rect 7055 24157 7064 24191
rect 7012 24148 7064 24157
rect 7104 24191 7156 24200
rect 7104 24157 7113 24191
rect 7113 24157 7147 24191
rect 7147 24157 7156 24191
rect 7104 24148 7156 24157
rect 7380 24191 7432 24200
rect 7380 24157 7389 24191
rect 7389 24157 7423 24191
rect 7423 24157 7432 24191
rect 7380 24148 7432 24157
rect 8668 24148 8720 24200
rect 12900 24216 12952 24268
rect 13084 24259 13136 24268
rect 13084 24225 13093 24259
rect 13093 24225 13127 24259
rect 13127 24225 13136 24259
rect 13084 24216 13136 24225
rect 17868 24327 17920 24336
rect 17868 24293 17877 24327
rect 17877 24293 17911 24327
rect 17911 24293 17920 24327
rect 17868 24284 17920 24293
rect 18512 24327 18564 24336
rect 18512 24293 18521 24327
rect 18521 24293 18555 24327
rect 18555 24293 18564 24327
rect 18512 24284 18564 24293
rect 21364 24284 21416 24336
rect 21640 24327 21692 24336
rect 21640 24293 21649 24327
rect 21649 24293 21683 24327
rect 21683 24293 21692 24327
rect 21640 24284 21692 24293
rect 25320 24327 25372 24336
rect 12992 24191 13044 24200
rect 12992 24157 13001 24191
rect 13001 24157 13035 24191
rect 13035 24157 13044 24191
rect 12992 24148 13044 24157
rect 1768 24080 1820 24132
rect 8852 24080 8904 24132
rect 9312 24080 9364 24132
rect 12624 24080 12676 24132
rect 12716 24080 12768 24132
rect 16488 24148 16540 24200
rect 16948 24148 17000 24200
rect 20444 24148 20496 24200
rect 21456 24216 21508 24268
rect 25320 24293 25329 24327
rect 25329 24293 25363 24327
rect 25363 24293 25372 24327
rect 25320 24284 25372 24293
rect 25412 24284 25464 24336
rect 24676 24259 24728 24268
rect 24676 24225 24685 24259
rect 24685 24225 24719 24259
rect 24719 24225 24728 24259
rect 24676 24216 24728 24225
rect 17132 24080 17184 24132
rect 17592 24080 17644 24132
rect 22468 24148 22520 24200
rect 23204 24148 23256 24200
rect 23388 24191 23440 24200
rect 23388 24157 23397 24191
rect 23397 24157 23431 24191
rect 23431 24157 23440 24191
rect 23388 24148 23440 24157
rect 23480 24191 23532 24200
rect 23480 24157 23489 24191
rect 23489 24157 23523 24191
rect 23523 24157 23532 24191
rect 23480 24148 23532 24157
rect 23756 24191 23808 24200
rect 23756 24157 23765 24191
rect 23765 24157 23799 24191
rect 23799 24157 23808 24191
rect 23756 24148 23808 24157
rect 23940 24148 23992 24200
rect 24860 24191 24912 24200
rect 24860 24157 24869 24191
rect 24869 24157 24903 24191
rect 24903 24157 24912 24191
rect 24860 24148 24912 24157
rect 25596 24191 25648 24200
rect 25596 24157 25605 24191
rect 25605 24157 25639 24191
rect 25639 24157 25648 24191
rect 25596 24148 25648 24157
rect 25688 24191 25740 24200
rect 26240 24216 26292 24268
rect 27528 24259 27580 24268
rect 27528 24225 27537 24259
rect 27537 24225 27571 24259
rect 27571 24225 27580 24259
rect 27528 24216 27580 24225
rect 27988 24216 28040 24268
rect 28172 24216 28224 24268
rect 32220 24284 32272 24336
rect 25688 24157 25722 24191
rect 25722 24157 25740 24191
rect 25688 24148 25740 24157
rect 6644 24055 6696 24064
rect 6644 24021 6653 24055
rect 6653 24021 6687 24055
rect 6687 24021 6696 24055
rect 6644 24012 6696 24021
rect 6736 24012 6788 24064
rect 9864 24012 9916 24064
rect 21732 24012 21784 24064
rect 23020 24012 23072 24064
rect 24032 24012 24084 24064
rect 26792 24191 26844 24200
rect 26792 24157 26801 24191
rect 26801 24157 26835 24191
rect 26835 24157 26844 24191
rect 26792 24148 26844 24157
rect 27804 24191 27856 24200
rect 27804 24157 27813 24191
rect 27813 24157 27847 24191
rect 27847 24157 27856 24191
rect 27804 24148 27856 24157
rect 32128 24148 32180 24200
rect 36084 24148 36136 24200
rect 26976 24012 27028 24064
rect 28264 24012 28316 24064
rect 36360 24055 36412 24064
rect 36360 24021 36369 24055
rect 36369 24021 36403 24055
rect 36403 24021 36412 24055
rect 36360 24012 36412 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 1768 23851 1820 23860
rect 1768 23817 1777 23851
rect 1777 23817 1811 23851
rect 1811 23817 1820 23851
rect 1768 23808 1820 23817
rect 2504 23851 2556 23860
rect 2504 23817 2513 23851
rect 2513 23817 2547 23851
rect 2547 23817 2556 23851
rect 2504 23808 2556 23817
rect 7288 23808 7340 23860
rect 7564 23851 7616 23860
rect 7564 23817 7573 23851
rect 7573 23817 7607 23851
rect 7607 23817 7616 23851
rect 7564 23808 7616 23817
rect 8852 23808 8904 23860
rect 3148 23740 3200 23792
rect 2872 23672 2924 23724
rect 2964 23715 3016 23724
rect 2964 23681 2973 23715
rect 2973 23681 3007 23715
rect 3007 23681 3016 23715
rect 2964 23672 3016 23681
rect 3792 23672 3844 23724
rect 8392 23783 8444 23792
rect 8392 23749 8401 23783
rect 8401 23749 8435 23783
rect 8435 23749 8444 23783
rect 8392 23740 8444 23749
rect 11520 23808 11572 23860
rect 13820 23808 13872 23860
rect 2688 23647 2740 23656
rect 2688 23613 2697 23647
rect 2697 23613 2731 23647
rect 2731 23613 2740 23647
rect 2688 23604 2740 23613
rect 6644 23604 6696 23656
rect 6184 23536 6236 23588
rect 8576 23715 8628 23724
rect 8576 23681 8585 23715
rect 8585 23681 8619 23715
rect 8619 23681 8628 23715
rect 8576 23672 8628 23681
rect 12716 23740 12768 23792
rect 14464 23851 14516 23860
rect 14464 23817 14473 23851
rect 14473 23817 14507 23851
rect 14507 23817 14516 23851
rect 14464 23808 14516 23817
rect 17776 23808 17828 23860
rect 17868 23808 17920 23860
rect 20444 23808 20496 23860
rect 21456 23808 21508 23860
rect 21640 23851 21692 23860
rect 21640 23817 21649 23851
rect 21649 23817 21683 23851
rect 21683 23817 21692 23851
rect 21640 23808 21692 23817
rect 21732 23808 21784 23860
rect 19984 23740 20036 23792
rect 23388 23808 23440 23860
rect 24860 23808 24912 23860
rect 26148 23808 26200 23860
rect 27988 23808 28040 23860
rect 29920 23808 29972 23860
rect 23204 23740 23256 23792
rect 9128 23715 9180 23724
rect 9128 23681 9137 23715
rect 9137 23681 9171 23715
rect 9171 23681 9180 23715
rect 9128 23672 9180 23681
rect 9864 23672 9916 23724
rect 11612 23715 11664 23724
rect 11612 23681 11621 23715
rect 11621 23681 11655 23715
rect 11655 23681 11664 23715
rect 11612 23672 11664 23681
rect 11888 23715 11940 23724
rect 11888 23681 11897 23715
rect 11897 23681 11931 23715
rect 11931 23681 11940 23715
rect 11888 23672 11940 23681
rect 12532 23672 12584 23724
rect 12992 23672 13044 23724
rect 13820 23715 13872 23724
rect 13820 23681 13829 23715
rect 13829 23681 13863 23715
rect 13863 23681 13872 23715
rect 13820 23672 13872 23681
rect 15016 23672 15068 23724
rect 15660 23672 15712 23724
rect 17592 23715 17644 23724
rect 17592 23681 17601 23715
rect 17601 23681 17635 23715
rect 17635 23681 17644 23715
rect 17592 23672 17644 23681
rect 17868 23715 17920 23724
rect 17868 23681 17877 23715
rect 17877 23681 17911 23715
rect 17911 23681 17920 23715
rect 17868 23672 17920 23681
rect 10048 23604 10100 23656
rect 10416 23647 10468 23656
rect 10416 23613 10425 23647
rect 10425 23613 10459 23647
rect 10459 23613 10468 23647
rect 10416 23604 10468 23613
rect 10600 23604 10652 23656
rect 10692 23647 10744 23656
rect 10692 23613 10701 23647
rect 10701 23613 10735 23647
rect 10735 23613 10744 23647
rect 10692 23604 10744 23613
rect 11060 23604 11112 23656
rect 12900 23604 12952 23656
rect 13176 23604 13228 23656
rect 13636 23647 13688 23656
rect 13636 23613 13670 23647
rect 13670 23613 13688 23647
rect 13636 23604 13688 23613
rect 16212 23604 16264 23656
rect 16764 23604 16816 23656
rect 9312 23536 9364 23588
rect 10232 23536 10284 23588
rect 4712 23468 4764 23520
rect 5816 23468 5868 23520
rect 8576 23468 8628 23520
rect 8944 23468 8996 23520
rect 10416 23468 10468 23520
rect 10784 23468 10836 23520
rect 10876 23468 10928 23520
rect 16948 23536 17000 23588
rect 16212 23468 16264 23520
rect 17224 23468 17276 23520
rect 18972 23511 19024 23520
rect 18972 23477 18981 23511
rect 18981 23477 19015 23511
rect 19015 23477 19024 23511
rect 18972 23468 19024 23477
rect 19708 23672 19760 23724
rect 19800 23715 19852 23724
rect 19800 23681 19809 23715
rect 19809 23681 19843 23715
rect 19843 23681 19852 23715
rect 19800 23672 19852 23681
rect 20720 23715 20772 23724
rect 20720 23681 20729 23715
rect 20729 23681 20763 23715
rect 20763 23681 20772 23715
rect 20720 23672 20772 23681
rect 22468 23672 22520 23724
rect 22836 23672 22888 23724
rect 19616 23647 19668 23656
rect 19616 23613 19625 23647
rect 19625 23613 19659 23647
rect 19659 23613 19668 23647
rect 19616 23604 19668 23613
rect 20076 23604 20128 23656
rect 20812 23647 20864 23656
rect 19892 23536 19944 23588
rect 20812 23613 20846 23647
rect 20846 23613 20864 23647
rect 20812 23604 20864 23613
rect 20444 23579 20496 23588
rect 20444 23545 20453 23579
rect 20453 23545 20487 23579
rect 20487 23545 20496 23579
rect 20444 23536 20496 23545
rect 23940 23604 23992 23656
rect 24676 23715 24728 23724
rect 24676 23681 24685 23715
rect 24685 23681 24719 23715
rect 24719 23681 24728 23715
rect 24676 23672 24728 23681
rect 26792 23740 26844 23792
rect 33232 23808 33284 23860
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 25688 23715 25740 23724
rect 25688 23681 25722 23715
rect 25722 23681 25740 23715
rect 25688 23672 25740 23681
rect 26976 23715 27028 23724
rect 26976 23681 26985 23715
rect 26985 23681 27019 23715
rect 27019 23681 27028 23715
rect 26976 23672 27028 23681
rect 33048 23740 33100 23792
rect 26056 23604 26108 23656
rect 27896 23715 27948 23724
rect 27896 23681 27905 23715
rect 27905 23681 27939 23715
rect 27939 23681 27948 23715
rect 27896 23672 27948 23681
rect 27988 23715 28040 23724
rect 27988 23681 28022 23715
rect 28022 23681 28040 23715
rect 27988 23672 28040 23681
rect 28908 23715 28960 23724
rect 28908 23681 28917 23715
rect 28917 23681 28951 23715
rect 28951 23681 28960 23715
rect 28908 23672 28960 23681
rect 29184 23715 29236 23724
rect 29184 23681 29218 23715
rect 29218 23681 29236 23715
rect 29184 23672 29236 23681
rect 23388 23579 23440 23588
rect 23388 23545 23397 23579
rect 23397 23545 23431 23579
rect 23431 23545 23440 23579
rect 23388 23536 23440 23545
rect 24032 23579 24084 23588
rect 24032 23545 24041 23579
rect 24041 23545 24075 23579
rect 24075 23545 24084 23579
rect 24032 23536 24084 23545
rect 25320 23579 25372 23588
rect 25320 23545 25329 23579
rect 25329 23545 25363 23579
rect 25363 23545 25372 23579
rect 25320 23536 25372 23545
rect 21548 23468 21600 23520
rect 22284 23468 22336 23520
rect 25136 23468 25188 23520
rect 27528 23604 27580 23656
rect 27620 23579 27672 23588
rect 27620 23545 27629 23579
rect 27629 23545 27663 23579
rect 27663 23545 27672 23579
rect 27620 23536 27672 23545
rect 27988 23468 28040 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 3792 23307 3844 23316
rect 3792 23273 3801 23307
rect 3801 23273 3835 23307
rect 3835 23273 3844 23307
rect 3792 23264 3844 23273
rect 3608 23196 3660 23248
rect 4068 23196 4120 23248
rect 4344 23196 4396 23248
rect 5448 23196 5500 23248
rect 4160 23128 4212 23180
rect 9864 23171 9916 23180
rect 9864 23137 9873 23171
rect 9873 23137 9907 23171
rect 9907 23137 9916 23171
rect 9864 23128 9916 23137
rect 10048 23171 10100 23180
rect 10048 23137 10057 23171
rect 10057 23137 10091 23171
rect 10091 23137 10100 23171
rect 10048 23128 10100 23137
rect 10968 23264 11020 23316
rect 11060 23264 11112 23316
rect 11520 23264 11572 23316
rect 11704 23307 11756 23316
rect 11704 23273 11713 23307
rect 11713 23273 11747 23307
rect 11747 23273 11756 23307
rect 11704 23264 11756 23273
rect 13176 23264 13228 23316
rect 13452 23264 13504 23316
rect 15660 23307 15712 23316
rect 15660 23273 15669 23307
rect 15669 23273 15703 23307
rect 15703 23273 15712 23307
rect 15660 23264 15712 23273
rect 11888 23196 11940 23248
rect 18604 23196 18656 23248
rect 20260 23196 20312 23248
rect 10600 23128 10652 23180
rect 16120 23128 16172 23180
rect 16488 23171 16540 23180
rect 16488 23137 16497 23171
rect 16497 23137 16531 23171
rect 16531 23137 16540 23171
rect 16488 23128 16540 23137
rect 19800 23171 19852 23180
rect 19800 23137 19809 23171
rect 19809 23137 19843 23171
rect 19843 23137 19852 23171
rect 19800 23128 19852 23137
rect 20076 23128 20128 23180
rect 20720 23171 20772 23180
rect 20720 23137 20729 23171
rect 20729 23137 20763 23171
rect 20763 23137 20772 23171
rect 20720 23128 20772 23137
rect 20812 23171 20864 23180
rect 20812 23137 20846 23171
rect 20846 23137 20864 23171
rect 21456 23264 21508 23316
rect 20812 23128 20864 23137
rect 5448 23060 5500 23112
rect 10784 23103 10836 23112
rect 10784 23069 10793 23103
rect 10793 23069 10827 23103
rect 10827 23069 10836 23103
rect 10784 23060 10836 23069
rect 11060 23103 11112 23112
rect 11060 23069 11069 23103
rect 11069 23069 11103 23103
rect 11103 23069 11112 23103
rect 11060 23060 11112 23069
rect 14464 23103 14516 23112
rect 14464 23069 14473 23103
rect 14473 23069 14507 23103
rect 14507 23069 14516 23103
rect 14464 23060 14516 23069
rect 4712 22992 4764 23044
rect 7564 22992 7616 23044
rect 4068 22924 4120 22976
rect 7104 22924 7156 22976
rect 8116 22924 8168 22976
rect 14280 22967 14332 22976
rect 14280 22933 14289 22967
rect 14289 22933 14323 22967
rect 14323 22933 14332 22967
rect 14280 22924 14332 22933
rect 18972 23103 19024 23112
rect 18972 23069 18981 23103
rect 18981 23069 19015 23103
rect 19015 23069 19024 23103
rect 18972 23060 19024 23069
rect 19616 23060 19668 23112
rect 20996 23103 21048 23112
rect 20996 23069 21005 23103
rect 21005 23069 21039 23103
rect 21039 23069 21048 23103
rect 20996 23060 21048 23069
rect 16488 22992 16540 23044
rect 16212 22924 16264 22976
rect 18788 22967 18840 22976
rect 18788 22933 18797 22967
rect 18797 22933 18831 22967
rect 18831 22933 18840 22967
rect 18788 22924 18840 22933
rect 19616 22924 19668 22976
rect 21456 22924 21508 22976
rect 21640 22967 21692 22976
rect 21640 22933 21649 22967
rect 21649 22933 21683 22967
rect 21683 22933 21692 22967
rect 21640 22924 21692 22933
rect 23756 22967 23808 22976
rect 23756 22933 23765 22967
rect 23765 22933 23799 22967
rect 23799 22933 23808 22967
rect 23756 22924 23808 22933
rect 26424 23128 26476 23180
rect 26516 23171 26568 23180
rect 26516 23137 26525 23171
rect 26525 23137 26559 23171
rect 26559 23137 26568 23171
rect 26516 23128 26568 23137
rect 29184 23307 29236 23316
rect 29184 23273 29193 23307
rect 29193 23273 29227 23307
rect 29227 23273 29236 23307
rect 29184 23264 29236 23273
rect 31668 23196 31720 23248
rect 32864 23196 32916 23248
rect 24860 23060 24912 23112
rect 25688 23060 25740 23112
rect 27620 23103 27672 23112
rect 27620 23069 27629 23103
rect 27629 23069 27663 23103
rect 27663 23069 27672 23103
rect 27620 23060 27672 23069
rect 27804 23060 27856 23112
rect 28908 23060 28960 23112
rect 25320 22992 25372 23044
rect 24676 22924 24728 22976
rect 25504 22924 25556 22976
rect 26240 22967 26292 22976
rect 26240 22933 26249 22967
rect 26249 22933 26283 22967
rect 26283 22933 26292 22967
rect 26240 22924 26292 22933
rect 28356 22924 28408 22976
rect 29920 23103 29972 23112
rect 29920 23069 29929 23103
rect 29929 23069 29963 23103
rect 29963 23069 29972 23103
rect 29920 23060 29972 23069
rect 32404 23171 32456 23180
rect 32404 23137 32413 23171
rect 32413 23137 32447 23171
rect 32447 23137 32456 23171
rect 32404 23128 32456 23137
rect 30656 23060 30708 23112
rect 30196 22924 30248 22976
rect 30564 22967 30616 22976
rect 30564 22933 30573 22967
rect 30573 22933 30607 22967
rect 30607 22933 30616 22967
rect 30564 22924 30616 22933
rect 30656 22924 30708 22976
rect 30932 22967 30984 22976
rect 30932 22933 30941 22967
rect 30941 22933 30975 22967
rect 30975 22933 30984 22967
rect 30932 22924 30984 22933
rect 31852 22992 31904 23044
rect 31392 22924 31444 22976
rect 32220 22924 32272 22976
rect 33232 23060 33284 23112
rect 33784 22992 33836 23044
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 4344 22720 4396 22772
rect 4804 22720 4856 22772
rect 5448 22763 5500 22772
rect 5448 22729 5457 22763
rect 5457 22729 5491 22763
rect 5491 22729 5500 22763
rect 5448 22720 5500 22729
rect 19892 22763 19944 22772
rect 19892 22729 19901 22763
rect 19901 22729 19935 22763
rect 19935 22729 19944 22763
rect 19892 22720 19944 22729
rect 20812 22720 20864 22772
rect 21088 22720 21140 22772
rect 24860 22720 24912 22772
rect 27620 22720 27672 22772
rect 30472 22720 30524 22772
rect 30932 22720 30984 22772
rect 32312 22763 32364 22772
rect 32312 22729 32321 22763
rect 32321 22729 32355 22763
rect 32355 22729 32364 22763
rect 32312 22720 32364 22729
rect 32404 22720 32456 22772
rect 33784 22763 33836 22772
rect 33784 22729 33793 22763
rect 33793 22729 33827 22763
rect 33827 22729 33836 22763
rect 33784 22720 33836 22729
rect 7656 22652 7708 22704
rect 2964 22584 3016 22636
rect 4068 22627 4120 22636
rect 4068 22593 4077 22627
rect 4077 22593 4111 22627
rect 4111 22593 4120 22627
rect 4068 22584 4120 22593
rect 4620 22584 4672 22636
rect 7564 22627 7616 22636
rect 7564 22593 7573 22627
rect 7573 22593 7607 22627
rect 7607 22593 7616 22627
rect 8576 22652 8628 22704
rect 7564 22584 7616 22593
rect 7840 22627 7892 22636
rect 7840 22593 7874 22627
rect 7874 22593 7892 22627
rect 7840 22584 7892 22593
rect 8392 22584 8444 22636
rect 10600 22584 10652 22636
rect 14280 22652 14332 22704
rect 18788 22695 18840 22704
rect 18788 22661 18822 22695
rect 18822 22661 18840 22695
rect 18788 22652 18840 22661
rect 23756 22652 23808 22704
rect 12532 22627 12584 22636
rect 12532 22593 12541 22627
rect 12541 22593 12575 22627
rect 12575 22593 12584 22627
rect 12532 22584 12584 22593
rect 13452 22627 13504 22636
rect 13452 22593 13461 22627
rect 13461 22593 13495 22627
rect 13495 22593 13504 22627
rect 13452 22584 13504 22593
rect 13636 22584 13688 22636
rect 15016 22584 15068 22636
rect 22836 22584 22888 22636
rect 27712 22652 27764 22704
rect 28356 22695 28408 22704
rect 28356 22661 28365 22695
rect 28365 22661 28399 22695
rect 28399 22661 28408 22695
rect 28356 22652 28408 22661
rect 25964 22584 26016 22636
rect 26516 22584 26568 22636
rect 940 22448 992 22500
rect 12624 22516 12676 22568
rect 12900 22516 12952 22568
rect 13176 22491 13228 22500
rect 13176 22457 13185 22491
rect 13185 22457 13219 22491
rect 13219 22457 13228 22491
rect 13176 22448 13228 22457
rect 3884 22380 3936 22432
rect 4436 22380 4488 22432
rect 9036 22423 9088 22432
rect 9036 22389 9045 22423
rect 9045 22389 9079 22423
rect 9079 22389 9088 22423
rect 9036 22380 9088 22389
rect 13728 22559 13780 22568
rect 13728 22525 13737 22559
rect 13737 22525 13771 22559
rect 13771 22525 13780 22559
rect 13728 22516 13780 22525
rect 14280 22448 14332 22500
rect 14372 22423 14424 22432
rect 14372 22389 14381 22423
rect 14381 22389 14415 22423
rect 14415 22389 14424 22423
rect 14372 22380 14424 22389
rect 16764 22380 16816 22432
rect 17408 22380 17460 22432
rect 17868 22380 17920 22432
rect 23112 22516 23164 22568
rect 28448 22559 28500 22568
rect 28448 22525 28457 22559
rect 28457 22525 28491 22559
rect 28491 22525 28500 22559
rect 28448 22516 28500 22525
rect 30840 22584 30892 22636
rect 30564 22516 30616 22568
rect 30932 22516 30984 22568
rect 32220 22584 32272 22636
rect 32312 22627 32364 22636
rect 32312 22593 32321 22627
rect 32321 22593 32355 22627
rect 32355 22593 32364 22627
rect 32312 22584 32364 22593
rect 32496 22584 32548 22636
rect 32864 22627 32916 22636
rect 32864 22593 32873 22627
rect 32873 22593 32907 22627
rect 32907 22593 32916 22627
rect 32864 22584 32916 22593
rect 33232 22584 33284 22636
rect 33140 22559 33192 22568
rect 33140 22525 33149 22559
rect 33149 22525 33183 22559
rect 33183 22525 33192 22559
rect 33140 22516 33192 22525
rect 31852 22448 31904 22500
rect 32496 22448 32548 22500
rect 21180 22380 21232 22432
rect 25596 22380 25648 22432
rect 31668 22423 31720 22432
rect 31668 22389 31677 22423
rect 31677 22389 31711 22423
rect 31711 22389 31720 22423
rect 31668 22380 31720 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 4620 22219 4672 22228
rect 4620 22185 4629 22219
rect 4629 22185 4663 22219
rect 4663 22185 4672 22219
rect 4620 22176 4672 22185
rect 7840 22176 7892 22228
rect 10140 22176 10192 22228
rect 2964 22108 3016 22160
rect 6920 22151 6972 22160
rect 6920 22117 6929 22151
rect 6929 22117 6963 22151
rect 6963 22117 6972 22151
rect 6920 22108 6972 22117
rect 1492 21972 1544 22024
rect 4160 22040 4212 22092
rect 4804 22015 4856 22024
rect 4804 21981 4813 22015
rect 4813 21981 4847 22015
rect 4847 21981 4856 22015
rect 4804 21972 4856 21981
rect 8300 22040 8352 22092
rect 8576 22040 8628 22092
rect 12624 22176 12676 22228
rect 14464 22176 14516 22228
rect 14740 22176 14792 22228
rect 17868 22176 17920 22228
rect 26240 22176 26292 22228
rect 31392 22176 31444 22228
rect 32312 22176 32364 22228
rect 11980 21972 12032 22024
rect 16488 22108 16540 22160
rect 32680 22108 32732 22160
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 16212 22083 16264 22092
rect 16212 22049 16221 22083
rect 16221 22049 16255 22083
rect 16255 22049 16264 22083
rect 16212 22040 16264 22049
rect 16764 22040 16816 22092
rect 16948 22040 17000 22092
rect 17132 22083 17184 22092
rect 17132 22049 17141 22083
rect 17141 22049 17175 22083
rect 17175 22049 17184 22083
rect 17132 22040 17184 22049
rect 17224 22083 17276 22092
rect 17224 22049 17258 22083
rect 17258 22049 17276 22083
rect 17224 22040 17276 22049
rect 17592 22040 17644 22092
rect 20168 22040 20220 22092
rect 21180 22040 21232 22092
rect 23112 22040 23164 22092
rect 25596 22083 25648 22092
rect 25596 22049 25605 22083
rect 25605 22049 25639 22083
rect 25639 22049 25648 22083
rect 25596 22040 25648 22049
rect 30748 22040 30800 22092
rect 13636 21972 13688 22024
rect 14280 21972 14332 22024
rect 21272 22015 21324 22024
rect 21272 21981 21281 22015
rect 21281 21981 21315 22015
rect 21315 21981 21324 22015
rect 21272 21972 21324 21981
rect 25504 22015 25556 22024
rect 25504 21981 25513 22015
rect 25513 21981 25547 22015
rect 25547 21981 25556 22015
rect 25504 21972 25556 21981
rect 30472 22015 30524 22024
rect 30472 21981 30481 22015
rect 30481 21981 30515 22015
rect 30515 21981 30524 22015
rect 30472 21972 30524 21981
rect 1952 21904 2004 21956
rect 7380 21904 7432 21956
rect 9036 21904 9088 21956
rect 9312 21904 9364 21956
rect 9680 21904 9732 21956
rect 11796 21904 11848 21956
rect 13084 21904 13136 21956
rect 2964 21879 3016 21888
rect 2964 21845 2973 21879
rect 2973 21845 3007 21879
rect 3007 21845 3016 21879
rect 2964 21836 3016 21845
rect 4804 21836 4856 21888
rect 5264 21836 5316 21888
rect 7012 21836 7064 21888
rect 7840 21836 7892 21888
rect 8484 21836 8536 21888
rect 10784 21879 10836 21888
rect 10784 21845 10793 21879
rect 10793 21845 10827 21879
rect 10827 21845 10836 21879
rect 10784 21836 10836 21845
rect 12900 21879 12952 21888
rect 12900 21845 12909 21879
rect 12909 21845 12943 21879
rect 12943 21845 12952 21879
rect 12900 21836 12952 21845
rect 13268 21836 13320 21888
rect 13452 21836 13504 21888
rect 15016 21836 15068 21888
rect 17040 21836 17092 21888
rect 17132 21836 17184 21888
rect 22192 21836 22244 21888
rect 30656 21904 30708 21956
rect 30748 21904 30800 21956
rect 32404 21972 32456 22024
rect 33140 21972 33192 22024
rect 30564 21879 30616 21888
rect 30564 21845 30573 21879
rect 30573 21845 30607 21879
rect 30607 21845 30616 21879
rect 30564 21836 30616 21845
rect 30840 21879 30892 21888
rect 30840 21845 30849 21879
rect 30849 21845 30883 21879
rect 30883 21845 30892 21879
rect 30840 21836 30892 21845
rect 32128 21879 32180 21888
rect 32128 21845 32137 21879
rect 32137 21845 32171 21879
rect 32171 21845 32180 21879
rect 32128 21836 32180 21845
rect 32588 21879 32640 21888
rect 32588 21845 32597 21879
rect 32597 21845 32631 21879
rect 32631 21845 32640 21879
rect 32588 21836 32640 21845
rect 33232 21836 33284 21888
rect 33416 21879 33468 21888
rect 33416 21845 33425 21879
rect 33425 21845 33459 21879
rect 33459 21845 33468 21879
rect 33416 21836 33468 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 1952 21675 2004 21684
rect 1952 21641 1961 21675
rect 1961 21641 1995 21675
rect 1995 21641 2004 21675
rect 1952 21632 2004 21641
rect 2780 21632 2832 21684
rect 3240 21632 3292 21684
rect 6184 21675 6236 21684
rect 6184 21641 6193 21675
rect 6193 21641 6227 21675
rect 6227 21641 6236 21675
rect 6184 21632 6236 21641
rect 7288 21632 7340 21684
rect 11796 21675 11848 21684
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 11980 21632 12032 21684
rect 15016 21632 15068 21684
rect 4068 21564 4120 21616
rect 2964 21496 3016 21548
rect 3148 21428 3200 21480
rect 5264 21539 5316 21548
rect 5264 21505 5273 21539
rect 5273 21505 5307 21539
rect 5307 21505 5316 21539
rect 5264 21496 5316 21505
rect 7196 21539 7248 21548
rect 7196 21505 7205 21539
rect 7205 21505 7239 21539
rect 7239 21505 7248 21539
rect 7196 21496 7248 21505
rect 7380 21496 7432 21548
rect 5448 21428 5500 21480
rect 6184 21428 6236 21480
rect 8024 21539 8076 21548
rect 8024 21505 8033 21539
rect 8033 21505 8067 21539
rect 8067 21505 8076 21539
rect 8024 21496 8076 21505
rect 8668 21428 8720 21480
rect 10784 21564 10836 21616
rect 8944 21496 8996 21548
rect 9128 21496 9180 21548
rect 9680 21496 9732 21548
rect 14740 21564 14792 21616
rect 17776 21632 17828 21684
rect 21272 21632 21324 21684
rect 22192 21675 22244 21684
rect 20076 21564 20128 21616
rect 22192 21641 22201 21675
rect 22201 21641 22235 21675
rect 22235 21641 22244 21675
rect 22192 21632 22244 21641
rect 22284 21675 22336 21684
rect 22284 21641 22293 21675
rect 22293 21641 22327 21675
rect 22327 21641 22336 21675
rect 22284 21632 22336 21641
rect 26332 21632 26384 21684
rect 28448 21632 28500 21684
rect 12900 21496 12952 21548
rect 16856 21496 16908 21548
rect 16948 21539 17000 21548
rect 16948 21505 16957 21539
rect 16957 21505 16991 21539
rect 16991 21505 17000 21539
rect 16948 21496 17000 21505
rect 17040 21539 17092 21548
rect 17040 21505 17049 21539
rect 17049 21505 17083 21539
rect 17083 21505 17092 21539
rect 17040 21496 17092 21505
rect 11520 21428 11572 21480
rect 14280 21428 14332 21480
rect 4620 21360 4672 21412
rect 4804 21360 4856 21412
rect 6000 21360 6052 21412
rect 9312 21403 9364 21412
rect 9312 21369 9321 21403
rect 9321 21369 9355 21403
rect 9355 21369 9364 21403
rect 9312 21360 9364 21369
rect 14188 21360 14240 21412
rect 16028 21471 16080 21480
rect 16028 21437 16037 21471
rect 16037 21437 16071 21471
rect 16071 21437 16080 21471
rect 16028 21428 16080 21437
rect 16488 21428 16540 21480
rect 19708 21496 19760 21548
rect 5448 21292 5500 21344
rect 5632 21292 5684 21344
rect 6920 21292 6972 21344
rect 7564 21335 7616 21344
rect 7564 21301 7573 21335
rect 7573 21301 7607 21335
rect 7607 21301 7616 21335
rect 7564 21292 7616 21301
rect 9772 21292 9824 21344
rect 13728 21292 13780 21344
rect 15476 21292 15528 21344
rect 22008 21496 22060 21548
rect 20720 21471 20772 21480
rect 20720 21437 20729 21471
rect 20729 21437 20763 21471
rect 20763 21437 20772 21471
rect 20720 21428 20772 21437
rect 20996 21471 21048 21480
rect 20996 21437 21005 21471
rect 21005 21437 21039 21471
rect 21039 21437 21048 21471
rect 20996 21428 21048 21437
rect 25320 21564 25372 21616
rect 23112 21539 23164 21548
rect 23112 21505 23121 21539
rect 23121 21505 23155 21539
rect 23155 21505 23164 21539
rect 23112 21496 23164 21505
rect 23388 21539 23440 21548
rect 23388 21505 23422 21539
rect 23422 21505 23440 21539
rect 23388 21496 23440 21505
rect 24492 21496 24544 21548
rect 26976 21496 27028 21548
rect 28632 21539 28684 21548
rect 28632 21505 28641 21539
rect 28641 21505 28675 21539
rect 28675 21505 28684 21539
rect 28632 21496 28684 21505
rect 33324 21539 33376 21548
rect 33324 21505 33333 21539
rect 33333 21505 33367 21539
rect 33367 21505 33376 21539
rect 33324 21496 33376 21505
rect 18144 21360 18196 21412
rect 22836 21428 22888 21480
rect 21640 21360 21692 21412
rect 20352 21292 20404 21344
rect 21456 21335 21508 21344
rect 21456 21301 21465 21335
rect 21465 21301 21499 21335
rect 21499 21301 21508 21335
rect 21456 21292 21508 21301
rect 22928 21292 22980 21344
rect 30840 21428 30892 21480
rect 24492 21335 24544 21344
rect 24492 21301 24501 21335
rect 24501 21301 24535 21335
rect 24535 21301 24544 21335
rect 24492 21292 24544 21301
rect 24584 21335 24636 21344
rect 24584 21301 24593 21335
rect 24593 21301 24627 21335
rect 24627 21301 24636 21335
rect 24584 21292 24636 21301
rect 29736 21292 29788 21344
rect 31024 21292 31076 21344
rect 31392 21292 31444 21344
rect 33232 21292 33284 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2688 21088 2740 21140
rect 8668 21088 8720 21140
rect 9864 21131 9916 21140
rect 9864 21097 9873 21131
rect 9873 21097 9907 21131
rect 9907 21097 9916 21131
rect 9864 21088 9916 21097
rect 9680 21020 9732 21072
rect 2964 20884 3016 20936
rect 3976 20952 4028 21004
rect 4620 20995 4672 21004
rect 4620 20961 4629 20995
rect 4629 20961 4663 20995
rect 4663 20961 4672 20995
rect 4620 20952 4672 20961
rect 5264 20995 5316 21004
rect 5264 20961 5273 20995
rect 5273 20961 5307 20995
rect 5307 20961 5316 20995
rect 5264 20952 5316 20961
rect 5356 20952 5408 21004
rect 5632 20995 5684 21004
rect 5632 20961 5666 20995
rect 5666 20961 5684 20995
rect 5632 20952 5684 20961
rect 7196 20995 7248 21004
rect 7196 20961 7205 20995
rect 7205 20961 7239 20995
rect 7239 20961 7248 20995
rect 7196 20952 7248 20961
rect 9588 20952 9640 21004
rect 10876 21063 10928 21072
rect 10876 21029 10885 21063
rect 10885 21029 10919 21063
rect 10919 21029 10928 21063
rect 10876 21020 10928 21029
rect 2688 20859 2740 20868
rect 2688 20825 2697 20859
rect 2697 20825 2731 20859
rect 2731 20825 2740 20859
rect 2688 20816 2740 20825
rect 2780 20816 2832 20868
rect 2044 20748 2096 20800
rect 3424 20791 3476 20800
rect 3424 20757 3433 20791
rect 3433 20757 3467 20791
rect 3467 20757 3476 20791
rect 3424 20748 3476 20757
rect 4068 20884 4120 20936
rect 5816 20927 5868 20936
rect 5816 20893 5825 20927
rect 5825 20893 5859 20927
rect 5859 20893 5868 20927
rect 5816 20884 5868 20893
rect 6920 20927 6972 20936
rect 6920 20893 6929 20927
rect 6929 20893 6963 20927
rect 6963 20893 6972 20927
rect 6920 20884 6972 20893
rect 7012 20927 7064 20936
rect 7012 20893 7021 20927
rect 7021 20893 7055 20927
rect 7055 20893 7064 20927
rect 7012 20884 7064 20893
rect 7564 20884 7616 20936
rect 8024 20884 8076 20936
rect 11244 20952 11296 21004
rect 9864 20884 9916 20936
rect 11428 20995 11480 21004
rect 11428 20961 11437 20995
rect 11437 20961 11471 20995
rect 11471 20961 11480 20995
rect 11428 20952 11480 20961
rect 11520 20995 11572 21004
rect 11520 20961 11529 20995
rect 11529 20961 11563 20995
rect 11563 20961 11572 20995
rect 14372 21020 14424 21072
rect 14188 20995 14240 21004
rect 11520 20952 11572 20961
rect 12072 20884 12124 20936
rect 14188 20961 14197 20995
rect 14197 20961 14231 20995
rect 14231 20961 14240 20995
rect 14188 20952 14240 20961
rect 14280 20884 14332 20936
rect 14556 21088 14608 21140
rect 4436 20816 4488 20868
rect 3884 20748 3936 20800
rect 4620 20748 4672 20800
rect 7380 20859 7432 20868
rect 7380 20825 7389 20859
rect 7389 20825 7423 20859
rect 7423 20825 7432 20859
rect 7380 20816 7432 20825
rect 9312 20816 9364 20868
rect 9772 20859 9824 20868
rect 9772 20825 9781 20859
rect 9781 20825 9815 20859
rect 9815 20825 9824 20859
rect 9772 20816 9824 20825
rect 10508 20859 10560 20868
rect 10508 20825 10517 20859
rect 10517 20825 10551 20859
rect 10551 20825 10560 20859
rect 10508 20816 10560 20825
rect 11888 20816 11940 20868
rect 13452 20859 13504 20868
rect 13452 20825 13461 20859
rect 13461 20825 13495 20859
rect 13495 20825 13504 20859
rect 13452 20816 13504 20825
rect 14556 20816 14608 20868
rect 14924 20927 14976 20936
rect 14924 20893 14933 20927
rect 14933 20893 14967 20927
rect 14967 20893 14976 20927
rect 14924 20884 14976 20893
rect 15752 20884 15804 20936
rect 16856 21088 16908 21140
rect 16948 21088 17000 21140
rect 17408 21088 17460 21140
rect 17776 21088 17828 21140
rect 19708 21131 19760 21140
rect 19708 21097 19717 21131
rect 19717 21097 19751 21131
rect 19751 21097 19760 21131
rect 19708 21088 19760 21097
rect 20352 21131 20404 21140
rect 20352 21097 20361 21131
rect 20361 21097 20395 21131
rect 20395 21097 20404 21131
rect 20352 21088 20404 21097
rect 20996 21088 21048 21140
rect 17132 21063 17184 21072
rect 17132 21029 17141 21063
rect 17141 21029 17175 21063
rect 17175 21029 17184 21063
rect 17132 21020 17184 21029
rect 19432 21020 19484 21072
rect 20720 21020 20772 21072
rect 21180 21020 21232 21072
rect 17592 20952 17644 21004
rect 17868 20995 17920 21004
rect 17868 20961 17877 20995
rect 17877 20961 17911 20995
rect 17911 20961 17920 20995
rect 17868 20952 17920 20961
rect 18696 20952 18748 21004
rect 17408 20884 17460 20936
rect 5632 20748 5684 20800
rect 7288 20748 7340 20800
rect 8484 20748 8536 20800
rect 9588 20791 9640 20800
rect 9588 20757 9597 20791
rect 9597 20757 9631 20791
rect 9631 20757 9640 20791
rect 9588 20748 9640 20757
rect 11704 20791 11756 20800
rect 11704 20757 11713 20791
rect 11713 20757 11747 20791
rect 11747 20757 11756 20791
rect 11704 20748 11756 20757
rect 11796 20791 11848 20800
rect 11796 20757 11805 20791
rect 11805 20757 11839 20791
rect 11839 20757 11848 20791
rect 11796 20748 11848 20757
rect 13912 20791 13964 20800
rect 13912 20757 13921 20791
rect 13921 20757 13955 20791
rect 13955 20757 13964 20791
rect 13912 20748 13964 20757
rect 14832 20791 14884 20800
rect 14832 20757 14841 20791
rect 14841 20757 14875 20791
rect 14875 20757 14884 20791
rect 14832 20748 14884 20757
rect 15292 20816 15344 20868
rect 19708 20884 19760 20936
rect 19892 20927 19944 20936
rect 19892 20893 19901 20927
rect 19901 20893 19935 20927
rect 19935 20893 19944 20927
rect 19892 20884 19944 20893
rect 20076 20927 20128 20936
rect 20076 20893 20085 20927
rect 20085 20893 20119 20927
rect 20119 20893 20128 20927
rect 20076 20884 20128 20893
rect 21456 20952 21508 21004
rect 23388 21131 23440 21140
rect 23388 21097 23397 21131
rect 23397 21097 23431 21131
rect 23431 21097 23440 21131
rect 23388 21088 23440 21097
rect 27068 21088 27120 21140
rect 27988 21088 28040 21140
rect 28632 21088 28684 21140
rect 31208 21088 31260 21140
rect 31668 21088 31720 21140
rect 32036 21088 32088 21140
rect 25136 21063 25188 21072
rect 25136 21029 25145 21063
rect 25145 21029 25179 21063
rect 25179 21029 25188 21063
rect 25136 21020 25188 21029
rect 27160 21020 27212 21072
rect 31024 21020 31076 21072
rect 31760 21020 31812 21072
rect 33048 21020 33100 21072
rect 25964 20952 26016 21004
rect 17960 20816 18012 20868
rect 19616 20859 19668 20868
rect 19616 20825 19625 20859
rect 19625 20825 19659 20859
rect 19659 20825 19668 20859
rect 19616 20816 19668 20825
rect 20812 20884 20864 20936
rect 21180 20884 21232 20936
rect 24584 20884 24636 20936
rect 26608 20952 26660 21004
rect 26332 20884 26384 20936
rect 26792 20884 26844 20936
rect 27804 20952 27856 21004
rect 30748 20952 30800 21004
rect 30932 20995 30984 21004
rect 30932 20961 30941 20995
rect 30941 20961 30975 20995
rect 30975 20961 30984 20995
rect 30932 20952 30984 20961
rect 17592 20748 17644 20800
rect 17868 20748 17920 20800
rect 18144 20791 18196 20800
rect 18144 20757 18153 20791
rect 18153 20757 18187 20791
rect 18187 20757 18196 20791
rect 18144 20748 18196 20757
rect 18420 20748 18472 20800
rect 24308 20816 24360 20868
rect 24860 20816 24912 20868
rect 25228 20791 25280 20800
rect 25228 20757 25237 20791
rect 25237 20757 25271 20791
rect 25271 20757 25280 20791
rect 25228 20748 25280 20757
rect 25320 20791 25372 20800
rect 25320 20757 25329 20791
rect 25329 20757 25363 20791
rect 25363 20757 25372 20791
rect 25320 20748 25372 20757
rect 26148 20748 26200 20800
rect 26516 20748 26568 20800
rect 29736 20927 29788 20936
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 29736 20884 29788 20893
rect 30564 20884 30616 20936
rect 31208 20884 31260 20936
rect 32128 20927 32180 20936
rect 32128 20893 32137 20927
rect 32137 20893 32171 20927
rect 32171 20893 32180 20927
rect 32128 20884 32180 20893
rect 33140 20995 33192 21004
rect 33140 20961 33149 20995
rect 33149 20961 33183 20995
rect 33183 20961 33192 20995
rect 33140 20952 33192 20961
rect 27160 20816 27212 20868
rect 28080 20748 28132 20800
rect 32036 20816 32088 20868
rect 33232 20884 33284 20936
rect 30380 20748 30432 20800
rect 31300 20748 31352 20800
rect 31944 20791 31996 20800
rect 31944 20757 31953 20791
rect 31953 20757 31987 20791
rect 31987 20757 31996 20791
rect 31944 20748 31996 20757
rect 36268 20816 36320 20868
rect 36360 20791 36412 20800
rect 36360 20757 36369 20791
rect 36369 20757 36403 20791
rect 36403 20757 36412 20791
rect 36360 20748 36412 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 2964 20544 3016 20596
rect 4436 20587 4488 20596
rect 4436 20553 4445 20587
rect 4445 20553 4479 20587
rect 4479 20553 4488 20587
rect 4436 20544 4488 20553
rect 7656 20544 7708 20596
rect 8760 20587 8812 20596
rect 8760 20553 8769 20587
rect 8769 20553 8803 20587
rect 8803 20553 8812 20587
rect 8760 20544 8812 20553
rect 15200 20544 15252 20596
rect 15292 20587 15344 20596
rect 15292 20553 15301 20587
rect 15301 20553 15335 20587
rect 15335 20553 15344 20587
rect 15292 20544 15344 20553
rect 18880 20544 18932 20596
rect 19340 20544 19392 20596
rect 19432 20587 19484 20596
rect 19432 20553 19441 20587
rect 19441 20553 19475 20587
rect 19475 20553 19484 20587
rect 19432 20544 19484 20553
rect 20076 20544 20128 20596
rect 22284 20587 22336 20596
rect 22284 20553 22293 20587
rect 22293 20553 22327 20587
rect 22327 20553 22336 20587
rect 22284 20544 22336 20553
rect 25872 20544 25924 20596
rect 27160 20544 27212 20596
rect 28080 20587 28132 20596
rect 28080 20553 28089 20587
rect 28089 20553 28123 20587
rect 28123 20553 28132 20587
rect 28080 20544 28132 20553
rect 29276 20544 29328 20596
rect 30656 20587 30708 20596
rect 30656 20553 30665 20587
rect 30665 20553 30699 20587
rect 30699 20553 30708 20587
rect 30656 20544 30708 20553
rect 32128 20544 32180 20596
rect 1492 20451 1544 20460
rect 1492 20417 1501 20451
rect 1501 20417 1535 20451
rect 1535 20417 1544 20451
rect 1492 20408 1544 20417
rect 1768 20451 1820 20460
rect 1768 20417 1802 20451
rect 1802 20417 1820 20451
rect 1768 20408 1820 20417
rect 3424 20476 3476 20528
rect 7288 20408 7340 20460
rect 8208 20408 8260 20460
rect 9312 20451 9364 20460
rect 9312 20417 9321 20451
rect 9321 20417 9355 20451
rect 9355 20417 9364 20451
rect 9312 20408 9364 20417
rect 10876 20451 10928 20460
rect 10876 20417 10885 20451
rect 10885 20417 10919 20451
rect 10919 20417 10928 20451
rect 10876 20408 10928 20417
rect 11796 20476 11848 20528
rect 11888 20476 11940 20528
rect 11244 20451 11296 20460
rect 11244 20417 11253 20451
rect 11253 20417 11287 20451
rect 11287 20417 11296 20451
rect 11244 20408 11296 20417
rect 12716 20451 12768 20460
rect 10508 20340 10560 20392
rect 11704 20340 11756 20392
rect 12716 20417 12725 20451
rect 12725 20417 12759 20451
rect 12759 20417 12768 20451
rect 12716 20408 12768 20417
rect 13360 20408 13412 20460
rect 14372 20451 14424 20460
rect 14372 20417 14381 20451
rect 14381 20417 14415 20451
rect 14415 20417 14424 20451
rect 14372 20408 14424 20417
rect 21824 20476 21876 20528
rect 15476 20451 15528 20460
rect 15476 20417 15485 20451
rect 15485 20417 15519 20451
rect 15519 20417 15528 20451
rect 15476 20408 15528 20417
rect 17408 20451 17460 20460
rect 17408 20417 17417 20451
rect 17417 20417 17451 20451
rect 17451 20417 17460 20451
rect 17408 20408 17460 20417
rect 14740 20340 14792 20392
rect 17132 20272 17184 20324
rect 17776 20451 17828 20460
rect 17776 20417 17785 20451
rect 17785 20417 17819 20451
rect 17819 20417 17828 20451
rect 17776 20408 17828 20417
rect 18236 20451 18288 20460
rect 18236 20417 18245 20451
rect 18245 20417 18279 20451
rect 18279 20417 18288 20451
rect 18236 20408 18288 20417
rect 19616 20408 19668 20460
rect 18604 20340 18656 20392
rect 21180 20272 21232 20324
rect 8300 20247 8352 20256
rect 8300 20213 8309 20247
rect 8309 20213 8343 20247
rect 8343 20213 8352 20247
rect 8300 20204 8352 20213
rect 9680 20204 9732 20256
rect 10416 20204 10468 20256
rect 10784 20204 10836 20256
rect 13728 20247 13780 20256
rect 13728 20213 13737 20247
rect 13737 20213 13771 20247
rect 13771 20213 13780 20247
rect 13728 20204 13780 20213
rect 13820 20204 13872 20256
rect 17500 20204 17552 20256
rect 17592 20204 17644 20256
rect 17868 20247 17920 20256
rect 17868 20213 17877 20247
rect 17877 20213 17911 20247
rect 17911 20213 17920 20247
rect 17868 20204 17920 20213
rect 21364 20204 21416 20256
rect 22284 20340 22336 20392
rect 22928 20340 22980 20392
rect 23572 20408 23624 20460
rect 24216 20408 24268 20460
rect 24308 20451 24360 20460
rect 24308 20417 24317 20451
rect 24317 20417 24351 20451
rect 24351 20417 24360 20451
rect 24308 20408 24360 20417
rect 24860 20408 24912 20460
rect 26240 20476 26292 20528
rect 26332 20519 26384 20528
rect 26332 20485 26341 20519
rect 26341 20485 26375 20519
rect 26375 20485 26384 20519
rect 26332 20476 26384 20485
rect 29184 20476 29236 20528
rect 30564 20476 30616 20528
rect 23296 20315 23348 20324
rect 23296 20281 23305 20315
rect 23305 20281 23339 20315
rect 23339 20281 23348 20315
rect 23296 20272 23348 20281
rect 30472 20408 30524 20460
rect 30932 20408 30984 20460
rect 31668 20451 31720 20460
rect 31668 20417 31677 20451
rect 31677 20417 31711 20451
rect 31711 20417 31720 20451
rect 31668 20408 31720 20417
rect 31852 20451 31904 20460
rect 31852 20417 31861 20451
rect 31861 20417 31895 20451
rect 31895 20417 31904 20451
rect 31852 20408 31904 20417
rect 32036 20408 32088 20460
rect 33140 20408 33192 20460
rect 30748 20383 30800 20392
rect 30748 20349 30757 20383
rect 30757 20349 30791 20383
rect 30791 20349 30800 20383
rect 30748 20340 30800 20349
rect 32128 20272 32180 20324
rect 24124 20247 24176 20256
rect 24124 20213 24133 20247
rect 24133 20213 24167 20247
rect 24167 20213 24176 20247
rect 24124 20204 24176 20213
rect 25228 20204 25280 20256
rect 30656 20204 30708 20256
rect 31852 20204 31904 20256
rect 34796 20204 34848 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 1768 20000 1820 20052
rect 7196 20000 7248 20052
rect 8484 20043 8536 20052
rect 8484 20009 8493 20043
rect 8493 20009 8527 20043
rect 8527 20009 8536 20043
rect 8484 20000 8536 20009
rect 10876 20000 10928 20052
rect 13360 20043 13412 20052
rect 13360 20009 13369 20043
rect 13369 20009 13403 20043
rect 13403 20009 13412 20043
rect 13360 20000 13412 20009
rect 13912 20000 13964 20052
rect 6644 19975 6696 19984
rect 6644 19941 6653 19975
rect 6653 19941 6687 19975
rect 6687 19941 6696 19975
rect 6644 19932 6696 19941
rect 7380 19932 7432 19984
rect 1584 19864 1636 19916
rect 11244 19932 11296 19984
rect 2044 19839 2096 19848
rect 2044 19805 2053 19839
rect 2053 19805 2087 19839
rect 2087 19805 2096 19839
rect 2044 19796 2096 19805
rect 7380 19796 7432 19848
rect 8300 19839 8352 19848
rect 8300 19805 8309 19839
rect 8309 19805 8343 19839
rect 8343 19805 8352 19839
rect 8300 19796 8352 19805
rect 9588 19796 9640 19848
rect 9680 19728 9732 19780
rect 4344 19660 4396 19712
rect 4620 19660 4672 19712
rect 5908 19660 5960 19712
rect 8116 19660 8168 19712
rect 13452 19864 13504 19916
rect 10416 19796 10468 19848
rect 14740 19864 14792 19916
rect 15200 19864 15252 19916
rect 23572 20043 23624 20052
rect 23572 20009 23581 20043
rect 23581 20009 23615 20043
rect 23615 20009 23624 20043
rect 23572 20000 23624 20009
rect 33324 20000 33376 20052
rect 30840 19932 30892 19984
rect 13820 19796 13872 19848
rect 14832 19796 14884 19848
rect 15108 19796 15160 19848
rect 16120 19796 16172 19848
rect 20996 19864 21048 19916
rect 21272 19796 21324 19848
rect 23664 19864 23716 19916
rect 30932 19864 30984 19916
rect 31668 19864 31720 19916
rect 32680 19864 32732 19916
rect 21364 19839 21416 19844
rect 21364 19805 21373 19839
rect 21373 19805 21407 19839
rect 21407 19805 21416 19839
rect 21364 19792 21416 19805
rect 12440 19728 12492 19780
rect 16028 19728 16080 19780
rect 20996 19728 21048 19780
rect 21548 19728 21600 19780
rect 22008 19728 22060 19780
rect 23388 19839 23440 19848
rect 23388 19805 23397 19839
rect 23397 19805 23431 19839
rect 23431 19805 23440 19839
rect 23388 19796 23440 19805
rect 28632 19796 28684 19848
rect 29920 19839 29972 19848
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 33048 19839 33100 19848
rect 33048 19805 33057 19839
rect 33057 19805 33091 19839
rect 33091 19805 33100 19839
rect 33048 19796 33100 19805
rect 34704 19728 34756 19780
rect 13728 19660 13780 19712
rect 15384 19660 15436 19712
rect 16304 19703 16356 19712
rect 16304 19669 16313 19703
rect 16313 19669 16347 19703
rect 16347 19669 16356 19703
rect 16304 19660 16356 19669
rect 20076 19703 20128 19712
rect 20076 19669 20085 19703
rect 20085 19669 20119 19703
rect 20119 19669 20128 19703
rect 20076 19660 20128 19669
rect 21272 19660 21324 19712
rect 21824 19660 21876 19712
rect 23112 19703 23164 19712
rect 23112 19669 23121 19703
rect 23121 19669 23155 19703
rect 23155 19669 23164 19703
rect 23112 19660 23164 19669
rect 26332 19660 26384 19712
rect 29736 19703 29788 19712
rect 29736 19669 29745 19703
rect 29745 19669 29779 19703
rect 29779 19669 29788 19703
rect 29736 19660 29788 19669
rect 33140 19703 33192 19712
rect 33140 19669 33149 19703
rect 33149 19669 33183 19703
rect 33183 19669 33192 19703
rect 33140 19660 33192 19669
rect 34612 19660 34664 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 12440 19456 12492 19508
rect 13084 19456 13136 19508
rect 14372 19456 14424 19508
rect 16028 19456 16080 19508
rect 16212 19456 16264 19508
rect 21272 19456 21324 19508
rect 21548 19456 21600 19508
rect 22008 19499 22060 19508
rect 22008 19465 22017 19499
rect 22017 19465 22051 19499
rect 22051 19465 22060 19499
rect 22008 19456 22060 19465
rect 25044 19456 25096 19508
rect 26056 19499 26108 19508
rect 26056 19465 26065 19499
rect 26065 19465 26099 19499
rect 26099 19465 26108 19499
rect 26056 19456 26108 19465
rect 35440 19456 35492 19508
rect 2964 19431 3016 19440
rect 2964 19397 2973 19431
rect 2973 19397 3007 19431
rect 3007 19397 3016 19431
rect 2964 19388 3016 19397
rect 2872 19363 2924 19372
rect 2872 19329 2881 19363
rect 2881 19329 2915 19363
rect 2915 19329 2924 19363
rect 2872 19320 2924 19329
rect 3608 19320 3660 19372
rect 14832 19388 14884 19440
rect 4344 19363 4396 19372
rect 4344 19329 4353 19363
rect 4353 19329 4387 19363
rect 4387 19329 4396 19363
rect 4344 19320 4396 19329
rect 4620 19320 4672 19372
rect 8300 19363 8352 19372
rect 8300 19329 8334 19363
rect 8334 19329 8352 19363
rect 8300 19320 8352 19329
rect 12900 19363 12952 19372
rect 12900 19329 12909 19363
rect 12909 19329 12943 19363
rect 12943 19329 12952 19363
rect 12900 19320 12952 19329
rect 2964 19252 3016 19304
rect 940 19116 992 19168
rect 2136 19116 2188 19168
rect 2688 19116 2740 19168
rect 4712 19116 4764 19168
rect 8024 19295 8076 19304
rect 8024 19261 8033 19295
rect 8033 19261 8067 19295
rect 8067 19261 8076 19295
rect 8024 19252 8076 19261
rect 9220 19252 9272 19304
rect 9036 19184 9088 19236
rect 12624 19184 12676 19236
rect 9220 19116 9272 19168
rect 9404 19159 9456 19168
rect 9404 19125 9413 19159
rect 9413 19125 9447 19159
rect 9447 19125 9456 19159
rect 9404 19116 9456 19125
rect 9864 19116 9916 19168
rect 10600 19116 10652 19168
rect 11980 19116 12032 19168
rect 12072 19159 12124 19168
rect 12072 19125 12081 19159
rect 12081 19125 12115 19159
rect 12115 19125 12124 19159
rect 12072 19116 12124 19125
rect 13084 19295 13136 19304
rect 13084 19261 13093 19295
rect 13093 19261 13127 19295
rect 13127 19261 13136 19295
rect 13084 19252 13136 19261
rect 13452 19252 13504 19304
rect 13820 19295 13872 19304
rect 13820 19261 13829 19295
rect 13829 19261 13863 19295
rect 13863 19261 13872 19295
rect 13820 19252 13872 19261
rect 13912 19295 13964 19304
rect 13912 19261 13946 19295
rect 13946 19261 13964 19295
rect 13912 19252 13964 19261
rect 14280 19252 14332 19304
rect 14648 19252 14700 19304
rect 15108 19252 15160 19304
rect 18144 19320 18196 19372
rect 19892 19320 19944 19372
rect 20812 19388 20864 19440
rect 20996 19388 21048 19440
rect 20076 19320 20128 19372
rect 16764 19252 16816 19304
rect 17040 19252 17092 19304
rect 17408 19252 17460 19304
rect 21548 19320 21600 19372
rect 24768 19388 24820 19440
rect 26332 19431 26384 19440
rect 26332 19397 26341 19431
rect 26341 19397 26375 19431
rect 26375 19397 26384 19431
rect 26332 19388 26384 19397
rect 29736 19431 29788 19440
rect 29736 19397 29770 19431
rect 29770 19397 29788 19431
rect 29736 19388 29788 19397
rect 34612 19388 34664 19440
rect 23388 19363 23440 19372
rect 23388 19329 23397 19363
rect 23397 19329 23431 19363
rect 23431 19329 23440 19363
rect 23388 19320 23440 19329
rect 24860 19320 24912 19372
rect 25412 19363 25464 19372
rect 25412 19329 25421 19363
rect 25421 19329 25455 19363
rect 25455 19329 25464 19363
rect 25412 19320 25464 19329
rect 25872 19363 25924 19372
rect 25872 19329 25881 19363
rect 25881 19329 25915 19363
rect 25915 19329 25924 19363
rect 25872 19320 25924 19329
rect 26976 19363 27028 19372
rect 26976 19329 26985 19363
rect 26985 19329 27019 19363
rect 27019 19329 27028 19363
rect 26976 19320 27028 19329
rect 27344 19320 27396 19372
rect 29552 19320 29604 19372
rect 21732 19252 21784 19304
rect 19340 19184 19392 19236
rect 21824 19184 21876 19236
rect 15200 19116 15252 19168
rect 17592 19116 17644 19168
rect 18052 19116 18104 19168
rect 20076 19116 20128 19168
rect 20168 19159 20220 19168
rect 20168 19125 20177 19159
rect 20177 19125 20211 19159
rect 20211 19125 20220 19159
rect 20168 19116 20220 19125
rect 20260 19116 20312 19168
rect 23296 19252 23348 19304
rect 25688 19252 25740 19304
rect 27068 19252 27120 19304
rect 27528 19252 27580 19304
rect 22008 19116 22060 19168
rect 23664 19159 23716 19168
rect 23664 19125 23673 19159
rect 23673 19125 23707 19159
rect 23707 19125 23716 19159
rect 23664 19116 23716 19125
rect 24952 19159 25004 19168
rect 24952 19125 24961 19159
rect 24961 19125 24995 19159
rect 24995 19125 25004 19159
rect 24952 19116 25004 19125
rect 25596 19116 25648 19168
rect 26424 19159 26476 19168
rect 26424 19125 26433 19159
rect 26433 19125 26467 19159
rect 26467 19125 26476 19159
rect 26424 19116 26476 19125
rect 28080 19252 28132 19304
rect 28540 19252 28592 19304
rect 28816 19295 28868 19304
rect 28816 19261 28825 19295
rect 28825 19261 28859 19295
rect 28859 19261 28868 19295
rect 28816 19252 28868 19261
rect 34152 19363 34204 19372
rect 34152 19329 34161 19363
rect 34161 19329 34195 19363
rect 34195 19329 34204 19363
rect 34152 19320 34204 19329
rect 35348 19320 35400 19372
rect 32404 19252 32456 19304
rect 28264 19116 28316 19168
rect 28356 19116 28408 19168
rect 30380 19116 30432 19168
rect 30840 19159 30892 19168
rect 30840 19125 30849 19159
rect 30849 19125 30883 19159
rect 30883 19125 30892 19159
rect 30840 19116 30892 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2872 18912 2924 18964
rect 4068 18776 4120 18828
rect 5264 18912 5316 18964
rect 6644 18912 6696 18964
rect 8024 18912 8076 18964
rect 8300 18912 8352 18964
rect 11244 18955 11296 18964
rect 11244 18921 11253 18955
rect 11253 18921 11287 18955
rect 11287 18921 11296 18955
rect 11244 18912 11296 18921
rect 7564 18776 7616 18828
rect 7932 18776 7984 18828
rect 9036 18776 9088 18828
rect 9404 18819 9456 18828
rect 9404 18785 9413 18819
rect 9413 18785 9447 18819
rect 9447 18785 9456 18819
rect 9404 18776 9456 18785
rect 9680 18776 9732 18828
rect 12900 18955 12952 18964
rect 12900 18921 12909 18955
rect 12909 18921 12943 18955
rect 12943 18921 12952 18955
rect 12900 18912 12952 18921
rect 16304 18912 16356 18964
rect 13176 18844 13228 18896
rect 14832 18819 14884 18828
rect 14832 18785 14841 18819
rect 14841 18785 14875 18819
rect 14875 18785 14884 18819
rect 14832 18776 14884 18785
rect 18236 18955 18288 18964
rect 18236 18921 18245 18955
rect 18245 18921 18279 18955
rect 18279 18921 18288 18955
rect 18236 18912 18288 18921
rect 16488 18844 16540 18896
rect 17040 18819 17092 18828
rect 17040 18785 17049 18819
rect 17049 18785 17083 18819
rect 17083 18785 17092 18819
rect 17040 18776 17092 18785
rect 1492 18708 1544 18760
rect 2136 18751 2188 18760
rect 2136 18717 2170 18751
rect 2170 18717 2188 18751
rect 2136 18708 2188 18717
rect 4528 18751 4580 18760
rect 4528 18717 4537 18751
rect 4537 18717 4571 18751
rect 4571 18717 4580 18751
rect 4528 18708 4580 18717
rect 5264 18751 5316 18760
rect 5264 18717 5273 18751
rect 5273 18717 5307 18751
rect 5307 18717 5316 18751
rect 5264 18708 5316 18717
rect 5448 18708 5500 18760
rect 5540 18751 5592 18760
rect 5540 18717 5549 18751
rect 5549 18717 5583 18751
rect 5583 18717 5592 18751
rect 5540 18708 5592 18717
rect 6184 18708 6236 18760
rect 9128 18751 9180 18760
rect 9128 18717 9137 18751
rect 9137 18717 9171 18751
rect 9171 18717 9180 18751
rect 9128 18708 9180 18717
rect 9220 18751 9272 18760
rect 9220 18717 9229 18751
rect 9229 18717 9263 18751
rect 9263 18717 9272 18751
rect 9220 18708 9272 18717
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 10508 18708 10560 18760
rect 10600 18751 10652 18760
rect 10600 18717 10609 18751
rect 10609 18717 10643 18751
rect 10643 18717 10652 18751
rect 10600 18708 10652 18717
rect 11520 18751 11572 18760
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 7932 18640 7984 18692
rect 9036 18640 9088 18692
rect 5540 18572 5592 18624
rect 5816 18572 5868 18624
rect 10600 18572 10652 18624
rect 13636 18708 13688 18760
rect 16580 18751 16632 18760
rect 16580 18717 16589 18751
rect 16589 18717 16623 18751
rect 16623 18717 16632 18751
rect 16580 18708 16632 18717
rect 17408 18751 17460 18760
rect 17408 18717 17442 18751
rect 17442 18717 17460 18751
rect 17408 18708 17460 18717
rect 17592 18751 17644 18760
rect 17592 18717 17601 18751
rect 17601 18717 17635 18751
rect 17635 18717 17644 18751
rect 17592 18708 17644 18717
rect 11888 18640 11940 18692
rect 11980 18640 12032 18692
rect 14280 18640 14332 18692
rect 15200 18640 15252 18692
rect 11704 18572 11756 18624
rect 18880 18844 18932 18896
rect 20260 18887 20312 18896
rect 20260 18853 20269 18887
rect 20269 18853 20303 18887
rect 20303 18853 20312 18887
rect 20260 18844 20312 18853
rect 21456 18955 21508 18964
rect 21456 18921 21465 18955
rect 21465 18921 21499 18955
rect 21499 18921 21508 18955
rect 21456 18912 21508 18921
rect 24216 18912 24268 18964
rect 26240 18955 26292 18964
rect 26240 18921 26249 18955
rect 26249 18921 26283 18955
rect 26283 18921 26292 18955
rect 26240 18912 26292 18921
rect 23848 18844 23900 18896
rect 20352 18776 20404 18828
rect 20812 18819 20864 18828
rect 20812 18785 20821 18819
rect 20821 18785 20855 18819
rect 20855 18785 20864 18819
rect 20812 18776 20864 18785
rect 23112 18776 23164 18828
rect 25044 18819 25096 18828
rect 25044 18785 25053 18819
rect 25053 18785 25087 18819
rect 25087 18785 25096 18819
rect 25044 18776 25096 18785
rect 25596 18819 25648 18828
rect 25596 18785 25605 18819
rect 25605 18785 25639 18819
rect 25639 18785 25648 18819
rect 25596 18776 25648 18785
rect 19340 18708 19392 18760
rect 19708 18708 19760 18760
rect 20536 18751 20588 18760
rect 20536 18717 20545 18751
rect 20545 18717 20579 18751
rect 20579 18717 20588 18751
rect 20536 18708 20588 18717
rect 21548 18708 21600 18760
rect 23572 18708 23624 18760
rect 24492 18708 24544 18760
rect 23204 18640 23256 18692
rect 24768 18708 24820 18760
rect 25320 18751 25372 18760
rect 25320 18717 25329 18751
rect 25329 18717 25363 18751
rect 25363 18717 25372 18751
rect 25320 18708 25372 18717
rect 26976 18751 27028 18760
rect 26976 18717 26985 18751
rect 26985 18717 27019 18751
rect 27019 18717 27028 18751
rect 26976 18708 27028 18717
rect 26148 18640 26200 18692
rect 27896 18776 27948 18828
rect 28080 18776 28132 18828
rect 29184 18955 29236 18964
rect 29184 18921 29193 18955
rect 29193 18921 29227 18955
rect 29227 18921 29236 18955
rect 29184 18912 29236 18921
rect 29920 18912 29972 18964
rect 30472 18912 30524 18964
rect 30380 18819 30432 18828
rect 30380 18785 30389 18819
rect 30389 18785 30423 18819
rect 30423 18785 30432 18819
rect 30380 18776 30432 18785
rect 32404 18819 32456 18828
rect 32404 18785 32413 18819
rect 32413 18785 32447 18819
rect 32447 18785 32456 18819
rect 32404 18776 32456 18785
rect 34152 18776 34204 18828
rect 27344 18751 27396 18760
rect 27344 18717 27353 18751
rect 27353 18717 27387 18751
rect 27387 18717 27396 18751
rect 27344 18708 27396 18717
rect 27528 18751 27580 18760
rect 27528 18717 27537 18751
rect 27537 18717 27571 18751
rect 27571 18717 27580 18751
rect 27528 18708 27580 18717
rect 28264 18751 28316 18760
rect 28264 18717 28273 18751
rect 28273 18717 28307 18751
rect 28307 18717 28316 18751
rect 28264 18708 28316 18717
rect 28356 18751 28408 18760
rect 28356 18717 28390 18751
rect 28390 18717 28408 18751
rect 28356 18708 28408 18717
rect 29828 18708 29880 18760
rect 20260 18572 20312 18624
rect 20536 18572 20588 18624
rect 23940 18572 23992 18624
rect 25320 18572 25372 18624
rect 30840 18708 30892 18760
rect 31576 18708 31628 18760
rect 34612 18708 34664 18760
rect 31208 18683 31260 18692
rect 31208 18649 31242 18683
rect 31242 18649 31260 18683
rect 31208 18640 31260 18649
rect 32220 18640 32272 18692
rect 31024 18572 31076 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 4988 18368 5040 18420
rect 5632 18368 5684 18420
rect 6368 18368 6420 18420
rect 2872 18300 2924 18352
rect 6092 18300 6144 18352
rect 7196 18368 7248 18420
rect 8208 18411 8260 18420
rect 8208 18377 8217 18411
rect 8217 18377 8251 18411
rect 8251 18377 8260 18411
rect 8208 18368 8260 18377
rect 9036 18411 9088 18420
rect 9036 18377 9045 18411
rect 9045 18377 9079 18411
rect 9079 18377 9088 18411
rect 9036 18368 9088 18377
rect 9128 18368 9180 18420
rect 10508 18368 10560 18420
rect 11152 18368 11204 18420
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 14004 18368 14056 18420
rect 15200 18411 15252 18420
rect 15200 18377 15209 18411
rect 15209 18377 15243 18411
rect 15243 18377 15252 18411
rect 15200 18368 15252 18377
rect 16488 18368 16540 18420
rect 17592 18368 17644 18420
rect 18512 18411 18564 18420
rect 18512 18377 18521 18411
rect 18521 18377 18555 18411
rect 18555 18377 18564 18411
rect 18512 18368 18564 18377
rect 8852 18300 8904 18352
rect 4068 18232 4120 18284
rect 4528 18275 4580 18284
rect 4528 18241 4537 18275
rect 4537 18241 4571 18275
rect 4571 18241 4580 18275
rect 4528 18232 4580 18241
rect 9220 18300 9272 18352
rect 9404 18232 9456 18284
rect 2688 18164 2740 18216
rect 2964 18207 3016 18216
rect 2964 18173 2973 18207
rect 2973 18173 3007 18207
rect 3007 18173 3016 18207
rect 2964 18164 3016 18173
rect 5080 18164 5132 18216
rect 5264 18207 5316 18216
rect 5264 18173 5273 18207
rect 5273 18173 5307 18207
rect 5307 18173 5316 18207
rect 5264 18164 5316 18173
rect 5448 18164 5500 18216
rect 6092 18164 6144 18216
rect 6368 18207 6420 18216
rect 6368 18173 6377 18207
rect 6377 18173 6411 18207
rect 6411 18173 6420 18207
rect 6368 18164 6420 18173
rect 6552 18207 6604 18216
rect 6552 18173 6561 18207
rect 6561 18173 6595 18207
rect 6595 18173 6604 18207
rect 6552 18164 6604 18173
rect 6920 18164 6972 18216
rect 7380 18207 7432 18216
rect 7380 18173 7414 18207
rect 7414 18173 7432 18207
rect 7380 18164 7432 18173
rect 9864 18232 9916 18284
rect 10416 18275 10468 18284
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10416 18232 10468 18241
rect 10508 18275 10560 18284
rect 10508 18241 10542 18275
rect 10542 18241 10560 18275
rect 10508 18232 10560 18241
rect 10692 18275 10744 18284
rect 10692 18241 10701 18275
rect 10701 18241 10735 18275
rect 10735 18241 10744 18275
rect 10692 18232 10744 18241
rect 12072 18275 12124 18284
rect 12072 18241 12081 18275
rect 12081 18241 12115 18275
rect 12115 18241 12124 18275
rect 12072 18232 12124 18241
rect 12900 18275 12952 18284
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 13820 18275 13872 18284
rect 13820 18241 13829 18275
rect 13829 18241 13863 18275
rect 13863 18241 13872 18275
rect 13820 18232 13872 18241
rect 13912 18275 13964 18284
rect 13912 18241 13946 18275
rect 13946 18241 13964 18275
rect 13912 18232 13964 18241
rect 15384 18275 15436 18284
rect 15384 18241 15393 18275
rect 15393 18241 15427 18275
rect 15427 18241 15436 18275
rect 15384 18232 15436 18241
rect 16304 18232 16356 18284
rect 17592 18275 17644 18284
rect 17592 18241 17601 18275
rect 17601 18241 17635 18275
rect 17635 18241 17644 18275
rect 17592 18232 17644 18241
rect 17868 18275 17920 18284
rect 17868 18241 17877 18275
rect 17877 18241 17911 18275
rect 17911 18241 17920 18275
rect 17868 18232 17920 18241
rect 21180 18411 21232 18420
rect 21180 18377 21189 18411
rect 21189 18377 21223 18411
rect 21223 18377 21232 18411
rect 21180 18368 21232 18377
rect 21640 18368 21692 18420
rect 25136 18368 25188 18420
rect 25412 18368 25464 18420
rect 28448 18368 28500 18420
rect 31208 18411 31260 18420
rect 31208 18377 31217 18411
rect 31217 18377 31251 18411
rect 31251 18377 31260 18411
rect 31208 18368 31260 18377
rect 32220 18411 32272 18420
rect 32220 18377 32229 18411
rect 32229 18377 32263 18411
rect 32263 18377 32272 18411
rect 32220 18368 32272 18377
rect 32404 18368 32456 18420
rect 35348 18411 35400 18420
rect 35348 18377 35357 18411
rect 35357 18377 35391 18411
rect 35391 18377 35400 18411
rect 35348 18368 35400 18377
rect 19340 18275 19392 18284
rect 19340 18241 19349 18275
rect 19349 18241 19383 18275
rect 19383 18241 19392 18275
rect 19340 18232 19392 18241
rect 20260 18275 20312 18284
rect 20260 18241 20269 18275
rect 20269 18241 20303 18275
rect 20303 18241 20312 18275
rect 20260 18232 20312 18241
rect 20536 18275 20588 18284
rect 20536 18241 20545 18275
rect 20545 18241 20579 18275
rect 20579 18241 20588 18275
rect 20536 18232 20588 18241
rect 9680 18207 9732 18216
rect 9680 18173 9689 18207
rect 9689 18173 9723 18207
rect 9723 18173 9732 18207
rect 9680 18164 9732 18173
rect 13176 18164 13228 18216
rect 14464 18164 14516 18216
rect 16580 18164 16632 18216
rect 16856 18207 16908 18216
rect 16856 18173 16865 18207
rect 16865 18173 16899 18207
rect 16899 18173 16908 18207
rect 16856 18164 16908 18173
rect 17408 18164 17460 18216
rect 19432 18164 19484 18216
rect 19708 18164 19760 18216
rect 4988 18139 5040 18148
rect 4988 18105 4997 18139
rect 4997 18105 5031 18139
rect 5031 18105 5040 18139
rect 4988 18096 5040 18105
rect 7012 18139 7064 18148
rect 7012 18105 7021 18139
rect 7021 18105 7055 18139
rect 7055 18105 7064 18139
rect 7012 18096 7064 18105
rect 10140 18139 10192 18148
rect 10140 18105 10149 18139
rect 10149 18105 10183 18139
rect 10183 18105 10192 18139
rect 10140 18096 10192 18105
rect 2044 18028 2096 18080
rect 4804 18028 4856 18080
rect 13636 18096 13688 18148
rect 12624 18028 12676 18080
rect 14556 18028 14608 18080
rect 18880 18096 18932 18148
rect 19984 18139 20036 18148
rect 19984 18105 19993 18139
rect 19993 18105 20027 18139
rect 20027 18105 20036 18139
rect 19984 18096 20036 18105
rect 18788 18071 18840 18080
rect 18788 18037 18797 18071
rect 18797 18037 18831 18071
rect 18831 18037 18840 18071
rect 18788 18028 18840 18037
rect 20352 18207 20404 18216
rect 20352 18173 20386 18207
rect 20386 18173 20404 18207
rect 20352 18164 20404 18173
rect 22100 18164 22152 18216
rect 22928 18275 22980 18284
rect 22928 18241 22937 18275
rect 22937 18241 22971 18275
rect 22971 18241 22980 18275
rect 22928 18232 22980 18241
rect 23204 18275 23256 18284
rect 23204 18241 23213 18275
rect 23213 18241 23247 18275
rect 23247 18241 23256 18275
rect 23204 18232 23256 18241
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 24216 18275 24268 18284
rect 24216 18241 24225 18275
rect 24225 18241 24259 18275
rect 24259 18241 24268 18275
rect 24216 18232 24268 18241
rect 25044 18232 25096 18284
rect 25964 18232 26016 18284
rect 21824 18071 21876 18080
rect 21824 18037 21833 18071
rect 21833 18037 21867 18071
rect 21867 18037 21876 18071
rect 21824 18028 21876 18037
rect 22744 18071 22796 18080
rect 22744 18037 22753 18071
rect 22753 18037 22787 18071
rect 22787 18037 22796 18071
rect 22744 18028 22796 18037
rect 23572 18164 23624 18216
rect 23664 18207 23716 18216
rect 23664 18173 23673 18207
rect 23673 18173 23707 18207
rect 23707 18173 23716 18207
rect 23664 18164 23716 18173
rect 23756 18164 23808 18216
rect 24032 18207 24084 18216
rect 24032 18173 24066 18207
rect 24066 18173 24084 18207
rect 24032 18164 24084 18173
rect 24860 18164 24912 18216
rect 26884 18164 26936 18216
rect 28540 18343 28592 18352
rect 28540 18309 28549 18343
rect 28549 18309 28583 18343
rect 28583 18309 28592 18343
rect 28540 18300 28592 18309
rect 31300 18300 31352 18352
rect 30380 18232 30432 18284
rect 25688 18028 25740 18080
rect 28632 18164 28684 18216
rect 27896 18096 27948 18148
rect 30564 18164 30616 18216
rect 30932 18207 30984 18216
rect 30932 18173 30941 18207
rect 30941 18173 30975 18207
rect 30975 18173 30984 18207
rect 30932 18164 30984 18173
rect 31392 18275 31444 18284
rect 31392 18241 31401 18275
rect 31401 18241 31435 18275
rect 31435 18241 31444 18275
rect 31392 18232 31444 18241
rect 32404 18275 32456 18284
rect 32404 18241 32413 18275
rect 32413 18241 32447 18275
rect 32447 18241 32456 18275
rect 32404 18232 32456 18241
rect 34704 18300 34756 18352
rect 33324 18275 33376 18284
rect 33324 18241 33358 18275
rect 33358 18241 33376 18275
rect 33324 18232 33376 18241
rect 35440 18232 35492 18284
rect 34520 18164 34572 18216
rect 34796 18164 34848 18216
rect 31392 18096 31444 18148
rect 28632 18028 28684 18080
rect 34704 18028 34756 18080
rect 35348 18028 35400 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 5080 17824 5132 17876
rect 5264 17824 5316 17876
rect 1492 17620 1544 17672
rect 2780 17620 2832 17672
rect 5632 17756 5684 17808
rect 6644 17799 6696 17808
rect 6644 17765 6653 17799
rect 6653 17765 6687 17799
rect 6687 17765 6696 17799
rect 6644 17756 6696 17765
rect 7748 17824 7800 17876
rect 9496 17824 9548 17876
rect 8024 17756 8076 17808
rect 10416 17824 10468 17876
rect 14648 17824 14700 17876
rect 22100 17867 22152 17876
rect 22100 17833 22109 17867
rect 22109 17833 22143 17867
rect 22143 17833 22152 17867
rect 22100 17824 22152 17833
rect 23848 17867 23900 17876
rect 23848 17833 23857 17867
rect 23857 17833 23891 17867
rect 23891 17833 23900 17867
rect 23848 17824 23900 17833
rect 25044 17824 25096 17876
rect 25136 17824 25188 17876
rect 1860 17552 1912 17604
rect 4068 17595 4120 17604
rect 4068 17561 4102 17595
rect 4102 17561 4120 17595
rect 4068 17552 4120 17561
rect 2872 17484 2924 17536
rect 6368 17688 6420 17740
rect 6920 17731 6972 17740
rect 6920 17697 6929 17731
rect 6929 17697 6963 17731
rect 6963 17697 6972 17731
rect 6920 17688 6972 17697
rect 7380 17688 7432 17740
rect 7012 17663 7064 17672
rect 7012 17629 7046 17663
rect 7046 17629 7064 17663
rect 7012 17620 7064 17629
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 7932 17620 7984 17672
rect 13084 17688 13136 17740
rect 14556 17731 14608 17740
rect 14556 17697 14565 17731
rect 14565 17697 14599 17731
rect 14599 17697 14608 17731
rect 14556 17688 14608 17697
rect 9588 17663 9640 17672
rect 9588 17629 9597 17663
rect 9597 17629 9631 17663
rect 9631 17629 9640 17663
rect 9588 17620 9640 17629
rect 10416 17620 10468 17672
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 10876 17620 10928 17629
rect 18788 17688 18840 17740
rect 17316 17620 17368 17672
rect 18880 17620 18932 17672
rect 19248 17663 19300 17672
rect 19248 17629 19257 17663
rect 19257 17629 19291 17663
rect 19291 17629 19300 17663
rect 19248 17620 19300 17629
rect 20812 17620 20864 17672
rect 22744 17663 22796 17672
rect 22744 17629 22778 17663
rect 22778 17629 22796 17663
rect 13544 17552 13596 17604
rect 16856 17552 16908 17604
rect 6552 17484 6604 17536
rect 6828 17484 6880 17536
rect 9312 17527 9364 17536
rect 9312 17493 9321 17527
rect 9321 17493 9355 17527
rect 9355 17493 9364 17527
rect 9312 17484 9364 17493
rect 9956 17484 10008 17536
rect 13452 17484 13504 17536
rect 17040 17527 17092 17536
rect 17040 17493 17049 17527
rect 17049 17493 17083 17527
rect 17083 17493 17092 17527
rect 17040 17484 17092 17493
rect 17592 17484 17644 17536
rect 20996 17595 21048 17604
rect 20996 17561 21030 17595
rect 21030 17561 21048 17595
rect 20996 17552 21048 17561
rect 22744 17620 22796 17629
rect 24952 17620 25004 17672
rect 25872 17663 25924 17672
rect 25872 17629 25881 17663
rect 25881 17629 25915 17663
rect 25915 17629 25924 17663
rect 25872 17620 25924 17629
rect 30472 17824 30524 17876
rect 33324 17824 33376 17876
rect 22652 17552 22704 17604
rect 24860 17552 24912 17604
rect 28356 17620 28408 17672
rect 29184 17688 29236 17740
rect 29552 17731 29604 17740
rect 29552 17697 29561 17731
rect 29561 17697 29595 17731
rect 29595 17697 29604 17731
rect 29552 17688 29604 17697
rect 30656 17620 30708 17672
rect 33600 17620 33652 17672
rect 20628 17527 20680 17536
rect 20628 17493 20637 17527
rect 20637 17493 20671 17527
rect 20671 17493 20680 17527
rect 20628 17484 20680 17493
rect 26240 17595 26292 17604
rect 26240 17561 26274 17595
rect 26274 17561 26292 17595
rect 26240 17552 26292 17561
rect 26424 17552 26476 17604
rect 29460 17552 29512 17604
rect 28172 17484 28224 17536
rect 30196 17484 30248 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 1860 17323 1912 17332
rect 1860 17289 1869 17323
rect 1869 17289 1903 17323
rect 1903 17289 1912 17323
rect 1860 17280 1912 17289
rect 4068 17280 4120 17332
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 4712 17280 4764 17332
rect 5264 17280 5316 17332
rect 7104 17280 7156 17332
rect 9680 17280 9732 17332
rect 10876 17280 10928 17332
rect 13176 17280 13228 17332
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 9588 17212 9640 17264
rect 14556 17280 14608 17332
rect 17592 17280 17644 17332
rect 18880 17323 18932 17332
rect 18880 17289 18889 17323
rect 18889 17289 18923 17323
rect 18923 17289 18932 17323
rect 18880 17280 18932 17289
rect 20352 17280 20404 17332
rect 20628 17280 20680 17332
rect 20996 17323 21048 17332
rect 20996 17289 21005 17323
rect 21005 17289 21039 17323
rect 21039 17289 21048 17323
rect 20996 17280 21048 17289
rect 22928 17280 22980 17332
rect 23848 17280 23900 17332
rect 26240 17323 26292 17332
rect 26240 17289 26249 17323
rect 26249 17289 26283 17323
rect 26283 17289 26292 17323
rect 26240 17280 26292 17289
rect 9956 17187 10008 17196
rect 9956 17153 9990 17187
rect 9990 17153 10008 17187
rect 9956 17144 10008 17153
rect 11520 17187 11572 17196
rect 11520 17153 11529 17187
rect 11529 17153 11563 17187
rect 11563 17153 11572 17187
rect 11520 17144 11572 17153
rect 11796 17187 11848 17196
rect 11796 17153 11830 17187
rect 11830 17153 11848 17187
rect 11796 17144 11848 17153
rect 13452 17187 13504 17196
rect 13452 17153 13461 17187
rect 13461 17153 13495 17187
rect 13495 17153 13504 17187
rect 13452 17144 13504 17153
rect 8852 17076 8904 17128
rect 9312 17076 9364 17128
rect 5264 17008 5316 17060
rect 6552 16940 6604 16992
rect 6828 17008 6880 17060
rect 8392 16940 8444 16992
rect 11520 16940 11572 16992
rect 12532 16940 12584 16992
rect 14832 17144 14884 17196
rect 16580 17144 16632 17196
rect 16764 17144 16816 17196
rect 17224 17144 17276 17196
rect 21824 17144 21876 17196
rect 23664 17212 23716 17264
rect 24676 17212 24728 17264
rect 28264 17280 28316 17332
rect 29460 17323 29512 17332
rect 29460 17289 29469 17323
rect 29469 17289 29503 17323
rect 29503 17289 29512 17323
rect 29460 17280 29512 17289
rect 32404 17280 32456 17332
rect 33600 17323 33652 17332
rect 33600 17289 33609 17323
rect 33609 17289 33643 17323
rect 33643 17289 33652 17323
rect 33600 17280 33652 17289
rect 27712 17212 27764 17264
rect 26424 17187 26476 17196
rect 26424 17153 26433 17187
rect 26433 17153 26467 17187
rect 26467 17153 26476 17187
rect 26424 17144 26476 17153
rect 29644 17187 29696 17196
rect 29644 17153 29653 17187
rect 29653 17153 29687 17187
rect 29687 17153 29696 17187
rect 29644 17144 29696 17153
rect 32496 17187 32548 17196
rect 32496 17153 32505 17187
rect 32505 17153 32539 17187
rect 32539 17153 32548 17187
rect 32496 17144 32548 17153
rect 34428 17144 34480 17196
rect 36452 17187 36504 17196
rect 36452 17153 36461 17187
rect 36461 17153 36495 17187
rect 36495 17153 36504 17187
rect 36452 17144 36504 17153
rect 18236 17008 18288 17060
rect 25136 17076 25188 17128
rect 19800 17008 19852 17060
rect 16396 16983 16448 16992
rect 16396 16949 16405 16983
rect 16405 16949 16439 16983
rect 16439 16949 16448 16983
rect 16396 16940 16448 16949
rect 32680 17076 32732 17128
rect 30288 17008 30340 17060
rect 34060 17119 34112 17128
rect 34060 17085 34069 17119
rect 34069 17085 34103 17119
rect 34103 17085 34112 17119
rect 34060 17076 34112 17085
rect 34336 17076 34388 17128
rect 29184 16940 29236 16992
rect 36176 16940 36228 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 4712 16668 4764 16720
rect 5264 16600 5316 16652
rect 8852 16736 8904 16788
rect 11796 16779 11848 16788
rect 11796 16745 11805 16779
rect 11805 16745 11839 16779
rect 11839 16745 11848 16779
rect 11796 16736 11848 16745
rect 9128 16668 9180 16720
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 8392 16532 8444 16584
rect 16396 16736 16448 16788
rect 17224 16779 17276 16788
rect 17224 16745 17233 16779
rect 17233 16745 17267 16779
rect 17267 16745 17276 16779
rect 17224 16736 17276 16745
rect 14832 16600 14884 16652
rect 16396 16600 16448 16652
rect 22192 16600 22244 16652
rect 23664 16600 23716 16652
rect 23940 16643 23992 16652
rect 23940 16609 23949 16643
rect 23949 16609 23983 16643
rect 23983 16609 23992 16643
rect 27712 16779 27764 16788
rect 27712 16745 27721 16779
rect 27721 16745 27755 16779
rect 27755 16745 27764 16779
rect 27712 16736 27764 16745
rect 29644 16736 29696 16788
rect 23940 16600 23992 16609
rect 27804 16600 27856 16652
rect 28172 16643 28224 16652
rect 28172 16609 28181 16643
rect 28181 16609 28215 16643
rect 28215 16609 28224 16643
rect 28172 16600 28224 16609
rect 31944 16736 31996 16788
rect 32496 16736 32548 16788
rect 30104 16668 30156 16720
rect 30288 16643 30340 16652
rect 30288 16609 30297 16643
rect 30297 16609 30331 16643
rect 30331 16609 30340 16643
rect 30288 16600 30340 16609
rect 31116 16643 31168 16652
rect 31116 16609 31125 16643
rect 31125 16609 31159 16643
rect 31159 16609 31168 16643
rect 31116 16600 31168 16609
rect 31576 16643 31628 16652
rect 31576 16609 31585 16643
rect 31585 16609 31619 16643
rect 31619 16609 31628 16643
rect 34152 16736 34204 16788
rect 34428 16736 34480 16788
rect 31576 16600 31628 16609
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 5448 16464 5500 16516
rect 6368 16464 6420 16516
rect 8024 16464 8076 16516
rect 3056 16396 3108 16448
rect 4160 16439 4212 16448
rect 4160 16405 4169 16439
rect 4169 16405 4203 16439
rect 4203 16405 4212 16439
rect 4160 16396 4212 16405
rect 4620 16439 4672 16448
rect 4620 16405 4629 16439
rect 4629 16405 4663 16439
rect 4663 16405 4672 16439
rect 4620 16396 4672 16405
rect 6828 16396 6880 16448
rect 9036 16439 9088 16448
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 13176 16532 13228 16584
rect 17040 16532 17092 16584
rect 20812 16532 20864 16584
rect 24860 16575 24912 16584
rect 24860 16541 24869 16575
rect 24869 16541 24903 16575
rect 24903 16541 24912 16575
rect 24860 16532 24912 16541
rect 28264 16532 28316 16584
rect 29552 16532 29604 16584
rect 33784 16532 33836 16584
rect 15292 16464 15344 16516
rect 13360 16396 13412 16448
rect 17316 16464 17368 16516
rect 23664 16507 23716 16516
rect 23664 16473 23673 16507
rect 23673 16473 23707 16507
rect 23707 16473 23716 16507
rect 23664 16464 23716 16473
rect 26332 16464 26384 16516
rect 30196 16507 30248 16516
rect 30196 16473 30205 16507
rect 30205 16473 30239 16507
rect 30239 16473 30248 16507
rect 30196 16464 30248 16473
rect 31852 16507 31904 16516
rect 31852 16473 31886 16507
rect 31886 16473 31904 16507
rect 31852 16464 31904 16473
rect 16396 16439 16448 16448
rect 16396 16405 16405 16439
rect 16405 16405 16439 16439
rect 16439 16405 16448 16439
rect 16396 16396 16448 16405
rect 16948 16396 17000 16448
rect 22836 16396 22888 16448
rect 26056 16396 26108 16448
rect 30104 16439 30156 16448
rect 30104 16405 30113 16439
rect 30113 16405 30147 16439
rect 30147 16405 30156 16439
rect 30104 16396 30156 16405
rect 30564 16439 30616 16448
rect 30564 16405 30573 16439
rect 30573 16405 30607 16439
rect 30607 16405 30616 16439
rect 30564 16396 30616 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 4160 16192 4212 16244
rect 6368 16235 6420 16244
rect 6368 16201 6377 16235
rect 6377 16201 6411 16235
rect 6411 16201 6420 16235
rect 6368 16192 6420 16201
rect 7840 16192 7892 16244
rect 9220 16192 9272 16244
rect 10324 16192 10376 16244
rect 1860 16056 1912 16108
rect 2780 16124 2832 16176
rect 4620 16167 4672 16176
rect 2688 16099 2740 16108
rect 2688 16065 2722 16099
rect 2722 16065 2740 16099
rect 2688 16056 2740 16065
rect 4620 16133 4654 16167
rect 4654 16133 4672 16167
rect 4620 16124 4672 16133
rect 9036 16124 9088 16176
rect 13820 16192 13872 16244
rect 15292 16235 15344 16244
rect 15292 16201 15301 16235
rect 15301 16201 15335 16235
rect 15335 16201 15344 16235
rect 15292 16192 15344 16201
rect 19616 16192 19668 16244
rect 20260 16192 20312 16244
rect 21548 16235 21600 16244
rect 21548 16201 21557 16235
rect 21557 16201 21591 16235
rect 21591 16201 21600 16235
rect 21548 16192 21600 16201
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 8392 16056 8444 16108
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 9128 16099 9180 16108
rect 9128 16065 9162 16099
rect 9162 16065 9180 16099
rect 9128 16056 9180 16065
rect 10232 16056 10284 16108
rect 12440 16099 12492 16108
rect 12440 16065 12449 16099
rect 12449 16065 12483 16099
rect 12483 16065 12492 16099
rect 12440 16056 12492 16065
rect 12532 16099 12584 16108
rect 12532 16065 12541 16099
rect 12541 16065 12575 16099
rect 12575 16065 12584 16099
rect 12532 16056 12584 16065
rect 16396 16056 16448 16108
rect 17592 16099 17644 16108
rect 17592 16065 17601 16099
rect 17601 16065 17635 16099
rect 17635 16065 17644 16099
rect 17592 16056 17644 16065
rect 19248 16124 19300 16176
rect 23756 16192 23808 16244
rect 24860 16192 24912 16244
rect 25872 16192 25924 16244
rect 26332 16235 26384 16244
rect 26332 16201 26341 16235
rect 26341 16201 26375 16235
rect 26375 16201 26384 16235
rect 26332 16192 26384 16201
rect 18696 16099 18748 16108
rect 18696 16065 18730 16099
rect 18730 16065 18748 16099
rect 18696 16056 18748 16065
rect 26148 16124 26200 16176
rect 30104 16192 30156 16244
rect 31852 16192 31904 16244
rect 20076 16056 20128 16108
rect 22836 16099 22888 16108
rect 22836 16065 22845 16099
rect 22845 16065 22879 16099
rect 22879 16065 22888 16099
rect 22836 16056 22888 16065
rect 25872 16056 25924 16108
rect 26976 16056 27028 16108
rect 29736 16056 29788 16108
rect 32496 16235 32548 16244
rect 32496 16201 32505 16235
rect 32505 16201 32539 16235
rect 32539 16201 32548 16235
rect 32496 16192 32548 16201
rect 32588 16192 32640 16244
rect 33784 16235 33836 16244
rect 33784 16201 33793 16235
rect 33793 16201 33827 16235
rect 33827 16201 33836 16235
rect 33784 16192 33836 16201
rect 34428 16192 34480 16244
rect 33508 16124 33560 16176
rect 34060 16124 34112 16176
rect 8024 15963 8076 15972
rect 8024 15929 8033 15963
rect 8033 15929 8067 15963
rect 8067 15929 8076 15963
rect 8024 15920 8076 15929
rect 940 15852 992 15904
rect 5724 15895 5776 15904
rect 5724 15861 5733 15895
rect 5733 15861 5767 15895
rect 5767 15861 5776 15895
rect 5724 15852 5776 15861
rect 7012 15852 7064 15904
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 10508 15852 10560 15904
rect 12716 15852 12768 15904
rect 15476 15852 15528 15904
rect 16764 15852 16816 15904
rect 22652 15988 22704 16040
rect 29184 16031 29236 16040
rect 29184 15997 29193 16031
rect 29193 15997 29227 16031
rect 29227 15997 29236 16031
rect 29184 15988 29236 15997
rect 32588 16031 32640 16040
rect 32588 15997 32597 16031
rect 32597 15997 32631 16031
rect 32631 15997 32640 16031
rect 32588 15988 32640 15997
rect 32680 16031 32732 16040
rect 32680 15997 32689 16031
rect 32689 15997 32723 16031
rect 32723 15997 32732 16031
rect 32680 15988 32732 15997
rect 33692 15988 33744 16040
rect 34336 16031 34388 16040
rect 34336 15997 34345 16031
rect 34345 15997 34379 16031
rect 34379 15997 34388 16031
rect 34336 15988 34388 15997
rect 20812 15852 20864 15904
rect 25412 15852 25464 15904
rect 28448 15852 28500 15904
rect 31116 15852 31168 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2688 15648 2740 15700
rect 4804 15691 4856 15700
rect 4804 15657 4813 15691
rect 4813 15657 4847 15691
rect 4847 15657 4856 15691
rect 4804 15648 4856 15657
rect 9128 15648 9180 15700
rect 12440 15648 12492 15700
rect 18696 15691 18748 15700
rect 18696 15657 18705 15691
rect 18705 15657 18739 15691
rect 18739 15657 18748 15691
rect 18696 15648 18748 15657
rect 20076 15691 20128 15700
rect 20076 15657 20085 15691
rect 20085 15657 20119 15691
rect 20119 15657 20128 15691
rect 20076 15648 20128 15657
rect 16856 15580 16908 15632
rect 5264 15512 5316 15564
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 5724 15444 5776 15496
rect 10324 15512 10376 15564
rect 7748 15376 7800 15428
rect 10232 15444 10284 15496
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 10784 15487 10836 15496
rect 10784 15453 10793 15487
rect 10793 15453 10827 15487
rect 10827 15453 10836 15487
rect 10784 15444 10836 15453
rect 16764 15555 16816 15564
rect 16764 15521 16773 15555
rect 16773 15521 16807 15555
rect 16807 15521 16816 15555
rect 16764 15512 16816 15521
rect 17592 15512 17644 15564
rect 13820 15444 13872 15496
rect 13360 15419 13412 15428
rect 13360 15385 13369 15419
rect 13369 15385 13403 15419
rect 13403 15385 13412 15419
rect 13360 15376 13412 15385
rect 18972 15376 19024 15428
rect 6000 15308 6052 15360
rect 6644 15308 6696 15360
rect 9220 15351 9272 15360
rect 9220 15317 9229 15351
rect 9229 15317 9263 15351
rect 9263 15317 9272 15351
rect 9220 15308 9272 15317
rect 12164 15308 12216 15360
rect 16488 15351 16540 15360
rect 16488 15317 16497 15351
rect 16497 15317 16531 15351
rect 16531 15317 16540 15351
rect 16488 15308 16540 15317
rect 16948 15308 17000 15360
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 20260 15487 20312 15496
rect 20260 15453 20269 15487
rect 20269 15453 20303 15487
rect 20303 15453 20312 15487
rect 20260 15444 20312 15453
rect 20720 15580 20772 15632
rect 22560 15648 22612 15700
rect 23388 15648 23440 15700
rect 26976 15691 27028 15700
rect 26976 15657 26985 15691
rect 26985 15657 27019 15691
rect 27019 15657 27028 15691
rect 26976 15648 27028 15657
rect 20812 15444 20864 15496
rect 22100 15444 22152 15496
rect 27252 15512 27304 15564
rect 29552 15648 29604 15700
rect 29736 15691 29788 15700
rect 29736 15657 29745 15691
rect 29745 15657 29779 15691
rect 29779 15657 29788 15691
rect 29736 15648 29788 15657
rect 33416 15580 33468 15632
rect 28448 15555 28500 15564
rect 28448 15521 28457 15555
rect 28457 15521 28491 15555
rect 28491 15521 28500 15555
rect 28448 15512 28500 15521
rect 30196 15555 30248 15564
rect 30196 15521 30205 15555
rect 30205 15521 30239 15555
rect 30239 15521 30248 15555
rect 30196 15512 30248 15521
rect 23940 15444 23992 15496
rect 24492 15444 24544 15496
rect 26148 15444 26200 15496
rect 27436 15444 27488 15496
rect 19800 15376 19852 15428
rect 22376 15376 22428 15428
rect 25136 15376 25188 15428
rect 28632 15487 28684 15496
rect 28632 15453 28641 15487
rect 28641 15453 28675 15487
rect 28675 15453 28684 15487
rect 28632 15444 28684 15453
rect 30104 15487 30156 15496
rect 30104 15453 30113 15487
rect 30113 15453 30147 15487
rect 30147 15453 30156 15487
rect 30104 15444 30156 15453
rect 32680 15512 32732 15564
rect 24400 15308 24452 15360
rect 25872 15308 25924 15360
rect 27528 15308 27580 15360
rect 28264 15351 28316 15360
rect 28264 15317 28273 15351
rect 28273 15317 28307 15351
rect 28307 15317 28316 15351
rect 28264 15308 28316 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 4620 15036 4672 15088
rect 5356 15036 5408 15088
rect 4804 14968 4856 15020
rect 6920 15104 6972 15156
rect 16488 15147 16540 15156
rect 16488 15113 16497 15147
rect 16497 15113 16531 15147
rect 16531 15113 16540 15147
rect 16488 15104 16540 15113
rect 10508 15036 10560 15088
rect 8116 15011 8168 15020
rect 8116 14977 8125 15011
rect 8125 14977 8159 15011
rect 8159 14977 8168 15011
rect 8116 14968 8168 14977
rect 15200 15036 15252 15088
rect 18420 15104 18472 15156
rect 24124 15104 24176 15156
rect 25136 15147 25188 15156
rect 25136 15113 25145 15147
rect 25145 15113 25179 15147
rect 25179 15113 25188 15147
rect 25136 15104 25188 15113
rect 17224 15036 17276 15088
rect 23020 15036 23072 15088
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 16304 14968 16356 15020
rect 16580 14968 16632 15020
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 17500 14968 17552 15020
rect 22284 14968 22336 15020
rect 27252 15104 27304 15156
rect 34060 15104 34112 15156
rect 25688 15036 25740 15088
rect 25412 14968 25464 15020
rect 6644 14900 6696 14952
rect 7748 14900 7800 14952
rect 17316 14943 17368 14952
rect 17316 14909 17325 14943
rect 17325 14909 17359 14943
rect 17359 14909 17368 14943
rect 17316 14900 17368 14909
rect 24860 14900 24912 14952
rect 27436 15011 27488 15020
rect 27436 14977 27445 15011
rect 27445 14977 27479 15011
rect 27479 14977 27488 15011
rect 27436 14968 27488 14977
rect 27528 14943 27580 14952
rect 27528 14909 27537 14943
rect 27537 14909 27571 14943
rect 27571 14909 27580 14943
rect 27528 14900 27580 14909
rect 28632 15036 28684 15088
rect 30748 14968 30800 15020
rect 34244 15011 34296 15020
rect 34244 14977 34253 15011
rect 34253 14977 34287 15011
rect 34287 14977 34296 15011
rect 34244 14968 34296 14977
rect 36176 14968 36228 15020
rect 33416 14900 33468 14952
rect 3976 14764 4028 14816
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 9864 14764 9916 14816
rect 14832 14807 14884 14816
rect 14832 14773 14841 14807
rect 14841 14773 14875 14807
rect 14875 14773 14884 14807
rect 14832 14764 14884 14773
rect 17960 14764 18012 14816
rect 27988 14832 28040 14884
rect 30288 14832 30340 14884
rect 22376 14807 22428 14816
rect 22376 14773 22385 14807
rect 22385 14773 22419 14807
rect 22419 14773 22428 14807
rect 22376 14764 22428 14773
rect 27160 14764 27212 14816
rect 31852 14764 31904 14816
rect 33232 14807 33284 14816
rect 33232 14773 33241 14807
rect 33241 14773 33275 14807
rect 33275 14773 33284 14807
rect 33232 14764 33284 14773
rect 33324 14764 33376 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 6920 14560 6972 14612
rect 9864 14603 9916 14612
rect 9864 14569 9873 14603
rect 9873 14569 9907 14603
rect 9907 14569 9916 14603
rect 9864 14560 9916 14569
rect 17224 14560 17276 14612
rect 20260 14560 20312 14612
rect 22284 14603 22336 14612
rect 22284 14569 22293 14603
rect 22293 14569 22327 14603
rect 22327 14569 22336 14603
rect 22284 14560 22336 14569
rect 27436 14560 27488 14612
rect 27988 14560 28040 14612
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 4712 14356 4764 14408
rect 5356 14399 5408 14408
rect 5356 14365 5390 14399
rect 5390 14365 5408 14399
rect 5356 14356 5408 14365
rect 6828 14356 6880 14408
rect 11704 14535 11756 14544
rect 11704 14501 11713 14535
rect 11713 14501 11747 14535
rect 11747 14501 11756 14535
rect 11704 14492 11756 14501
rect 17316 14492 17368 14544
rect 18144 14492 18196 14544
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 10968 14424 11020 14476
rect 13912 14424 13964 14476
rect 19524 14424 19576 14476
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 10784 14356 10836 14408
rect 7932 14288 7984 14340
rect 11520 14288 11572 14340
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 13728 14356 13780 14408
rect 12532 14288 12584 14340
rect 14096 14399 14148 14408
rect 14096 14365 14105 14399
rect 14105 14365 14139 14399
rect 14139 14365 14148 14399
rect 14096 14356 14148 14365
rect 14832 14356 14884 14408
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 18420 14356 18472 14408
rect 18512 14399 18564 14408
rect 18512 14365 18521 14399
rect 18521 14365 18555 14399
rect 18555 14365 18564 14399
rect 18512 14356 18564 14365
rect 17776 14288 17828 14340
rect 19984 14492 20036 14544
rect 25412 14492 25464 14544
rect 30196 14492 30248 14544
rect 30748 14535 30800 14544
rect 30748 14501 30757 14535
rect 30757 14501 30791 14535
rect 30791 14501 30800 14535
rect 30748 14492 30800 14501
rect 34060 14492 34112 14544
rect 20996 14467 21048 14476
rect 20996 14433 21005 14467
rect 21005 14433 21039 14467
rect 21039 14433 21048 14467
rect 20996 14424 21048 14433
rect 21364 14424 21416 14476
rect 23020 14424 23072 14476
rect 26148 14424 26200 14476
rect 28172 14424 28224 14476
rect 30288 14424 30340 14476
rect 32864 14424 32916 14476
rect 33324 14467 33376 14476
rect 33324 14433 33333 14467
rect 33333 14433 33367 14467
rect 33367 14433 33376 14467
rect 33324 14424 33376 14433
rect 25412 14399 25464 14408
rect 25412 14365 25421 14399
rect 25421 14365 25455 14399
rect 25455 14365 25464 14399
rect 25412 14356 25464 14365
rect 26424 14356 26476 14408
rect 29368 14399 29420 14408
rect 29368 14365 29377 14399
rect 29377 14365 29411 14399
rect 29411 14365 29420 14399
rect 29368 14356 29420 14365
rect 21364 14288 21416 14340
rect 22744 14331 22796 14340
rect 22744 14297 22753 14331
rect 22753 14297 22787 14331
rect 22787 14297 22796 14331
rect 22744 14288 22796 14297
rect 24492 14331 24544 14340
rect 24492 14297 24501 14331
rect 24501 14297 24535 14331
rect 24535 14297 24544 14331
rect 24492 14288 24544 14297
rect 26976 14288 27028 14340
rect 3792 14263 3844 14272
rect 3792 14229 3801 14263
rect 3801 14229 3835 14263
rect 3835 14229 3844 14263
rect 3792 14220 3844 14229
rect 8208 14220 8260 14272
rect 11796 14220 11848 14272
rect 11888 14263 11940 14272
rect 11888 14229 11897 14263
rect 11897 14229 11931 14263
rect 11931 14229 11940 14263
rect 11888 14220 11940 14229
rect 12348 14263 12400 14272
rect 12348 14229 12357 14263
rect 12357 14229 12391 14263
rect 12391 14229 12400 14263
rect 12348 14220 12400 14229
rect 13268 14220 13320 14272
rect 13728 14263 13780 14272
rect 13728 14229 13737 14263
rect 13737 14229 13771 14263
rect 13771 14229 13780 14263
rect 13728 14220 13780 14229
rect 14556 14220 14608 14272
rect 16488 14263 16540 14272
rect 16488 14229 16497 14263
rect 16497 14229 16531 14263
rect 16531 14229 16540 14263
rect 16488 14220 16540 14229
rect 18604 14220 18656 14272
rect 19616 14263 19668 14272
rect 19616 14229 19625 14263
rect 19625 14229 19659 14263
rect 19659 14229 19668 14263
rect 19616 14220 19668 14229
rect 20444 14263 20496 14272
rect 20444 14229 20453 14263
rect 20453 14229 20487 14263
rect 20487 14229 20496 14263
rect 20444 14220 20496 14229
rect 20812 14263 20864 14272
rect 20812 14229 20821 14263
rect 20821 14229 20855 14263
rect 20855 14229 20864 14263
rect 20812 14220 20864 14229
rect 21180 14220 21232 14272
rect 22652 14263 22704 14272
rect 22652 14229 22661 14263
rect 22661 14229 22695 14263
rect 22695 14229 22704 14263
rect 22652 14220 22704 14229
rect 24124 14220 24176 14272
rect 26424 14263 26476 14272
rect 26424 14229 26433 14263
rect 26433 14229 26467 14263
rect 26467 14229 26476 14263
rect 26424 14220 26476 14229
rect 31852 14399 31904 14408
rect 31852 14365 31861 14399
rect 31861 14365 31895 14399
rect 31895 14365 31904 14399
rect 31852 14356 31904 14365
rect 33232 14399 33284 14408
rect 33232 14365 33241 14399
rect 33241 14365 33275 14399
rect 33275 14365 33284 14399
rect 33232 14356 33284 14365
rect 29276 14220 29328 14272
rect 30012 14220 30064 14272
rect 31208 14263 31260 14272
rect 31208 14229 31217 14263
rect 31217 14229 31251 14263
rect 31251 14229 31260 14263
rect 31208 14220 31260 14229
rect 32864 14288 32916 14340
rect 32588 14263 32640 14272
rect 32588 14229 32597 14263
rect 32597 14229 32631 14263
rect 32631 14229 32640 14263
rect 32588 14220 32640 14229
rect 36360 14263 36412 14272
rect 36360 14229 36369 14263
rect 36369 14229 36403 14263
rect 36403 14229 36412 14263
rect 36360 14220 36412 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 4620 14016 4672 14068
rect 3792 13948 3844 14000
rect 6736 13948 6788 14000
rect 4712 13880 4764 13932
rect 6828 13880 6880 13932
rect 10692 14016 10744 14068
rect 10968 14016 11020 14068
rect 9772 13948 9824 14000
rect 9864 13880 9916 13932
rect 10232 13880 10284 13932
rect 12072 14016 12124 14068
rect 12532 13991 12584 14000
rect 12532 13957 12541 13991
rect 12541 13957 12575 13991
rect 12575 13957 12584 13991
rect 12532 13948 12584 13957
rect 11612 13880 11664 13932
rect 12348 13923 12400 13932
rect 12348 13889 12357 13923
rect 12357 13889 12391 13923
rect 12391 13889 12400 13923
rect 12348 13880 12400 13889
rect 13176 13991 13228 14000
rect 13176 13957 13185 13991
rect 13185 13957 13219 13991
rect 13219 13957 13228 13991
rect 13176 13948 13228 13957
rect 11520 13855 11572 13864
rect 11520 13821 11529 13855
rect 11529 13821 11563 13855
rect 11563 13821 11572 13855
rect 11520 13812 11572 13821
rect 11704 13855 11756 13864
rect 11704 13821 11713 13855
rect 11713 13821 11747 13855
rect 11747 13821 11756 13855
rect 11704 13812 11756 13821
rect 11796 13812 11848 13864
rect 13268 13923 13320 13932
rect 13268 13889 13277 13923
rect 13277 13889 13311 13923
rect 13311 13889 13320 13923
rect 13268 13880 13320 13889
rect 14096 14016 14148 14068
rect 15476 14016 15528 14068
rect 13728 13923 13780 13932
rect 13728 13889 13752 13923
rect 13752 13889 13780 13923
rect 13728 13880 13780 13889
rect 2320 13676 2372 13728
rect 10600 13744 10652 13796
rect 8392 13676 8444 13728
rect 9772 13676 9824 13728
rect 10784 13744 10836 13796
rect 13912 13923 13964 13932
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 14188 13948 14240 14000
rect 19616 14016 19668 14068
rect 19984 14016 20036 14068
rect 20812 14016 20864 14068
rect 22652 14016 22704 14068
rect 14096 13880 14148 13932
rect 14556 13923 14608 13932
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 16304 13880 16356 13932
rect 18604 13880 18656 13932
rect 21272 13948 21324 14000
rect 21548 13948 21600 14000
rect 22284 13991 22336 14000
rect 22284 13957 22318 13991
rect 22318 13957 22336 13991
rect 22284 13948 22336 13957
rect 25412 14016 25464 14068
rect 26976 14059 27028 14068
rect 26976 14025 26985 14059
rect 26985 14025 27019 14059
rect 27019 14025 27028 14059
rect 26976 14016 27028 14025
rect 29368 14016 29420 14068
rect 30196 14016 30248 14068
rect 28172 13948 28224 14000
rect 33140 14059 33192 14068
rect 33140 14025 33149 14059
rect 33149 14025 33183 14059
rect 33183 14025 33192 14059
rect 33140 14016 33192 14025
rect 34060 14016 34112 14068
rect 20260 13923 20312 13932
rect 20260 13889 20294 13923
rect 20294 13889 20312 13923
rect 20260 13880 20312 13889
rect 15200 13812 15252 13864
rect 21824 13812 21876 13864
rect 22008 13855 22060 13864
rect 22008 13821 22017 13855
rect 22017 13821 22051 13855
rect 22051 13821 22060 13855
rect 24032 13923 24084 13932
rect 24032 13889 24041 13923
rect 24041 13889 24075 13923
rect 24075 13889 24084 13923
rect 24032 13880 24084 13889
rect 24124 13923 24176 13932
rect 24124 13889 24133 13923
rect 24133 13889 24167 13923
rect 24167 13889 24176 13923
rect 24124 13880 24176 13889
rect 24216 13880 24268 13932
rect 25872 13923 25924 13932
rect 25872 13889 25881 13923
rect 25881 13889 25915 13923
rect 25915 13889 25924 13923
rect 25872 13880 25924 13889
rect 27160 13923 27212 13932
rect 27160 13889 27169 13923
rect 27169 13889 27203 13923
rect 27203 13889 27212 13923
rect 27160 13880 27212 13889
rect 28448 13923 28500 13932
rect 28448 13889 28457 13923
rect 28457 13889 28491 13923
rect 28491 13889 28500 13923
rect 28448 13880 28500 13889
rect 29276 13923 29328 13932
rect 29276 13889 29285 13923
rect 29285 13889 29319 13923
rect 29319 13889 29328 13923
rect 29276 13880 29328 13889
rect 22008 13812 22060 13821
rect 10876 13676 10928 13728
rect 12072 13744 12124 13796
rect 12348 13744 12400 13796
rect 17960 13744 18012 13796
rect 25504 13787 25556 13796
rect 25504 13753 25513 13787
rect 25513 13753 25547 13787
rect 25547 13753 25556 13787
rect 25504 13744 25556 13753
rect 13912 13676 13964 13728
rect 14004 13676 14056 13728
rect 22284 13676 22336 13728
rect 23848 13676 23900 13728
rect 27988 13676 28040 13728
rect 28172 13855 28224 13864
rect 28172 13821 28181 13855
rect 28181 13821 28215 13855
rect 28215 13821 28224 13855
rect 28172 13812 28224 13821
rect 28540 13676 28592 13728
rect 29920 13744 29972 13796
rect 30288 13812 30340 13864
rect 30748 13923 30800 13932
rect 30748 13889 30757 13923
rect 30757 13889 30791 13923
rect 30791 13889 30800 13923
rect 30748 13880 30800 13889
rect 31944 13923 31996 13932
rect 31944 13889 31953 13923
rect 31953 13889 31987 13923
rect 31987 13889 31996 13923
rect 31944 13880 31996 13889
rect 33508 13880 33560 13932
rect 30656 13676 30708 13728
rect 33600 13855 33652 13864
rect 33600 13821 33609 13855
rect 33609 13821 33643 13855
rect 33643 13821 33652 13855
rect 33600 13812 33652 13821
rect 33692 13855 33744 13864
rect 33692 13821 33701 13855
rect 33701 13821 33735 13855
rect 33735 13821 33744 13855
rect 33692 13812 33744 13821
rect 32956 13676 33008 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4620 13268 4672 13320
rect 7196 13404 7248 13456
rect 9404 13472 9456 13524
rect 10048 13404 10100 13456
rect 10968 13404 11020 13456
rect 16672 13472 16724 13524
rect 17684 13472 17736 13524
rect 18512 13472 18564 13524
rect 20260 13515 20312 13524
rect 20260 13481 20269 13515
rect 20269 13481 20303 13515
rect 20303 13481 20312 13515
rect 20260 13472 20312 13481
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 21824 13472 21876 13524
rect 24032 13472 24084 13524
rect 28448 13472 28500 13524
rect 30748 13472 30800 13524
rect 6644 13336 6696 13388
rect 6276 13311 6328 13320
rect 6276 13277 6285 13311
rect 6285 13277 6319 13311
rect 6319 13277 6328 13311
rect 6276 13268 6328 13277
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 10692 13336 10744 13388
rect 11796 13336 11848 13388
rect 13084 13336 13136 13388
rect 15292 13336 15344 13388
rect 6828 13200 6880 13252
rect 8852 13200 8904 13252
rect 11060 13268 11112 13320
rect 11888 13268 11940 13320
rect 16304 13336 16356 13388
rect 23848 13404 23900 13456
rect 19064 13336 19116 13388
rect 19524 13336 19576 13388
rect 14924 13200 14976 13252
rect 17592 13268 17644 13320
rect 16764 13243 16816 13252
rect 16764 13209 16798 13243
rect 16798 13209 16816 13243
rect 16764 13200 16816 13209
rect 18052 13200 18104 13252
rect 19616 13311 19668 13320
rect 19616 13277 19625 13311
rect 19625 13277 19659 13311
rect 19659 13277 19668 13311
rect 19616 13268 19668 13277
rect 21180 13379 21232 13388
rect 21180 13345 21189 13379
rect 21189 13345 21223 13379
rect 21223 13345 21232 13379
rect 21180 13336 21232 13345
rect 21364 13379 21416 13388
rect 21364 13345 21373 13379
rect 21373 13345 21407 13379
rect 21407 13345 21416 13379
rect 21364 13336 21416 13345
rect 22928 13379 22980 13388
rect 20444 13311 20496 13320
rect 20444 13277 20453 13311
rect 20453 13277 20487 13311
rect 20487 13277 20496 13311
rect 20444 13268 20496 13277
rect 20812 13268 20864 13320
rect 20996 13200 21048 13252
rect 22928 13345 22937 13379
rect 22937 13345 22971 13379
rect 22971 13345 22980 13379
rect 22928 13336 22980 13345
rect 22652 13311 22704 13320
rect 22652 13277 22661 13311
rect 22661 13277 22695 13311
rect 22695 13277 22704 13311
rect 22652 13268 22704 13277
rect 22744 13311 22796 13320
rect 22744 13277 22753 13311
rect 22753 13277 22787 13311
rect 22787 13277 22796 13311
rect 22744 13268 22796 13277
rect 24032 13336 24084 13388
rect 25504 13336 25556 13388
rect 26332 13379 26384 13388
rect 26332 13345 26341 13379
rect 26341 13345 26375 13379
rect 26375 13345 26384 13379
rect 26332 13336 26384 13345
rect 29092 13404 29144 13456
rect 27160 13311 27212 13320
rect 27160 13277 27169 13311
rect 27169 13277 27203 13311
rect 27203 13277 27212 13311
rect 27160 13268 27212 13277
rect 32036 13336 32088 13388
rect 32956 13336 33008 13388
rect 29000 13268 29052 13320
rect 29092 13311 29144 13320
rect 29092 13277 29101 13311
rect 29101 13277 29135 13311
rect 29135 13277 29144 13311
rect 29092 13268 29144 13277
rect 32864 13268 32916 13320
rect 5448 13175 5500 13184
rect 5448 13141 5457 13175
rect 5457 13141 5491 13175
rect 5491 13141 5500 13175
rect 5448 13132 5500 13141
rect 7380 13132 7432 13184
rect 8300 13175 8352 13184
rect 8300 13141 8309 13175
rect 8309 13141 8343 13175
rect 8343 13141 8352 13175
rect 8300 13132 8352 13141
rect 10416 13132 10468 13184
rect 10600 13132 10652 13184
rect 15016 13132 15068 13184
rect 15292 13132 15344 13184
rect 16396 13132 16448 13184
rect 19064 13132 19116 13184
rect 24308 13200 24360 13252
rect 31944 13200 31996 13252
rect 22100 13132 22152 13184
rect 22744 13132 22796 13184
rect 23388 13132 23440 13184
rect 24768 13175 24820 13184
rect 24768 13141 24777 13175
rect 24777 13141 24811 13175
rect 24811 13141 24820 13175
rect 24768 13132 24820 13141
rect 25596 13132 25648 13184
rect 26148 13175 26200 13184
rect 26148 13141 26157 13175
rect 26157 13141 26191 13175
rect 26191 13141 26200 13175
rect 26148 13132 26200 13141
rect 26240 13175 26292 13184
rect 26240 13141 26249 13175
rect 26249 13141 26283 13175
rect 26283 13141 26292 13175
rect 26240 13132 26292 13141
rect 27252 13132 27304 13184
rect 27988 13132 28040 13184
rect 28448 13175 28500 13184
rect 28448 13141 28457 13175
rect 28457 13141 28491 13175
rect 28491 13141 28500 13175
rect 28448 13132 28500 13141
rect 28540 13175 28592 13184
rect 28540 13141 28549 13175
rect 28549 13141 28583 13175
rect 28583 13141 28592 13175
rect 28540 13132 28592 13141
rect 29000 13132 29052 13184
rect 30104 13132 30156 13184
rect 31116 13132 31168 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 7748 12928 7800 12980
rect 5356 12860 5408 12912
rect 8852 12971 8904 12980
rect 8852 12937 8861 12971
rect 8861 12937 8895 12971
rect 8895 12937 8904 12971
rect 8852 12928 8904 12937
rect 9772 12903 9824 12912
rect 5448 12792 5500 12844
rect 6828 12792 6880 12844
rect 7104 12792 7156 12844
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 5908 12724 5960 12776
rect 6368 12767 6420 12776
rect 6368 12733 6377 12767
rect 6377 12733 6411 12767
rect 6411 12733 6420 12767
rect 6368 12724 6420 12733
rect 7656 12767 7708 12776
rect 7656 12733 7665 12767
rect 7665 12733 7699 12767
rect 7699 12733 7708 12767
rect 7656 12724 7708 12733
rect 8576 12835 8628 12844
rect 8576 12801 8585 12835
rect 8585 12801 8619 12835
rect 8619 12801 8628 12835
rect 8576 12792 8628 12801
rect 9772 12869 9781 12903
rect 9781 12869 9815 12903
rect 9815 12869 9824 12903
rect 9772 12860 9824 12869
rect 8024 12724 8076 12776
rect 8944 12767 8996 12776
rect 8944 12733 8953 12767
rect 8953 12733 8987 12767
rect 8987 12733 8996 12767
rect 8944 12724 8996 12733
rect 9128 12792 9180 12844
rect 9404 12835 9456 12844
rect 9404 12801 9413 12835
rect 9413 12801 9447 12835
rect 9447 12801 9456 12835
rect 9404 12792 9456 12801
rect 10876 12792 10928 12844
rect 15384 12860 15436 12912
rect 16764 12928 16816 12980
rect 21180 12928 21232 12980
rect 24584 12928 24636 12980
rect 24768 12928 24820 12980
rect 11060 12792 11112 12844
rect 12164 12656 12216 12708
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 13912 12792 13964 12844
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 15016 12792 15068 12844
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 14004 12767 14056 12776
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 14096 12767 14148 12776
rect 14096 12733 14105 12767
rect 14105 12733 14139 12767
rect 14139 12733 14148 12767
rect 14096 12724 14148 12733
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 15752 12835 15804 12844
rect 15752 12801 15761 12835
rect 15761 12801 15795 12835
rect 15795 12801 15804 12835
rect 15752 12792 15804 12801
rect 16120 12792 16172 12844
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 18328 12792 18380 12844
rect 24308 12792 24360 12844
rect 25596 12835 25648 12844
rect 25596 12801 25605 12835
rect 25605 12801 25639 12835
rect 25639 12801 25648 12835
rect 25596 12792 25648 12801
rect 26148 12792 26200 12844
rect 28264 12928 28316 12980
rect 28448 12928 28500 12980
rect 29276 12928 29328 12980
rect 29644 12928 29696 12980
rect 17132 12724 17184 12776
rect 15752 12656 15804 12708
rect 18420 12724 18472 12776
rect 25412 12724 25464 12776
rect 28172 12860 28224 12912
rect 33324 12928 33376 12980
rect 33600 12928 33652 12980
rect 35992 12971 36044 12980
rect 35992 12937 36001 12971
rect 36001 12937 36035 12971
rect 36035 12937 36044 12971
rect 35992 12928 36044 12937
rect 27252 12835 27304 12844
rect 27252 12801 27261 12835
rect 27261 12801 27295 12835
rect 27295 12801 27304 12835
rect 27252 12792 27304 12801
rect 29184 12835 29236 12844
rect 29184 12801 29218 12835
rect 29218 12801 29236 12835
rect 29184 12792 29236 12801
rect 32956 12835 33008 12844
rect 32956 12801 32965 12835
rect 32965 12801 32999 12835
rect 32999 12801 33008 12835
rect 32956 12792 33008 12801
rect 33048 12835 33100 12844
rect 33048 12801 33057 12835
rect 33057 12801 33091 12835
rect 33091 12801 33100 12835
rect 33048 12792 33100 12801
rect 34704 12792 34756 12844
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 8300 12588 8352 12640
rect 14004 12588 14056 12640
rect 15660 12588 15712 12640
rect 18604 12699 18656 12708
rect 18604 12665 18613 12699
rect 18613 12665 18647 12699
rect 18647 12665 18656 12699
rect 18604 12656 18656 12665
rect 18880 12588 18932 12640
rect 22744 12588 22796 12640
rect 24216 12588 24268 12640
rect 27620 12588 27672 12640
rect 27988 12631 28040 12640
rect 27988 12597 27997 12631
rect 27997 12597 28031 12631
rect 28031 12597 28040 12631
rect 27988 12588 28040 12597
rect 34612 12588 34664 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 8944 12384 8996 12436
rect 7748 12291 7800 12300
rect 7748 12257 7757 12291
rect 7757 12257 7791 12291
rect 7791 12257 7800 12291
rect 7748 12248 7800 12257
rect 11428 12384 11480 12436
rect 11612 12427 11664 12436
rect 11612 12393 11621 12427
rect 11621 12393 11655 12427
rect 11655 12393 11664 12427
rect 11612 12384 11664 12393
rect 9588 12359 9640 12368
rect 9588 12325 9597 12359
rect 9597 12325 9631 12359
rect 9631 12325 9640 12359
rect 9588 12316 9640 12325
rect 10324 12316 10376 12368
rect 16948 12384 17000 12436
rect 19248 12384 19300 12436
rect 21088 12384 21140 12436
rect 22928 12427 22980 12436
rect 22928 12393 22937 12427
rect 22937 12393 22971 12427
rect 22971 12393 22980 12427
rect 22928 12384 22980 12393
rect 27160 12384 27212 12436
rect 29184 12427 29236 12436
rect 29184 12393 29193 12427
rect 29193 12393 29227 12427
rect 29227 12393 29236 12427
rect 29184 12384 29236 12393
rect 29276 12384 29328 12436
rect 29920 12384 29972 12436
rect 30012 12384 30064 12436
rect 5724 12223 5776 12232
rect 5724 12189 5733 12223
rect 5733 12189 5767 12223
rect 5767 12189 5776 12223
rect 5724 12180 5776 12189
rect 4712 12112 4764 12164
rect 6828 12180 6880 12232
rect 7104 12223 7156 12232
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 7104 12180 7156 12189
rect 7380 12180 7432 12232
rect 7564 12180 7616 12232
rect 8576 12180 8628 12232
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 6920 12112 6972 12164
rect 7840 12112 7892 12164
rect 8208 12112 8260 12164
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 10876 12248 10928 12300
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 5356 12044 5408 12096
rect 8944 12044 8996 12096
rect 10324 12044 10376 12096
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 11888 12112 11940 12164
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 12532 12112 12584 12164
rect 13452 12112 13504 12164
rect 14096 12112 14148 12164
rect 15384 12180 15436 12232
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 16120 12180 16172 12232
rect 18604 12248 18656 12300
rect 24032 12316 24084 12368
rect 24124 12316 24176 12368
rect 18328 12223 18380 12232
rect 18328 12189 18338 12223
rect 18338 12189 18372 12223
rect 18372 12189 18380 12223
rect 18328 12180 18380 12189
rect 17960 12155 18012 12164
rect 17960 12121 17969 12155
rect 17969 12121 18003 12155
rect 18003 12121 18012 12155
rect 17960 12112 18012 12121
rect 18972 12180 19024 12232
rect 19524 12223 19576 12232
rect 19524 12189 19533 12223
rect 19533 12189 19567 12223
rect 19567 12189 19576 12223
rect 19524 12180 19576 12189
rect 19984 12223 20036 12232
rect 19984 12189 19998 12223
rect 19998 12189 20032 12223
rect 20032 12189 20036 12223
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 19984 12180 20036 12189
rect 21916 12180 21968 12232
rect 22008 12180 22060 12232
rect 22468 12180 22520 12232
rect 22744 12223 22796 12232
rect 22744 12189 22753 12223
rect 22753 12189 22787 12223
rect 22787 12189 22796 12223
rect 22744 12180 22796 12189
rect 23112 12180 23164 12232
rect 18512 12155 18564 12164
rect 18512 12121 18521 12155
rect 18521 12121 18555 12155
rect 18555 12121 18564 12155
rect 18512 12112 18564 12121
rect 19156 12112 19208 12164
rect 13728 12044 13780 12096
rect 14924 12044 14976 12096
rect 15292 12044 15344 12096
rect 16120 12087 16172 12096
rect 16120 12053 16129 12087
rect 16129 12053 16163 12087
rect 16163 12053 16172 12087
rect 16120 12044 16172 12053
rect 19708 12044 19760 12096
rect 19892 12155 19944 12164
rect 19892 12121 19901 12155
rect 19901 12121 19935 12155
rect 19935 12121 19944 12155
rect 19892 12112 19944 12121
rect 21824 12112 21876 12164
rect 22652 12087 22704 12096
rect 22652 12053 22661 12087
rect 22661 12053 22695 12087
rect 22695 12053 22704 12087
rect 22652 12044 22704 12053
rect 23756 12112 23808 12164
rect 24124 12223 24176 12232
rect 24124 12189 24133 12223
rect 24133 12189 24167 12223
rect 24167 12189 24176 12223
rect 24124 12180 24176 12189
rect 24216 12223 24268 12232
rect 24216 12189 24225 12223
rect 24225 12189 24259 12223
rect 24259 12189 24268 12223
rect 24216 12180 24268 12189
rect 29276 12248 29328 12300
rect 29552 12248 29604 12300
rect 30104 12291 30156 12300
rect 30104 12257 30113 12291
rect 30113 12257 30147 12291
rect 30147 12257 30156 12291
rect 30104 12248 30156 12257
rect 30656 12316 30708 12368
rect 31576 12316 31628 12368
rect 32036 12384 32088 12436
rect 32956 12427 33008 12436
rect 32956 12393 32965 12427
rect 32965 12393 32999 12427
rect 32999 12393 33008 12427
rect 32956 12384 33008 12393
rect 34704 12427 34756 12436
rect 34704 12393 34713 12427
rect 34713 12393 34747 12427
rect 34747 12393 34756 12427
rect 34704 12384 34756 12393
rect 30932 12248 30984 12300
rect 27988 12180 28040 12232
rect 24400 12112 24452 12164
rect 27804 12112 27856 12164
rect 26240 12044 26292 12096
rect 27988 12044 28040 12096
rect 29644 12180 29696 12232
rect 31116 12180 31168 12232
rect 31300 12223 31352 12232
rect 31300 12189 31309 12223
rect 31309 12189 31343 12223
rect 31343 12189 31352 12223
rect 31300 12180 31352 12189
rect 33324 12248 33376 12300
rect 33416 12291 33468 12300
rect 33416 12257 33425 12291
rect 33425 12257 33459 12291
rect 33459 12257 33468 12291
rect 33416 12248 33468 12257
rect 31576 12180 31628 12232
rect 32128 12223 32180 12232
rect 32128 12189 32137 12223
rect 32137 12189 32171 12223
rect 32171 12189 32180 12223
rect 32128 12180 32180 12189
rect 34888 12223 34940 12232
rect 34888 12189 34897 12223
rect 34897 12189 34931 12223
rect 34931 12189 34940 12223
rect 34888 12180 34940 12189
rect 35992 12180 36044 12232
rect 29920 12087 29972 12096
rect 29920 12053 29929 12087
rect 29929 12053 29963 12087
rect 29963 12053 29972 12087
rect 29920 12044 29972 12053
rect 30288 12044 30340 12096
rect 31944 12044 31996 12096
rect 32036 12087 32088 12096
rect 32036 12053 32045 12087
rect 32045 12053 32079 12087
rect 32079 12053 32088 12087
rect 32036 12044 32088 12053
rect 34796 12044 34848 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 7748 11840 7800 11892
rect 4620 11772 4672 11824
rect 7564 11815 7616 11824
rect 7564 11781 7573 11815
rect 7573 11781 7607 11815
rect 7607 11781 7616 11815
rect 7564 11772 7616 11781
rect 8208 11772 8260 11824
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 7380 11704 7432 11756
rect 7748 11704 7800 11756
rect 7932 11747 7984 11756
rect 7932 11713 7941 11747
rect 7941 11713 7975 11747
rect 7975 11713 7984 11747
rect 7932 11704 7984 11713
rect 8392 11840 8444 11892
rect 11704 11840 11756 11892
rect 12256 11840 12308 11892
rect 12348 11840 12400 11892
rect 12624 11840 12676 11892
rect 12808 11840 12860 11892
rect 9128 11772 9180 11824
rect 10416 11747 10468 11756
rect 10416 11713 10425 11747
rect 10425 11713 10459 11747
rect 10459 11713 10468 11747
rect 10416 11704 10468 11713
rect 10508 11704 10560 11756
rect 8208 11679 8260 11688
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 8576 11636 8628 11688
rect 10324 11679 10376 11688
rect 10324 11645 10333 11679
rect 10333 11645 10367 11679
rect 10367 11645 10376 11679
rect 10324 11636 10376 11645
rect 9128 11568 9180 11620
rect 12440 11747 12492 11756
rect 12440 11713 12449 11747
rect 12449 11713 12483 11747
rect 12483 11713 12492 11747
rect 12440 11704 12492 11713
rect 12532 11747 12584 11756
rect 12532 11713 12541 11747
rect 12541 11713 12575 11747
rect 12575 11713 12584 11747
rect 12532 11704 12584 11713
rect 13084 11747 13136 11756
rect 13084 11713 13093 11747
rect 13093 11713 13127 11747
rect 13127 11713 13136 11747
rect 13084 11704 13136 11713
rect 14280 11840 14332 11892
rect 17960 11840 18012 11892
rect 18236 11772 18288 11824
rect 18512 11840 18564 11892
rect 19064 11840 19116 11892
rect 21824 11883 21876 11892
rect 21824 11849 21833 11883
rect 21833 11849 21867 11883
rect 21867 11849 21876 11883
rect 21824 11840 21876 11849
rect 21916 11840 21968 11892
rect 22100 11840 22152 11892
rect 23756 11840 23808 11892
rect 18696 11772 18748 11824
rect 18880 11815 18932 11824
rect 18880 11781 18889 11815
rect 18889 11781 18923 11815
rect 18923 11781 18932 11815
rect 18880 11772 18932 11781
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 12808 11636 12860 11688
rect 13912 11636 13964 11688
rect 11336 11568 11388 11620
rect 12440 11568 12492 11620
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 16120 11704 16172 11756
rect 17408 11747 17460 11756
rect 17408 11713 17417 11747
rect 17417 11713 17451 11747
rect 17451 11713 17460 11747
rect 17408 11704 17460 11713
rect 17960 11747 18012 11756
rect 17960 11713 17969 11747
rect 17969 11713 18003 11747
rect 18003 11713 18012 11747
rect 17960 11704 18012 11713
rect 18604 11704 18656 11756
rect 19248 11704 19300 11756
rect 19708 11747 19760 11756
rect 19708 11713 19717 11747
rect 19717 11713 19751 11747
rect 19751 11713 19760 11747
rect 19708 11704 19760 11713
rect 19800 11747 19852 11756
rect 19800 11713 19809 11747
rect 19809 11713 19843 11747
rect 19843 11713 19852 11747
rect 19800 11704 19852 11713
rect 19984 11704 20036 11756
rect 20444 11704 20496 11756
rect 18420 11636 18472 11688
rect 22284 11747 22336 11756
rect 22284 11713 22293 11747
rect 22293 11713 22327 11747
rect 22327 11713 22336 11747
rect 22284 11704 22336 11713
rect 22652 11704 22704 11756
rect 23020 11747 23072 11756
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 4620 11500 4672 11552
rect 7288 11543 7340 11552
rect 7288 11509 7297 11543
rect 7297 11509 7331 11543
rect 7331 11509 7340 11543
rect 7288 11500 7340 11509
rect 8024 11543 8076 11552
rect 8024 11509 8033 11543
rect 8033 11509 8067 11543
rect 8067 11509 8076 11543
rect 8024 11500 8076 11509
rect 9404 11500 9456 11552
rect 11612 11500 11664 11552
rect 11980 11543 12032 11552
rect 11980 11509 11989 11543
rect 11989 11509 12023 11543
rect 12023 11509 12032 11543
rect 11980 11500 12032 11509
rect 12072 11500 12124 11552
rect 19524 11568 19576 11620
rect 22836 11679 22888 11688
rect 22836 11645 22845 11679
rect 22845 11645 22879 11679
rect 22879 11645 22888 11679
rect 22836 11636 22888 11645
rect 22928 11679 22980 11688
rect 22928 11645 22937 11679
rect 22937 11645 22971 11679
rect 22971 11645 22980 11679
rect 22928 11636 22980 11645
rect 23020 11568 23072 11620
rect 18696 11543 18748 11552
rect 18696 11509 18705 11543
rect 18705 11509 18739 11543
rect 18739 11509 18748 11543
rect 18696 11500 18748 11509
rect 18972 11500 19024 11552
rect 19984 11500 20036 11552
rect 24400 11772 24452 11824
rect 23756 11747 23808 11756
rect 23756 11713 23765 11747
rect 23765 11713 23799 11747
rect 23799 11713 23808 11747
rect 23756 11704 23808 11713
rect 23848 11747 23900 11756
rect 23848 11713 23857 11747
rect 23857 11713 23891 11747
rect 23891 11713 23900 11747
rect 23848 11704 23900 11713
rect 24032 11704 24084 11756
rect 24584 11747 24636 11756
rect 24584 11713 24593 11747
rect 24593 11713 24627 11747
rect 24627 11713 24636 11747
rect 24584 11704 24636 11713
rect 24124 11679 24176 11688
rect 24124 11645 24133 11679
rect 24133 11645 24167 11679
rect 24167 11645 24176 11679
rect 34888 11840 34940 11892
rect 30288 11747 30340 11756
rect 30288 11713 30297 11747
rect 30297 11713 30331 11747
rect 30331 11713 30340 11747
rect 30288 11704 30340 11713
rect 31300 11772 31352 11824
rect 30656 11704 30708 11756
rect 31760 11772 31812 11824
rect 31668 11704 31720 11756
rect 24124 11636 24176 11645
rect 31392 11636 31444 11688
rect 30380 11568 30432 11620
rect 31760 11679 31812 11688
rect 31760 11645 31769 11679
rect 31769 11645 31803 11679
rect 31803 11645 31812 11679
rect 31760 11636 31812 11645
rect 32128 11636 32180 11688
rect 33140 11747 33192 11756
rect 33140 11713 33149 11747
rect 33149 11713 33183 11747
rect 33183 11713 33192 11747
rect 33140 11704 33192 11713
rect 34612 11704 34664 11756
rect 36268 11704 36320 11756
rect 31576 11568 31628 11620
rect 31944 11568 31996 11620
rect 33508 11679 33560 11688
rect 33508 11645 33517 11679
rect 33517 11645 33551 11679
rect 33551 11645 33560 11679
rect 33508 11636 33560 11645
rect 29920 11500 29972 11552
rect 31024 11500 31076 11552
rect 32220 11500 32272 11552
rect 33600 11500 33652 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 7288 11296 7340 11348
rect 12072 11296 12124 11348
rect 12532 11296 12584 11348
rect 16856 11296 16908 11348
rect 17960 11296 18012 11348
rect 22284 11339 22336 11348
rect 22284 11305 22293 11339
rect 22293 11305 22327 11339
rect 22327 11305 22336 11339
rect 22284 11296 22336 11305
rect 22744 11296 22796 11348
rect 23756 11296 23808 11348
rect 24124 11296 24176 11348
rect 29276 11296 29328 11348
rect 31300 11339 31352 11348
rect 31300 11305 31309 11339
rect 31309 11305 31343 11339
rect 31343 11305 31352 11339
rect 31300 11296 31352 11305
rect 31392 11296 31444 11348
rect 33140 11296 33192 11348
rect 36268 11339 36320 11348
rect 36268 11305 36277 11339
rect 36277 11305 36311 11339
rect 36311 11305 36320 11339
rect 36268 11296 36320 11305
rect 9036 11228 9088 11280
rect 11796 11228 11848 11280
rect 19248 11228 19300 11280
rect 7196 11092 7248 11144
rect 5724 10956 5776 11008
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 11336 11160 11388 11212
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 16856 11160 16908 11212
rect 17776 11160 17828 11212
rect 18604 11160 18656 11212
rect 19984 11228 20036 11280
rect 25044 11228 25096 11280
rect 25688 11228 25740 11280
rect 34796 11228 34848 11280
rect 7840 11024 7892 11076
rect 10324 11092 10376 11144
rect 11796 11135 11848 11144
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 11796 11092 11848 11101
rect 12808 11092 12860 11144
rect 14648 11135 14700 11144
rect 14648 11101 14657 11135
rect 14657 11101 14691 11135
rect 14691 11101 14700 11135
rect 14648 11092 14700 11101
rect 10416 11024 10468 11076
rect 14096 11024 14148 11076
rect 14924 11135 14976 11144
rect 14924 11101 14933 11135
rect 14933 11101 14967 11135
rect 14967 11101 14976 11135
rect 14924 11092 14976 11101
rect 15200 11135 15252 11144
rect 15200 11101 15209 11135
rect 15209 11101 15243 11135
rect 15243 11101 15252 11135
rect 15200 11092 15252 11101
rect 18788 11135 18840 11144
rect 18788 11101 18797 11135
rect 18797 11101 18831 11135
rect 18831 11101 18840 11135
rect 18788 11092 18840 11101
rect 18972 11092 19024 11144
rect 19248 11067 19300 11076
rect 19248 11033 19257 11067
rect 19257 11033 19291 11067
rect 19291 11033 19300 11067
rect 19248 11024 19300 11033
rect 15016 10999 15068 11008
rect 15016 10965 15025 10999
rect 15025 10965 15059 10999
rect 15059 10965 15068 10999
rect 15016 10956 15068 10965
rect 17132 10999 17184 11008
rect 17132 10965 17141 10999
rect 17141 10965 17175 10999
rect 17175 10965 17184 10999
rect 17132 10956 17184 10965
rect 17500 10956 17552 11008
rect 19064 10999 19116 11008
rect 19064 10965 19073 10999
rect 19073 10965 19107 10999
rect 19107 10965 19116 10999
rect 19064 10956 19116 10965
rect 19524 11067 19576 11076
rect 19524 11033 19533 11067
rect 19533 11033 19567 11067
rect 19567 11033 19576 11067
rect 19524 11024 19576 11033
rect 19984 11135 20036 11144
rect 19984 11101 19993 11135
rect 19993 11101 20027 11135
rect 20027 11101 20036 11135
rect 19984 11092 20036 11101
rect 20260 11135 20312 11144
rect 20260 11101 20269 11135
rect 20269 11101 20303 11135
rect 20303 11101 20312 11135
rect 20260 11092 20312 11101
rect 20444 11135 20496 11144
rect 20444 11101 20453 11135
rect 20453 11101 20487 11135
rect 20487 11101 20496 11135
rect 20444 11092 20496 11101
rect 22192 11160 22244 11212
rect 23020 11160 23072 11212
rect 24584 11160 24636 11212
rect 20812 11092 20864 11144
rect 22928 11092 22980 11144
rect 21180 11024 21232 11076
rect 22100 11067 22152 11076
rect 22100 11033 22109 11067
rect 22109 11033 22143 11067
rect 22143 11033 22152 11067
rect 22100 11024 22152 11033
rect 22836 11024 22888 11076
rect 26884 11092 26936 11144
rect 27988 11092 28040 11144
rect 25412 11024 25464 11076
rect 28172 11092 28224 11144
rect 31484 11160 31536 11212
rect 31668 11160 31720 11212
rect 28724 11092 28776 11144
rect 31392 11092 31444 11144
rect 31944 11135 31996 11144
rect 31944 11101 31953 11135
rect 31953 11101 31987 11135
rect 31987 11101 31996 11135
rect 31944 11092 31996 11101
rect 32036 11135 32088 11144
rect 32036 11101 32045 11135
rect 32045 11101 32079 11135
rect 32079 11101 32088 11135
rect 32036 11092 32088 11101
rect 32220 11135 32272 11144
rect 32220 11101 32229 11135
rect 32229 11101 32263 11135
rect 32263 11101 32272 11135
rect 32220 11092 32272 11101
rect 35348 11092 35400 11144
rect 36452 11135 36504 11144
rect 36452 11101 36461 11135
rect 36461 11101 36495 11135
rect 36495 11101 36504 11135
rect 36452 11092 36504 11101
rect 31300 11024 31352 11076
rect 32128 11024 32180 11076
rect 22376 10956 22428 11008
rect 24308 10956 24360 11008
rect 26332 10956 26384 11008
rect 28540 10956 28592 11008
rect 28632 10956 28684 11008
rect 29000 10956 29052 11008
rect 34520 10956 34572 11008
rect 34704 10956 34756 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 7472 10795 7524 10804
rect 7472 10761 7481 10795
rect 7481 10761 7515 10795
rect 7515 10761 7524 10795
rect 7472 10752 7524 10761
rect 9220 10752 9272 10804
rect 14096 10795 14148 10804
rect 14096 10761 14105 10795
rect 14105 10761 14139 10795
rect 14139 10761 14148 10795
rect 14096 10752 14148 10761
rect 14648 10752 14700 10804
rect 15016 10752 15068 10804
rect 4988 10659 5040 10668
rect 4988 10625 4997 10659
rect 4997 10625 5031 10659
rect 5031 10625 5040 10659
rect 4988 10616 5040 10625
rect 5080 10659 5132 10668
rect 5080 10625 5089 10659
rect 5089 10625 5123 10659
rect 5123 10625 5132 10659
rect 5080 10616 5132 10625
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 5908 10659 5960 10668
rect 5908 10625 5917 10659
rect 5917 10625 5951 10659
rect 5951 10625 5960 10659
rect 5908 10616 5960 10625
rect 6920 10616 6972 10668
rect 8024 10684 8076 10736
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 10324 10659 10376 10668
rect 10324 10625 10333 10659
rect 10333 10625 10367 10659
rect 10367 10625 10376 10659
rect 10324 10616 10376 10625
rect 13636 10684 13688 10736
rect 16396 10752 16448 10804
rect 17132 10752 17184 10804
rect 21272 10684 21324 10736
rect 27896 10752 27948 10804
rect 28816 10752 28868 10804
rect 29000 10684 29052 10736
rect 31484 10795 31536 10804
rect 31484 10761 31493 10795
rect 31493 10761 31527 10795
rect 31527 10761 31536 10795
rect 31484 10752 31536 10761
rect 29368 10684 29420 10736
rect 34244 10752 34296 10804
rect 7564 10548 7616 10600
rect 7932 10548 7984 10600
rect 6368 10412 6420 10464
rect 13544 10616 13596 10668
rect 14648 10616 14700 10668
rect 10968 10591 11020 10600
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 11980 10548 12032 10600
rect 13268 10548 13320 10600
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 16764 10616 16816 10668
rect 20628 10616 20680 10668
rect 21916 10659 21968 10668
rect 21916 10625 21925 10659
rect 21925 10625 21959 10659
rect 21959 10625 21968 10659
rect 21916 10616 21968 10625
rect 22284 10616 22336 10668
rect 23940 10616 23992 10668
rect 24216 10616 24268 10668
rect 25044 10659 25096 10668
rect 25044 10625 25053 10659
rect 25053 10625 25087 10659
rect 25087 10625 25096 10659
rect 25044 10616 25096 10625
rect 12348 10480 12400 10532
rect 21364 10548 21416 10600
rect 25136 10548 25188 10600
rect 25412 10591 25464 10600
rect 25412 10557 25421 10591
rect 25421 10557 25455 10591
rect 25455 10557 25464 10591
rect 25412 10548 25464 10557
rect 27712 10548 27764 10600
rect 28172 10616 28224 10668
rect 27988 10548 28040 10600
rect 13452 10412 13504 10464
rect 13820 10412 13872 10464
rect 19248 10480 19300 10532
rect 21272 10480 21324 10532
rect 17776 10412 17828 10464
rect 24768 10480 24820 10532
rect 25044 10480 25096 10532
rect 27620 10480 27672 10532
rect 28632 10616 28684 10668
rect 28816 10659 28868 10668
rect 28816 10625 28825 10659
rect 28825 10625 28859 10659
rect 28859 10625 28868 10659
rect 28816 10616 28868 10625
rect 29644 10659 29696 10668
rect 28540 10591 28592 10600
rect 28540 10557 28549 10591
rect 28549 10557 28583 10591
rect 28583 10557 28592 10591
rect 29644 10625 29653 10659
rect 29653 10625 29687 10659
rect 29687 10625 29696 10659
rect 29644 10616 29696 10625
rect 31300 10659 31352 10668
rect 31300 10625 31309 10659
rect 31309 10625 31343 10659
rect 31343 10625 31352 10659
rect 31300 10616 31352 10625
rect 31392 10659 31444 10668
rect 31392 10625 31401 10659
rect 31401 10625 31435 10659
rect 31435 10625 31444 10659
rect 31392 10616 31444 10625
rect 31668 10659 31720 10668
rect 31668 10625 31677 10659
rect 31677 10625 31711 10659
rect 31711 10625 31720 10659
rect 33232 10684 33284 10736
rect 33968 10684 34020 10736
rect 31668 10616 31720 10625
rect 32220 10659 32272 10668
rect 32220 10625 32229 10659
rect 32229 10625 32263 10659
rect 32263 10625 32272 10659
rect 32220 10616 32272 10625
rect 28540 10548 28592 10557
rect 31024 10548 31076 10600
rect 31944 10591 31996 10600
rect 31944 10557 31953 10591
rect 31953 10557 31987 10591
rect 31987 10557 31996 10591
rect 31944 10548 31996 10557
rect 32036 10548 32088 10600
rect 32864 10616 32916 10668
rect 33416 10616 33468 10668
rect 33600 10659 33652 10668
rect 33600 10625 33609 10659
rect 33609 10625 33643 10659
rect 33643 10625 33652 10659
rect 33600 10616 33652 10625
rect 33784 10659 33836 10668
rect 33784 10625 33793 10659
rect 33793 10625 33827 10659
rect 33827 10625 33836 10659
rect 33784 10616 33836 10625
rect 34152 10616 34204 10668
rect 35900 10752 35952 10804
rect 36360 10795 36412 10804
rect 36360 10761 36369 10795
rect 36369 10761 36403 10795
rect 36403 10761 36412 10795
rect 36360 10752 36412 10761
rect 34796 10616 34848 10668
rect 21824 10412 21876 10464
rect 23296 10412 23348 10464
rect 23848 10412 23900 10464
rect 24676 10412 24728 10464
rect 27160 10412 27212 10464
rect 27804 10412 27856 10464
rect 28908 10480 28960 10532
rect 28816 10412 28868 10464
rect 29092 10455 29144 10464
rect 29092 10421 29101 10455
rect 29101 10421 29135 10455
rect 29135 10421 29144 10455
rect 29092 10412 29144 10421
rect 30288 10480 30340 10532
rect 30104 10412 30156 10464
rect 32956 10591 33008 10600
rect 32956 10557 32965 10591
rect 32965 10557 32999 10591
rect 32999 10557 33008 10591
rect 32956 10548 33008 10557
rect 33232 10548 33284 10600
rect 33876 10591 33928 10600
rect 33876 10557 33885 10591
rect 33885 10557 33919 10591
rect 33919 10557 33928 10591
rect 33876 10548 33928 10557
rect 34704 10548 34756 10600
rect 33140 10480 33192 10532
rect 33508 10480 33560 10532
rect 31852 10455 31904 10464
rect 31852 10421 31861 10455
rect 31861 10421 31895 10455
rect 31895 10421 31904 10455
rect 31852 10412 31904 10421
rect 32680 10412 32732 10464
rect 33600 10412 33652 10464
rect 33784 10412 33836 10464
rect 33968 10412 34020 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4804 10208 4856 10260
rect 5632 10140 5684 10192
rect 7288 10208 7340 10260
rect 7380 10208 7432 10260
rect 9404 10208 9456 10260
rect 12348 10208 12400 10260
rect 12532 10251 12584 10260
rect 12532 10217 12541 10251
rect 12541 10217 12575 10251
rect 12575 10217 12584 10251
rect 12532 10208 12584 10217
rect 13912 10208 13964 10260
rect 14924 10208 14976 10260
rect 16764 10251 16816 10260
rect 16764 10217 16773 10251
rect 16773 10217 16807 10251
rect 16807 10217 16816 10251
rect 16764 10208 16816 10217
rect 17776 10208 17828 10260
rect 4160 10004 4212 10056
rect 4620 10072 4672 10124
rect 5080 10072 5132 10124
rect 4804 10004 4856 10056
rect 4988 10004 5040 10056
rect 1492 9979 1544 9988
rect 1492 9945 1501 9979
rect 1501 9945 1535 9979
rect 1535 9945 1544 9979
rect 1492 9936 1544 9945
rect 5724 9936 5776 9988
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 6920 10004 6972 10056
rect 7104 10115 7156 10124
rect 7104 10081 7113 10115
rect 7113 10081 7147 10115
rect 7147 10081 7156 10115
rect 7104 10072 7156 10081
rect 7380 10047 7432 10056
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 6460 9979 6512 9988
rect 6460 9945 6469 9979
rect 6469 9945 6503 9979
rect 6503 9945 6512 9979
rect 6460 9936 6512 9945
rect 7840 10047 7892 10056
rect 7840 10013 7849 10047
rect 7849 10013 7883 10047
rect 7883 10013 7892 10047
rect 7840 10004 7892 10013
rect 8944 10115 8996 10124
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 13360 10072 13412 10124
rect 13452 10072 13504 10124
rect 13636 10140 13688 10192
rect 12440 10047 12492 10056
rect 12440 10013 12449 10047
rect 12449 10013 12483 10047
rect 12483 10013 12492 10047
rect 12440 10004 12492 10013
rect 13636 10047 13688 10056
rect 13636 10013 13645 10047
rect 13645 10013 13679 10047
rect 13679 10013 13688 10047
rect 13636 10004 13688 10013
rect 9496 9936 9548 9988
rect 11612 9936 11664 9988
rect 11888 9979 11940 9988
rect 11888 9945 11897 9979
rect 11897 9945 11931 9979
rect 11931 9945 11940 9979
rect 11888 9936 11940 9945
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 6552 9868 6604 9920
rect 8576 9868 8628 9920
rect 8944 9868 8996 9920
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12072 9868 12124 9877
rect 15016 10072 15068 10124
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 17132 10047 17184 10056
rect 17132 10013 17141 10047
rect 17141 10013 17175 10047
rect 17175 10013 17184 10047
rect 17132 10004 17184 10013
rect 17316 10115 17368 10124
rect 17316 10081 17325 10115
rect 17325 10081 17359 10115
rect 17359 10081 17368 10115
rect 17316 10072 17368 10081
rect 17592 10072 17644 10124
rect 19248 10115 19300 10124
rect 19248 10081 19257 10115
rect 19257 10081 19291 10115
rect 19291 10081 19300 10115
rect 19248 10072 19300 10081
rect 12808 9868 12860 9920
rect 17408 9936 17460 9988
rect 17776 9979 17828 9988
rect 17776 9945 17785 9979
rect 17785 9945 17819 9979
rect 17819 9945 17828 9979
rect 17776 9936 17828 9945
rect 20812 10004 20864 10056
rect 22376 10208 22428 10260
rect 22100 10140 22152 10192
rect 22560 10140 22612 10192
rect 23204 10208 23256 10260
rect 27712 10208 27764 10260
rect 28632 10208 28684 10260
rect 28816 10208 28868 10260
rect 30656 10208 30708 10260
rect 34796 10208 34848 10260
rect 21824 10115 21876 10124
rect 21824 10081 21833 10115
rect 21833 10081 21867 10115
rect 21867 10081 21876 10115
rect 21824 10072 21876 10081
rect 22008 10072 22060 10124
rect 21364 10047 21416 10056
rect 21364 10013 21373 10047
rect 21373 10013 21407 10047
rect 21407 10013 21416 10047
rect 21364 10004 21416 10013
rect 24768 10115 24820 10124
rect 24768 10081 24777 10115
rect 24777 10081 24811 10115
rect 24811 10081 24820 10115
rect 24768 10072 24820 10081
rect 25964 10072 26016 10124
rect 29368 10140 29420 10192
rect 30196 10140 30248 10192
rect 15660 9868 15712 9920
rect 17500 9868 17552 9920
rect 17960 9868 18012 9920
rect 20628 9911 20680 9920
rect 20628 9877 20637 9911
rect 20637 9877 20671 9911
rect 20671 9877 20680 9911
rect 20628 9868 20680 9877
rect 21548 9936 21600 9988
rect 21732 9936 21784 9988
rect 21824 9868 21876 9920
rect 22468 9868 22520 9920
rect 23112 10047 23164 10056
rect 23112 10013 23121 10047
rect 23121 10013 23155 10047
rect 23155 10013 23164 10047
rect 23112 10004 23164 10013
rect 23204 10047 23256 10056
rect 23204 10013 23213 10047
rect 23213 10013 23247 10047
rect 23247 10013 23256 10047
rect 23204 10004 23256 10013
rect 23664 10004 23716 10056
rect 24400 10047 24452 10056
rect 24400 10013 24409 10047
rect 24409 10013 24443 10047
rect 24443 10013 24452 10047
rect 24400 10004 24452 10013
rect 27160 10047 27212 10056
rect 27160 10013 27169 10047
rect 27169 10013 27203 10047
rect 27203 10013 27212 10047
rect 27160 10004 27212 10013
rect 27252 10004 27304 10056
rect 23296 9936 23348 9988
rect 26056 9936 26108 9988
rect 22652 9868 22704 9920
rect 23020 9911 23072 9920
rect 23020 9877 23029 9911
rect 23029 9877 23063 9911
rect 23063 9877 23072 9911
rect 23020 9868 23072 9877
rect 23112 9868 23164 9920
rect 23940 9868 23992 9920
rect 24952 9868 25004 9920
rect 28540 10004 28592 10056
rect 28908 10115 28960 10124
rect 28908 10081 28917 10115
rect 28917 10081 28951 10115
rect 28951 10081 28960 10115
rect 28908 10072 28960 10081
rect 29092 10072 29144 10124
rect 32036 10140 32088 10192
rect 31668 10072 31720 10124
rect 29828 9979 29880 9988
rect 29828 9945 29837 9979
rect 29837 9945 29871 9979
rect 29871 9945 29880 9979
rect 29828 9936 29880 9945
rect 30104 10047 30156 10056
rect 30104 10013 30113 10047
rect 30113 10013 30147 10047
rect 30147 10013 30156 10047
rect 30104 10004 30156 10013
rect 30288 10004 30340 10056
rect 31024 10004 31076 10056
rect 31208 10004 31260 10056
rect 32220 10004 32272 10056
rect 33140 10072 33192 10124
rect 33784 10072 33836 10124
rect 33968 10115 34020 10124
rect 33968 10081 33977 10115
rect 33977 10081 34011 10115
rect 34011 10081 34020 10115
rect 33968 10072 34020 10081
rect 32680 10047 32732 10056
rect 32680 10013 32689 10047
rect 32689 10013 32723 10047
rect 32723 10013 32732 10047
rect 32680 10004 32732 10013
rect 32864 10004 32916 10056
rect 32956 10047 33008 10056
rect 32956 10013 32965 10047
rect 32965 10013 32999 10047
rect 32999 10013 33008 10047
rect 32956 10004 33008 10013
rect 30748 9936 30800 9988
rect 33692 10047 33744 10056
rect 33692 10013 33701 10047
rect 33701 10013 33735 10047
rect 33735 10013 33744 10047
rect 33692 10004 33744 10013
rect 34336 10004 34388 10056
rect 35900 10004 35952 10056
rect 29920 9868 29972 9920
rect 30012 9911 30064 9920
rect 30012 9877 30021 9911
rect 30021 9877 30055 9911
rect 30055 9877 30064 9911
rect 30012 9868 30064 9877
rect 30288 9868 30340 9920
rect 31392 9868 31444 9920
rect 31760 9911 31812 9920
rect 31760 9877 31769 9911
rect 31769 9877 31803 9911
rect 31803 9877 31812 9911
rect 31760 9868 31812 9877
rect 31944 9868 31996 9920
rect 33140 9911 33192 9920
rect 33140 9877 33149 9911
rect 33149 9877 33183 9911
rect 33183 9877 33192 9911
rect 33140 9868 33192 9877
rect 34888 9911 34940 9920
rect 34888 9877 34897 9911
rect 34897 9877 34931 9911
rect 34931 9877 34940 9911
rect 34888 9868 34940 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 6552 9664 6604 9716
rect 8944 9664 8996 9716
rect 5540 9596 5592 9648
rect 4804 9528 4856 9580
rect 5632 9528 5684 9580
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 7932 9596 7984 9648
rect 12072 9664 12124 9716
rect 14924 9664 14976 9716
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 9588 9571 9640 9580
rect 9588 9537 9597 9571
rect 9597 9537 9631 9571
rect 9631 9537 9640 9571
rect 9588 9528 9640 9537
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 5448 9460 5500 9512
rect 5908 9460 5960 9512
rect 6460 9460 6512 9512
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 7380 9392 7432 9444
rect 9588 9392 9640 9444
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 12532 9596 12584 9648
rect 14556 9596 14608 9648
rect 17776 9664 17828 9716
rect 18880 9596 18932 9648
rect 21548 9707 21600 9716
rect 21548 9673 21557 9707
rect 21557 9673 21591 9707
rect 21591 9673 21600 9707
rect 21548 9664 21600 9673
rect 22652 9664 22704 9716
rect 23664 9664 23716 9716
rect 26056 9664 26108 9716
rect 30012 9664 30064 9716
rect 23020 9596 23072 9648
rect 24952 9596 25004 9648
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 12992 9571 13044 9580
rect 12992 9537 13006 9571
rect 13006 9537 13040 9571
rect 13040 9537 13044 9571
rect 12992 9528 13044 9537
rect 14832 9528 14884 9580
rect 16672 9571 16724 9580
rect 16672 9537 16681 9571
rect 16681 9537 16715 9571
rect 16715 9537 16724 9571
rect 16672 9528 16724 9537
rect 17316 9528 17368 9580
rect 11888 9503 11940 9512
rect 11888 9469 11897 9503
rect 11897 9469 11931 9503
rect 11931 9469 11940 9503
rect 11888 9460 11940 9469
rect 15568 9460 15620 9512
rect 17960 9503 18012 9512
rect 17960 9469 17969 9503
rect 17969 9469 18003 9503
rect 18003 9469 18012 9503
rect 17960 9460 18012 9469
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 21732 9528 21784 9580
rect 20812 9460 20864 9512
rect 16856 9435 16908 9444
rect 16856 9401 16865 9435
rect 16865 9401 16899 9435
rect 16899 9401 16908 9435
rect 16856 9392 16908 9401
rect 17316 9392 17368 9444
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 9312 9367 9364 9376
rect 9312 9333 9321 9367
rect 9321 9333 9355 9367
rect 9355 9333 9364 9367
rect 9312 9324 9364 9333
rect 9496 9324 9548 9376
rect 11336 9324 11388 9376
rect 17224 9324 17276 9376
rect 22008 9392 22060 9444
rect 21088 9367 21140 9376
rect 21088 9333 21097 9367
rect 21097 9333 21131 9367
rect 21131 9333 21140 9367
rect 21088 9324 21140 9333
rect 23572 9571 23624 9580
rect 23572 9537 23581 9571
rect 23581 9537 23615 9571
rect 23615 9537 23624 9571
rect 23572 9528 23624 9537
rect 22560 9460 22612 9512
rect 23204 9460 23256 9512
rect 22928 9392 22980 9444
rect 24216 9571 24268 9580
rect 24216 9537 24225 9571
rect 24225 9537 24259 9571
rect 24259 9537 24268 9571
rect 24216 9528 24268 9537
rect 24676 9571 24728 9580
rect 24676 9537 24685 9571
rect 24685 9537 24719 9571
rect 24719 9537 24728 9571
rect 24676 9528 24728 9537
rect 25136 9571 25188 9580
rect 25136 9537 25145 9571
rect 25145 9537 25179 9571
rect 25179 9537 25188 9571
rect 25136 9528 25188 9537
rect 30104 9639 30156 9648
rect 30104 9605 30113 9639
rect 30113 9605 30147 9639
rect 30147 9605 30156 9639
rect 30104 9596 30156 9605
rect 31576 9664 31628 9716
rect 31944 9664 31996 9716
rect 33692 9664 33744 9716
rect 25964 9571 26016 9580
rect 25964 9537 25973 9571
rect 25973 9537 26007 9571
rect 26007 9537 26016 9571
rect 25964 9528 26016 9537
rect 29828 9528 29880 9580
rect 24032 9460 24084 9512
rect 29276 9460 29328 9512
rect 24860 9392 24912 9444
rect 27712 9392 27764 9444
rect 28908 9392 28960 9444
rect 30748 9571 30800 9580
rect 30748 9537 30757 9571
rect 30757 9537 30791 9571
rect 30791 9537 30800 9571
rect 30748 9528 30800 9537
rect 31760 9528 31812 9580
rect 33140 9596 33192 9648
rect 33600 9596 33652 9648
rect 33048 9528 33100 9580
rect 34888 9664 34940 9716
rect 33232 9460 33284 9512
rect 26424 9324 26476 9376
rect 30472 9324 30524 9376
rect 34244 9503 34296 9512
rect 34244 9469 34253 9503
rect 34253 9469 34287 9503
rect 34287 9469 34296 9503
rect 34244 9460 34296 9469
rect 34336 9503 34388 9512
rect 34336 9469 34345 9503
rect 34345 9469 34379 9503
rect 34379 9469 34388 9503
rect 34336 9460 34388 9469
rect 30932 9367 30984 9376
rect 30932 9333 30941 9367
rect 30941 9333 30975 9367
rect 30975 9333 30984 9367
rect 30932 9324 30984 9333
rect 32312 9324 32364 9376
rect 33140 9324 33192 9376
rect 33416 9367 33468 9376
rect 33416 9333 33425 9367
rect 33425 9333 33459 9367
rect 33459 9333 33468 9367
rect 33416 9324 33468 9333
rect 33876 9324 33928 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 10968 9163 11020 9172
rect 10968 9129 10977 9163
rect 10977 9129 11011 9163
rect 11011 9129 11020 9163
rect 10968 9120 11020 9129
rect 11336 9120 11388 9172
rect 13176 9120 13228 9172
rect 14280 9120 14332 9172
rect 14464 9163 14516 9172
rect 14464 9129 14473 9163
rect 14473 9129 14507 9163
rect 14507 9129 14516 9163
rect 14464 9120 14516 9129
rect 14832 9163 14884 9172
rect 14832 9129 14841 9163
rect 14841 9129 14875 9163
rect 14875 9129 14884 9163
rect 14832 9120 14884 9129
rect 22100 9120 22152 9172
rect 11888 9052 11940 9104
rect 11980 9052 12032 9104
rect 12164 9052 12216 9104
rect 16856 9052 16908 9104
rect 20996 9052 21048 9104
rect 22008 9052 22060 9104
rect 7932 8984 7984 9036
rect 4160 8916 4212 8968
rect 10416 8959 10468 8968
rect 10416 8925 10425 8959
rect 10425 8925 10459 8959
rect 10459 8925 10468 8959
rect 10416 8916 10468 8925
rect 11520 8984 11572 9036
rect 10508 8848 10560 8900
rect 5264 8780 5316 8832
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 11428 8959 11480 8968
rect 11428 8925 11437 8959
rect 11437 8925 11471 8959
rect 11471 8925 11480 8959
rect 11428 8916 11480 8925
rect 11612 8959 11664 8968
rect 11612 8925 11621 8959
rect 11621 8925 11655 8959
rect 11655 8925 11664 8959
rect 11612 8916 11664 8925
rect 12716 8916 12768 8968
rect 11980 8848 12032 8900
rect 12440 8848 12492 8900
rect 12624 8848 12676 8900
rect 16212 8848 16264 8900
rect 16488 8848 16540 8900
rect 17224 8916 17276 8968
rect 17316 8959 17368 8968
rect 17316 8925 17325 8959
rect 17325 8925 17359 8959
rect 17359 8925 17368 8959
rect 17316 8916 17368 8925
rect 20904 8916 20956 8968
rect 21272 8916 21324 8968
rect 21916 8984 21968 9036
rect 22928 9027 22980 9036
rect 22928 8993 22937 9027
rect 22937 8993 22971 9027
rect 22971 8993 22980 9027
rect 22928 8984 22980 8993
rect 22560 8959 22612 8968
rect 22560 8925 22569 8959
rect 22569 8925 22603 8959
rect 22603 8925 22612 8959
rect 22560 8916 22612 8925
rect 23572 9163 23624 9172
rect 23572 9129 23581 9163
rect 23581 9129 23615 9163
rect 23615 9129 23624 9163
rect 23572 9120 23624 9129
rect 23204 9052 23256 9104
rect 24032 9163 24084 9172
rect 24032 9129 24041 9163
rect 24041 9129 24075 9163
rect 24075 9129 24084 9163
rect 24032 9120 24084 9129
rect 26424 9120 26476 9172
rect 27344 9052 27396 9104
rect 29920 9120 29972 9172
rect 34244 9120 34296 9172
rect 23572 8916 23624 8968
rect 26792 8984 26844 9036
rect 23940 8916 23992 8968
rect 25136 8916 25188 8968
rect 27804 8959 27856 8968
rect 27804 8925 27813 8959
rect 27813 8925 27847 8959
rect 27847 8925 27856 8959
rect 27804 8916 27856 8925
rect 27896 8959 27948 8968
rect 27896 8925 27905 8959
rect 27905 8925 27939 8959
rect 27939 8925 27948 8959
rect 27896 8916 27948 8925
rect 36176 8984 36228 9036
rect 30932 8916 30984 8968
rect 12348 8780 12400 8832
rect 15200 8780 15252 8832
rect 15292 8780 15344 8832
rect 16028 8780 16080 8832
rect 16396 8823 16448 8832
rect 16396 8789 16405 8823
rect 16405 8789 16439 8823
rect 16439 8789 16448 8823
rect 16396 8780 16448 8789
rect 18696 8823 18748 8832
rect 18696 8789 18705 8823
rect 18705 8789 18739 8823
rect 18739 8789 18748 8823
rect 18696 8780 18748 8789
rect 27896 8780 27948 8832
rect 28264 8891 28316 8900
rect 28264 8857 28273 8891
rect 28273 8857 28307 8891
rect 28307 8857 28316 8891
rect 28264 8848 28316 8857
rect 31852 8848 31904 8900
rect 29184 8780 29236 8832
rect 30564 8780 30616 8832
rect 32128 8780 32180 8832
rect 33048 8780 33100 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 8576 8508 8628 8560
rect 12624 8576 12676 8628
rect 12900 8576 12952 8628
rect 14004 8576 14056 8628
rect 16028 8576 16080 8628
rect 16580 8576 16632 8628
rect 7196 8440 7248 8492
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 9312 8440 9364 8492
rect 5816 8372 5868 8424
rect 12624 8440 12676 8492
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 13728 8440 13780 8492
rect 16396 8508 16448 8560
rect 20076 8508 20128 8560
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 12440 8372 12492 8424
rect 14188 8372 14240 8424
rect 14648 8440 14700 8492
rect 15108 8440 15160 8492
rect 15200 8440 15252 8492
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 20996 8440 21048 8492
rect 21272 8483 21324 8492
rect 21272 8449 21281 8483
rect 21281 8449 21315 8483
rect 21315 8449 21324 8483
rect 21272 8440 21324 8449
rect 21732 8440 21784 8492
rect 22560 8576 22612 8628
rect 23940 8619 23992 8628
rect 23940 8585 23949 8619
rect 23949 8585 23983 8619
rect 23983 8585 23992 8619
rect 23940 8576 23992 8585
rect 26792 8619 26844 8628
rect 26792 8585 26801 8619
rect 26801 8585 26835 8619
rect 26835 8585 26844 8619
rect 26792 8576 26844 8585
rect 28448 8576 28500 8628
rect 32036 8576 32088 8628
rect 22100 8440 22152 8492
rect 14556 8415 14608 8424
rect 14556 8381 14565 8415
rect 14565 8381 14599 8415
rect 14599 8381 14608 8415
rect 14556 8372 14608 8381
rect 17776 8372 17828 8424
rect 22836 8440 22888 8492
rect 26516 8483 26568 8492
rect 26516 8449 26525 8483
rect 26525 8449 26559 8483
rect 26559 8449 26568 8483
rect 26516 8440 26568 8449
rect 12532 8304 12584 8356
rect 13636 8347 13688 8356
rect 13636 8313 13645 8347
rect 13645 8313 13679 8347
rect 13679 8313 13688 8347
rect 13636 8304 13688 8313
rect 19064 8304 19116 8356
rect 23572 8372 23624 8424
rect 27620 8508 27672 8560
rect 27344 8483 27396 8492
rect 27344 8449 27353 8483
rect 27353 8449 27387 8483
rect 27387 8449 27396 8483
rect 27344 8440 27396 8449
rect 27712 8483 27764 8492
rect 27712 8449 27721 8483
rect 27721 8449 27755 8483
rect 27755 8449 27764 8483
rect 27712 8440 27764 8449
rect 1492 8236 1544 8288
rect 7012 8236 7064 8288
rect 7656 8236 7708 8288
rect 11888 8236 11940 8288
rect 13544 8236 13596 8288
rect 20720 8236 20772 8288
rect 21088 8347 21140 8356
rect 21088 8313 21097 8347
rect 21097 8313 21131 8347
rect 21131 8313 21140 8347
rect 21088 8304 21140 8313
rect 24216 8304 24268 8356
rect 27528 8372 27580 8424
rect 28356 8483 28408 8492
rect 28356 8449 28365 8483
rect 28365 8449 28399 8483
rect 28399 8449 28408 8483
rect 28356 8440 28408 8449
rect 29184 8551 29236 8560
rect 29184 8517 29193 8551
rect 29193 8517 29227 8551
rect 29227 8517 29236 8551
rect 29184 8508 29236 8517
rect 32128 8551 32180 8560
rect 32128 8517 32137 8551
rect 32137 8517 32171 8551
rect 32171 8517 32180 8551
rect 32128 8508 32180 8517
rect 31852 8440 31904 8492
rect 32956 8576 33008 8628
rect 34336 8576 34388 8628
rect 33048 8508 33100 8560
rect 34244 8508 34296 8560
rect 32864 8483 32916 8492
rect 32864 8449 32873 8483
rect 32873 8449 32907 8483
rect 32907 8449 32916 8483
rect 32864 8440 32916 8449
rect 32404 8372 32456 8424
rect 27436 8347 27488 8356
rect 27436 8313 27445 8347
rect 27445 8313 27479 8347
rect 27479 8313 27488 8347
rect 27436 8304 27488 8313
rect 31668 8304 31720 8356
rect 34612 8347 34664 8356
rect 34612 8313 34621 8347
rect 34621 8313 34655 8347
rect 34655 8313 34664 8347
rect 34612 8304 34664 8313
rect 26332 8236 26384 8288
rect 27252 8236 27304 8288
rect 29184 8236 29236 8288
rect 29368 8279 29420 8288
rect 29368 8245 29377 8279
rect 29377 8245 29411 8279
rect 29411 8245 29420 8279
rect 29368 8236 29420 8245
rect 30012 8236 30064 8288
rect 31944 8236 31996 8288
rect 32404 8236 32456 8288
rect 32496 8279 32548 8288
rect 32496 8245 32505 8279
rect 32505 8245 32539 8279
rect 32539 8245 32548 8279
rect 32496 8236 32548 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 5356 8032 5408 8084
rect 5448 7964 5500 8016
rect 6368 8032 6420 8084
rect 7012 8032 7064 8084
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 5356 7828 5408 7880
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 7288 7896 7340 7948
rect 6736 7828 6788 7880
rect 4620 7735 4672 7744
rect 4620 7701 4629 7735
rect 4629 7701 4663 7735
rect 4663 7701 4672 7735
rect 4620 7692 4672 7701
rect 5448 7803 5500 7812
rect 5448 7769 5457 7803
rect 5457 7769 5491 7803
rect 5491 7769 5500 7803
rect 5448 7760 5500 7769
rect 6920 7828 6972 7880
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 11428 8032 11480 8084
rect 12164 8032 12216 8084
rect 13820 8075 13872 8084
rect 13820 8041 13829 8075
rect 13829 8041 13863 8075
rect 13863 8041 13872 8075
rect 13820 8032 13872 8041
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 17224 8032 17276 8084
rect 18880 8075 18932 8084
rect 18880 8041 18889 8075
rect 18889 8041 18923 8075
rect 18923 8041 18932 8075
rect 18880 8032 18932 8041
rect 7472 7896 7524 7948
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 17132 7964 17184 8016
rect 7932 7828 7984 7880
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 8392 7828 8444 7837
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10324 7828 10376 7880
rect 10784 7828 10836 7880
rect 7840 7692 7892 7744
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 12164 7939 12216 7948
rect 12164 7905 12173 7939
rect 12173 7905 12207 7939
rect 12207 7905 12216 7939
rect 12164 7896 12216 7905
rect 13544 7896 13596 7948
rect 13636 7896 13688 7948
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 18236 7896 18288 7948
rect 19064 7896 19116 7948
rect 26332 8032 26384 8084
rect 26516 8032 26568 8084
rect 28356 8032 28408 8084
rect 30564 8032 30616 8084
rect 31760 8032 31812 8084
rect 21916 7964 21968 8016
rect 27712 7964 27764 8016
rect 14280 7828 14332 7880
rect 13176 7760 13228 7812
rect 14464 7828 14516 7880
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 18420 7871 18472 7880
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 18604 7828 18656 7880
rect 19248 7871 19300 7880
rect 19248 7837 19257 7871
rect 19257 7837 19291 7871
rect 19291 7837 19300 7871
rect 19248 7828 19300 7837
rect 20812 7871 20864 7880
rect 20812 7837 20821 7871
rect 20821 7837 20855 7871
rect 20855 7837 20864 7871
rect 20812 7828 20864 7837
rect 21272 7896 21324 7948
rect 26608 7896 26660 7948
rect 27620 7939 27672 7948
rect 27620 7905 27629 7939
rect 27629 7905 27663 7939
rect 27663 7905 27672 7939
rect 27620 7896 27672 7905
rect 27896 7896 27948 7948
rect 18696 7760 18748 7812
rect 21088 7760 21140 7812
rect 21364 7828 21416 7880
rect 21640 7871 21692 7880
rect 21640 7837 21649 7871
rect 21649 7837 21683 7871
rect 21683 7837 21692 7871
rect 21640 7828 21692 7837
rect 21824 7871 21876 7880
rect 21824 7837 21833 7871
rect 21833 7837 21867 7871
rect 21867 7837 21876 7871
rect 21824 7828 21876 7837
rect 22744 7871 22796 7880
rect 22744 7837 22753 7871
rect 22753 7837 22787 7871
rect 22787 7837 22796 7871
rect 22744 7828 22796 7837
rect 22836 7871 22888 7880
rect 22836 7837 22845 7871
rect 22845 7837 22879 7871
rect 22879 7837 22888 7871
rect 22836 7828 22888 7837
rect 12532 7692 12584 7744
rect 17592 7735 17644 7744
rect 17592 7701 17601 7735
rect 17601 7701 17635 7735
rect 17635 7701 17644 7735
rect 17592 7692 17644 7701
rect 18420 7692 18472 7744
rect 22376 7760 22428 7812
rect 23480 7828 23532 7880
rect 25044 7828 25096 7880
rect 26792 7828 26844 7880
rect 21456 7692 21508 7744
rect 22192 7692 22244 7744
rect 24124 7760 24176 7812
rect 25964 7760 26016 7812
rect 27528 7871 27580 7880
rect 27528 7837 27537 7871
rect 27537 7837 27571 7871
rect 27571 7837 27580 7871
rect 27528 7828 27580 7837
rect 30196 7896 30248 7948
rect 30472 7896 30524 7948
rect 32956 7964 33008 8016
rect 33600 7964 33652 8016
rect 34060 7964 34112 8016
rect 29184 7803 29236 7812
rect 29184 7769 29193 7803
rect 29193 7769 29227 7803
rect 29227 7769 29236 7803
rect 29184 7760 29236 7769
rect 30012 7871 30064 7880
rect 30012 7837 30021 7871
rect 30021 7837 30055 7871
rect 30055 7837 30064 7871
rect 30012 7828 30064 7837
rect 30472 7803 30524 7812
rect 30472 7769 30493 7803
rect 30493 7769 30524 7803
rect 30472 7760 30524 7769
rect 30748 7871 30800 7880
rect 30748 7837 30757 7871
rect 30757 7837 30791 7871
rect 30791 7837 30800 7871
rect 30748 7828 30800 7837
rect 30840 7828 30892 7880
rect 31116 7871 31168 7880
rect 31116 7837 31125 7871
rect 31125 7837 31159 7871
rect 31159 7837 31168 7871
rect 31116 7828 31168 7837
rect 31208 7871 31260 7880
rect 31208 7837 31217 7871
rect 31217 7837 31251 7871
rect 31251 7837 31260 7871
rect 31208 7828 31260 7837
rect 31576 7828 31628 7880
rect 31392 7760 31444 7812
rect 31852 7828 31904 7880
rect 32036 7871 32088 7880
rect 32036 7837 32045 7871
rect 32045 7837 32079 7871
rect 32079 7837 32088 7871
rect 32036 7828 32088 7837
rect 28172 7692 28224 7744
rect 28448 7692 28500 7744
rect 29092 7692 29144 7744
rect 29736 7735 29788 7744
rect 29736 7701 29745 7735
rect 29745 7701 29779 7735
rect 29779 7701 29788 7735
rect 29736 7692 29788 7701
rect 31484 7692 31536 7744
rect 32220 7803 32272 7812
rect 32220 7769 32229 7803
rect 32229 7769 32263 7803
rect 32263 7769 32272 7803
rect 32220 7760 32272 7769
rect 31944 7735 31996 7744
rect 31944 7701 31953 7735
rect 31953 7701 31987 7735
rect 31987 7701 31996 7735
rect 31944 7692 31996 7701
rect 32036 7692 32088 7744
rect 32680 7760 32732 7812
rect 32956 7760 33008 7812
rect 33324 7871 33376 7880
rect 33324 7837 33333 7871
rect 33333 7837 33367 7871
rect 33367 7837 33376 7871
rect 33324 7828 33376 7837
rect 34520 7828 34572 7880
rect 34704 7871 34756 7880
rect 34704 7837 34713 7871
rect 34713 7837 34747 7871
rect 34747 7837 34756 7871
rect 34704 7828 34756 7837
rect 36452 7871 36504 7880
rect 36452 7837 36461 7871
rect 36461 7837 36495 7871
rect 36495 7837 36504 7871
rect 36452 7828 36504 7837
rect 33692 7760 33744 7812
rect 34060 7760 34112 7812
rect 32864 7692 32916 7744
rect 34520 7692 34572 7744
rect 36268 7735 36320 7744
rect 36268 7701 36277 7735
rect 36277 7701 36311 7735
rect 36311 7701 36320 7735
rect 36268 7692 36320 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 7104 7488 7156 7540
rect 7564 7488 7616 7540
rect 9956 7488 10008 7540
rect 10324 7531 10376 7540
rect 10324 7497 10333 7531
rect 10333 7497 10367 7531
rect 10367 7497 10376 7531
rect 10324 7488 10376 7497
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 12808 7488 12860 7540
rect 19984 7531 20036 7540
rect 19984 7497 19993 7531
rect 19993 7497 20027 7531
rect 20027 7497 20036 7531
rect 19984 7488 20036 7497
rect 20996 7531 21048 7540
rect 20996 7497 21005 7531
rect 21005 7497 21039 7531
rect 21039 7497 21048 7531
rect 20996 7488 21048 7497
rect 21272 7488 21324 7540
rect 5448 7352 5500 7404
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 5816 7284 5868 7336
rect 7196 7352 7248 7404
rect 7564 7352 7616 7404
rect 16580 7420 16632 7472
rect 20444 7420 20496 7472
rect 8116 7352 8168 7404
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 11980 7352 12032 7361
rect 12532 7352 12584 7404
rect 12716 7352 12768 7404
rect 13820 7352 13872 7404
rect 14280 7352 14332 7404
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 14188 7284 14240 7336
rect 16580 7284 16632 7336
rect 17316 7352 17368 7404
rect 19892 7395 19944 7404
rect 19892 7361 19901 7395
rect 19901 7361 19935 7395
rect 19935 7361 19944 7395
rect 19892 7352 19944 7361
rect 20076 7395 20128 7404
rect 20076 7361 20085 7395
rect 20085 7361 20119 7395
rect 20119 7361 20128 7395
rect 20076 7352 20128 7361
rect 20536 7352 20588 7404
rect 21272 7352 21324 7404
rect 21456 7395 21508 7404
rect 21456 7361 21465 7395
rect 21465 7361 21499 7395
rect 21499 7361 21508 7395
rect 21456 7352 21508 7361
rect 22008 7420 22060 7472
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 22744 7488 22796 7540
rect 23480 7531 23532 7540
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 24124 7531 24176 7540
rect 24124 7497 24133 7531
rect 24133 7497 24167 7531
rect 24167 7497 24176 7531
rect 24124 7488 24176 7497
rect 27528 7488 27580 7540
rect 30472 7488 30524 7540
rect 30748 7531 30800 7540
rect 30748 7497 30757 7531
rect 30757 7497 30791 7531
rect 30791 7497 30800 7531
rect 30748 7488 30800 7497
rect 33324 7488 33376 7540
rect 33692 7488 33744 7540
rect 23848 7420 23900 7472
rect 29736 7420 29788 7472
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 4620 7216 4672 7268
rect 9864 7216 9916 7268
rect 23572 7284 23624 7336
rect 24308 7352 24360 7404
rect 24216 7327 24268 7336
rect 24216 7293 24225 7327
rect 24225 7293 24259 7327
rect 24259 7293 24268 7327
rect 24216 7284 24268 7293
rect 12808 7148 12860 7200
rect 17592 7148 17644 7200
rect 18512 7148 18564 7200
rect 22376 7216 22428 7268
rect 24952 7327 25004 7336
rect 24952 7293 24961 7327
rect 24961 7293 24995 7327
rect 24995 7293 25004 7327
rect 24952 7284 25004 7293
rect 26608 7284 26660 7336
rect 29092 7395 29144 7404
rect 29092 7361 29101 7395
rect 29101 7361 29135 7395
rect 29135 7361 29144 7395
rect 29092 7352 29144 7361
rect 21640 7148 21692 7200
rect 21916 7148 21968 7200
rect 22008 7148 22060 7200
rect 26700 7216 26752 7268
rect 29920 7284 29972 7336
rect 30380 7352 30432 7404
rect 30564 7352 30616 7404
rect 30840 7352 30892 7404
rect 30748 7327 30800 7336
rect 30748 7293 30757 7327
rect 30757 7293 30791 7327
rect 30791 7293 30800 7327
rect 30748 7284 30800 7293
rect 31208 7395 31260 7404
rect 31208 7361 31217 7395
rect 31217 7361 31251 7395
rect 31251 7361 31260 7395
rect 31208 7352 31260 7361
rect 31392 7352 31444 7404
rect 31944 7395 31996 7404
rect 31944 7361 31953 7395
rect 31953 7361 31987 7395
rect 31987 7361 31996 7395
rect 31944 7352 31996 7361
rect 33876 7463 33928 7472
rect 33876 7429 33885 7463
rect 33885 7429 33919 7463
rect 33919 7429 33928 7463
rect 33876 7420 33928 7429
rect 32404 7395 32456 7404
rect 32404 7361 32413 7395
rect 32413 7361 32447 7395
rect 32447 7361 32456 7395
rect 32404 7352 32456 7361
rect 32680 7395 32732 7404
rect 32680 7361 32689 7395
rect 32689 7361 32723 7395
rect 32723 7361 32732 7395
rect 32680 7352 32732 7361
rect 31668 7284 31720 7336
rect 33784 7395 33836 7404
rect 33784 7361 33793 7395
rect 33793 7361 33827 7395
rect 33827 7361 33836 7395
rect 33784 7352 33836 7361
rect 34612 7488 34664 7540
rect 34796 7488 34848 7540
rect 33968 7284 34020 7336
rect 34336 7352 34388 7404
rect 34520 7395 34572 7404
rect 34520 7361 34529 7395
rect 34529 7361 34563 7395
rect 34563 7361 34572 7395
rect 34520 7352 34572 7361
rect 31760 7259 31812 7268
rect 31760 7225 31769 7259
rect 31769 7225 31803 7259
rect 31803 7225 31812 7259
rect 31760 7216 31812 7225
rect 32496 7216 32548 7268
rect 34796 7284 34848 7336
rect 23940 7148 23992 7200
rect 25964 7148 26016 7200
rect 29460 7148 29512 7200
rect 30564 7191 30616 7200
rect 30564 7157 30573 7191
rect 30573 7157 30607 7191
rect 30607 7157 30616 7191
rect 30564 7148 30616 7157
rect 31300 7148 31352 7200
rect 32312 7148 32364 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 5816 6876 5868 6928
rect 10232 6944 10284 6996
rect 11980 6944 12032 6996
rect 11796 6876 11848 6928
rect 5448 6808 5500 6860
rect 12716 6808 12768 6860
rect 14464 6808 14516 6860
rect 19248 6944 19300 6996
rect 20904 6944 20956 6996
rect 22008 6944 22060 6996
rect 23572 6987 23624 6996
rect 23572 6953 23581 6987
rect 23581 6953 23615 6987
rect 23615 6953 23624 6987
rect 23572 6944 23624 6953
rect 31024 6944 31076 6996
rect 33600 6944 33652 6996
rect 17132 6876 17184 6928
rect 25964 6876 26016 6928
rect 29368 6876 29420 6928
rect 33784 6876 33836 6928
rect 1952 6672 2004 6724
rect 11060 6740 11112 6792
rect 16672 6808 16724 6860
rect 18236 6808 18288 6860
rect 20444 6808 20496 6860
rect 22100 6808 22152 6860
rect 22376 6851 22428 6860
rect 22376 6817 22385 6851
rect 22385 6817 22419 6851
rect 22419 6817 22428 6851
rect 22376 6808 22428 6817
rect 14464 6672 14516 6724
rect 5264 6604 5316 6656
rect 6368 6604 6420 6656
rect 7288 6604 7340 6656
rect 7840 6604 7892 6656
rect 8576 6604 8628 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 18328 6783 18380 6792
rect 18328 6749 18337 6783
rect 18337 6749 18371 6783
rect 18371 6749 18380 6783
rect 18328 6740 18380 6749
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 18972 6783 19024 6792
rect 18972 6749 18981 6783
rect 18981 6749 19015 6783
rect 19015 6749 19024 6783
rect 18972 6740 19024 6749
rect 20812 6740 20864 6792
rect 18696 6715 18748 6724
rect 18696 6681 18705 6715
rect 18705 6681 18739 6715
rect 18739 6681 18748 6715
rect 18696 6672 18748 6681
rect 21916 6783 21968 6792
rect 21916 6749 21925 6783
rect 21925 6749 21959 6783
rect 21959 6749 21968 6783
rect 21916 6740 21968 6749
rect 22468 6740 22520 6792
rect 30564 6808 30616 6860
rect 31760 6808 31812 6860
rect 28908 6783 28960 6792
rect 28908 6749 28917 6783
rect 28917 6749 28951 6783
rect 28951 6749 28960 6783
rect 28908 6740 28960 6749
rect 29092 6783 29144 6792
rect 29092 6749 29101 6783
rect 29101 6749 29135 6783
rect 29135 6749 29144 6783
rect 29092 6740 29144 6749
rect 31208 6740 31260 6792
rect 31484 6783 31536 6792
rect 31484 6749 31493 6783
rect 31493 6749 31527 6783
rect 31527 6749 31536 6783
rect 31484 6740 31536 6749
rect 31668 6740 31720 6792
rect 33876 6783 33928 6792
rect 33876 6749 33885 6783
rect 33885 6749 33919 6783
rect 33919 6749 33928 6783
rect 33876 6740 33928 6749
rect 34796 6740 34848 6792
rect 22008 6715 22060 6724
rect 22008 6681 22017 6715
rect 22017 6681 22051 6715
rect 22051 6681 22060 6715
rect 22008 6672 22060 6681
rect 22560 6672 22612 6724
rect 26700 6672 26752 6724
rect 30380 6672 30432 6724
rect 18328 6604 18380 6656
rect 21824 6647 21876 6656
rect 21824 6613 21833 6647
rect 21833 6613 21867 6647
rect 21867 6613 21876 6647
rect 21824 6604 21876 6613
rect 22100 6604 22152 6656
rect 29000 6604 29052 6656
rect 29368 6604 29420 6656
rect 31392 6604 31444 6656
rect 33968 6647 34020 6656
rect 33968 6613 33977 6647
rect 33977 6613 34011 6647
rect 34011 6613 34020 6647
rect 33968 6604 34020 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 5356 6400 5408 6452
rect 1676 6375 1728 6384
rect 1676 6341 1710 6375
rect 1710 6341 1728 6375
rect 1676 6332 1728 6341
rect 4068 6264 4120 6316
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 10508 6400 10560 6452
rect 14188 6400 14240 6452
rect 7380 6264 7432 6316
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 7840 6307 7892 6316
rect 7840 6273 7849 6307
rect 7849 6273 7883 6307
rect 7883 6273 7892 6307
rect 7840 6264 7892 6273
rect 8024 6264 8076 6316
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 8484 6264 8536 6316
rect 11060 6264 11112 6316
rect 11336 6264 11388 6316
rect 14096 6332 14148 6384
rect 14464 6332 14516 6384
rect 15660 6400 15712 6452
rect 16304 6400 16356 6452
rect 19984 6400 20036 6452
rect 22008 6400 22060 6452
rect 22100 6400 22152 6452
rect 24216 6400 24268 6452
rect 28172 6400 28224 6452
rect 15568 6332 15620 6384
rect 16764 6332 16816 6384
rect 18696 6332 18748 6384
rect 14556 6264 14608 6316
rect 15384 6264 15436 6316
rect 16212 6264 16264 6316
rect 17316 6264 17368 6316
rect 6092 6171 6144 6180
rect 6092 6137 6101 6171
rect 6101 6137 6135 6171
rect 6135 6137 6144 6171
rect 6092 6128 6144 6137
rect 11796 6239 11848 6248
rect 11796 6205 11805 6239
rect 11805 6205 11839 6239
rect 11839 6205 11848 6239
rect 11796 6196 11848 6205
rect 8576 6171 8628 6180
rect 8576 6137 8585 6171
rect 8585 6137 8619 6171
rect 8619 6137 8628 6171
rect 8576 6128 8628 6137
rect 8668 6128 8720 6180
rect 7564 6060 7616 6112
rect 10232 6103 10284 6112
rect 10232 6069 10241 6103
rect 10241 6069 10275 6103
rect 10275 6069 10284 6103
rect 10232 6060 10284 6069
rect 16580 6196 16632 6248
rect 17132 6196 17184 6248
rect 18236 6264 18288 6316
rect 18880 6307 18932 6316
rect 18880 6273 18889 6307
rect 18889 6273 18923 6307
rect 18923 6273 18932 6307
rect 18880 6264 18932 6273
rect 19064 6264 19116 6316
rect 20720 6264 20772 6316
rect 18788 6239 18840 6248
rect 18788 6205 18797 6239
rect 18797 6205 18831 6239
rect 18831 6205 18840 6239
rect 18788 6196 18840 6205
rect 19248 6196 19300 6248
rect 21824 6264 21876 6316
rect 21916 6264 21968 6316
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 22560 6307 22612 6316
rect 22560 6273 22569 6307
rect 22569 6273 22603 6307
rect 22603 6273 22612 6307
rect 22560 6264 22612 6273
rect 22652 6264 22704 6316
rect 23940 6307 23992 6316
rect 23940 6273 23949 6307
rect 23949 6273 23983 6307
rect 23983 6273 23992 6307
rect 23940 6264 23992 6273
rect 25044 6264 25096 6316
rect 25688 6264 25740 6316
rect 27528 6264 27580 6316
rect 24216 6196 24268 6248
rect 28448 6264 28500 6316
rect 29092 6332 29144 6384
rect 33140 6400 33192 6452
rect 33968 6400 34020 6452
rect 28908 6264 28960 6316
rect 29460 6307 29512 6316
rect 29460 6273 29469 6307
rect 29469 6273 29503 6307
rect 29503 6273 29512 6307
rect 29460 6264 29512 6273
rect 31116 6264 31168 6316
rect 31300 6307 31352 6316
rect 31300 6273 31309 6307
rect 31309 6273 31343 6307
rect 31343 6273 31352 6307
rect 31300 6264 31352 6273
rect 31392 6307 31444 6316
rect 31392 6273 31401 6307
rect 31401 6273 31435 6307
rect 31435 6273 31444 6307
rect 31392 6264 31444 6273
rect 31576 6264 31628 6316
rect 14556 6128 14608 6180
rect 24860 6128 24912 6180
rect 26700 6128 26752 6180
rect 30840 6128 30892 6180
rect 31852 6128 31904 6180
rect 16304 6060 16356 6112
rect 18328 6060 18380 6112
rect 19340 6103 19392 6112
rect 19340 6069 19349 6103
rect 19349 6069 19383 6103
rect 19383 6069 19392 6103
rect 19340 6060 19392 6069
rect 20628 6103 20680 6112
rect 20628 6069 20637 6103
rect 20637 6069 20671 6103
rect 20671 6069 20680 6103
rect 20628 6060 20680 6069
rect 21180 6060 21232 6112
rect 23664 6060 23716 6112
rect 25872 6060 25924 6112
rect 27620 6103 27672 6112
rect 27620 6069 27629 6103
rect 27629 6069 27663 6103
rect 27663 6069 27672 6103
rect 27620 6060 27672 6069
rect 27712 6060 27764 6112
rect 29644 6060 29696 6112
rect 31024 6103 31076 6112
rect 31024 6069 31033 6103
rect 31033 6069 31067 6103
rect 31067 6069 31076 6103
rect 31024 6060 31076 6069
rect 31300 6060 31352 6112
rect 31944 6060 31996 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1308 5856 1360 5908
rect 7472 5856 7524 5908
rect 8024 5856 8076 5908
rect 1860 5788 1912 5840
rect 10876 5856 10928 5908
rect 11796 5856 11848 5908
rect 12808 5856 12860 5908
rect 12992 5856 13044 5908
rect 18512 5856 18564 5908
rect 18788 5856 18840 5908
rect 21364 5856 21416 5908
rect 8576 5720 8628 5772
rect 5816 5652 5868 5704
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 7380 5652 7432 5704
rect 7932 5652 7984 5704
rect 8668 5695 8720 5704
rect 8668 5661 8677 5695
rect 8677 5661 8711 5695
rect 8711 5661 8720 5695
rect 9220 5720 9272 5772
rect 12532 5720 12584 5772
rect 8668 5652 8720 5661
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 7748 5559 7800 5568
rect 7748 5525 7757 5559
rect 7757 5525 7791 5559
rect 7791 5525 7800 5559
rect 11060 5652 11112 5704
rect 7748 5516 7800 5525
rect 8300 5559 8352 5568
rect 8300 5525 8309 5559
rect 8309 5525 8343 5559
rect 8343 5525 8352 5559
rect 8300 5516 8352 5525
rect 9680 5516 9732 5568
rect 9864 5516 9916 5568
rect 12256 5695 12308 5704
rect 12256 5661 12265 5695
rect 12265 5661 12299 5695
rect 12299 5661 12308 5695
rect 12256 5652 12308 5661
rect 12440 5695 12492 5704
rect 12440 5661 12449 5695
rect 12449 5661 12483 5695
rect 12483 5661 12492 5695
rect 12440 5652 12492 5661
rect 14924 5695 14976 5704
rect 14924 5661 14933 5695
rect 14933 5661 14967 5695
rect 14967 5661 14976 5695
rect 14924 5652 14976 5661
rect 12624 5584 12676 5636
rect 15476 5652 15528 5704
rect 15568 5695 15620 5704
rect 20168 5788 20220 5840
rect 17224 5720 17276 5772
rect 18880 5720 18932 5772
rect 18972 5720 19024 5772
rect 15568 5661 15602 5695
rect 15602 5661 15620 5695
rect 15568 5652 15620 5661
rect 18328 5652 18380 5704
rect 19340 5652 19392 5704
rect 19708 5695 19760 5704
rect 19708 5661 19717 5695
rect 19717 5661 19751 5695
rect 19751 5661 19760 5695
rect 19708 5652 19760 5661
rect 19984 5695 20036 5704
rect 19984 5661 19993 5695
rect 19993 5661 20027 5695
rect 20027 5661 20036 5695
rect 19984 5652 20036 5661
rect 20076 5652 20128 5704
rect 20260 5695 20312 5704
rect 20260 5661 20270 5695
rect 20270 5661 20304 5695
rect 20304 5661 20312 5695
rect 20260 5652 20312 5661
rect 20628 5695 20680 5704
rect 20628 5661 20642 5695
rect 20642 5661 20676 5695
rect 20676 5661 20680 5695
rect 20628 5652 20680 5661
rect 21180 5695 21232 5704
rect 21180 5661 21189 5695
rect 21189 5661 21223 5695
rect 21223 5661 21232 5695
rect 21180 5652 21232 5661
rect 22468 5856 22520 5908
rect 22560 5856 22612 5908
rect 24216 5899 24268 5908
rect 24216 5865 24225 5899
rect 24225 5865 24259 5899
rect 24259 5865 24268 5899
rect 24216 5856 24268 5865
rect 25044 5788 25096 5840
rect 25872 5788 25924 5840
rect 26608 5763 26660 5772
rect 26608 5729 26617 5763
rect 26617 5729 26651 5763
rect 26651 5729 26660 5763
rect 26608 5720 26660 5729
rect 31300 5856 31352 5908
rect 31852 5899 31904 5908
rect 31852 5865 31861 5899
rect 31861 5865 31895 5899
rect 31895 5865 31904 5899
rect 31852 5856 31904 5865
rect 33600 5899 33652 5908
rect 33600 5865 33609 5899
rect 33609 5865 33643 5899
rect 33643 5865 33652 5899
rect 33600 5856 33652 5865
rect 21548 5695 21600 5704
rect 21548 5661 21557 5695
rect 21557 5661 21591 5695
rect 21591 5661 21600 5695
rect 21548 5652 21600 5661
rect 21824 5695 21876 5704
rect 21824 5661 21833 5695
rect 21833 5661 21867 5695
rect 21867 5661 21876 5695
rect 21824 5652 21876 5661
rect 15384 5559 15436 5568
rect 15384 5525 15393 5559
rect 15393 5525 15427 5559
rect 15427 5525 15436 5559
rect 15384 5516 15436 5525
rect 15660 5516 15712 5568
rect 16212 5584 16264 5636
rect 17132 5627 17184 5636
rect 17132 5593 17141 5627
rect 17141 5593 17175 5627
rect 17175 5593 17184 5627
rect 17132 5584 17184 5593
rect 17408 5584 17460 5636
rect 18420 5584 18472 5636
rect 19064 5584 19116 5636
rect 16764 5516 16816 5568
rect 20904 5584 20956 5636
rect 21732 5584 21784 5636
rect 22192 5695 22244 5704
rect 22192 5661 22199 5695
rect 22199 5661 22233 5695
rect 22233 5661 22244 5695
rect 22192 5652 22244 5661
rect 22008 5584 22060 5636
rect 22284 5584 22336 5636
rect 22836 5584 22888 5636
rect 23664 5652 23716 5704
rect 23848 5652 23900 5704
rect 24860 5652 24912 5704
rect 25872 5695 25924 5704
rect 25872 5661 25881 5695
rect 25881 5661 25915 5695
rect 25915 5661 25924 5695
rect 25872 5652 25924 5661
rect 25964 5695 26016 5704
rect 25964 5661 25973 5695
rect 25973 5661 26007 5695
rect 26007 5661 26016 5695
rect 25964 5652 26016 5661
rect 27528 5720 27580 5772
rect 27252 5652 27304 5704
rect 27712 5652 27764 5704
rect 31024 5720 31076 5772
rect 31668 5788 31720 5840
rect 31760 5788 31812 5840
rect 26700 5627 26752 5636
rect 26700 5593 26709 5627
rect 26709 5593 26743 5627
rect 26743 5593 26752 5627
rect 26700 5584 26752 5593
rect 22192 5516 22244 5568
rect 27436 5584 27488 5636
rect 28540 5652 28592 5704
rect 29460 5652 29512 5704
rect 29644 5652 29696 5704
rect 34704 5720 34756 5772
rect 31944 5652 31996 5704
rect 32220 5695 32272 5704
rect 32220 5661 32229 5695
rect 32229 5661 32263 5695
rect 32263 5661 32272 5695
rect 32220 5652 32272 5661
rect 32312 5652 32364 5704
rect 31852 5627 31904 5636
rect 31852 5593 31861 5627
rect 31861 5593 31895 5627
rect 31895 5593 31904 5627
rect 31852 5584 31904 5593
rect 27804 5559 27856 5568
rect 27804 5525 27813 5559
rect 27813 5525 27847 5559
rect 27847 5525 27856 5559
rect 27804 5516 27856 5525
rect 30656 5516 30708 5568
rect 31116 5559 31168 5568
rect 31116 5525 31125 5559
rect 31125 5525 31159 5559
rect 31159 5525 31168 5559
rect 31116 5516 31168 5525
rect 31208 5516 31260 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 8668 5312 8720 5364
rect 9864 5312 9916 5364
rect 9956 5312 10008 5364
rect 12440 5312 12492 5364
rect 12624 5312 12676 5364
rect 15384 5312 15436 5364
rect 14924 5244 14976 5296
rect 15660 5244 15712 5296
rect 7656 5176 7708 5228
rect 7748 5219 7800 5228
rect 7748 5185 7757 5219
rect 7757 5185 7791 5219
rect 7791 5185 7800 5219
rect 7748 5176 7800 5185
rect 8300 5176 8352 5228
rect 9680 5176 9732 5228
rect 11060 5176 11112 5228
rect 12532 5176 12584 5228
rect 17316 5312 17368 5364
rect 19892 5312 19944 5364
rect 19708 5244 19760 5296
rect 20260 5312 20312 5364
rect 21824 5312 21876 5364
rect 22100 5312 22152 5364
rect 23940 5312 23992 5364
rect 25964 5312 26016 5364
rect 27436 5355 27488 5364
rect 27436 5321 27445 5355
rect 27445 5321 27479 5355
rect 27479 5321 27488 5355
rect 27436 5312 27488 5321
rect 31484 5312 31536 5364
rect 31944 5312 31996 5364
rect 13084 5108 13136 5160
rect 15016 5151 15068 5160
rect 15016 5117 15025 5151
rect 15025 5117 15059 5151
rect 15059 5117 15068 5151
rect 15016 5108 15068 5117
rect 15476 5151 15528 5160
rect 15476 5117 15485 5151
rect 15485 5117 15519 5151
rect 15519 5117 15528 5151
rect 15476 5108 15528 5117
rect 16212 5219 16264 5228
rect 16212 5185 16221 5219
rect 16221 5185 16255 5219
rect 16255 5185 16264 5219
rect 16212 5176 16264 5185
rect 16304 5219 16356 5228
rect 16304 5185 16313 5219
rect 16313 5185 16347 5219
rect 16347 5185 16356 5219
rect 16304 5176 16356 5185
rect 16764 5219 16816 5228
rect 16764 5185 16773 5219
rect 16773 5185 16807 5219
rect 16807 5185 16816 5219
rect 16764 5176 16816 5185
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 17224 5219 17276 5228
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 17408 5219 17460 5228
rect 17408 5185 17417 5219
rect 17417 5185 17451 5219
rect 17451 5185 17460 5219
rect 17408 5176 17460 5185
rect 17500 5176 17552 5228
rect 18604 5176 18656 5228
rect 20168 5287 20220 5296
rect 20168 5253 20177 5287
rect 20177 5253 20211 5287
rect 20211 5253 20220 5287
rect 20168 5244 20220 5253
rect 7380 5040 7432 5092
rect 12256 5040 12308 5092
rect 19984 5176 20036 5228
rect 20628 5244 20680 5296
rect 24216 5244 24268 5296
rect 27252 5287 27304 5296
rect 27252 5253 27261 5287
rect 27261 5253 27295 5287
rect 27295 5253 27304 5287
rect 27252 5244 27304 5253
rect 30196 5244 30248 5296
rect 31300 5244 31352 5296
rect 36544 5312 36596 5364
rect 20444 5176 20496 5228
rect 21548 5176 21600 5228
rect 24860 5176 24912 5228
rect 27804 5176 27856 5228
rect 30656 5176 30708 5228
rect 32220 5176 32272 5228
rect 32772 5219 32824 5228
rect 32772 5185 32781 5219
rect 32781 5185 32815 5219
rect 32815 5185 32824 5219
rect 32772 5176 32824 5185
rect 20076 5040 20128 5092
rect 22008 5108 22060 5160
rect 22652 5151 22704 5160
rect 22652 5117 22661 5151
rect 22661 5117 22695 5151
rect 22695 5117 22704 5151
rect 22652 5108 22704 5117
rect 23940 5151 23992 5160
rect 23940 5117 23949 5151
rect 23949 5117 23983 5151
rect 23983 5117 23992 5151
rect 23940 5108 23992 5117
rect 24124 5151 24176 5160
rect 24124 5117 24133 5151
rect 24133 5117 24167 5151
rect 24167 5117 24176 5151
rect 24124 5108 24176 5117
rect 21088 5040 21140 5092
rect 31116 5108 31168 5160
rect 36176 5219 36228 5228
rect 36176 5185 36185 5219
rect 36185 5185 36219 5219
rect 36219 5185 36228 5219
rect 36176 5176 36228 5185
rect 25688 5040 25740 5092
rect 10232 4972 10284 5024
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 20444 4972 20496 5024
rect 26240 4972 26292 5024
rect 31300 4972 31352 5024
rect 36360 5015 36412 5024
rect 36360 4981 36369 5015
rect 36369 4981 36403 5015
rect 36403 4981 36412 5015
rect 36360 4972 36412 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 10140 4768 10192 4820
rect 18328 4768 18380 4820
rect 25044 4768 25096 4820
rect 27620 4768 27672 4820
rect 16764 4632 16816 4684
rect 25688 4700 25740 4752
rect 16948 4607 17000 4616
rect 16948 4573 16957 4607
rect 16957 4573 16991 4607
rect 16991 4573 17000 4607
rect 16948 4564 17000 4573
rect 21364 4564 21416 4616
rect 22008 4564 22060 4616
rect 26700 4632 26752 4684
rect 25228 4564 25280 4616
rect 23848 4496 23900 4548
rect 25688 4607 25740 4616
rect 25688 4573 25697 4607
rect 25697 4573 25731 4607
rect 25731 4573 25740 4607
rect 25688 4564 25740 4573
rect 27252 4564 27304 4616
rect 28264 4700 28316 4752
rect 27804 4632 27856 4684
rect 28356 4632 28408 4684
rect 15016 4428 15068 4480
rect 25044 4428 25096 4480
rect 27436 4496 27488 4548
rect 27896 4539 27948 4548
rect 27896 4505 27905 4539
rect 27905 4505 27939 4539
rect 27939 4505 27948 4539
rect 27896 4496 27948 4505
rect 26516 4428 26568 4480
rect 28172 4564 28224 4616
rect 28264 4607 28316 4616
rect 28264 4573 28273 4607
rect 28273 4573 28307 4607
rect 28307 4573 28316 4607
rect 28264 4564 28316 4573
rect 28448 4564 28500 4616
rect 31116 4700 31168 4752
rect 31668 4700 31720 4752
rect 31300 4564 31352 4616
rect 29000 4539 29052 4548
rect 29000 4505 29009 4539
rect 29009 4505 29043 4539
rect 29043 4505 29052 4539
rect 29000 4496 29052 4505
rect 29736 4428 29788 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 19432 4224 19484 4276
rect 19984 4267 20036 4276
rect 19984 4233 19993 4267
rect 19993 4233 20027 4267
rect 20027 4233 20036 4267
rect 19984 4224 20036 4233
rect 21364 4224 21416 4276
rect 22928 4224 22980 4276
rect 5908 4088 5960 4140
rect 9128 4088 9180 4140
rect 4068 4020 4120 4072
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 18604 4131 18656 4140
rect 18604 4097 18613 4131
rect 18613 4097 18647 4131
rect 18647 4097 18656 4131
rect 18604 4088 18656 4097
rect 21824 4088 21876 4140
rect 23480 4156 23532 4208
rect 27896 4156 27948 4208
rect 28448 4156 28500 4208
rect 23940 4088 23992 4140
rect 25044 4131 25096 4140
rect 25044 4097 25053 4131
rect 25053 4097 25087 4131
rect 25087 4097 25096 4131
rect 25044 4088 25096 4097
rect 25228 4131 25280 4140
rect 25228 4097 25237 4131
rect 25237 4097 25271 4131
rect 25271 4097 25280 4131
rect 25228 4088 25280 4097
rect 25688 4088 25740 4140
rect 26240 4131 26292 4140
rect 26240 4097 26249 4131
rect 26249 4097 26283 4131
rect 26283 4097 26292 4131
rect 26240 4088 26292 4097
rect 18696 4063 18748 4072
rect 18696 4029 18705 4063
rect 18705 4029 18739 4063
rect 18739 4029 18748 4063
rect 18696 4020 18748 4029
rect 19340 4020 19392 4072
rect 22468 4020 22520 4072
rect 26516 4131 26568 4140
rect 26516 4097 26525 4131
rect 26525 4097 26559 4131
rect 26559 4097 26568 4131
rect 26516 4088 26568 4097
rect 26700 4131 26752 4140
rect 26700 4097 26709 4131
rect 26709 4097 26743 4131
rect 26743 4097 26752 4131
rect 26700 4088 26752 4097
rect 30288 4131 30340 4140
rect 30288 4097 30297 4131
rect 30297 4097 30331 4131
rect 30331 4097 30340 4131
rect 30288 4088 30340 4097
rect 30564 4156 30616 4208
rect 31116 4156 31168 4208
rect 26608 4063 26660 4072
rect 26608 4029 26617 4063
rect 26617 4029 26651 4063
rect 26651 4029 26660 4063
rect 26608 4020 26660 4029
rect 30932 4088 30984 4140
rect 27988 3952 28040 4004
rect 30380 3952 30432 4004
rect 31208 4020 31260 4072
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 19616 3927 19668 3936
rect 19616 3893 19625 3927
rect 19625 3893 19659 3927
rect 19659 3893 19668 3927
rect 19616 3884 19668 3893
rect 21548 3884 21600 3936
rect 22836 3884 22888 3936
rect 26148 3884 26200 3936
rect 30748 3884 30800 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 18696 3680 18748 3732
rect 19248 3587 19300 3596
rect 16580 3476 16632 3528
rect 17592 3476 17644 3528
rect 16212 3408 16264 3460
rect 17132 3383 17184 3392
rect 17132 3349 17141 3383
rect 17141 3349 17175 3383
rect 17175 3349 17184 3383
rect 17132 3340 17184 3349
rect 17500 3383 17552 3392
rect 17500 3349 17509 3383
rect 17509 3349 17543 3383
rect 17543 3349 17552 3383
rect 17500 3340 17552 3349
rect 18052 3519 18104 3528
rect 18052 3485 18061 3519
rect 18061 3485 18095 3519
rect 18095 3485 18104 3519
rect 18052 3476 18104 3485
rect 19248 3553 19257 3587
rect 19257 3553 19291 3587
rect 19291 3553 19300 3587
rect 19248 3544 19300 3553
rect 22008 3680 22060 3732
rect 23480 3723 23532 3732
rect 23480 3689 23489 3723
rect 23489 3689 23523 3723
rect 23523 3689 23532 3723
rect 23480 3680 23532 3689
rect 24492 3680 24544 3732
rect 20904 3587 20956 3596
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 21088 3587 21140 3596
rect 21088 3553 21097 3587
rect 21097 3553 21131 3587
rect 21131 3553 21140 3587
rect 21088 3544 21140 3553
rect 22100 3544 22152 3596
rect 19432 3476 19484 3528
rect 19984 3476 20036 3528
rect 20536 3476 20588 3528
rect 21548 3519 21600 3528
rect 21548 3485 21557 3519
rect 21557 3485 21591 3519
rect 21591 3485 21600 3519
rect 21548 3476 21600 3485
rect 22652 3476 22704 3528
rect 25688 3476 25740 3528
rect 25964 3519 26016 3528
rect 25964 3485 25973 3519
rect 25973 3485 26007 3519
rect 26007 3485 26016 3519
rect 25964 3476 26016 3485
rect 18328 3408 18380 3460
rect 30288 3680 30340 3732
rect 30380 3680 30432 3732
rect 31300 3680 31352 3732
rect 31852 3680 31904 3732
rect 36084 3680 36136 3732
rect 26148 3587 26200 3596
rect 26148 3553 26157 3587
rect 26157 3553 26191 3587
rect 26191 3553 26200 3587
rect 26148 3544 26200 3553
rect 26240 3544 26292 3596
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 26608 3476 26660 3528
rect 27528 3544 27580 3596
rect 27068 3519 27120 3528
rect 27068 3485 27077 3519
rect 27077 3485 27111 3519
rect 27111 3485 27120 3519
rect 27068 3476 27120 3485
rect 32220 3612 32272 3664
rect 30472 3544 30524 3596
rect 30748 3544 30800 3596
rect 31668 3544 31720 3596
rect 29828 3476 29880 3528
rect 30196 3519 30248 3528
rect 30196 3485 30205 3519
rect 30205 3485 30239 3519
rect 30239 3485 30248 3519
rect 30196 3476 30248 3485
rect 30840 3519 30892 3528
rect 30840 3485 30849 3519
rect 30849 3485 30883 3519
rect 30883 3485 30892 3519
rect 30840 3476 30892 3485
rect 30932 3519 30984 3528
rect 30932 3485 30941 3519
rect 30941 3485 30975 3519
rect 30975 3485 30984 3519
rect 30932 3476 30984 3485
rect 31300 3519 31352 3528
rect 31300 3485 31309 3519
rect 31309 3485 31343 3519
rect 31343 3485 31352 3519
rect 31300 3476 31352 3485
rect 31392 3519 31444 3528
rect 31392 3485 31401 3519
rect 31401 3485 31435 3519
rect 31435 3485 31444 3519
rect 31392 3476 31444 3485
rect 31484 3519 31536 3528
rect 31484 3485 31493 3519
rect 31493 3485 31527 3519
rect 31527 3485 31536 3519
rect 31484 3476 31536 3485
rect 31852 3519 31904 3528
rect 31852 3485 31861 3519
rect 31861 3485 31895 3519
rect 31895 3485 31904 3519
rect 31852 3476 31904 3485
rect 32404 3519 32456 3528
rect 32404 3485 32413 3519
rect 32413 3485 32447 3519
rect 32447 3485 32456 3519
rect 32404 3476 32456 3485
rect 29000 3408 29052 3460
rect 32772 3519 32824 3528
rect 32772 3485 32781 3519
rect 32781 3485 32815 3519
rect 32815 3485 32824 3519
rect 32772 3476 32824 3485
rect 18236 3340 18288 3392
rect 18604 3340 18656 3392
rect 20076 3340 20128 3392
rect 20812 3383 20864 3392
rect 20812 3349 20821 3383
rect 20821 3349 20855 3383
rect 20855 3349 20864 3383
rect 20812 3340 20864 3349
rect 20904 3340 20956 3392
rect 23388 3340 23440 3392
rect 25136 3340 25188 3392
rect 29552 3383 29604 3392
rect 29552 3349 29561 3383
rect 29561 3349 29595 3383
rect 29595 3349 29604 3383
rect 29552 3340 29604 3349
rect 29736 3383 29788 3392
rect 29736 3349 29745 3383
rect 29745 3349 29779 3383
rect 29779 3349 29788 3383
rect 29736 3340 29788 3349
rect 31576 3408 31628 3460
rect 32220 3408 32272 3460
rect 30656 3383 30708 3392
rect 30656 3349 30665 3383
rect 30665 3349 30699 3383
rect 30699 3349 30708 3383
rect 30656 3340 30708 3349
rect 31116 3383 31168 3392
rect 31116 3349 31125 3383
rect 31125 3349 31159 3383
rect 31159 3349 31168 3383
rect 31116 3340 31168 3349
rect 31208 3383 31260 3392
rect 31208 3349 31217 3383
rect 31217 3349 31251 3383
rect 31251 3349 31260 3383
rect 31208 3340 31260 3349
rect 31300 3340 31352 3392
rect 31760 3340 31812 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 16212 3179 16264 3188
rect 16212 3145 16221 3179
rect 16221 3145 16255 3179
rect 16255 3145 16264 3179
rect 16212 3136 16264 3145
rect 18604 3136 18656 3188
rect 18696 3136 18748 3188
rect 19432 3179 19484 3188
rect 19432 3145 19441 3179
rect 19441 3145 19475 3179
rect 19475 3145 19484 3179
rect 19432 3136 19484 3145
rect 16028 3068 16080 3120
rect 17132 3111 17184 3120
rect 17132 3077 17141 3111
rect 17141 3077 17175 3111
rect 17175 3077 17184 3111
rect 17132 3068 17184 3077
rect 940 3000 992 3052
rect 4068 3000 4120 3052
rect 4252 2907 4304 2916
rect 4252 2873 4261 2907
rect 4261 2873 4295 2907
rect 4295 2873 4304 2907
rect 4252 2864 4304 2873
rect 17776 3068 17828 3120
rect 20812 3136 20864 3188
rect 21824 3179 21876 3188
rect 21824 3145 21833 3179
rect 21833 3145 21867 3179
rect 21867 3145 21876 3179
rect 21824 3136 21876 3145
rect 22008 3136 22060 3188
rect 22652 3179 22704 3188
rect 22652 3145 22661 3179
rect 22661 3145 22695 3179
rect 22695 3145 22704 3179
rect 22652 3136 22704 3145
rect 25044 3136 25096 3188
rect 17592 3043 17644 3052
rect 17592 3009 17601 3043
rect 17601 3009 17635 3043
rect 17635 3009 17644 3043
rect 17592 3000 17644 3009
rect 18144 3000 18196 3052
rect 19616 3043 19668 3052
rect 19616 3009 19625 3043
rect 19625 3009 19659 3043
rect 19659 3009 19668 3043
rect 19616 3000 19668 3009
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 19340 2932 19392 2984
rect 20352 3000 20404 3052
rect 23388 3068 23440 3120
rect 25688 3179 25740 3188
rect 25688 3145 25697 3179
rect 25697 3145 25731 3179
rect 25731 3145 25740 3179
rect 25688 3136 25740 3145
rect 26148 3136 26200 3188
rect 27068 3136 27120 3188
rect 27528 3179 27580 3188
rect 27528 3145 27537 3179
rect 27537 3145 27571 3179
rect 27571 3145 27580 3179
rect 27528 3136 27580 3145
rect 21088 2932 21140 2984
rect 22836 3043 22888 3052
rect 22836 3009 22845 3043
rect 22845 3009 22879 3043
rect 22879 3009 22888 3043
rect 22836 3000 22888 3009
rect 23940 3043 23992 3052
rect 23940 3009 23949 3043
rect 23949 3009 23983 3043
rect 23983 3009 23992 3043
rect 23940 3000 23992 3009
rect 26056 3000 26108 3052
rect 24308 2975 24360 2984
rect 24308 2941 24317 2975
rect 24317 2941 24351 2975
rect 24351 2941 24360 2975
rect 24308 2932 24360 2941
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 22928 2864 22980 2916
rect 25320 2864 25372 2916
rect 26240 3000 26292 3052
rect 30472 3136 30524 3188
rect 30564 3179 30616 3188
rect 30564 3145 30573 3179
rect 30573 3145 30607 3179
rect 30607 3145 30616 3179
rect 30564 3136 30616 3145
rect 30656 3136 30708 3188
rect 31576 3179 31628 3188
rect 31576 3145 31585 3179
rect 31585 3145 31619 3179
rect 31619 3145 31628 3179
rect 31576 3136 31628 3145
rect 34152 3179 34204 3188
rect 34152 3145 34161 3179
rect 34161 3145 34195 3179
rect 34195 3145 34204 3179
rect 34152 3136 34204 3145
rect 29552 3068 29604 3120
rect 28540 3043 28592 3052
rect 28540 3009 28549 3043
rect 28549 3009 28583 3043
rect 28583 3009 28592 3043
rect 28540 3000 28592 3009
rect 30380 3043 30432 3052
rect 30380 3009 30389 3043
rect 30389 3009 30423 3043
rect 30423 3009 30432 3043
rect 30380 3000 30432 3009
rect 31484 3068 31536 3120
rect 32404 3068 32456 3120
rect 30932 3000 30984 3052
rect 31392 3000 31444 3052
rect 31668 3043 31720 3052
rect 31668 3009 31677 3043
rect 31677 3009 31711 3043
rect 31711 3009 31720 3043
rect 31668 3000 31720 3009
rect 32772 3043 32824 3052
rect 32772 3009 32781 3043
rect 32781 3009 32815 3043
rect 32815 3009 32824 3043
rect 32772 3000 32824 3009
rect 33048 3043 33100 3052
rect 33048 3009 33082 3043
rect 33082 3009 33100 3043
rect 33048 3000 33100 3009
rect 24308 2796 24360 2848
rect 30196 2796 30248 2848
rect 30288 2796 30340 2848
rect 35440 2864 35492 2916
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 5908 2635 5960 2644
rect 5908 2601 5917 2635
rect 5917 2601 5951 2635
rect 5951 2601 5960 2635
rect 5908 2592 5960 2601
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 19524 2592 19576 2644
rect 25964 2592 26016 2644
rect 33048 2592 33100 2644
rect 29920 2524 29972 2576
rect 30472 2524 30524 2576
rect 31208 2524 31260 2576
rect 5816 2388 5868 2440
rect 9036 2388 9088 2440
rect 24308 2456 24360 2508
rect 25964 2499 26016 2508
rect 25964 2465 25973 2499
rect 25973 2465 26007 2499
rect 26007 2465 26016 2499
rect 25964 2456 26016 2465
rect 26148 2499 26200 2508
rect 26148 2465 26157 2499
rect 26157 2465 26191 2499
rect 26191 2465 26200 2499
rect 26148 2456 26200 2465
rect 36084 2456 36136 2508
rect 16028 2388 16080 2440
rect 18052 2388 18104 2440
rect 21272 2388 21324 2440
rect 23848 2388 23900 2440
rect 25320 2388 25372 2440
rect 26240 2388 26292 2440
rect 27068 2388 27120 2440
rect 29644 2388 29696 2440
rect 32864 2388 32916 2440
rect 35900 2431 35952 2440
rect 35900 2397 35909 2431
rect 35909 2397 35943 2431
rect 35943 2397 35952 2431
rect 35900 2388 35952 2397
rect 20 2320 72 2372
rect 19156 2320 19208 2372
rect 2228 2295 2280 2304
rect 2228 2261 2237 2295
rect 2237 2261 2271 2295
rect 2271 2261 2280 2295
rect 2228 2252 2280 2261
rect 2596 2295 2648 2304
rect 2596 2261 2605 2295
rect 2605 2261 2639 2295
rect 2639 2261 2648 2295
rect 2596 2252 2648 2261
rect 11612 2252 11664 2304
rect 14832 2252 14884 2304
rect 23848 2252 23900 2304
rect 30196 2363 30248 2372
rect 30196 2329 30205 2363
rect 30205 2329 30239 2363
rect 30239 2329 30248 2363
rect 30196 2320 30248 2329
rect 30380 2252 30432 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 2228 1980 2280 2032
rect 30748 1980 30800 2032
<< metal2 >>
rect 1306 39280 1362 40080
rect 4526 39386 4582 40080
rect 7102 39386 7158 40080
rect 10322 39386 10378 40080
rect 4526 39358 4660 39386
rect 4526 39280 4582 39358
rect 938 38176 994 38185
rect 938 38111 994 38120
rect 952 37466 980 38111
rect 940 37460 992 37466
rect 940 37402 992 37408
rect 1320 37194 1348 39280
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37330 4660 39358
rect 7102 39358 7420 39386
rect 7102 39280 7158 39358
rect 4620 37324 4672 37330
rect 4620 37266 4672 37272
rect 5448 37256 5500 37262
rect 5448 37198 5500 37204
rect 6828 37256 6880 37262
rect 6828 37198 6880 37204
rect 1308 37188 1360 37194
rect 1308 37130 1360 37136
rect 2320 37120 2372 37126
rect 2320 37062 2372 37068
rect 2136 35080 2188 35086
rect 2136 35022 2188 35028
rect 940 34944 992 34950
rect 940 34886 992 34892
rect 952 34785 980 34886
rect 938 34776 994 34785
rect 938 34711 994 34720
rect 1952 32836 2004 32842
rect 1952 32778 2004 32784
rect 1964 32570 1992 32778
rect 1952 32564 2004 32570
rect 1952 32506 2004 32512
rect 1492 32428 1544 32434
rect 1492 32370 1544 32376
rect 940 32224 992 32230
rect 940 32166 992 32172
rect 952 32065 980 32166
rect 938 32056 994 32065
rect 938 31991 994 32000
rect 1504 26234 1532 32370
rect 1768 31408 1820 31414
rect 1768 31350 1820 31356
rect 1780 29170 1808 31350
rect 1860 31340 1912 31346
rect 1860 31282 1912 31288
rect 1872 30938 1900 31282
rect 1860 30932 1912 30938
rect 1860 30874 1912 30880
rect 1584 29164 1636 29170
rect 1584 29106 1636 29112
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 2044 29164 2096 29170
rect 2044 29106 2096 29112
rect 1596 28665 1624 29106
rect 1676 29028 1728 29034
rect 1676 28970 1728 28976
rect 1582 28656 1638 28665
rect 1582 28591 1638 28600
rect 1504 26206 1624 26234
rect 1398 25256 1454 25265
rect 1398 25191 1454 25200
rect 1412 24818 1440 25191
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 938 22536 994 22545
rect 938 22471 940 22480
rect 992 22471 994 22480
rect 940 22442 992 22448
rect 1492 22024 1544 22030
rect 1492 21966 1544 21972
rect 1504 20466 1532 21966
rect 1492 20460 1544 20466
rect 1492 20402 1544 20408
rect 1596 19922 1624 26206
rect 1584 19916 1636 19922
rect 1584 19858 1636 19864
rect 940 19168 992 19174
rect 938 19136 940 19145
rect 992 19136 994 19145
rect 938 19071 994 19080
rect 1492 18760 1544 18766
rect 1492 18702 1544 18708
rect 1504 17678 1532 18702
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 940 15904 992 15910
rect 940 15846 992 15852
rect 952 15745 980 15846
rect 938 15736 994 15745
rect 938 15671 994 15680
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12345 1624 12582
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1492 9988 1544 9994
rect 1492 9930 1544 9936
rect 1504 8294 1532 9930
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1596 9625 1624 9862
rect 1582 9616 1638 9625
rect 1582 9551 1638 9560
rect 1492 8288 1544 8294
rect 1492 8230 1544 8236
rect 1688 6390 1716 28970
rect 2056 28762 2084 29106
rect 2044 28756 2096 28762
rect 2044 28698 2096 28704
rect 1768 27396 1820 27402
rect 1768 27338 1820 27344
rect 1780 27130 1808 27338
rect 1768 27124 1820 27130
rect 1768 27066 1820 27072
rect 2148 26234 2176 35022
rect 2056 26206 2176 26234
rect 1768 25696 1820 25702
rect 1768 25638 1820 25644
rect 1780 25294 1808 25638
rect 1768 25288 1820 25294
rect 1768 25230 1820 25236
rect 1860 24744 1912 24750
rect 1860 24686 1912 24692
rect 1768 24132 1820 24138
rect 1768 24074 1820 24080
rect 1780 23866 1808 24074
rect 1768 23860 1820 23866
rect 1768 23802 1820 23808
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1780 20058 1808 20402
rect 1768 20052 1820 20058
rect 1768 19994 1820 20000
rect 1872 19938 1900 24686
rect 1952 21956 2004 21962
rect 1952 21898 2004 21904
rect 1964 21690 1992 21898
rect 1952 21684 2004 21690
rect 1952 21626 2004 21632
rect 2056 21570 2084 26206
rect 1780 19910 1900 19938
rect 1964 21542 2084 21570
rect 1780 12209 1808 19910
rect 1860 17604 1912 17610
rect 1860 17546 1912 17552
rect 1872 17338 1900 17546
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1766 12200 1822 12209
rect 1766 12135 1822 12144
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 1306 6216 1362 6225
rect 1306 6151 1362 6160
rect 1320 5914 1348 6151
rect 1308 5908 1360 5914
rect 1308 5850 1360 5856
rect 1872 5846 1900 16050
rect 1964 6730 1992 21542
rect 2044 20800 2096 20806
rect 2044 20742 2096 20748
rect 2056 19854 2084 20742
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2148 18766 2176 19110
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 2056 17202 2084 18022
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2332 13734 2360 37062
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 3792 36168 3844 36174
rect 3792 36110 3844 36116
rect 3804 34542 3832 36110
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4620 34604 4672 34610
rect 4620 34546 4672 34552
rect 3792 34536 3844 34542
rect 3792 34478 3844 34484
rect 3804 34066 3832 34478
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4632 34202 4660 34546
rect 4712 34400 4764 34406
rect 4712 34342 4764 34348
rect 4620 34196 4672 34202
rect 4620 34138 4672 34144
rect 3792 34060 3844 34066
rect 3792 34002 3844 34008
rect 2688 33108 2740 33114
rect 2688 33050 2740 33056
rect 2700 32570 2728 33050
rect 3804 32978 3832 34002
rect 4724 33998 4752 34342
rect 4712 33992 4764 33998
rect 4712 33934 4764 33940
rect 5264 33924 5316 33930
rect 5264 33866 5316 33872
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 5276 33658 5304 33866
rect 5356 33856 5408 33862
rect 5356 33798 5408 33804
rect 5264 33652 5316 33658
rect 5264 33594 5316 33600
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 3792 32972 3844 32978
rect 3792 32914 3844 32920
rect 3608 32904 3660 32910
rect 3608 32846 3660 32852
rect 3620 32570 3648 32846
rect 4252 32768 4304 32774
rect 4252 32710 4304 32716
rect 4264 32570 4292 32710
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 2688 32564 2740 32570
rect 2688 32506 2740 32512
rect 3608 32564 3660 32570
rect 3608 32506 3660 32512
rect 4252 32564 4304 32570
rect 4252 32506 4304 32512
rect 3332 32496 3384 32502
rect 3332 32438 3384 32444
rect 2596 32428 2648 32434
rect 2596 32370 2648 32376
rect 2608 30802 2636 32370
rect 3344 31754 3372 32438
rect 4620 32224 4672 32230
rect 4620 32166 4672 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4632 31890 4660 32166
rect 4620 31884 4672 31890
rect 4620 31826 4672 31832
rect 5368 31822 5396 33798
rect 5356 31816 5408 31822
rect 5356 31758 5408 31764
rect 2780 31748 2832 31754
rect 2780 31690 2832 31696
rect 3252 31726 3372 31754
rect 2688 31136 2740 31142
rect 2688 31078 2740 31084
rect 2596 30796 2648 30802
rect 2596 30738 2648 30744
rect 2700 30734 2728 31078
rect 2792 30734 2820 31690
rect 2688 30728 2740 30734
rect 2688 30670 2740 30676
rect 2780 30728 2832 30734
rect 2780 30670 2832 30676
rect 2792 28994 2820 30670
rect 2792 28966 2912 28994
rect 2884 28422 2912 28966
rect 3148 28960 3200 28966
rect 3148 28902 3200 28908
rect 3160 28490 3188 28902
rect 3148 28484 3200 28490
rect 3148 28426 3200 28432
rect 2872 28416 2924 28422
rect 2872 28358 2924 28364
rect 2884 27418 2912 28358
rect 3056 28008 3108 28014
rect 3056 27950 3108 27956
rect 3068 27470 3096 27950
rect 3252 27470 3280 31726
rect 3424 31680 3476 31686
rect 3424 31622 3476 31628
rect 3436 31346 3464 31622
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 3424 31340 3476 31346
rect 3424 31282 3476 31288
rect 3516 31272 3568 31278
rect 3516 31214 3568 31220
rect 3528 30258 3556 31214
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 5368 30802 5396 31758
rect 5356 30796 5408 30802
rect 5356 30738 5408 30744
rect 5264 30660 5316 30666
rect 5264 30602 5316 30608
rect 4804 30592 4856 30598
rect 4804 30534 4856 30540
rect 4816 30326 4844 30534
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4804 30320 4856 30326
rect 4804 30262 4856 30268
rect 3516 30252 3568 30258
rect 3516 30194 3568 30200
rect 3528 29714 3556 30194
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 5276 29850 5304 30602
rect 5356 30048 5408 30054
rect 5356 29990 5408 29996
rect 5264 29844 5316 29850
rect 5264 29786 5316 29792
rect 3516 29708 3568 29714
rect 3516 29650 3568 29656
rect 5368 29646 5396 29990
rect 3608 29640 3660 29646
rect 3608 29582 3660 29588
rect 5356 29640 5408 29646
rect 5356 29582 5408 29588
rect 3620 29306 3648 29582
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 3608 29300 3660 29306
rect 3608 29242 3660 29248
rect 4712 29300 4764 29306
rect 4712 29242 4764 29248
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 3516 28620 3568 28626
rect 3516 28562 3568 28568
rect 3528 27538 3556 28562
rect 3884 28076 3936 28082
rect 3884 28018 3936 28024
rect 3896 27674 3924 28018
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3884 27668 3936 27674
rect 3884 27610 3936 27616
rect 3516 27532 3568 27538
rect 3516 27474 3568 27480
rect 2792 27390 2912 27418
rect 3056 27464 3108 27470
rect 3056 27406 3108 27412
rect 3240 27464 3292 27470
rect 3240 27406 3292 27412
rect 2792 25974 2820 27390
rect 2872 27328 2924 27334
rect 2872 27270 2924 27276
rect 2884 26994 2912 27270
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 2964 26988 3016 26994
rect 2964 26930 3016 26936
rect 2976 26586 3004 26930
rect 3068 26926 3096 27406
rect 3056 26920 3108 26926
rect 3056 26862 3108 26868
rect 2964 26580 3016 26586
rect 2964 26522 3016 26528
rect 2780 25968 2832 25974
rect 2780 25910 2832 25916
rect 2504 24336 2556 24342
rect 2504 24278 2556 24284
rect 2516 23866 2544 24278
rect 2504 23860 2556 23866
rect 2504 23802 2556 23808
rect 2792 23712 2820 25910
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 2884 25498 2912 25842
rect 2872 25492 2924 25498
rect 2872 25434 2924 25440
rect 3068 25378 3096 26862
rect 3148 25832 3200 25838
rect 3148 25774 3200 25780
rect 2884 25350 3096 25378
rect 2884 25226 2912 25350
rect 2872 25220 2924 25226
rect 2872 25162 2924 25168
rect 2884 24750 2912 25162
rect 2872 24744 2924 24750
rect 2872 24686 2924 24692
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 2976 23730 3004 24142
rect 3160 23798 3188 25774
rect 3148 23792 3200 23798
rect 3148 23734 3200 23740
rect 2872 23724 2924 23730
rect 2792 23684 2872 23712
rect 2872 23666 2924 23672
rect 2964 23724 3016 23730
rect 2964 23666 3016 23672
rect 2688 23656 2740 23662
rect 2688 23598 2740 23604
rect 2700 21146 2728 23598
rect 2780 21684 2832 21690
rect 2780 21626 2832 21632
rect 2688 21140 2740 21146
rect 2688 21082 2740 21088
rect 2792 20874 2820 21626
rect 2688 20868 2740 20874
rect 2688 20810 2740 20816
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2700 19174 2728 20810
rect 2884 20210 2912 23666
rect 2976 22642 3004 23666
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 2976 22166 3004 22578
rect 2964 22160 3016 22166
rect 2964 22102 3016 22108
rect 2964 21888 3016 21894
rect 2964 21830 3016 21836
rect 2976 21554 3004 21830
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 3160 21486 3188 23734
rect 3252 21690 3280 27406
rect 4252 27328 4304 27334
rect 4080 27276 4252 27282
rect 4080 27270 4304 27276
rect 4080 27254 4292 27270
rect 3792 25152 3844 25158
rect 3792 25094 3844 25100
rect 3804 24886 3832 25094
rect 3792 24880 3844 24886
rect 3792 24822 3844 24828
rect 3332 24744 3384 24750
rect 3332 24686 3384 24692
rect 3344 24410 3372 24686
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3804 23322 3832 23666
rect 3792 23316 3844 23322
rect 3792 23258 3844 23264
rect 4080 23254 4108 27254
rect 4620 26852 4672 26858
rect 4620 26794 4672 26800
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26450 4660 26794
rect 4620 26444 4672 26450
rect 4620 26386 4672 26392
rect 4620 26308 4672 26314
rect 4620 26250 4672 26256
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4528 25152 4580 25158
rect 4528 25094 4580 25100
rect 4540 24954 4568 25094
rect 4528 24948 4580 24954
rect 4528 24890 4580 24896
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3608 23248 3660 23254
rect 3608 23190 3660 23196
rect 4068 23248 4120 23254
rect 4068 23190 4120 23196
rect 4344 23248 4396 23254
rect 4344 23190 4396 23196
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3148 21480 3200 21486
rect 3148 21422 3200 21428
rect 2964 20936 3016 20942
rect 2964 20878 3016 20884
rect 2976 20602 3004 20878
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 3436 20534 3464 20742
rect 3424 20528 3476 20534
rect 3424 20470 3476 20476
rect 2884 20182 3004 20210
rect 2976 19446 3004 20182
rect 2964 19440 3016 19446
rect 2964 19382 3016 19388
rect 3620 19378 3648 23190
rect 4160 23180 4212 23186
rect 4160 23122 4212 23128
rect 4068 22976 4120 22982
rect 4068 22918 4120 22924
rect 4080 22642 4108 22918
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 4172 22522 4200 23122
rect 4356 22778 4384 23190
rect 4632 22794 4660 26250
rect 4724 25226 4752 29242
rect 5368 28694 5396 29582
rect 5460 28994 5488 37198
rect 6840 36922 6868 37198
rect 7392 37126 7420 39358
rect 10322 39358 10640 39386
rect 10322 39280 10378 39358
rect 10416 37256 10468 37262
rect 10416 37198 10468 37204
rect 7380 37120 7432 37126
rect 7380 37062 7432 37068
rect 6828 36916 6880 36922
rect 6828 36858 6880 36864
rect 6920 36780 6972 36786
rect 6920 36722 6972 36728
rect 6368 36100 6420 36106
rect 6368 36042 6420 36048
rect 6380 35834 6408 36042
rect 6368 35828 6420 35834
rect 6368 35770 6420 35776
rect 6184 35692 6236 35698
rect 6184 35634 6236 35640
rect 6196 35290 6224 35634
rect 6184 35284 6236 35290
rect 6184 35226 6236 35232
rect 6736 35148 6788 35154
rect 6736 35090 6788 35096
rect 6368 34740 6420 34746
rect 6368 34682 6420 34688
rect 5632 34604 5684 34610
rect 5632 34546 5684 34552
rect 5644 33998 5672 34546
rect 5632 33992 5684 33998
rect 5684 33952 5764 33980
rect 5632 33934 5684 33940
rect 5540 31680 5592 31686
rect 5540 31622 5592 31628
rect 5632 31680 5684 31686
rect 5632 31622 5684 31628
rect 5552 31210 5580 31622
rect 5540 31204 5592 31210
rect 5540 31146 5592 31152
rect 5644 31142 5672 31622
rect 5632 31136 5684 31142
rect 5632 31078 5684 31084
rect 5644 30802 5672 31078
rect 5632 30796 5684 30802
rect 5632 30738 5684 30744
rect 5736 29714 5764 33952
rect 6276 33856 6328 33862
rect 6276 33798 6328 33804
rect 6288 33522 6316 33798
rect 6276 33516 6328 33522
rect 6276 33458 6328 33464
rect 6380 31822 6408 34682
rect 6748 34542 6776 35090
rect 6932 34542 6960 36722
rect 10428 36650 10456 37198
rect 10612 37126 10640 39358
rect 13542 39280 13598 40080
rect 16118 39386 16174 40080
rect 19338 39386 19394 40080
rect 22558 39386 22614 40080
rect 25778 39386 25834 40080
rect 28354 39386 28410 40080
rect 31574 39386 31630 40080
rect 16118 39358 16436 39386
rect 16118 39280 16174 39358
rect 12808 37256 12860 37262
rect 12808 37198 12860 37204
rect 10600 37120 10652 37126
rect 10600 37062 10652 37068
rect 10416 36644 10468 36650
rect 10416 36586 10468 36592
rect 8484 36168 8536 36174
rect 8484 36110 8536 36116
rect 7196 36032 7248 36038
rect 7196 35974 7248 35980
rect 7208 35086 7236 35974
rect 7196 35080 7248 35086
rect 7196 35022 7248 35028
rect 7012 34604 7064 34610
rect 7012 34546 7064 34552
rect 6736 34536 6788 34542
rect 6736 34478 6788 34484
rect 6920 34536 6972 34542
rect 6920 34478 6972 34484
rect 7024 34202 7052 34546
rect 7104 34400 7156 34406
rect 7104 34342 7156 34348
rect 7012 34196 7064 34202
rect 7012 34138 7064 34144
rect 7012 34060 7064 34066
rect 7012 34002 7064 34008
rect 6828 33040 6880 33046
rect 7024 32994 7052 34002
rect 7116 33930 7144 34342
rect 7104 33924 7156 33930
rect 7104 33866 7156 33872
rect 6880 32988 7052 32994
rect 6828 32982 7052 32988
rect 6840 32966 7052 32982
rect 6828 32904 6880 32910
rect 6828 32846 6880 32852
rect 6840 32434 6868 32846
rect 6932 32570 6960 32966
rect 7116 32892 7144 33866
rect 7208 33046 7236 35022
rect 7288 35012 7340 35018
rect 7288 34954 7340 34960
rect 7300 33862 7328 34954
rect 8496 34610 8524 36110
rect 10324 35284 10376 35290
rect 10324 35226 10376 35232
rect 9864 35012 9916 35018
rect 9864 34954 9916 34960
rect 9220 34944 9272 34950
rect 9220 34886 9272 34892
rect 9232 34678 9260 34886
rect 9876 34746 9904 34954
rect 9864 34740 9916 34746
rect 9864 34682 9916 34688
rect 10048 34740 10100 34746
rect 10048 34682 10100 34688
rect 9220 34672 9272 34678
rect 9220 34614 9272 34620
rect 8484 34604 8536 34610
rect 8484 34546 8536 34552
rect 7564 34400 7616 34406
rect 7564 34342 7616 34348
rect 7576 34066 7604 34342
rect 8496 34202 8524 34546
rect 8484 34196 8536 34202
rect 8484 34138 8536 34144
rect 7564 34060 7616 34066
rect 7564 34002 7616 34008
rect 9772 33924 9824 33930
rect 9772 33866 9824 33872
rect 7288 33856 7340 33862
rect 7288 33798 7340 33804
rect 7196 33040 7248 33046
rect 7196 32982 7248 32988
rect 7024 32864 7144 32892
rect 6920 32564 6972 32570
rect 6920 32506 6972 32512
rect 6828 32428 6880 32434
rect 6828 32370 6880 32376
rect 6918 32328 6974 32337
rect 6918 32263 6920 32272
rect 6972 32263 6974 32272
rect 6920 32234 6972 32240
rect 6644 32020 6696 32026
rect 6644 31962 6696 31968
rect 6656 31822 6684 31962
rect 6368 31816 6420 31822
rect 6196 31764 6368 31770
rect 6196 31758 6420 31764
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6644 31816 6696 31822
rect 6644 31758 6696 31764
rect 6196 31742 6408 31758
rect 6196 30802 6224 31742
rect 6472 31210 6500 31758
rect 6460 31204 6512 31210
rect 6460 31146 6512 31152
rect 5816 30796 5868 30802
rect 5816 30738 5868 30744
rect 6184 30796 6236 30802
rect 6184 30738 6236 30744
rect 6368 30796 6420 30802
rect 6472 30784 6500 31146
rect 6644 30796 6696 30802
rect 6420 30756 6500 30784
rect 6564 30756 6644 30784
rect 6368 30738 6420 30744
rect 5724 29708 5776 29714
rect 5724 29650 5776 29656
rect 5736 29306 5764 29650
rect 5724 29300 5776 29306
rect 5724 29242 5776 29248
rect 5460 28966 5580 28994
rect 5828 28966 5856 30738
rect 5908 29776 5960 29782
rect 5908 29718 5960 29724
rect 5920 29170 5948 29718
rect 6368 29708 6420 29714
rect 6368 29650 6420 29656
rect 6184 29504 6236 29510
rect 6184 29446 6236 29452
rect 6196 29170 6224 29446
rect 5908 29164 5960 29170
rect 5908 29106 5960 29112
rect 6184 29164 6236 29170
rect 6184 29106 6236 29112
rect 5356 28688 5408 28694
rect 5276 28636 5356 28642
rect 5276 28630 5408 28636
rect 5276 28614 5396 28630
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5276 27554 5304 28614
rect 5356 28552 5408 28558
rect 5356 28494 5408 28500
rect 5368 28218 5396 28494
rect 5356 28212 5408 28218
rect 5356 28154 5408 28160
rect 4804 27532 4856 27538
rect 4804 27474 4856 27480
rect 5092 27526 5304 27554
rect 5368 27538 5396 28154
rect 5356 27532 5408 27538
rect 4816 26450 4844 27474
rect 5092 27470 5120 27526
rect 5356 27474 5408 27480
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4804 26444 4856 26450
rect 4804 26386 4856 26392
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4988 25968 5040 25974
rect 4988 25910 5040 25916
rect 5000 25362 5028 25910
rect 4988 25356 5040 25362
rect 4988 25298 5040 25304
rect 5448 25356 5500 25362
rect 5448 25298 5500 25304
rect 4804 25288 4856 25294
rect 4804 25230 4856 25236
rect 5264 25288 5316 25294
rect 5264 25230 5316 25236
rect 4712 25220 4764 25226
rect 4712 25162 4764 25168
rect 4724 24018 4752 25162
rect 4816 24206 4844 25230
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5276 24426 5304 25230
rect 5184 24398 5304 24426
rect 5184 24274 5212 24398
rect 5264 24336 5316 24342
rect 5264 24278 5316 24284
rect 5172 24268 5224 24274
rect 5172 24210 5224 24216
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4724 23990 4844 24018
rect 4712 23520 4764 23526
rect 4712 23462 4764 23468
rect 4724 23050 4752 23462
rect 4712 23044 4764 23050
rect 4712 22986 4764 22992
rect 4816 22930 4844 23990
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4344 22772 4396 22778
rect 4344 22714 4396 22720
rect 4448 22766 4660 22794
rect 4724 22902 4844 22930
rect 4080 22494 4200 22522
rect 3884 22432 3936 22438
rect 3884 22374 3936 22380
rect 3896 20806 3924 22374
rect 4080 22216 4108 22494
rect 4448 22438 4476 22766
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4436 22432 4488 22438
rect 4436 22374 4488 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22234 4660 22578
rect 4620 22228 4672 22234
rect 4080 22188 4200 22216
rect 4080 22094 4108 22188
rect 4172 22098 4200 22188
rect 4620 22170 4672 22176
rect 3988 22066 4108 22094
rect 4160 22092 4212 22098
rect 3988 21010 4016 22066
rect 4160 22034 4212 22040
rect 4068 21616 4120 21622
rect 4068 21558 4120 21564
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 4080 20942 4108 21558
rect 4620 21412 4672 21418
rect 4620 21354 4672 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21010 4660 21354
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 4436 20868 4488 20874
rect 4436 20810 4488 20816
rect 3884 20800 3936 20806
rect 3884 20742 3936 20748
rect 4448 20602 4476 20810
rect 4620 20800 4672 20806
rect 4620 20742 4672 20748
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4632 19718 4660 20742
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4356 19378 4384 19654
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2700 18222 2728 19110
rect 2884 18970 2912 19314
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2872 18352 2924 18358
rect 2872 18294 2924 18300
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2792 16182 2820 17614
rect 2884 17542 2912 18294
rect 2976 18222 3004 19246
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4080 18290 4108 18770
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4540 18290 4568 18702
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4528 18284 4580 18290
rect 4528 18226 4580 18232
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 4080 17338 4108 17546
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4632 17218 4660 19314
rect 4724 19174 4752 22902
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4804 22772 4856 22778
rect 4804 22714 4856 22720
rect 4816 22030 4844 22714
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 5276 21894 5304 24278
rect 5460 23254 5488 25298
rect 5448 23248 5500 23254
rect 5448 23190 5500 23196
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5460 22778 5488 23054
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 4804 21888 4856 21894
rect 4804 21830 4856 21836
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 4816 21418 4844 21830
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5460 21570 5488 22714
rect 5276 21554 5488 21570
rect 5264 21548 5488 21554
rect 5316 21542 5488 21548
rect 5264 21490 5316 21496
rect 4804 21412 4856 21418
rect 4804 21354 4856 21360
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4724 17338 4752 19110
rect 4816 18086 4844 21354
rect 5368 21010 5396 21542
rect 5448 21480 5500 21486
rect 5448 21422 5500 21428
rect 5460 21350 5488 21422
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5356 21004 5408 21010
rect 5356 20946 5408 20952
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5276 18970 5304 20946
rect 5552 19334 5580 28966
rect 5816 28960 5868 28966
rect 5816 28902 5868 28908
rect 5828 28694 5856 28902
rect 5816 28688 5868 28694
rect 5816 28630 5868 28636
rect 5920 28626 5948 29106
rect 6380 29102 6408 29650
rect 6368 29096 6420 29102
rect 6368 29038 6420 29044
rect 6564 28626 6592 30756
rect 6644 30738 6696 30744
rect 7024 30258 7052 32864
rect 7208 32366 7236 32982
rect 7196 32360 7248 32366
rect 7196 32302 7248 32308
rect 7104 32292 7156 32298
rect 7104 32234 7156 32240
rect 7116 31958 7144 32234
rect 7104 31952 7156 31958
rect 7104 31894 7156 31900
rect 7196 31884 7248 31890
rect 7196 31826 7248 31832
rect 7208 30818 7236 31826
rect 7300 31414 7328 33798
rect 7380 33108 7432 33114
rect 7380 33050 7432 33056
rect 9496 33108 9548 33114
rect 9496 33050 9548 33056
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 7392 31890 7420 33050
rect 8024 32972 8076 32978
rect 8024 32914 8076 32920
rect 7656 32904 7708 32910
rect 7656 32846 7708 32852
rect 7668 32774 7696 32846
rect 7656 32768 7708 32774
rect 7656 32710 7708 32716
rect 7564 32428 7616 32434
rect 7668 32416 7696 32710
rect 8036 32450 8064 32914
rect 9508 32570 9536 33050
rect 9588 32768 9640 32774
rect 9588 32710 9640 32716
rect 8208 32564 8260 32570
rect 8208 32506 8260 32512
rect 8944 32564 8996 32570
rect 8944 32506 8996 32512
rect 9496 32564 9548 32570
rect 9496 32506 9548 32512
rect 8036 32422 8156 32450
rect 7616 32388 7696 32416
rect 7564 32370 7616 32376
rect 7840 32360 7892 32366
rect 7840 32302 7892 32308
rect 7852 32026 7880 32302
rect 7840 32020 7892 32026
rect 7840 31962 7892 31968
rect 7380 31884 7432 31890
rect 7380 31826 7432 31832
rect 7472 31816 7524 31822
rect 8128 31793 8156 32422
rect 8220 32230 8248 32506
rect 8956 32434 8984 32506
rect 8484 32428 8536 32434
rect 8484 32370 8536 32376
rect 8944 32428 8996 32434
rect 8944 32370 8996 32376
rect 8392 32360 8444 32366
rect 8392 32302 8444 32308
rect 8208 32224 8260 32230
rect 8208 32166 8260 32172
rect 7472 31758 7524 31764
rect 8114 31784 8170 31793
rect 7288 31408 7340 31414
rect 7288 31350 7340 31356
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7392 30938 7420 31282
rect 7380 30932 7432 30938
rect 7380 30874 7432 30880
rect 7208 30790 7328 30818
rect 7196 30728 7248 30734
rect 7196 30670 7248 30676
rect 7104 30592 7156 30598
rect 7104 30534 7156 30540
rect 7116 30433 7144 30534
rect 7102 30424 7158 30433
rect 7102 30359 7158 30368
rect 7208 30326 7236 30670
rect 7196 30320 7248 30326
rect 7196 30262 7248 30268
rect 7012 30252 7064 30258
rect 7012 30194 7064 30200
rect 7300 30002 7328 30790
rect 7208 29974 7328 30002
rect 5908 28620 5960 28626
rect 5908 28562 5960 28568
rect 6552 28620 6604 28626
rect 6552 28562 6604 28568
rect 5920 27538 5948 28562
rect 6184 28552 6236 28558
rect 6104 28512 6184 28540
rect 6104 28422 6132 28512
rect 6184 28494 6236 28500
rect 6092 28416 6144 28422
rect 6092 28358 6144 28364
rect 7104 28416 7156 28422
rect 7104 28358 7156 28364
rect 6104 27538 6132 28358
rect 5908 27532 5960 27538
rect 5908 27474 5960 27480
rect 6092 27532 6144 27538
rect 6092 27474 6144 27480
rect 6920 27532 6972 27538
rect 6920 27474 6972 27480
rect 6184 27464 6236 27470
rect 6184 27406 6236 27412
rect 6196 26858 6224 27406
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6184 26852 6236 26858
rect 6184 26794 6236 26800
rect 6196 25514 6224 26794
rect 6840 26042 6868 27270
rect 6932 26926 6960 27474
rect 7012 27464 7064 27470
rect 7012 27406 7064 27412
rect 7024 26994 7052 27406
rect 7012 26988 7064 26994
rect 7012 26930 7064 26936
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 6368 25900 6420 25906
rect 6368 25842 6420 25848
rect 6104 25486 6224 25514
rect 5816 25356 5868 25362
rect 5816 25298 5868 25304
rect 5828 25158 5856 25298
rect 5908 25288 5960 25294
rect 5908 25230 5960 25236
rect 5816 25152 5868 25158
rect 5816 25094 5868 25100
rect 5828 24800 5856 25094
rect 5736 24772 5856 24800
rect 5736 24274 5764 24772
rect 5920 24698 5948 25230
rect 5828 24670 5948 24698
rect 5724 24268 5776 24274
rect 5724 24210 5776 24216
rect 5828 24206 5856 24670
rect 5816 24200 5868 24206
rect 5816 24142 5868 24148
rect 6000 24200 6052 24206
rect 6000 24142 6052 24148
rect 5828 23526 5856 24142
rect 5816 23520 5868 23526
rect 5816 23462 5868 23468
rect 6012 21418 6040 24142
rect 6000 21412 6052 21418
rect 6000 21354 6052 21360
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5644 21010 5672 21286
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5644 20806 5672 20946
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5368 19306 5580 19334
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 5000 18154 5028 18362
rect 5276 18222 5304 18702
rect 5368 18329 5396 19306
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5354 18320 5410 18329
rect 5354 18255 5410 18264
rect 5460 18222 5488 18702
rect 5552 18630 5580 18702
rect 5828 18630 5856 20878
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5538 18320 5594 18329
rect 5538 18255 5594 18264
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5264 18216 5316 18222
rect 5448 18216 5500 18222
rect 5316 18176 5396 18204
rect 5264 18158 5316 18164
rect 4988 18148 5040 18154
rect 4988 18090 5040 18096
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 5092 17882 5120 18158
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5276 17338 5304 17818
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 4632 17190 4752 17218
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4724 16726 4752 17190
rect 5264 17060 5316 17066
rect 5264 17002 5316 17008
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 2780 16176 2832 16182
rect 2780 16118 2832 16124
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2700 15706 2728 16050
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 3068 15502 3096 16390
rect 4172 16250 4200 16390
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4632 16182 4660 16390
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4724 15586 4752 16662
rect 5276 16658 5304 17002
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4816 15706 4844 16526
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4724 15558 4844 15586
rect 5276 15570 5304 16594
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3988 14414 4016 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3804 14006 3832 14214
rect 4632 14074 4660 15030
rect 4816 15026 4844 15558
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5368 15094 5396 18176
rect 5448 18158 5500 18164
rect 5460 16522 5488 18158
rect 5448 16516 5500 16522
rect 5448 16458 5500 16464
rect 5552 16402 5580 18255
rect 5644 17814 5672 18362
rect 5920 18034 5948 19654
rect 6104 18358 6132 25486
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 6184 23588 6236 23594
rect 6184 23530 6236 23536
rect 6196 21690 6224 23530
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6184 21480 6236 21486
rect 6184 21422 6236 21428
rect 6196 18766 6224 21422
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6092 18352 6144 18358
rect 6092 18294 6144 18300
rect 6104 18222 6132 18294
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 5920 18006 6040 18034
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 6012 17202 6040 18006
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 5460 16374 5580 16402
rect 5356 15088 5408 15094
rect 5356 15030 5408 15036
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 4724 13938 4752 14350
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12152 4660 13262
rect 4712 12164 4764 12170
rect 4632 12124 4712 12152
rect 4632 11830 4660 12124
rect 4712 12106 4764 12112
rect 4620 11824 4672 11830
rect 4158 11792 4214 11801
rect 4620 11766 4672 11772
rect 4158 11727 4160 11736
rect 4212 11727 4214 11736
rect 4160 11698 4212 11704
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10130 4660 11494
rect 4816 10266 4844 14962
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5368 14414 5396 14758
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5460 14226 5488 16374
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5736 15502 5764 15846
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 6012 15366 6040 17138
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 5368 14198 5488 14226
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5368 12918 5396 14198
rect 6288 13326 6316 24550
rect 6380 18426 6408 25842
rect 6644 25696 6696 25702
rect 6644 25638 6696 25644
rect 6656 24818 6684 25638
rect 7012 25220 7064 25226
rect 7012 25162 7064 25168
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 6644 24812 6696 24818
rect 6644 24754 6696 24760
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6656 23662 6684 24006
rect 6644 23656 6696 23662
rect 6644 23598 6696 23604
rect 6644 19984 6696 19990
rect 6644 19926 6696 19932
rect 6656 18970 6684 19926
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6368 18420 6420 18426
rect 6368 18362 6420 18368
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 6642 18184 6698 18193
rect 6380 17746 6408 18158
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 6564 17542 6592 18158
rect 6642 18119 6698 18128
rect 6656 17814 6684 18119
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6368 16516 6420 16522
rect 6368 16458 6420 16464
rect 6380 16250 6408 16458
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6564 16114 6592 16934
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6656 14958 6684 15302
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6656 13394 6684 14894
rect 6748 14006 6776 24006
rect 6932 22166 6960 25094
rect 7024 24750 7052 25162
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 7116 24698 7144 28358
rect 7208 25498 7236 29974
rect 7392 27606 7420 30874
rect 7288 27600 7340 27606
rect 7288 27542 7340 27548
rect 7380 27600 7432 27606
rect 7380 27542 7432 27548
rect 7300 26858 7328 27542
rect 7288 26852 7340 26858
rect 7288 26794 7340 26800
rect 7300 26518 7328 26794
rect 7288 26512 7340 26518
rect 7288 26454 7340 26460
rect 7288 25832 7340 25838
rect 7288 25774 7340 25780
rect 7196 25492 7248 25498
rect 7196 25434 7248 25440
rect 7300 25294 7328 25774
rect 7380 25696 7432 25702
rect 7380 25638 7432 25644
rect 7288 25288 7340 25294
rect 7288 25230 7340 25236
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 7208 24818 7236 25094
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 7024 24206 7052 24686
rect 7116 24670 7236 24698
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7116 24206 7144 24550
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7104 22976 7156 22982
rect 7104 22918 7156 22924
rect 6920 22160 6972 22166
rect 6920 22102 6972 22108
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6932 20942 6960 21286
rect 7024 20942 7052 21830
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7010 19272 7066 19281
rect 7010 19207 7066 19216
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6932 17746 6960 18158
rect 7024 18154 7052 19207
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6840 17066 6868 17478
rect 6828 17060 6880 17066
rect 6828 17002 6880 17008
rect 6840 16454 6868 17002
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6932 15162 6960 17682
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7024 15910 7052 17614
rect 7116 17338 7144 22918
rect 7208 22094 7236 24670
rect 7288 24268 7340 24274
rect 7288 24210 7340 24216
rect 7300 23866 7328 24210
rect 7392 24206 7420 25638
rect 7484 25362 7512 31758
rect 8114 31719 8170 31728
rect 7656 31340 7708 31346
rect 7656 31282 7708 31288
rect 7564 31272 7616 31278
rect 7564 31214 7616 31220
rect 7576 29782 7604 31214
rect 7564 29776 7616 29782
rect 7564 29718 7616 29724
rect 7576 29578 7604 29718
rect 7668 29646 7696 31282
rect 8024 31136 8076 31142
rect 8024 31078 8076 31084
rect 7840 30660 7892 30666
rect 7840 30602 7892 30608
rect 7852 30394 7880 30602
rect 7840 30388 7892 30394
rect 7840 30330 7892 30336
rect 8036 30258 8064 31078
rect 8024 30252 8076 30258
rect 8024 30194 8076 30200
rect 7656 29640 7708 29646
rect 7656 29582 7708 29588
rect 7564 29572 7616 29578
rect 7564 29514 7616 29520
rect 7840 29504 7892 29510
rect 7840 29446 7892 29452
rect 7852 29306 7880 29446
rect 7840 29300 7892 29306
rect 7840 29242 7892 29248
rect 7852 27470 7880 29242
rect 8128 28506 8156 31719
rect 8404 31278 8432 32302
rect 8496 32026 8524 32370
rect 8760 32224 8812 32230
rect 8760 32166 8812 32172
rect 8484 32020 8536 32026
rect 8484 31962 8536 31968
rect 8772 31754 8800 32166
rect 8956 31822 8984 32370
rect 9496 32360 9548 32366
rect 9496 32302 9548 32308
rect 9128 32224 9180 32230
rect 9128 32166 9180 32172
rect 9140 31822 9168 32166
rect 9312 31952 9364 31958
rect 9312 31894 9364 31900
rect 8944 31816 8996 31822
rect 8944 31758 8996 31764
rect 9128 31816 9180 31822
rect 9128 31758 9180 31764
rect 8680 31726 8800 31754
rect 8576 31680 8628 31686
rect 8576 31622 8628 31628
rect 8392 31272 8444 31278
rect 8392 31214 8444 31220
rect 8404 30190 8432 31214
rect 8392 30184 8444 30190
rect 8392 30126 8444 30132
rect 8208 29640 8260 29646
rect 8208 29582 8260 29588
rect 8036 28478 8156 28506
rect 7840 27464 7892 27470
rect 7576 27412 7840 27418
rect 7576 27406 7892 27412
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 7576 27390 7880 27406
rect 7576 26994 7604 27390
rect 7944 27334 7972 27406
rect 7656 27328 7708 27334
rect 7656 27270 7708 27276
rect 7932 27328 7984 27334
rect 7932 27270 7984 27276
rect 7668 26994 7696 27270
rect 7564 26988 7616 26994
rect 7564 26930 7616 26936
rect 7656 26988 7708 26994
rect 7656 26930 7708 26936
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 7564 25900 7616 25906
rect 7564 25842 7616 25848
rect 7576 25362 7604 25842
rect 7472 25356 7524 25362
rect 7472 25298 7524 25304
rect 7564 25356 7616 25362
rect 7564 25298 7616 25304
rect 7668 24818 7696 26726
rect 7932 26512 7984 26518
rect 7932 26454 7984 26460
rect 7748 24880 7800 24886
rect 7748 24822 7800 24828
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7564 24676 7616 24682
rect 7564 24618 7616 24624
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7576 23866 7604 24618
rect 7288 23860 7340 23866
rect 7288 23802 7340 23808
rect 7564 23860 7616 23866
rect 7564 23802 7616 23808
rect 7564 23044 7616 23050
rect 7564 22986 7616 22992
rect 7576 22642 7604 22986
rect 7656 22704 7708 22710
rect 7656 22646 7708 22652
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7208 22066 7328 22094
rect 7194 21856 7250 21865
rect 7194 21791 7250 21800
rect 7208 21554 7236 21791
rect 7300 21690 7328 22066
rect 7380 21956 7432 21962
rect 7380 21898 7432 21904
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 7392 21554 7420 21898
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 7208 20058 7236 20946
rect 7576 20942 7604 21286
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7380 20868 7432 20874
rect 7380 20810 7432 20816
rect 7288 20800 7340 20806
rect 7288 20742 7340 20748
rect 7300 20466 7328 20742
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7392 19990 7420 20810
rect 7668 20602 7696 22646
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7380 19984 7432 19990
rect 7380 19926 7432 19932
rect 7392 19854 7420 19926
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7208 17678 7236 18362
rect 7380 18216 7432 18222
rect 7576 18193 7604 18770
rect 7380 18158 7432 18164
rect 7562 18184 7618 18193
rect 7392 17746 7420 18158
rect 7562 18119 7618 18128
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6932 14618 6960 15098
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6840 13938 6868 14350
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6840 13258 6868 13874
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5460 12850 5488 13126
rect 6840 12850 6868 13194
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5356 12096 5408 12102
rect 5736 12073 5764 12174
rect 5356 12038 5408 12044
rect 5722 12064 5778 12073
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9364 4200 9998
rect 4080 9336 4200 9364
rect 4080 9058 4108 9336
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9178 4660 10066
rect 5000 10062 5028 10610
rect 5092 10130 5120 10610
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4816 9586 4844 9998
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4080 9030 4200 9058
rect 4172 8974 4200 9030
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 5276 7886 5304 8774
rect 5368 8090 5396 12038
rect 5722 11999 5778 12008
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5736 10674 5764 10950
rect 5920 10674 5948 12718
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5552 9654 5580 10610
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5644 9586 5672 10134
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5460 8022 5488 9454
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4632 7274 4660 7686
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5276 6322 5304 6598
rect 5368 6458 5396 7822
rect 5460 7818 5488 7958
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 6866 5488 7346
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5736 6322 5764 9930
rect 5920 9518 5948 10610
rect 6380 10470 6408 12718
rect 6840 12238 6868 12786
rect 7116 12238 7144 12786
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6932 11762 6960 12106
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 7208 11150 7236 13398
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12850 7420 13126
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7668 12782 7696 20538
rect 7760 17882 7788 24822
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7852 22234 7880 22578
rect 7840 22228 7892 22234
rect 7840 22170 7892 22176
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7852 16250 7880 21830
rect 7944 18834 7972 26454
rect 8036 25498 8064 28478
rect 8116 27464 8168 27470
rect 8116 27406 8168 27412
rect 8128 27334 8156 27406
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 8220 27146 8248 29582
rect 8404 29170 8432 30126
rect 8392 29164 8444 29170
rect 8392 29106 8444 29112
rect 8404 28082 8432 29106
rect 8588 28422 8616 31622
rect 8576 28416 8628 28422
rect 8576 28358 8628 28364
rect 8392 28076 8444 28082
rect 8392 28018 8444 28024
rect 8128 27118 8248 27146
rect 8024 25492 8076 25498
rect 8024 25434 8076 25440
rect 8128 22982 8156 27118
rect 8484 26988 8536 26994
rect 8484 26930 8536 26936
rect 8496 26314 8524 26930
rect 8588 26450 8616 28358
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 8208 25900 8260 25906
rect 8208 25842 8260 25848
rect 8220 25770 8248 25842
rect 8208 25764 8260 25770
rect 8208 25706 8260 25712
rect 8220 24954 8248 25706
rect 8208 24948 8260 24954
rect 8208 24890 8260 24896
rect 8220 24750 8248 24890
rect 8208 24744 8260 24750
rect 8208 24686 8260 24692
rect 8392 23792 8444 23798
rect 8390 23760 8392 23769
rect 8444 23760 8446 23769
rect 8390 23695 8446 23704
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 8300 22094 8352 22098
rect 8404 22094 8432 22578
rect 8300 22092 8432 22094
rect 8352 22066 8432 22092
rect 8300 22034 8352 22040
rect 8496 21894 8524 26250
rect 8588 23730 8616 26386
rect 8680 25838 8708 31726
rect 9324 31414 9352 31894
rect 9508 31754 9536 32302
rect 9416 31726 9536 31754
rect 9312 31408 9364 31414
rect 9312 31350 9364 31356
rect 9416 31346 9444 31726
rect 9404 31340 9456 31346
rect 9404 31282 9456 31288
rect 9128 30252 9180 30258
rect 9128 30194 9180 30200
rect 9140 29850 9168 30194
rect 9128 29844 9180 29850
rect 9128 29786 9180 29792
rect 9496 29640 9548 29646
rect 9496 29582 9548 29588
rect 9508 29306 9536 29582
rect 9496 29300 9548 29306
rect 9496 29242 9548 29248
rect 8944 28688 8996 28694
rect 8944 28630 8996 28636
rect 8956 28150 8984 28630
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 9324 28150 9352 28494
rect 8944 28144 8996 28150
rect 8944 28086 8996 28092
rect 9312 28144 9364 28150
rect 9312 28086 9364 28092
rect 8760 27328 8812 27334
rect 8760 27270 8812 27276
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8668 25696 8720 25702
rect 8668 25638 8720 25644
rect 8680 24206 8708 25638
rect 8668 24200 8720 24206
rect 8668 24142 8720 24148
rect 8576 23724 8628 23730
rect 8576 23666 8628 23672
rect 8588 23526 8616 23666
rect 8576 23520 8628 23526
rect 8576 23462 8628 23468
rect 8680 23338 8708 24142
rect 8588 23310 8708 23338
rect 8588 22710 8616 23310
rect 8576 22704 8628 22710
rect 8576 22646 8628 22652
rect 8588 22098 8616 22646
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 8036 20942 8064 21490
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8680 21146 8708 21422
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8024 20936 8076 20942
rect 8024 20878 8076 20884
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 8036 18970 8064 19246
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 7932 18692 7984 18698
rect 7932 18634 7984 18640
rect 7944 17678 7972 18634
rect 8036 17814 8064 18906
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7748 15428 7800 15434
rect 7748 15370 7800 15376
rect 7760 14958 7788 15370
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7944 14346 7972 17614
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 8036 15978 8064 16458
rect 8024 15972 8076 15978
rect 8024 15914 8076 15920
rect 8128 15026 8156 19654
rect 8220 18426 8248 20402
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8312 19854 8340 20198
rect 8496 20058 8524 20742
rect 8772 20602 8800 27270
rect 9508 26790 9536 29242
rect 9496 26784 9548 26790
rect 9496 26726 9548 26732
rect 9220 26376 9272 26382
rect 9220 26318 9272 26324
rect 9128 25900 9180 25906
rect 9128 25842 9180 25848
rect 9140 25498 9168 25842
rect 9232 25702 9260 26318
rect 9404 26036 9456 26042
rect 9404 25978 9456 25984
rect 9416 25906 9444 25978
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 9416 25514 9444 25842
rect 9128 25492 9180 25498
rect 9128 25434 9180 25440
rect 9324 25486 9444 25514
rect 9324 25362 9352 25486
rect 9312 25356 9364 25362
rect 9312 25298 9364 25304
rect 9508 25294 9536 26726
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 8852 24132 8904 24138
rect 8852 24074 8904 24080
rect 9312 24132 9364 24138
rect 9312 24074 9364 24080
rect 8864 23866 8892 24074
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 9126 23760 9182 23769
rect 9126 23695 9128 23704
rect 9180 23695 9182 23704
rect 9128 23666 9180 23672
rect 9324 23594 9352 24074
rect 9312 23588 9364 23594
rect 9312 23530 9364 23536
rect 8944 23520 8996 23526
rect 8944 23462 8996 23468
rect 8956 21554 8984 23462
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 9048 21962 9076 22374
rect 9036 21956 9088 21962
rect 9036 21898 9088 21904
rect 9312 21956 9364 21962
rect 9312 21898 9364 21904
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8312 18970 8340 19314
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 9048 18834 9076 19178
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 9140 18766 9168 21490
rect 9324 21418 9352 21898
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 9312 20868 9364 20874
rect 9312 20810 9364 20816
rect 9324 20466 9352 20810
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9232 19174 9260 19246
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9232 18766 9260 19110
rect 9416 18834 9444 19110
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 9048 18426 9076 18634
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 8852 18352 8904 18358
rect 8850 18320 8852 18329
rect 8904 18320 8906 18329
rect 8850 18255 8906 18264
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16590 8432 16934
rect 8864 16794 8892 17070
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8404 16114 8432 16526
rect 8864 16114 8892 16730
rect 9140 16726 9168 18362
rect 9232 18358 9260 18702
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 9416 18290 9444 18770
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9508 17882 9536 25230
rect 9600 21010 9628 32710
rect 9692 32337 9720 33050
rect 9784 32434 9812 33866
rect 9876 33046 9904 34682
rect 9864 33040 9916 33046
rect 9864 32982 9916 32988
rect 10060 32910 10088 34682
rect 10232 34604 10284 34610
rect 10232 34546 10284 34552
rect 10244 34202 10272 34546
rect 10232 34196 10284 34202
rect 10232 34138 10284 34144
rect 10336 34134 10364 35226
rect 11704 35148 11756 35154
rect 11704 35090 11756 35096
rect 11060 35080 11112 35086
rect 11060 35022 11112 35028
rect 11072 34134 11100 35022
rect 11716 34610 11744 35090
rect 11704 34604 11756 34610
rect 11704 34546 11756 34552
rect 12164 34604 12216 34610
rect 12164 34546 12216 34552
rect 11612 34400 11664 34406
rect 11612 34342 11664 34348
rect 10324 34128 10376 34134
rect 10324 34070 10376 34076
rect 11060 34128 11112 34134
rect 11060 34070 11112 34076
rect 10048 32904 10100 32910
rect 10048 32846 10100 32852
rect 10232 32904 10284 32910
rect 10232 32846 10284 32852
rect 9772 32428 9824 32434
rect 9772 32370 9824 32376
rect 9678 32328 9734 32337
rect 9678 32263 9734 32272
rect 9692 31822 9720 32263
rect 10060 31890 10088 32846
rect 10048 31884 10100 31890
rect 10048 31826 10100 31832
rect 10244 31822 10272 32846
rect 9680 31816 9732 31822
rect 9680 31758 9732 31764
rect 10232 31816 10284 31822
rect 10232 31758 10284 31764
rect 10244 31482 10272 31758
rect 10232 31476 10284 31482
rect 10232 31418 10284 31424
rect 10232 30252 10284 30258
rect 10232 30194 10284 30200
rect 9864 30048 9916 30054
rect 9864 29990 9916 29996
rect 10140 30048 10192 30054
rect 10140 29990 10192 29996
rect 9876 29578 9904 29990
rect 9864 29572 9916 29578
rect 9864 29514 9916 29520
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 10048 28552 10100 28558
rect 10152 28540 10180 29990
rect 10244 29850 10272 30194
rect 10232 29844 10284 29850
rect 10232 29786 10284 29792
rect 10336 29306 10364 34070
rect 11624 34066 11652 34342
rect 11612 34060 11664 34066
rect 11612 34002 11664 34008
rect 11716 33930 11744 34546
rect 12176 34202 12204 34546
rect 12164 34196 12216 34202
rect 12164 34138 12216 34144
rect 11704 33924 11756 33930
rect 11704 33866 11756 33872
rect 11796 33108 11848 33114
rect 11440 33068 11796 33096
rect 11440 32978 11468 33068
rect 11848 33068 11928 33096
rect 11796 33050 11848 33056
rect 10692 32972 10744 32978
rect 10692 32914 10744 32920
rect 11428 32972 11480 32978
rect 11428 32914 11480 32920
rect 10508 30252 10560 30258
rect 10508 30194 10560 30200
rect 10520 29510 10548 30194
rect 10600 29640 10652 29646
rect 10600 29582 10652 29588
rect 10508 29504 10560 29510
rect 10508 29446 10560 29452
rect 10612 29306 10640 29582
rect 10324 29300 10376 29306
rect 10324 29242 10376 29248
rect 10600 29300 10652 29306
rect 10600 29242 10652 29248
rect 10704 28966 10732 32914
rect 10968 32904 11020 32910
rect 10968 32846 11020 32852
rect 11060 32904 11112 32910
rect 11060 32846 11112 32852
rect 10980 31890 11008 32846
rect 11072 32230 11100 32846
rect 11520 32768 11572 32774
rect 11440 32728 11520 32756
rect 11244 32496 11296 32502
rect 11244 32438 11296 32444
rect 11060 32224 11112 32230
rect 11060 32166 11112 32172
rect 11072 31890 11100 32166
rect 11256 31890 11284 32438
rect 10968 31884 11020 31890
rect 10968 31826 11020 31832
rect 11060 31884 11112 31890
rect 11060 31826 11112 31832
rect 11244 31884 11296 31890
rect 11244 31826 11296 31832
rect 11336 30728 11388 30734
rect 11336 30670 11388 30676
rect 11348 30394 11376 30670
rect 11336 30388 11388 30394
rect 11336 30330 11388 30336
rect 10968 29572 11020 29578
rect 10968 29514 11020 29520
rect 10692 28960 10744 28966
rect 10692 28902 10744 28908
rect 10100 28512 10180 28540
rect 10416 28552 10468 28558
rect 10048 28494 10100 28500
rect 10416 28494 10468 28500
rect 9784 28218 9812 28494
rect 9772 28212 9824 28218
rect 9772 28154 9824 28160
rect 10060 27538 10088 28494
rect 10428 27538 10456 28494
rect 10704 27538 10732 28902
rect 10876 28620 10928 28626
rect 10876 28562 10928 28568
rect 10048 27532 10100 27538
rect 10048 27474 10100 27480
rect 10416 27532 10468 27538
rect 10416 27474 10468 27480
rect 10692 27532 10744 27538
rect 10692 27474 10744 27480
rect 10428 27130 10456 27474
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 10244 26586 10272 26930
rect 10232 26580 10284 26586
rect 10232 26522 10284 26528
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 10336 25702 10364 25842
rect 10324 25696 10376 25702
rect 10324 25638 10376 25644
rect 10416 25696 10468 25702
rect 10416 25638 10468 25644
rect 10692 25696 10744 25702
rect 10692 25638 10744 25644
rect 9956 25152 10008 25158
rect 9956 25094 10008 25100
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 9876 23730 9904 24006
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9876 23186 9904 23666
rect 9864 23180 9916 23186
rect 9864 23122 9916 23128
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9692 21554 9720 21898
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9692 21078 9720 21490
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9680 21072 9732 21078
rect 9680 21014 9732 21020
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 9784 20874 9812 21286
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9876 20942 9904 21082
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9600 19854 9628 20742
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9692 19786 9720 20198
rect 9680 19780 9732 19786
rect 9680 19722 9732 19728
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9692 18222 9720 18770
rect 9876 18290 9904 19110
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9324 17134 9352 17478
rect 9600 17270 9628 17614
rect 9692 17338 9720 18158
rect 9968 17762 9996 25094
rect 10048 23656 10100 23662
rect 10336 23644 10364 25638
rect 10428 25430 10456 25638
rect 10416 25424 10468 25430
rect 10416 25366 10468 25372
rect 10704 25294 10732 25638
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10888 24682 10916 28562
rect 10980 28540 11008 29514
rect 11244 28620 11296 28626
rect 11244 28562 11296 28568
rect 11152 28552 11204 28558
rect 10980 28512 11152 28540
rect 10980 27470 11008 28512
rect 11152 28494 11204 28500
rect 11256 27554 11284 28562
rect 11072 27538 11284 27554
rect 11060 27532 11284 27538
rect 11112 27526 11284 27532
rect 11060 27474 11112 27480
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 11244 27464 11296 27470
rect 11348 27418 11376 30330
rect 11296 27412 11376 27418
rect 11244 27406 11376 27412
rect 11256 27390 11376 27406
rect 11244 26988 11296 26994
rect 11244 26930 11296 26936
rect 10968 26852 11020 26858
rect 10968 26794 11020 26800
rect 10980 26518 11008 26794
rect 10968 26512 11020 26518
rect 10968 26454 11020 26460
rect 11256 26382 11284 26930
rect 11336 26920 11388 26926
rect 11336 26862 11388 26868
rect 11348 26790 11376 26862
rect 11336 26784 11388 26790
rect 11336 26726 11388 26732
rect 11348 26382 11376 26726
rect 11244 26376 11296 26382
rect 11244 26318 11296 26324
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 11152 25152 11204 25158
rect 11152 25094 11204 25100
rect 10876 24676 10928 24682
rect 10876 24618 10928 24624
rect 10416 23656 10468 23662
rect 10336 23616 10416 23644
rect 10048 23598 10100 23604
rect 10416 23598 10468 23604
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 10692 23656 10744 23662
rect 10692 23598 10744 23604
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 10060 23186 10088 23598
rect 10232 23588 10284 23594
rect 10232 23530 10284 23536
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 10060 22216 10088 23122
rect 10140 22228 10192 22234
rect 10060 22188 10140 22216
rect 10140 22170 10192 22176
rect 10244 19281 10272 23530
rect 10428 23526 10456 23598
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10612 23186 10640 23598
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10612 22642 10640 23122
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10704 22094 10732 23598
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10876 23520 10928 23526
rect 11072 23474 11100 23598
rect 10876 23462 10928 23468
rect 10796 23118 10824 23462
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10612 22066 10732 22094
rect 10508 20868 10560 20874
rect 10508 20810 10560 20816
rect 10520 20398 10548 20810
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10428 19854 10456 20198
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10230 19272 10286 19281
rect 10230 19207 10286 19216
rect 10612 19174 10640 22066
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10796 21622 10824 21830
rect 10784 21616 10836 21622
rect 10784 21558 10836 21564
rect 10888 21078 10916 23462
rect 10980 23446 11100 23474
rect 10980 23322 11008 23446
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 11072 23118 11100 23258
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10600 19168 10652 19174
rect 10600 19110 10652 19116
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10336 18306 10364 18702
rect 10520 18426 10548 18702
rect 10612 18630 10640 18702
rect 10600 18624 10652 18630
rect 10600 18566 10652 18572
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10336 18290 10456 18306
rect 10520 18290 10548 18362
rect 10690 18320 10746 18329
rect 10336 18284 10468 18290
rect 10336 18278 10416 18284
rect 10138 18184 10194 18193
rect 10138 18119 10140 18128
rect 10192 18119 10194 18128
rect 10140 18090 10192 18096
rect 9968 17734 10088 17762
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9968 17202 9996 17478
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 9140 16590 9168 16662
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 9048 16182 9076 16390
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9140 15706 9168 16050
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9232 15366 9260 16186
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7760 12306 7788 12922
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 8036 12434 8064 12718
rect 8220 12434 8248 14214
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 13326 8432 13670
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 12646 8340 13126
rect 8864 12986 8892 13194
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 7852 12406 8064 12434
rect 8128 12406 8248 12434
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7392 11762 7420 12174
rect 7576 11830 7604 12174
rect 7852 12170 7880 12406
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7564 11824 7616 11830
rect 7564 11766 7616 11772
rect 7760 11762 7788 11834
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7300 11354 7328 11494
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7208 10962 7236 11086
rect 7208 10934 7328 10962
rect 7300 10674 7328 10934
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6932 10062 6960 10610
rect 7300 10266 7328 10610
rect 7392 10266 7420 11698
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7484 10810 7512 11086
rect 7852 11082 7880 12106
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6380 9586 6408 9998
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5828 7886 5856 8366
rect 6380 8090 6408 9522
rect 6472 9518 6500 9930
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6564 9722 6592 9862
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 8090 7052 8230
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6736 7880 6788 7886
rect 6920 7880 6972 7886
rect 6788 7840 6920 7868
rect 6736 7822 6788 7828
rect 6920 7822 6972 7828
rect 5828 7342 5856 7822
rect 5920 7410 5948 7822
rect 7116 7546 7144 10066
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7392 9450 7420 9998
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7208 7886 7236 8434
rect 7300 7954 7328 8434
rect 7484 7954 7512 10746
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7208 7410 7236 7822
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7300 7342 7328 7890
rect 7576 7546 7604 10542
rect 7852 10062 7880 11018
rect 7944 10606 7972 11698
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 10742 8064 11494
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 7944 9042 7972 9590
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7886 7696 8230
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 5828 6934 5856 7278
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 4080 4078 4108 6258
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 5828 5710 5856 6870
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 6380 6322 6408 6598
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 6104 5817 6132 6122
rect 6090 5808 6146 5817
rect 6090 5743 6146 5752
rect 7300 5710 7328 6598
rect 7576 6458 7604 7346
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7392 5710 7420 6258
rect 7484 5914 7512 6258
rect 7576 6118 7604 6394
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7668 5692 7696 7822
rect 7852 7750 7880 7890
rect 7944 7886 7972 8978
rect 7932 7880 7984 7886
rect 8128 7868 8156 12406
rect 8588 12238 8616 12786
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 12442 8984 12718
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 9140 12238 9168 12786
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8220 11830 8248 12106
rect 8390 12064 8446 12073
rect 8390 11999 8446 12008
rect 8404 11898 8432 11999
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 8220 11694 8248 11766
rect 8588 11694 8616 12174
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8956 10130 8984 12038
rect 9140 11830 9168 12174
rect 9128 11824 9180 11830
rect 9128 11766 9180 11772
rect 9140 11626 9168 11766
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8588 9518 8616 9862
rect 8956 9722 8984 9862
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 8956 9586 8984 9658
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 9048 9518 9076 11222
rect 9232 10810 9260 15302
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9876 14618 9904 14758
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9784 14006 9812 14350
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9784 13734 9812 13942
rect 9876 13938 9904 14554
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9416 12850 9444 13466
rect 10060 13462 10088 17734
rect 10336 16250 10364 18278
rect 10416 18226 10468 18232
rect 10508 18284 10560 18290
rect 10690 18255 10692 18264
rect 10508 18226 10560 18232
rect 10744 18255 10746 18264
rect 10692 18226 10744 18232
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10428 17678 10456 17818
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10244 15502 10272 16050
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10336 15570 10364 15846
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10520 15502 10548 15846
rect 10796 15502 10824 20198
rect 10888 20058 10916 20402
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 11164 18426 11192 25094
rect 11256 24410 11284 25298
rect 11244 24404 11296 24410
rect 11244 24346 11296 24352
rect 11440 21010 11468 32728
rect 11520 32710 11572 32716
rect 11796 32020 11848 32026
rect 11796 31962 11848 31968
rect 11520 30048 11572 30054
rect 11520 29990 11572 29996
rect 11532 29714 11560 29990
rect 11520 29708 11572 29714
rect 11520 29650 11572 29656
rect 11612 28620 11664 28626
rect 11612 28562 11664 28568
rect 11520 26784 11572 26790
rect 11520 26726 11572 26732
rect 11532 26450 11560 26726
rect 11520 26444 11572 26450
rect 11520 26386 11572 26392
rect 11520 25832 11572 25838
rect 11520 25774 11572 25780
rect 11532 25498 11560 25774
rect 11520 25492 11572 25498
rect 11520 25434 11572 25440
rect 11520 25356 11572 25362
rect 11520 25298 11572 25304
rect 11532 24954 11560 25298
rect 11520 24948 11572 24954
rect 11520 24890 11572 24896
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11532 23322 11560 23802
rect 11624 23769 11652 28562
rect 11808 25906 11836 31962
rect 11900 30394 11928 33068
rect 12440 32904 12492 32910
rect 12440 32846 12492 32852
rect 12256 32768 12308 32774
rect 12256 32710 12308 32716
rect 12268 32502 12296 32710
rect 12256 32496 12308 32502
rect 12256 32438 12308 32444
rect 11980 32428 12032 32434
rect 11980 32370 12032 32376
rect 11992 31754 12020 32370
rect 12452 32026 12480 32846
rect 12440 32020 12492 32026
rect 12440 31962 12492 31968
rect 11992 31726 12112 31754
rect 12084 30734 12112 31726
rect 12072 30728 12124 30734
rect 12124 30688 12204 30716
rect 12072 30670 12124 30676
rect 11888 30388 11940 30394
rect 11888 30330 11940 30336
rect 12176 30326 12204 30688
rect 12348 30660 12400 30666
rect 12348 30602 12400 30608
rect 12360 30394 12388 30602
rect 12348 30388 12400 30394
rect 12348 30330 12400 30336
rect 12164 30320 12216 30326
rect 12164 30262 12216 30268
rect 12176 28626 12204 30262
rect 12532 29164 12584 29170
rect 12532 29106 12584 29112
rect 12440 29028 12492 29034
rect 12440 28970 12492 28976
rect 12164 28620 12216 28626
rect 12164 28562 12216 28568
rect 12452 28558 12480 28970
rect 12440 28552 12492 28558
rect 12440 28494 12492 28500
rect 12072 28416 12124 28422
rect 12072 28358 12124 28364
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 11888 26376 11940 26382
rect 11888 26318 11940 26324
rect 11796 25900 11848 25906
rect 11796 25842 11848 25848
rect 11900 24818 11928 26318
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 11888 24676 11940 24682
rect 11888 24618 11940 24624
rect 11704 24336 11756 24342
rect 11704 24278 11756 24284
rect 11610 23760 11666 23769
rect 11610 23695 11612 23704
rect 11664 23695 11666 23704
rect 11612 23666 11664 23672
rect 11716 23322 11744 24278
rect 11900 23730 11928 24618
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 11704 23316 11756 23322
rect 11704 23258 11756 23264
rect 11900 23254 11928 23666
rect 11888 23248 11940 23254
rect 11888 23190 11940 23196
rect 11992 22094 12020 27270
rect 12084 25226 12112 28358
rect 12544 28218 12572 29106
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12164 26784 12216 26790
rect 12164 26726 12216 26732
rect 12176 26382 12204 26726
rect 12164 26376 12216 26382
rect 12164 26318 12216 26324
rect 12452 26042 12480 26930
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12164 25832 12216 25838
rect 12164 25774 12216 25780
rect 12176 25430 12204 25774
rect 12164 25424 12216 25430
rect 12164 25366 12216 25372
rect 12072 25220 12124 25226
rect 12072 25162 12124 25168
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12624 24812 12676 24818
rect 12624 24754 12676 24760
rect 12360 24410 12388 24754
rect 12348 24404 12400 24410
rect 12348 24346 12400 24352
rect 12636 24138 12664 24754
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12716 24132 12768 24138
rect 12716 24074 12768 24080
rect 12728 23798 12756 24074
rect 12716 23792 12768 23798
rect 12716 23734 12768 23740
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12544 22642 12572 23666
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12624 22568 12676 22574
rect 12624 22510 12676 22516
rect 12636 22234 12664 22510
rect 12624 22228 12676 22234
rect 12624 22170 12676 22176
rect 11992 22066 12112 22094
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11796 21956 11848 21962
rect 11796 21898 11848 21904
rect 11808 21690 11836 21898
rect 11992 21690 12020 21966
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11520 21480 11572 21486
rect 11520 21422 11572 21428
rect 11532 21010 11560 21422
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11256 20466 11284 20946
rect 12084 20942 12112 22066
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 11888 20868 11940 20874
rect 11888 20810 11940 20816
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11716 20398 11744 20742
rect 11808 20534 11836 20742
rect 11900 20534 11928 20810
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11888 20528 11940 20534
rect 11888 20470 11940 20476
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 11704 20392 11756 20398
rect 11704 20334 11756 20340
rect 11244 19984 11296 19990
rect 11244 19926 11296 19932
rect 11256 18970 11284 19926
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12452 19514 12480 19722
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12624 19236 12676 19242
rect 12624 19178 12676 19184
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10888 17338 10916 17614
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 11532 17202 11560 18702
rect 11992 18698 12020 19110
rect 11888 18692 11940 18698
rect 11888 18634 11940 18640
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11716 18329 11744 18566
rect 11900 18426 11928 18634
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11702 18320 11758 18329
rect 12084 18290 12112 19110
rect 11702 18255 11758 18264
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12636 18086 12664 19178
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11532 16998 11560 17138
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11808 16794 11836 17138
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 12544 16114 12572 16934
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12452 15706 12480 16050
rect 12728 15910 12756 20402
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10520 15094 10548 15438
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10704 14074 10732 14350
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9416 11150 9444 11494
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 8392 7880 8444 7886
rect 7932 7822 7984 7828
rect 8036 7840 8392 7868
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7852 6322 7880 6598
rect 8036 6322 8064 7840
rect 8392 7822 8444 7828
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8128 6322 8156 7346
rect 8496 6322 8524 9318
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8588 7886 8616 8502
rect 9324 8498 9352 9318
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8588 6662 8616 7822
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8036 5914 8064 6258
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8588 5778 8616 6122
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8680 5710 8708 6122
rect 9218 5808 9274 5817
rect 9218 5743 9220 5752
rect 9272 5743 9274 5752
rect 9220 5714 9272 5720
rect 7932 5704 7984 5710
rect 7668 5664 7932 5692
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 7392 5098 7420 5646
rect 7668 5234 7696 5664
rect 7932 5646 7984 5652
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 7760 5234 7788 5510
rect 8312 5234 8340 5510
rect 8680 5370 8708 5646
rect 9416 5624 9444 10202
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9508 9382 9536 9930
rect 9600 9586 9628 12310
rect 9784 12238 9812 12854
rect 10244 12434 10272 13874
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10612 13190 10640 13738
rect 10704 13394 10732 14010
rect 10796 13802 10824 14350
rect 10980 14074 11008 14418
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10152 12406 10272 12434
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9600 9450 9628 9522
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9876 7274 9904 7822
rect 9968 7546 9996 8366
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9324 5596 9444 5624
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 7380 5092 7432 5098
rect 7380 5034 7432 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4080 3058 4108 4014
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 940 3052 992 3058
rect 940 2994 992 3000
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 952 2825 980 2994
rect 4250 2952 4306 2961
rect 4250 2887 4252 2896
rect 4304 2887 4306 2896
rect 4252 2858 4304 2864
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5920 2650 5948 4082
rect 9140 2650 9168 4082
rect 9324 4078 9352 5596
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9692 5234 9720 5510
rect 9876 5370 9904 5510
rect 9968 5370 9996 5646
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 10152 4826 10180 12406
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10336 12102 10364 12310
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10336 11694 10364 12038
rect 10428 11762 10456 13126
rect 10888 12850 10916 13670
rect 10980 13462 11008 14010
rect 11532 13870 11560 14282
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11520 13864 11572 13870
rect 11518 13832 11520 13841
rect 11572 13832 11574 13841
rect 11518 13767 11574 13776
rect 10968 13456 11020 13462
rect 10968 13398 11020 13404
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11072 12850 11100 13262
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10888 12306 10916 12786
rect 11624 12442 11652 13874
rect 11716 13870 11744 14486
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11808 13870 11836 14214
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11808 13394 11836 13806
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11900 13326 11928 14214
rect 12084 14074 12112 14350
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12084 13802 12112 14010
rect 12072 13796 12124 13802
rect 12072 13738 12124 13744
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 12176 12714 12204 15302
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12360 13938 12388 14214
rect 12544 14006 12572 14282
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 11440 12238 11468 12378
rect 11794 12336 11850 12345
rect 11794 12271 11796 12280
rect 11848 12271 11850 12280
rect 11796 12242 11848 12248
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 10520 11762 10548 12174
rect 11702 11928 11758 11937
rect 11702 11863 11704 11872
rect 11756 11863 11758 11872
rect 11704 11834 11756 11840
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10336 11150 10364 11630
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10428 11082 10456 11698
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 11348 11218 11376 11562
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11624 11218 11652 11494
rect 11808 11286 11836 12242
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10322 10704 10378 10713
rect 10322 10639 10324 10648
rect 10376 10639 10378 10648
rect 10324 10610 10376 10616
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10506 9616 10562 9625
rect 10506 9551 10508 9560
rect 10560 9551 10562 9560
rect 10784 9580 10836 9586
rect 10508 9522 10560 9528
rect 10784 9522 10836 9528
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10428 8634 10456 8910
rect 10520 8906 10548 9522
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10796 7886 10824 9522
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10336 7546 10364 7822
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10244 7002 10272 7346
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10520 6458 10548 7346
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5030 10272 6054
rect 10888 5914 10916 9522
rect 10980 9178 11008 10542
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 9178 11376 9318
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11348 8974 11376 9114
rect 11532 9042 11560 9522
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11624 8974 11652 9930
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11428 8968 11480 8974
rect 11612 8968 11664 8974
rect 11428 8910 11480 8916
rect 11610 8936 11612 8945
rect 11664 8936 11666 8945
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 6322 11100 6734
rect 11348 6322 11376 8910
rect 11440 8090 11468 8910
rect 11610 8871 11666 8880
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11808 7546 11836 11086
rect 11900 9994 11928 12106
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11992 10606 12020 11494
rect 12084 11354 12112 11494
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 12084 9722 12112 9862
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11900 9110 11928 9454
rect 12176 9110 12204 12650
rect 12360 11898 12388 13738
rect 12820 12434 12848 37198
rect 13556 37126 13584 39280
rect 16408 37126 16436 39358
rect 19338 39358 19656 39386
rect 19338 39280 19394 39358
rect 17040 37324 17092 37330
rect 17040 37266 17092 37272
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 16396 37120 16448 37126
rect 16396 37062 16448 37068
rect 17052 36854 17080 37266
rect 19628 37262 19656 39358
rect 22558 39358 22968 39386
rect 22558 39280 22614 39358
rect 21272 37460 21324 37466
rect 21272 37402 21324 37408
rect 17868 37256 17920 37262
rect 17868 37198 17920 37204
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19616 37256 19668 37262
rect 19616 37198 19668 37204
rect 17224 37188 17276 37194
rect 17224 37130 17276 37136
rect 17040 36848 17092 36854
rect 17040 36790 17092 36796
rect 16672 36780 16724 36786
rect 16672 36722 16724 36728
rect 16120 36576 16172 36582
rect 16120 36518 16172 36524
rect 16132 36174 16160 36518
rect 16120 36168 16172 36174
rect 16120 36110 16172 36116
rect 16684 35834 16712 36722
rect 17236 36378 17264 37130
rect 17408 36712 17460 36718
rect 17408 36654 17460 36660
rect 17224 36372 17276 36378
rect 17224 36314 17276 36320
rect 17236 35834 17264 36314
rect 17316 36168 17368 36174
rect 17316 36110 17368 36116
rect 16672 35828 16724 35834
rect 16672 35770 16724 35776
rect 17224 35828 17276 35834
rect 17224 35770 17276 35776
rect 16948 35692 17000 35698
rect 16948 35634 17000 35640
rect 12900 35012 12952 35018
rect 12900 34954 12952 34960
rect 12912 33998 12940 34954
rect 13820 34944 13872 34950
rect 13820 34886 13872 34892
rect 14556 34944 14608 34950
rect 14556 34886 14608 34892
rect 15568 34944 15620 34950
rect 15568 34886 15620 34892
rect 13728 34604 13780 34610
rect 13728 34546 13780 34552
rect 12992 34400 13044 34406
rect 12992 34342 13044 34348
rect 13004 34066 13032 34342
rect 13740 34202 13768 34546
rect 13728 34196 13780 34202
rect 13728 34138 13780 34144
rect 12992 34060 13044 34066
rect 12992 34002 13044 34008
rect 12900 33992 12952 33998
rect 12900 33934 12952 33940
rect 12900 32836 12952 32842
rect 12900 32778 12952 32784
rect 12912 31890 12940 32778
rect 13004 32366 13032 34002
rect 13832 33998 13860 34886
rect 14568 34746 14596 34886
rect 14004 34740 14056 34746
rect 14004 34682 14056 34688
rect 14556 34740 14608 34746
rect 14556 34682 14608 34688
rect 13084 33992 13136 33998
rect 13084 33934 13136 33940
rect 13820 33992 13872 33998
rect 13820 33934 13872 33940
rect 12992 32360 13044 32366
rect 12992 32302 13044 32308
rect 12992 32224 13044 32230
rect 12992 32166 13044 32172
rect 13004 31890 13032 32166
rect 12900 31884 12952 31890
rect 12900 31826 12952 31832
rect 12992 31884 13044 31890
rect 12992 31826 13044 31832
rect 12912 28082 12940 31826
rect 13096 31754 13124 33934
rect 13176 32768 13228 32774
rect 13176 32710 13228 32716
rect 13188 31822 13216 32710
rect 13820 32564 13872 32570
rect 13820 32506 13872 32512
rect 13268 32224 13320 32230
rect 13268 32166 13320 32172
rect 13280 32026 13308 32166
rect 13268 32020 13320 32026
rect 13268 31962 13320 31968
rect 13176 31816 13228 31822
rect 13176 31758 13228 31764
rect 13004 31726 13124 31754
rect 13004 30258 13032 31726
rect 13176 31680 13228 31686
rect 13280 31634 13308 31962
rect 13832 31929 13860 32506
rect 14016 32366 14044 34682
rect 14096 34672 14148 34678
rect 14096 34614 14148 34620
rect 14108 33998 14136 34614
rect 14096 33992 14148 33998
rect 14096 33934 14148 33940
rect 14372 33924 14424 33930
rect 14372 33866 14424 33872
rect 14384 33658 14412 33866
rect 15200 33856 15252 33862
rect 15200 33798 15252 33804
rect 14372 33652 14424 33658
rect 14372 33594 14424 33600
rect 14464 33516 14516 33522
rect 14464 33458 14516 33464
rect 14186 33144 14242 33153
rect 14476 33114 14504 33458
rect 14186 33079 14188 33088
rect 14240 33079 14242 33088
rect 14464 33108 14516 33114
rect 14188 33050 14240 33056
rect 14464 33050 14516 33056
rect 15212 32910 15240 33798
rect 15200 32904 15252 32910
rect 15200 32846 15252 32852
rect 15476 32904 15528 32910
rect 15580 32858 15608 34886
rect 16856 34604 16908 34610
rect 16856 34546 16908 34552
rect 16672 34400 16724 34406
rect 16672 34342 16724 34348
rect 16684 34066 16712 34342
rect 16868 34202 16896 34546
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 16672 34060 16724 34066
rect 16672 34002 16724 34008
rect 15528 32852 15608 32858
rect 15476 32846 15608 32852
rect 15212 32570 15240 32846
rect 15488 32830 15608 32846
rect 14280 32564 14332 32570
rect 14280 32506 14332 32512
rect 15200 32564 15252 32570
rect 15200 32506 15252 32512
rect 14004 32360 14056 32366
rect 14004 32302 14056 32308
rect 13818 31920 13874 31929
rect 14016 31890 14044 32302
rect 14292 31890 14320 32506
rect 15476 32496 15528 32502
rect 15304 32456 15476 32484
rect 15304 32450 15332 32456
rect 14740 32428 14792 32434
rect 14740 32370 14792 32376
rect 15120 32422 15332 32450
rect 15476 32438 15528 32444
rect 14648 32360 14700 32366
rect 14648 32302 14700 32308
rect 13818 31855 13874 31864
rect 14004 31884 14056 31890
rect 14004 31826 14056 31832
rect 14280 31884 14332 31890
rect 14280 31826 14332 31832
rect 14660 31770 14688 32302
rect 14752 32042 14780 32370
rect 14752 32026 14872 32042
rect 14740 32020 14872 32026
rect 14792 32014 14872 32020
rect 14740 31962 14792 31968
rect 14738 31920 14794 31929
rect 14844 31890 14872 32014
rect 14738 31855 14740 31864
rect 14792 31855 14794 31864
rect 14832 31884 14884 31890
rect 14740 31826 14792 31832
rect 14832 31826 14884 31832
rect 15016 31816 15068 31822
rect 14660 31764 15016 31770
rect 14660 31758 15068 31764
rect 14660 31742 15056 31758
rect 15120 31686 15148 32422
rect 15580 32314 15608 32830
rect 16028 32836 16080 32842
rect 16028 32778 16080 32784
rect 16212 32836 16264 32842
rect 16212 32778 16264 32784
rect 15488 32286 15608 32314
rect 15292 31816 15344 31822
rect 15290 31784 15292 31793
rect 15344 31784 15346 31793
rect 15290 31719 15346 31728
rect 13228 31628 13308 31634
rect 13176 31622 13308 31628
rect 15108 31680 15160 31686
rect 15108 31622 15160 31628
rect 13188 31606 13308 31622
rect 15488 30734 15516 32286
rect 15568 32224 15620 32230
rect 15568 32166 15620 32172
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 13360 30592 13412 30598
rect 13360 30534 13412 30540
rect 14096 30592 14148 30598
rect 14096 30534 14148 30540
rect 13372 30394 13400 30534
rect 13360 30388 13412 30394
rect 13360 30330 13412 30336
rect 12992 30252 13044 30258
rect 12992 30194 13044 30200
rect 13004 29510 13032 30194
rect 13268 30184 13320 30190
rect 13268 30126 13320 30132
rect 13280 29782 13308 30126
rect 13268 29776 13320 29782
rect 13268 29718 13320 29724
rect 12992 29504 13044 29510
rect 12992 29446 13044 29452
rect 12900 28076 12952 28082
rect 12900 28018 12952 28024
rect 12912 26586 12940 28018
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12912 24274 12940 26522
rect 13004 26042 13032 29446
rect 13372 28422 13400 30330
rect 14108 30326 14136 30534
rect 14096 30320 14148 30326
rect 14096 30262 14148 30268
rect 14292 29850 14320 30670
rect 15488 30054 15516 30670
rect 14556 30048 14608 30054
rect 14556 29990 14608 29996
rect 15476 30048 15528 30054
rect 15476 29990 15528 29996
rect 14280 29844 14332 29850
rect 14280 29786 14332 29792
rect 14568 29646 14596 29990
rect 14556 29640 14608 29646
rect 14556 29582 14608 29588
rect 14372 28688 14424 28694
rect 14372 28630 14424 28636
rect 14096 28620 14148 28626
rect 14096 28562 14148 28568
rect 13912 28552 13964 28558
rect 13912 28494 13964 28500
rect 13360 28416 13412 28422
rect 13360 28358 13412 28364
rect 13924 27946 13952 28494
rect 14108 28014 14136 28562
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 14292 28082 14320 28358
rect 14384 28218 14412 28630
rect 14464 28620 14516 28626
rect 14568 28608 14596 29582
rect 14516 28580 14596 28608
rect 14464 28562 14516 28568
rect 15016 28552 15068 28558
rect 15016 28494 15068 28500
rect 15028 28422 15056 28494
rect 15016 28416 15068 28422
rect 15016 28358 15068 28364
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 14372 28212 14424 28218
rect 14372 28154 14424 28160
rect 14384 28082 14412 28154
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 14372 28076 14424 28082
rect 14372 28018 14424 28024
rect 14096 28008 14148 28014
rect 14096 27950 14148 27956
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 13912 27940 13964 27946
rect 13912 27882 13964 27888
rect 14004 27940 14056 27946
rect 14004 27882 14056 27888
rect 13636 27396 13688 27402
rect 13636 27338 13688 27344
rect 13648 26926 13676 27338
rect 13924 27146 13952 27882
rect 14016 27674 14044 27882
rect 14004 27668 14056 27674
rect 14004 27610 14056 27616
rect 14568 27538 14596 27950
rect 15200 27872 15252 27878
rect 15200 27814 15252 27820
rect 14556 27532 14608 27538
rect 14556 27474 14608 27480
rect 14280 27464 14332 27470
rect 14280 27406 14332 27412
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 13924 27130 14044 27146
rect 13924 27124 14056 27130
rect 13924 27118 14004 27124
rect 14004 27066 14056 27072
rect 14108 27062 14136 27270
rect 14096 27056 14148 27062
rect 14096 26998 14148 27004
rect 13636 26920 13688 26926
rect 13636 26862 13688 26868
rect 14292 26586 14320 27406
rect 14740 27328 14792 27334
rect 14740 27270 14792 27276
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14476 26382 14504 27066
rect 14648 26852 14700 26858
rect 14648 26794 14700 26800
rect 14660 26450 14688 26794
rect 14648 26444 14700 26450
rect 14648 26386 14700 26392
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 13360 26308 13412 26314
rect 13360 26250 13412 26256
rect 13176 26240 13228 26246
rect 13176 26182 13228 26188
rect 12992 26036 13044 26042
rect 12992 25978 13044 25984
rect 13188 25770 13216 26182
rect 13372 25906 13400 26250
rect 13544 26036 13596 26042
rect 13544 25978 13596 25984
rect 13360 25900 13412 25906
rect 13360 25842 13412 25848
rect 13176 25764 13228 25770
rect 13176 25706 13228 25712
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12900 24268 12952 24274
rect 12900 24210 12952 24216
rect 13004 24206 13032 24550
rect 13084 24268 13136 24274
rect 13084 24210 13136 24216
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 13004 23730 13032 24142
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12900 23656 12952 23662
rect 12900 23598 12952 23604
rect 12912 22574 12940 23598
rect 12900 22568 12952 22574
rect 12900 22510 12952 22516
rect 13096 21962 13124 24210
rect 13188 23662 13216 25706
rect 13176 23656 13228 23662
rect 13176 23598 13228 23604
rect 13188 23322 13216 23598
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 13176 22500 13228 22506
rect 13176 22442 13228 22448
rect 13084 21956 13136 21962
rect 13084 21898 13136 21904
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12912 21554 12940 21830
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 13096 19514 13124 21898
rect 13188 21729 13216 22442
rect 13372 22094 13400 25842
rect 13556 25702 13584 25978
rect 14752 25838 14780 27270
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 15016 26988 15068 26994
rect 15016 26930 15068 26936
rect 14740 25832 14792 25838
rect 14924 25832 14976 25838
rect 14740 25774 14792 25780
rect 14922 25800 14924 25809
rect 14976 25800 14978 25809
rect 14922 25735 14978 25744
rect 13544 25696 13596 25702
rect 13544 25638 13596 25644
rect 14648 25696 14700 25702
rect 14648 25638 14700 25644
rect 13452 23316 13504 23322
rect 13452 23258 13504 23264
rect 13464 22642 13492 23258
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13372 22066 13492 22094
rect 13464 21894 13492 22066
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13174 21720 13230 21729
rect 13174 21655 13230 21664
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12912 18970 12940 19314
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 12912 18290 12940 18906
rect 13096 18290 13124 19246
rect 13188 18902 13216 21655
rect 13280 19802 13308 21830
rect 13452 20868 13504 20874
rect 13452 20810 13504 20816
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13372 20058 13400 20402
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13464 19922 13492 20810
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 13280 19774 13400 19802
rect 13176 18896 13228 18902
rect 13176 18838 13228 18844
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13096 17746 13124 18226
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 13188 17338 13216 18158
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13188 16590 13216 17274
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13372 16454 13400 19774
rect 13452 19304 13504 19310
rect 13450 19272 13452 19281
rect 13504 19272 13506 19281
rect 13450 19207 13506 19216
rect 13556 17610 13584 25638
rect 14464 25152 14516 25158
rect 14464 25094 14516 25100
rect 14476 24818 14504 25094
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14660 24750 14688 25638
rect 14936 25294 14964 25735
rect 14924 25288 14976 25294
rect 14924 25230 14976 25236
rect 14648 24744 14700 24750
rect 14648 24686 14700 24692
rect 14832 24744 14884 24750
rect 14832 24686 14884 24692
rect 14004 24676 14056 24682
rect 14004 24618 14056 24624
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13832 23730 13860 23802
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13636 23656 13688 23662
rect 13688 23604 13860 23610
rect 13636 23598 13860 23604
rect 13648 23582 13860 23598
rect 13832 23202 13860 23582
rect 13648 23174 13860 23202
rect 13648 22642 13676 23174
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 13648 22030 13676 22578
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13740 22273 13768 22510
rect 13726 22264 13782 22273
rect 13726 22199 13782 22208
rect 13636 22024 13688 22030
rect 13636 21966 13688 21972
rect 13740 21468 13768 22199
rect 13648 21440 13768 21468
rect 13648 18766 13676 21440
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13740 20913 13768 21286
rect 13726 20904 13782 20913
rect 13726 20839 13782 20848
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13740 19718 13768 20198
rect 13832 19854 13860 20198
rect 13924 20058 13952 20742
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13636 18148 13688 18154
rect 13636 18090 13688 18096
rect 13648 18057 13676 18090
rect 13634 18048 13690 18057
rect 13634 17983 13690 17992
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 17202 13492 17478
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 15434 13400 16390
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13740 14414 13768 19654
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13832 18290 13860 19246
rect 13924 18290 13952 19246
rect 14016 18426 14044 24618
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13832 16250 13860 18226
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13832 15502 13860 16186
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 14108 15026 14136 24550
rect 14476 23866 14504 24618
rect 14844 24410 14872 24686
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 15028 23730 15056 26930
rect 15120 26790 15148 27066
rect 15108 26784 15160 26790
rect 15108 26726 15160 26732
rect 15120 25906 15148 26726
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 15016 23724 15068 23730
rect 15016 23666 15068 23672
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14292 22710 14320 22918
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14280 22500 14332 22506
rect 14280 22442 14332 22448
rect 14292 22030 14320 22442
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14188 21412 14240 21418
rect 14188 21354 14240 21360
rect 14200 21010 14228 21354
rect 14188 21004 14240 21010
rect 14188 20946 14240 20952
rect 14292 20942 14320 21422
rect 14384 21078 14412 22374
rect 14476 22234 14504 23054
rect 15028 22642 15056 23666
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14752 22098 14780 22170
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14752 21622 14780 22034
rect 15028 21894 15056 22578
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 15028 21690 15056 21830
rect 15016 21684 15068 21690
rect 15016 21626 15068 21632
rect 14740 21616 14792 21622
rect 14740 21558 14792 21564
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14568 20874 14596 21082
rect 14924 20936 14976 20942
rect 15028 20924 15056 21626
rect 14976 20896 15056 20924
rect 14924 20878 14976 20884
rect 14556 20868 14608 20874
rect 14556 20810 14608 20816
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14384 19514 14412 20402
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14752 19922 14780 20334
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14844 19854 14872 20742
rect 15212 20602 15240 27814
rect 15304 25226 15332 28358
rect 15476 27872 15528 27878
rect 15476 27814 15528 27820
rect 15488 27470 15516 27814
rect 15476 27464 15528 27470
rect 15476 27406 15528 27412
rect 15580 27334 15608 32166
rect 15752 31952 15804 31958
rect 15752 31894 15804 31900
rect 15568 27328 15620 27334
rect 15568 27270 15620 27276
rect 15292 25220 15344 25226
rect 15292 25162 15344 25168
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15672 23322 15700 23666
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 15304 20602 15332 20810
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15488 20466 15516 21286
rect 15764 20942 15792 31894
rect 16040 31822 16068 32778
rect 16224 32502 16252 32778
rect 16856 32768 16908 32774
rect 16856 32710 16908 32716
rect 16868 32570 16896 32710
rect 16856 32564 16908 32570
rect 16856 32506 16908 32512
rect 16212 32496 16264 32502
rect 16132 32456 16212 32484
rect 16028 31816 16080 31822
rect 16028 31758 16080 31764
rect 16132 28218 16160 32456
rect 16212 32438 16264 32444
rect 16304 32360 16356 32366
rect 16304 32302 16356 32308
rect 16212 32224 16264 32230
rect 16212 32166 16264 32172
rect 16224 31822 16252 32166
rect 16316 31822 16344 32302
rect 16684 32298 16896 32314
rect 16684 32292 16908 32298
rect 16684 32286 16856 32292
rect 16684 32230 16712 32286
rect 16856 32234 16908 32240
rect 16672 32224 16724 32230
rect 16672 32166 16724 32172
rect 16212 31816 16264 31822
rect 16212 31758 16264 31764
rect 16304 31816 16356 31822
rect 16304 31758 16356 31764
rect 16960 31754 16988 35634
rect 17132 35080 17184 35086
rect 17132 35022 17184 35028
rect 17040 35012 17092 35018
rect 17040 34954 17092 34960
rect 17052 34746 17080 34954
rect 17040 34740 17092 34746
rect 17040 34682 17092 34688
rect 17144 34542 17172 35022
rect 17328 34950 17356 36110
rect 17420 36038 17448 36654
rect 17880 36174 17908 37198
rect 17960 36780 18012 36786
rect 17960 36722 18012 36728
rect 19156 36780 19208 36786
rect 19156 36722 19208 36728
rect 17972 36378 18000 36722
rect 18328 36576 18380 36582
rect 18328 36518 18380 36524
rect 17960 36372 18012 36378
rect 17960 36314 18012 36320
rect 17868 36168 17920 36174
rect 17868 36110 17920 36116
rect 18340 36038 18368 36518
rect 19168 36378 19196 36722
rect 19248 36712 19300 36718
rect 19248 36654 19300 36660
rect 19156 36372 19208 36378
rect 19156 36314 19208 36320
rect 19064 36236 19116 36242
rect 19064 36178 19116 36184
rect 18420 36168 18472 36174
rect 18420 36110 18472 36116
rect 17408 36032 17460 36038
rect 17408 35974 17460 35980
rect 18328 36032 18380 36038
rect 18328 35974 18380 35980
rect 17316 34944 17368 34950
rect 17316 34886 17368 34892
rect 17328 34542 17356 34886
rect 17132 34536 17184 34542
rect 17132 34478 17184 34484
rect 17316 34536 17368 34542
rect 17316 34478 17368 34484
rect 17420 33522 17448 35974
rect 18328 34740 18380 34746
rect 18328 34682 18380 34688
rect 17684 34536 17736 34542
rect 17684 34478 17736 34484
rect 17696 33930 17724 34478
rect 17868 34128 17920 34134
rect 17868 34070 17920 34076
rect 17684 33924 17736 33930
rect 17684 33866 17736 33872
rect 17316 33516 17368 33522
rect 17316 33458 17368 33464
rect 17408 33516 17460 33522
rect 17408 33458 17460 33464
rect 17328 33114 17356 33458
rect 17316 33108 17368 33114
rect 17316 33050 17368 33056
rect 17040 33040 17092 33046
rect 17040 32982 17092 32988
rect 17052 32434 17080 32982
rect 17040 32428 17092 32434
rect 17040 32370 17092 32376
rect 17224 32428 17276 32434
rect 17224 32370 17276 32376
rect 17052 31890 17080 32370
rect 17236 31890 17264 32370
rect 17500 32292 17552 32298
rect 17500 32234 17552 32240
rect 17040 31884 17092 31890
rect 17040 31826 17092 31832
rect 17224 31884 17276 31890
rect 17224 31826 17276 31832
rect 16960 31726 17080 31754
rect 16856 30252 16908 30258
rect 16856 30194 16908 30200
rect 16580 30048 16632 30054
rect 16580 29990 16632 29996
rect 16592 29714 16620 29990
rect 16868 29850 16896 30194
rect 16856 29844 16908 29850
rect 16856 29786 16908 29792
rect 16580 29708 16632 29714
rect 16580 29650 16632 29656
rect 16592 28694 16620 29650
rect 16948 29572 17000 29578
rect 16948 29514 17000 29520
rect 16580 28688 16632 28694
rect 16580 28630 16632 28636
rect 16960 28626 16988 29514
rect 16948 28620 17000 28626
rect 16948 28562 17000 28568
rect 16120 28212 16172 28218
rect 16120 28154 16172 28160
rect 16132 26586 16160 28154
rect 16488 28144 16540 28150
rect 16488 28086 16540 28092
rect 16500 27946 16528 28086
rect 16960 28082 16988 28562
rect 16580 28076 16632 28082
rect 16580 28018 16632 28024
rect 16948 28076 17000 28082
rect 16948 28018 17000 28024
rect 16488 27940 16540 27946
rect 16488 27882 16540 27888
rect 16592 27334 16620 28018
rect 16672 27872 16724 27878
rect 16672 27814 16724 27820
rect 16684 27674 16712 27814
rect 16672 27668 16724 27674
rect 16672 27610 16724 27616
rect 16580 27328 16632 27334
rect 16580 27270 16632 27276
rect 16120 26580 16172 26586
rect 16120 26522 16172 26528
rect 15844 25900 15896 25906
rect 15844 25842 15896 25848
rect 15856 25226 15884 25842
rect 15844 25220 15896 25226
rect 15844 25162 15896 25168
rect 16132 23186 16160 26522
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 16672 25696 16724 25702
rect 16672 25638 16724 25644
rect 16684 25294 16712 25638
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 16488 24676 16540 24682
rect 16488 24618 16540 24624
rect 16500 24206 16528 24618
rect 16672 24608 16724 24614
rect 16672 24550 16724 24556
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 16224 23526 16252 23598
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 16120 23180 16172 23186
rect 16120 23122 16172 23128
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 16040 21049 16068 21422
rect 16132 21185 16160 23122
rect 16224 22982 16252 23462
rect 16500 23186 16528 24142
rect 16488 23180 16540 23186
rect 16488 23122 16540 23128
rect 16488 23044 16540 23050
rect 16488 22986 16540 22992
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 16224 22098 16252 22918
rect 16500 22166 16528 22986
rect 16488 22160 16540 22166
rect 16488 22102 16540 22108
rect 16212 22092 16264 22098
rect 16212 22034 16264 22040
rect 16500 21486 16528 22102
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16118 21176 16174 21185
rect 16118 21111 16174 21120
rect 16026 21040 16082 21049
rect 16026 20975 16082 20984
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 14292 19009 14320 19246
rect 14278 19000 14334 19009
rect 14278 18935 14334 18944
rect 14292 18698 14320 18935
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14462 18320 14518 18329
rect 14462 18255 14518 18264
rect 14476 18222 14504 18255
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14556 18080 14608 18086
rect 14554 18048 14556 18057
rect 14608 18048 14610 18057
rect 14554 17983 14610 17992
rect 14660 17882 14688 19246
rect 14844 18834 14872 19382
rect 15120 19310 15148 19790
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15212 19174 15240 19858
rect 16132 19854 16160 21111
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14568 17338 14596 17682
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13176 14000 13228 14006
rect 13174 13968 13176 13977
rect 13228 13968 13230 13977
rect 13280 13938 13308 14214
rect 13740 13938 13768 14214
rect 13924 13938 13952 14418
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 14074 14136 14350
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14188 14000 14240 14006
rect 14186 13968 14188 13977
rect 14240 13968 14242 13977
rect 13174 13903 13230 13912
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13912 13932 13964 13938
rect 14096 13932 14148 13938
rect 13964 13892 14096 13920
rect 13912 13874 13964 13880
rect 14568 13938 14596 14214
rect 14186 13903 14242 13912
rect 14556 13932 14608 13938
rect 14096 13874 14148 13880
rect 14556 13874 14608 13880
rect 13280 13841 13308 13874
rect 13266 13832 13322 13841
rect 13266 13767 13322 13776
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 12820 12406 12940 12434
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12544 12050 12572 12106
rect 12452 12022 12572 12050
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 11992 8906 12020 9046
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 12268 8786 12296 11834
rect 12452 11762 12480 12022
rect 12636 11898 12664 12174
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12360 10266 12388 10474
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12452 10062 12480 11562
rect 12544 11354 12572 11698
rect 12820 11694 12848 11834
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12820 11150 12848 11630
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12544 9654 12572 10202
rect 12820 9926 12848 11086
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 12348 8832 12400 8838
rect 12268 8780 12348 8786
rect 12268 8774 12400 8780
rect 12268 8758 12388 8774
rect 12452 8430 12480 8842
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12544 8362 12572 9590
rect 12820 9586 12848 9862
rect 12912 9704 12940 12406
rect 13096 11762 13124 13330
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13280 10606 13308 13767
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 13924 12850 13952 13670
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13464 10470 13492 12106
rect 13740 12102 13768 12786
rect 14016 12782 14044 13670
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14016 12646 14044 12718
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14002 12336 14058 12345
rect 14108 12288 14136 12718
rect 14058 12280 14136 12288
rect 14002 12271 14136 12280
rect 14016 12260 14136 12271
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13464 10130 13492 10406
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13372 10010 13400 10066
rect 13556 10010 13584 10610
rect 13648 10198 13676 10678
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13636 10056 13688 10062
rect 13372 10004 13636 10010
rect 13372 9998 13688 10004
rect 13372 9982 13676 9998
rect 12912 9676 13124 9704
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12636 8906 12664 9522
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12898 8936 12954 8945
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12636 8634 12664 8842
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12622 8528 12678 8537
rect 12622 8463 12624 8472
rect 12676 8463 12678 8472
rect 12624 8434 12676 8440
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11900 7886 11928 8230
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12176 7954 12204 8026
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 12544 7750 12572 8298
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 12544 7410 12572 7686
rect 12728 7410 12756 8910
rect 12898 8871 12954 8880
rect 12912 8634 12940 8871
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12820 7546 12848 8434
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 11992 7002 12020 7346
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 11072 5710 11100 6258
rect 11808 6254 11836 6870
rect 12728 6866 12756 7346
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11808 5914 11836 6190
rect 12820 5914 12848 7142
rect 13004 5914 13032 9522
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11072 5234 11100 5646
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11808 5030 11836 5850
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12268 5098 12296 5646
rect 12452 5370 12480 5646
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12544 5234 12572 5714
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 12636 5370 12664 5578
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 13096 5166 13124 9676
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13188 7818 13216 9114
rect 13648 8362 13676 9982
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13556 7954 13584 8230
rect 13648 7954 13676 8298
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13740 7886 13768 8434
rect 13832 8090 13860 10406
rect 13924 10266 13952 11630
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14016 8634 14044 12260
rect 14096 12164 14148 12170
rect 14096 12106 14148 12112
rect 14108 11762 14136 12106
rect 14292 11898 14320 12718
rect 14660 12434 14688 17818
rect 14844 17202 14872 18770
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 15212 18426 15240 18634
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15396 18290 15424 19654
rect 16040 19514 16068 19722
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 15384 18284 15436 18290
rect 15384 18226 15436 18232
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14844 16658 14872 17138
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15304 16250 15332 16458
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14844 14414 14872 14758
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 15212 13954 15240 15030
rect 15488 14414 15516 15846
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15488 14074 15516 14350
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15212 13926 15332 13954
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14936 12850 14964 13194
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 15028 12850 15056 13126
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 14568 12406 14688 12434
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14108 10810 14136 11018
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14292 9178 14320 9998
rect 14568 9654 14596 12406
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14936 11150 14964 12038
rect 15212 11150 15240 13806
rect 15304 13394 15332 13926
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15304 13190 15332 13330
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15304 12102 15332 12786
rect 15396 12238 15424 12854
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 15764 12714 15792 12786
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 14660 10810 14688 11086
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15028 10810 15056 10950
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13832 7410 13860 8026
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 14200 7342 14228 8366
rect 14476 7886 14504 9114
rect 14568 8430 14596 9590
rect 14660 8498 14688 10610
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14936 10266 14964 10542
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 15028 10130 15056 10746
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14936 9722 14964 9998
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14844 9178 14872 9522
rect 15580 9518 15608 11698
rect 15672 9926 15700 12582
rect 15764 12238 15792 12650
rect 16132 12238 16160 12786
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16132 11762 16160 12038
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 16224 9625 16252 19450
rect 16316 18970 16344 19654
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16316 18290 16344 18906
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 16500 18426 16528 18838
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16488 18420 16540 18426
rect 16488 18362 16540 18368
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16408 16794 16436 16934
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 16408 16658 16436 16730
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16408 16114 16436 16390
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16500 15366 16528 18362
rect 16592 18222 16620 18702
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 15162 16528 15302
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16592 15026 16620 17138
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16316 13938 16344 14962
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16316 13394 16344 13874
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16408 10810 16436 13126
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16210 9616 16266 9625
rect 16210 9551 16266 9560
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 16224 8906 16252 9551
rect 16500 8906 16528 14214
rect 16684 13530 16712 24550
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16776 22438 16804 23598
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16776 22098 16804 22374
rect 16764 22092 16816 22098
rect 16764 22034 16816 22040
rect 16868 21978 16896 26250
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16960 23594 16988 24142
rect 16948 23588 17000 23594
rect 16948 23530 17000 23536
rect 16948 22092 17000 22098
rect 16948 22034 17000 22040
rect 16776 21950 16896 21978
rect 16776 21049 16804 21950
rect 16854 21856 16910 21865
rect 16854 21791 16910 21800
rect 16868 21554 16896 21791
rect 16960 21729 16988 22034
rect 17052 21978 17080 31726
rect 17224 30592 17276 30598
rect 17224 30534 17276 30540
rect 17132 30252 17184 30258
rect 17132 30194 17184 30200
rect 17144 29850 17172 30194
rect 17236 30190 17264 30534
rect 17224 30184 17276 30190
rect 17224 30126 17276 30132
rect 17132 29844 17184 29850
rect 17132 29786 17184 29792
rect 17316 29504 17368 29510
rect 17316 29446 17368 29452
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 17144 28014 17172 28494
rect 17132 28008 17184 28014
rect 17132 27950 17184 27956
rect 17144 27674 17172 27950
rect 17132 27668 17184 27674
rect 17132 27610 17184 27616
rect 17328 26450 17356 29446
rect 17512 28762 17540 32234
rect 17696 29510 17724 33866
rect 17880 32450 17908 34070
rect 18340 34066 18368 34682
rect 18328 34060 18380 34066
rect 18328 34002 18380 34008
rect 18052 32972 18104 32978
rect 18052 32914 18104 32920
rect 17960 32904 18012 32910
rect 17960 32846 18012 32852
rect 17972 32570 18000 32846
rect 18064 32570 18092 32914
rect 18328 32768 18380 32774
rect 18328 32710 18380 32716
rect 17960 32564 18012 32570
rect 17960 32506 18012 32512
rect 18052 32564 18104 32570
rect 18052 32506 18104 32512
rect 17880 32434 18000 32450
rect 17880 32428 18012 32434
rect 17880 32422 17960 32428
rect 17960 32370 18012 32376
rect 17776 31952 17828 31958
rect 17774 31920 17776 31929
rect 17828 31920 17830 31929
rect 17972 31890 18000 32370
rect 18052 32360 18104 32366
rect 18052 32302 18104 32308
rect 18064 31890 18092 32302
rect 17774 31855 17830 31864
rect 17960 31884 18012 31890
rect 17960 31826 18012 31832
rect 18052 31884 18104 31890
rect 18052 31826 18104 31832
rect 18236 31816 18288 31822
rect 18234 31784 18236 31793
rect 18288 31784 18290 31793
rect 18234 31719 18290 31728
rect 17868 30048 17920 30054
rect 17868 29990 17920 29996
rect 17880 29594 17908 29990
rect 17788 29578 17908 29594
rect 17776 29572 17908 29578
rect 17828 29566 17908 29572
rect 17776 29514 17828 29520
rect 17684 29504 17736 29510
rect 17684 29446 17736 29452
rect 17500 28756 17552 28762
rect 17500 28698 17552 28704
rect 17512 28014 17540 28698
rect 17592 28620 17644 28626
rect 17592 28562 17644 28568
rect 17684 28620 17736 28626
rect 17736 28580 17816 28608
rect 17684 28562 17736 28568
rect 17500 28008 17552 28014
rect 17500 27950 17552 27956
rect 17500 27872 17552 27878
rect 17500 27814 17552 27820
rect 17512 27554 17540 27814
rect 17604 27554 17632 28562
rect 17788 28082 17816 28580
rect 17960 28552 18012 28558
rect 17880 28500 17960 28506
rect 17880 28494 18012 28500
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 17880 28478 18000 28494
rect 17880 28082 17908 28478
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 18064 28082 18092 28358
rect 17776 28076 17828 28082
rect 17776 28018 17828 28024
rect 17868 28076 17920 28082
rect 17868 28018 17920 28024
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 17512 27526 17632 27554
rect 17408 27396 17460 27402
rect 17408 27338 17460 27344
rect 17420 26994 17448 27338
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17316 26444 17368 26450
rect 17316 26386 17368 26392
rect 17328 26042 17356 26386
rect 17316 26036 17368 26042
rect 17316 25978 17368 25984
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 17144 24138 17172 25774
rect 17132 24132 17184 24138
rect 17132 24074 17184 24080
rect 17144 22098 17172 24074
rect 17224 23520 17276 23526
rect 17224 23462 17276 23468
rect 17236 22137 17264 23462
rect 17222 22128 17278 22137
rect 17132 22092 17184 22098
rect 17222 22063 17224 22072
rect 17132 22034 17184 22040
rect 17276 22063 17278 22072
rect 17224 22034 17276 22040
rect 17052 21950 17264 21978
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 16946 21720 17002 21729
rect 16946 21655 17002 21664
rect 17052 21554 17080 21830
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 17040 21548 17092 21554
rect 17040 21490 17092 21496
rect 16868 21146 16896 21490
rect 16960 21146 16988 21490
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 17144 21078 17172 21830
rect 17132 21072 17184 21078
rect 16762 21040 16818 21049
rect 16762 20975 16818 20984
rect 16946 21040 17002 21049
rect 17132 21014 17184 21020
rect 16946 20975 17002 20984
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16776 17202 16804 19246
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16868 17610 16896 18158
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16960 16454 16988 20975
rect 17130 20360 17186 20369
rect 17130 20295 17132 20304
rect 17184 20295 17186 20304
rect 17132 20266 17184 20272
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 17052 18873 17080 19246
rect 17038 18864 17094 18873
rect 17038 18799 17040 18808
rect 17092 18799 17094 18808
rect 17040 18770 17092 18776
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 17052 16590 17080 17478
rect 17236 17354 17264 21950
rect 17328 17678 17356 25978
rect 17408 22432 17460 22438
rect 17408 22374 17460 22380
rect 17420 21146 17448 22374
rect 17408 21140 17460 21146
rect 17408 21082 17460 21088
rect 17420 20942 17448 21082
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17406 20496 17462 20505
rect 17406 20431 17408 20440
rect 17460 20431 17462 20440
rect 17408 20402 17460 20408
rect 17512 20346 17540 27526
rect 17592 27396 17644 27402
rect 17592 27338 17644 27344
rect 17604 26586 17632 27338
rect 17880 27334 17908 28018
rect 18156 27878 18184 28494
rect 18236 28008 18288 28014
rect 18236 27950 18288 27956
rect 18144 27872 18196 27878
rect 18144 27814 18196 27820
rect 17868 27328 17920 27334
rect 17868 27270 17920 27276
rect 17684 26920 17736 26926
rect 17684 26862 17736 26868
rect 17592 26580 17644 26586
rect 17592 26522 17644 26528
rect 17696 26314 17724 26862
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 17788 26382 17816 26726
rect 17776 26376 17828 26382
rect 17776 26318 17828 26324
rect 17684 26308 17736 26314
rect 17684 26250 17736 26256
rect 17868 26308 17920 26314
rect 17868 26250 17920 26256
rect 17880 25838 17908 26250
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 17682 25528 17738 25537
rect 17682 25463 17684 25472
rect 17736 25463 17738 25472
rect 17684 25434 17736 25440
rect 17592 24132 17644 24138
rect 17592 24074 17644 24080
rect 17604 23730 17632 24074
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 17590 22264 17646 22273
rect 17590 22199 17646 22208
rect 17604 22098 17632 22199
rect 17592 22092 17644 22098
rect 17592 22034 17644 22040
rect 17590 21176 17646 21185
rect 17590 21111 17646 21120
rect 17604 21010 17632 21111
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17420 20318 17540 20346
rect 17420 19310 17448 20318
rect 17604 20262 17632 20742
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17420 18222 17448 18702
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17144 17326 17264 17354
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16776 15570 16804 15846
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16868 15026 16896 15574
rect 16960 15366 16988 16390
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16776 12986 16804 13194
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16868 11354 16896 12786
rect 16960 12442 16988 15302
rect 17144 12782 17172 17326
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17236 16794 17264 17138
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17316 16516 17368 16522
rect 17420 16504 17448 18158
rect 17368 16476 17448 16504
rect 17316 16458 17368 16464
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17236 14618 17264 15030
rect 17512 15026 17540 20198
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17604 18766 17632 19110
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 17604 18290 17632 18362
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17604 17338 17632 17478
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17604 15570 17632 16050
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17328 14550 17356 14894
rect 17316 14544 17368 14550
rect 17316 14486 17368 14492
rect 17696 13530 17724 25434
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 17972 24410 18000 24754
rect 17960 24404 18012 24410
rect 17960 24346 18012 24352
rect 17868 24336 17920 24342
rect 17868 24278 17920 24284
rect 17880 23866 17908 24278
rect 17776 23860 17828 23866
rect 17776 23802 17828 23808
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 17788 23746 17816 23802
rect 17788 23730 17908 23746
rect 17788 23724 17920 23730
rect 17788 23718 17868 23724
rect 17868 23666 17920 23672
rect 17868 22432 17920 22438
rect 17868 22374 17920 22380
rect 17880 22234 17908 22374
rect 17868 22228 17920 22234
rect 17868 22170 17920 22176
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17788 21146 17816 21626
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 17880 21010 17908 22170
rect 18156 22094 18184 27814
rect 18248 27130 18276 27950
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 18340 25974 18368 32710
rect 18328 25968 18380 25974
rect 18328 25910 18380 25916
rect 18328 25832 18380 25838
rect 18326 25800 18328 25809
rect 18380 25800 18382 25809
rect 18326 25735 18382 25744
rect 18432 22094 18460 36110
rect 19076 35630 19104 36178
rect 19260 35766 19288 36654
rect 19248 35760 19300 35766
rect 19248 35702 19300 35708
rect 19064 35624 19116 35630
rect 19064 35566 19116 35572
rect 18788 35080 18840 35086
rect 18788 35022 18840 35028
rect 18696 34944 18748 34950
rect 18696 34886 18748 34892
rect 18708 34678 18736 34886
rect 18696 34672 18748 34678
rect 18696 34614 18748 34620
rect 18708 33046 18736 34614
rect 18800 34542 18828 35022
rect 18788 34536 18840 34542
rect 18788 34478 18840 34484
rect 18880 33516 18932 33522
rect 18880 33458 18932 33464
rect 18788 33312 18840 33318
rect 18788 33254 18840 33260
rect 18696 33040 18748 33046
rect 18696 32982 18748 32988
rect 18800 32910 18828 33254
rect 18892 33114 18920 33458
rect 18880 33108 18932 33114
rect 18880 33050 18932 33056
rect 18788 32904 18840 32910
rect 18788 32846 18840 32852
rect 18880 32768 18932 32774
rect 18880 32710 18932 32716
rect 18892 32502 18920 32710
rect 18880 32496 18932 32502
rect 18880 32438 18932 32444
rect 18604 32360 18656 32366
rect 18604 32302 18656 32308
rect 18512 31680 18564 31686
rect 18616 31634 18644 32302
rect 18788 31884 18840 31890
rect 18788 31826 18840 31832
rect 18564 31628 18644 31634
rect 18512 31622 18644 31628
rect 18524 31606 18644 31622
rect 18616 28608 18644 31606
rect 18696 28620 18748 28626
rect 18616 28580 18696 28608
rect 18616 28422 18644 28580
rect 18696 28562 18748 28568
rect 18604 28416 18656 28422
rect 18604 28358 18656 28364
rect 18696 27872 18748 27878
rect 18696 27814 18748 27820
rect 18604 27668 18656 27674
rect 18604 27610 18656 27616
rect 18616 27130 18644 27610
rect 18604 27124 18656 27130
rect 18604 27066 18656 27072
rect 18708 26042 18736 27814
rect 18696 26036 18748 26042
rect 18696 25978 18748 25984
rect 18800 25922 18828 31826
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18892 29714 18920 29990
rect 18880 29708 18932 29714
rect 18880 29650 18932 29656
rect 18880 28416 18932 28422
rect 18880 28358 18932 28364
rect 18708 25894 18828 25922
rect 18512 25696 18564 25702
rect 18512 25638 18564 25644
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 18524 24750 18552 25638
rect 18616 24886 18644 25638
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18512 24744 18564 24750
rect 18512 24686 18564 24692
rect 18604 24676 18656 24682
rect 18604 24618 18656 24624
rect 18616 24410 18644 24618
rect 18604 24404 18656 24410
rect 18604 24346 18656 24352
rect 18512 24336 18564 24342
rect 18512 24278 18564 24284
rect 18064 22066 18184 22094
rect 18340 22066 18460 22094
rect 17868 21004 17920 21010
rect 17868 20946 17920 20952
rect 17866 20904 17922 20913
rect 17866 20839 17922 20848
rect 17960 20868 18012 20874
rect 17880 20806 17908 20839
rect 17960 20810 18012 20816
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 17776 20460 17828 20466
rect 17972 20448 18000 20810
rect 17828 20420 18000 20448
rect 17776 20402 17828 20408
rect 17866 20360 17922 20369
rect 17866 20295 17922 20304
rect 17880 20262 17908 20295
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 18064 19174 18092 22066
rect 18144 21412 18196 21418
rect 18144 21354 18196 21360
rect 18156 20806 18184 21354
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 17866 18320 17922 18329
rect 17866 18255 17868 18264
rect 17920 18255 17922 18264
rect 17868 18226 17920 18232
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17776 14340 17828 14346
rect 17776 14282 17828 14288
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16776 10266 16804 10610
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 15212 8498 15240 8774
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 15120 8090 15148 8434
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15304 7886 15332 8774
rect 16040 8634 16068 8774
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16408 8566 16436 8774
rect 16396 8560 16448 8566
rect 16500 8537 16528 8842
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16396 8502 16448 8508
rect 16486 8528 16542 8537
rect 16486 8463 16542 8472
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 14292 7410 14320 7822
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6390 14136 6598
rect 14200 6458 14228 7278
rect 14476 6866 14504 7822
rect 16592 7478 16620 8570
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14476 6390 14504 6666
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14464 6384 14516 6390
rect 14464 6326 14516 6332
rect 15568 6384 15620 6390
rect 15568 6326 15620 6332
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 14568 6186 14596 6258
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14936 5302 14964 5646
rect 15396 5574 15424 6258
rect 15580 5710 15608 6326
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15396 5370 15424 5510
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 14924 5296 14976 5302
rect 14924 5238 14976 5244
rect 15488 5166 15516 5646
rect 15672 5574 15700 6394
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16224 5642 16252 6258
rect 16316 6118 16344 6394
rect 16592 6254 16620 7278
rect 16684 6866 16712 9522
rect 16868 9450 16896 11154
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10810 17172 10950
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17144 10062 17172 10746
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 17328 9586 17356 10066
rect 17420 9994 17448 11698
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17512 9926 17540 10950
rect 17604 10130 17632 13262
rect 17788 11218 17816 14282
rect 17972 13802 18000 14758
rect 18156 14550 18184 19314
rect 18248 18970 18276 20402
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 18144 14544 18196 14550
rect 18144 14486 18196 14492
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 18064 12434 18092 13194
rect 17880 12406 18092 12434
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 10266 17816 10406
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 16856 9444 16908 9450
rect 16856 9386 16908 9392
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 16868 9110 16896 9386
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 17236 8974 17264 9318
rect 17328 8974 17356 9386
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17236 8090 17264 8434
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 17144 6934 17172 7958
rect 17328 7410 17356 8910
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17132 6928 17184 6934
rect 17132 6870 17184 6876
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15672 5302 15700 5510
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 16224 5234 16252 5578
rect 16316 5234 16344 6054
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 15028 4486 15056 5102
rect 15016 4480 15068 4486
rect 15016 4422 15068 4428
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 16592 3534 16620 6190
rect 16776 5574 16804 6326
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17144 5642 17172 6190
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16776 5234 16804 5510
rect 17236 5234 17264 5714
rect 17328 5370 17356 6258
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17420 5234 17448 5578
rect 17512 5234 17540 9862
rect 17788 9722 17816 9930
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17880 9602 17908 12406
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 17972 11898 18000 12106
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 18248 11830 18276 17002
rect 18340 14260 18368 22066
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 18432 20505 18460 20742
rect 18418 20496 18474 20505
rect 18418 20431 18474 20440
rect 18524 18426 18552 24278
rect 18604 23248 18656 23254
rect 18604 23190 18656 23196
rect 18616 20398 18644 23190
rect 18708 21010 18736 25894
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18800 22710 18828 22918
rect 18788 22704 18840 22710
rect 18788 22646 18840 22652
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18892 20602 18920 28358
rect 18972 27872 19024 27878
rect 18972 27814 19024 27820
rect 18984 27062 19012 27814
rect 18972 27056 19024 27062
rect 18972 26998 19024 27004
rect 18972 25900 19024 25906
rect 18972 25842 19024 25848
rect 18984 25362 19012 25842
rect 18972 25356 19024 25362
rect 18972 25298 19024 25304
rect 18972 25152 19024 25158
rect 18972 25094 19024 25100
rect 18984 24954 19012 25094
rect 18972 24948 19024 24954
rect 18972 24890 19024 24896
rect 18972 23520 19024 23526
rect 18972 23462 19024 23468
rect 18984 23118 19012 23462
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18512 18420 18564 18426
rect 18512 18362 18564 18368
rect 18892 18154 18920 18838
rect 18880 18148 18932 18154
rect 18880 18090 18932 18096
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18800 17746 18828 18022
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18892 17338 18920 17614
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18708 15706 18736 16050
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18972 15428 19024 15434
rect 18972 15370 19024 15376
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18432 14414 18460 15098
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18340 14232 18460 14260
rect 18432 13818 18460 14232
rect 18340 13790 18460 13818
rect 18340 12850 18368 13790
rect 18524 13530 18552 14350
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18616 13938 18644 14214
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18984 13002 19012 15370
rect 19076 13394 19104 35566
rect 19260 35442 19288 35702
rect 19168 35414 19288 35442
rect 19168 33454 19196 35414
rect 19156 33448 19208 33454
rect 19156 33390 19208 33396
rect 19156 32836 19208 32842
rect 19156 32778 19208 32784
rect 19168 31958 19196 32778
rect 19156 31952 19208 31958
rect 19156 31894 19208 31900
rect 19156 29164 19208 29170
rect 19156 29106 19208 29112
rect 19168 28762 19196 29106
rect 19156 28756 19208 28762
rect 19156 28698 19208 28704
rect 19352 28082 19380 37198
rect 20628 37188 20680 37194
rect 20628 37130 20680 37136
rect 20168 37120 20220 37126
rect 20168 37062 20220 37068
rect 20180 36854 20208 37062
rect 20640 36922 20668 37130
rect 20628 36916 20680 36922
rect 20628 36858 20680 36864
rect 20168 36848 20220 36854
rect 20168 36790 20220 36796
rect 20640 36310 20668 36858
rect 20628 36304 20680 36310
rect 20628 36246 20680 36252
rect 21284 36242 21312 37402
rect 22284 37256 22336 37262
rect 22284 37198 22336 37204
rect 22296 36922 22324 37198
rect 22940 37126 22968 39358
rect 25778 39358 26096 39386
rect 25778 39280 25834 39358
rect 25872 37256 25924 37262
rect 25872 37198 25924 37204
rect 25136 37188 25188 37194
rect 25136 37130 25188 37136
rect 22928 37120 22980 37126
rect 22928 37062 22980 37068
rect 22284 36916 22336 36922
rect 22284 36858 22336 36864
rect 21548 36576 21600 36582
rect 21548 36518 21600 36524
rect 21272 36236 21324 36242
rect 21272 36178 21324 36184
rect 19524 36032 19576 36038
rect 19524 35974 19576 35980
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 19444 29238 19472 30670
rect 19432 29232 19484 29238
rect 19432 29174 19484 29180
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19352 26382 19380 27610
rect 19432 27328 19484 27334
rect 19432 27270 19484 27276
rect 19444 26926 19472 27270
rect 19432 26920 19484 26926
rect 19432 26862 19484 26868
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19352 25378 19380 26318
rect 19260 25350 19380 25378
rect 19260 25294 19288 25350
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19352 24954 19380 25230
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 19338 21448 19394 21457
rect 19338 21383 19394 21392
rect 19352 20602 19380 21383
rect 19432 21072 19484 21078
rect 19432 21014 19484 21020
rect 19444 20602 19472 21014
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19352 18766 19380 19178
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19352 18290 19380 18702
rect 19430 18320 19486 18329
rect 19340 18284 19392 18290
rect 19430 18255 19486 18264
rect 19340 18226 19392 18232
rect 19444 18222 19472 18255
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19260 16182 19288 17614
rect 19248 16176 19300 16182
rect 19248 16118 19300 16124
rect 19536 14482 19564 35974
rect 21284 35766 21312 36178
rect 21560 36174 21588 36518
rect 22296 36378 22324 36858
rect 22560 36780 22612 36786
rect 22560 36722 22612 36728
rect 22836 36780 22888 36786
rect 22836 36722 22888 36728
rect 22284 36372 22336 36378
rect 22284 36314 22336 36320
rect 21548 36168 21600 36174
rect 21548 36110 21600 36116
rect 21272 35760 21324 35766
rect 21272 35702 21324 35708
rect 19708 35692 19760 35698
rect 19708 35634 19760 35640
rect 19720 35290 19748 35634
rect 20996 35488 21048 35494
rect 20996 35430 21048 35436
rect 19708 35284 19760 35290
rect 19708 35226 19760 35232
rect 19800 35148 19852 35154
rect 19800 35090 19852 35096
rect 19812 34610 19840 35090
rect 21008 35086 21036 35430
rect 21284 35086 21312 35702
rect 20996 35080 21048 35086
rect 20996 35022 21048 35028
rect 21088 35080 21140 35086
rect 21088 35022 21140 35028
rect 21272 35080 21324 35086
rect 21272 35022 21324 35028
rect 20352 34944 20404 34950
rect 20352 34886 20404 34892
rect 20364 34678 20392 34886
rect 20352 34672 20404 34678
rect 20352 34614 20404 34620
rect 21008 34626 21036 35022
rect 21100 34746 21128 35022
rect 21088 34740 21140 34746
rect 21088 34682 21140 34688
rect 19800 34604 19852 34610
rect 19800 34546 19852 34552
rect 20260 33312 20312 33318
rect 20260 33254 20312 33260
rect 20272 33046 20300 33254
rect 20260 33040 20312 33046
rect 19982 33008 20038 33017
rect 20260 32982 20312 32988
rect 19982 32943 19984 32952
rect 20036 32943 20038 32952
rect 19984 32914 20036 32920
rect 19892 32768 19944 32774
rect 19892 32710 19944 32716
rect 19904 32502 19932 32710
rect 19892 32496 19944 32502
rect 19892 32438 19944 32444
rect 19904 31754 19932 32438
rect 19996 32434 20024 32914
rect 20272 32910 20300 32982
rect 20260 32904 20312 32910
rect 20260 32846 20312 32852
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 20364 31754 20392 34614
rect 21008 34598 21128 34626
rect 20994 33144 21050 33153
rect 20994 33079 21050 33088
rect 20812 32972 20864 32978
rect 20812 32914 20864 32920
rect 19904 31726 20024 31754
rect 19892 31340 19944 31346
rect 19892 31282 19944 31288
rect 19708 31136 19760 31142
rect 19708 31078 19760 31084
rect 19720 30734 19748 31078
rect 19708 30728 19760 30734
rect 19708 30670 19760 30676
rect 19904 30394 19932 31282
rect 19892 30388 19944 30394
rect 19892 30330 19944 30336
rect 19708 30048 19760 30054
rect 19708 29990 19760 29996
rect 19720 29782 19748 29990
rect 19708 29776 19760 29782
rect 19708 29718 19760 29724
rect 19892 28960 19944 28966
rect 19892 28902 19944 28908
rect 19904 28558 19932 28902
rect 19996 28626 20024 31726
rect 20272 31726 20392 31754
rect 20272 30258 20300 31726
rect 20720 30592 20772 30598
rect 20720 30534 20772 30540
rect 20732 30394 20760 30534
rect 20720 30388 20772 30394
rect 20720 30330 20772 30336
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20260 30252 20312 30258
rect 20260 30194 20312 30200
rect 20272 30054 20300 30194
rect 20260 30048 20312 30054
rect 20260 29990 20312 29996
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 20456 29034 20484 29446
rect 20640 29306 20668 30262
rect 20628 29300 20680 29306
rect 20628 29242 20680 29248
rect 20536 29096 20588 29102
rect 20536 29038 20588 29044
rect 20444 29028 20496 29034
rect 20444 28970 20496 28976
rect 19984 28620 20036 28626
rect 19984 28562 20036 28568
rect 20168 28620 20220 28626
rect 20168 28562 20220 28568
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19996 27946 20024 28562
rect 20180 28082 20208 28562
rect 20456 28218 20484 28970
rect 20548 28404 20576 29038
rect 20640 28558 20668 29242
rect 20732 29102 20760 30330
rect 20824 29510 20852 32914
rect 20904 30048 20956 30054
rect 20904 29990 20956 29996
rect 20812 29504 20864 29510
rect 20812 29446 20864 29452
rect 20720 29096 20772 29102
rect 20720 29038 20772 29044
rect 20812 29096 20864 29102
rect 20812 29038 20864 29044
rect 20732 28694 20760 29038
rect 20824 28966 20852 29038
rect 20812 28960 20864 28966
rect 20812 28902 20864 28908
rect 20720 28688 20772 28694
rect 20720 28630 20772 28636
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20720 28552 20772 28558
rect 20720 28494 20772 28500
rect 20732 28404 20760 28494
rect 20548 28376 20760 28404
rect 20444 28212 20496 28218
rect 20444 28154 20496 28160
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 20352 28076 20404 28082
rect 20352 28018 20404 28024
rect 20364 27985 20392 28018
rect 20350 27976 20406 27985
rect 19984 27940 20036 27946
rect 20350 27911 20406 27920
rect 19984 27882 20036 27888
rect 20732 27878 20760 28376
rect 20812 27940 20864 27946
rect 20812 27882 20864 27888
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20732 27402 20760 27814
rect 20720 27396 20772 27402
rect 20720 27338 20772 27344
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 20640 27062 20668 27270
rect 19708 27056 19760 27062
rect 19708 26998 19760 27004
rect 20628 27056 20680 27062
rect 20628 26998 20680 27004
rect 19616 26784 19668 26790
rect 19616 26726 19668 26732
rect 19628 26382 19656 26726
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 19720 23730 19748 26998
rect 20824 26994 20852 27882
rect 19892 26988 19944 26994
rect 19892 26930 19944 26936
rect 20812 26988 20864 26994
rect 20812 26930 20864 26936
rect 19904 26042 19932 26930
rect 20720 26240 20772 26246
rect 20720 26182 20772 26188
rect 20732 26042 20760 26182
rect 19892 26036 19944 26042
rect 19892 25978 19944 25984
rect 20720 26036 20772 26042
rect 20720 25978 20772 25984
rect 20168 25832 20220 25838
rect 20168 25774 20220 25780
rect 20536 25832 20588 25838
rect 20536 25774 20588 25780
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19996 24954 20024 25094
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 19996 23798 20024 24890
rect 20180 24818 20208 25774
rect 20548 25362 20576 25774
rect 20536 25356 20588 25362
rect 20536 25298 20588 25304
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20456 23866 20484 24142
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19708 23724 19760 23730
rect 19708 23666 19760 23672
rect 19800 23724 19852 23730
rect 19800 23666 19852 23672
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19628 23118 19656 23598
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19628 22982 19656 23054
rect 19616 22976 19668 22982
rect 19616 22918 19668 22924
rect 19720 22094 19748 23666
rect 19812 23186 19840 23666
rect 20076 23656 20128 23662
rect 20076 23598 20128 23604
rect 19892 23588 19944 23594
rect 19892 23530 19944 23536
rect 19800 23180 19852 23186
rect 19800 23122 19852 23128
rect 19904 22778 19932 23530
rect 20088 23186 20116 23598
rect 20456 23594 20484 23802
rect 20732 23730 20760 25978
rect 20824 25786 20852 26930
rect 20916 26772 20944 29990
rect 21008 29170 21036 33079
rect 21100 32910 21128 34598
rect 21284 33522 21312 35022
rect 22100 34944 22152 34950
rect 22100 34886 22152 34892
rect 22112 34542 22140 34886
rect 22100 34536 22152 34542
rect 22100 34478 22152 34484
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 21362 33144 21418 33153
rect 22112 33114 22140 34478
rect 22284 33312 22336 33318
rect 22284 33254 22336 33260
rect 21362 33079 21418 33088
rect 22100 33108 22152 33114
rect 21376 32910 21404 33079
rect 22100 33050 22152 33056
rect 22192 33108 22244 33114
rect 22192 33050 22244 33056
rect 22112 32978 22140 33050
rect 22100 32972 22152 32978
rect 22100 32914 22152 32920
rect 21088 32904 21140 32910
rect 21088 32846 21140 32852
rect 21364 32904 21416 32910
rect 22204 32858 22232 33050
rect 22296 32978 22324 33254
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 21364 32846 21416 32852
rect 21100 32570 21128 32846
rect 21836 32830 22232 32858
rect 22296 32842 22324 32914
rect 22284 32836 22336 32842
rect 21088 32564 21140 32570
rect 21088 32506 21140 32512
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 21192 30394 21220 30670
rect 21180 30388 21232 30394
rect 21180 30330 21232 30336
rect 21088 29640 21140 29646
rect 21088 29582 21140 29588
rect 20996 29164 21048 29170
rect 20996 29106 21048 29112
rect 21008 28218 21036 29106
rect 21100 28626 21128 29582
rect 21180 29096 21232 29102
rect 21180 29038 21232 29044
rect 21088 28620 21140 28626
rect 21088 28562 21140 28568
rect 20996 28212 21048 28218
rect 20996 28154 21048 28160
rect 20996 26784 21048 26790
rect 20916 26744 20996 26772
rect 20996 26726 21048 26732
rect 21008 25906 21036 26726
rect 21192 26466 21220 29038
rect 21548 28960 21600 28966
rect 21548 28902 21600 28908
rect 21560 28626 21588 28902
rect 21548 28620 21600 28626
rect 21548 28562 21600 28568
rect 21732 28552 21784 28558
rect 21732 28494 21784 28500
rect 21744 28422 21772 28494
rect 21732 28416 21784 28422
rect 21732 28358 21784 28364
rect 21732 28144 21784 28150
rect 21652 28092 21732 28098
rect 21652 28086 21784 28092
rect 21548 28076 21600 28082
rect 21548 28018 21600 28024
rect 21652 28070 21772 28086
rect 21560 27674 21588 28018
rect 21652 27946 21680 28070
rect 21640 27940 21692 27946
rect 21640 27882 21692 27888
rect 21732 27940 21784 27946
rect 21732 27882 21784 27888
rect 21744 27674 21772 27882
rect 21548 27668 21600 27674
rect 21548 27610 21600 27616
rect 21732 27668 21784 27674
rect 21732 27610 21784 27616
rect 21272 26580 21324 26586
rect 21272 26522 21324 26528
rect 21100 26438 21220 26466
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 20824 25758 20944 25786
rect 20812 25696 20864 25702
rect 20812 25638 20864 25644
rect 20824 25498 20852 25638
rect 20812 25492 20864 25498
rect 20812 25434 20864 25440
rect 20916 24954 20944 25758
rect 20904 24948 20956 24954
rect 20904 24890 20956 24896
rect 20916 24698 20944 24890
rect 20916 24670 21036 24698
rect 21008 24614 21036 24670
rect 20904 24608 20956 24614
rect 20904 24550 20956 24556
rect 20996 24608 21048 24614
rect 20996 24550 21048 24556
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20444 23588 20496 23594
rect 20444 23530 20496 23536
rect 20260 23248 20312 23254
rect 20260 23190 20312 23196
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19892 22772 19944 22778
rect 19892 22714 19944 22720
rect 19720 22066 19840 22094
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 19720 21146 19748 21490
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19706 21040 19762 21049
rect 19706 20975 19762 20984
rect 19720 20942 19748 20975
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19616 20868 19668 20874
rect 19616 20810 19668 20816
rect 19628 20466 19656 20810
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19720 18222 19748 18702
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 19812 17066 19840 22066
rect 19982 21720 20038 21729
rect 19982 21655 20038 21664
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19904 19378 19932 20878
rect 19996 19666 20024 21655
rect 20088 21622 20116 23122
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 20076 21616 20128 21622
rect 20076 21558 20128 21564
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 20088 20602 20116 20878
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 20076 19712 20128 19718
rect 19996 19660 20076 19666
rect 19996 19654 20128 19660
rect 19996 19638 20116 19654
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19996 18154 20024 19638
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20088 19174 20116 19314
rect 20180 19258 20208 22034
rect 20272 19417 20300 23190
rect 20732 23186 20760 23666
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20824 23186 20852 23598
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20364 21146 20392 21286
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20732 21078 20760 21422
rect 20720 21072 20772 21078
rect 20720 21014 20772 21020
rect 20824 20942 20852 22714
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20812 19440 20864 19446
rect 20258 19408 20314 19417
rect 20258 19343 20314 19352
rect 20810 19408 20812 19417
rect 20864 19408 20866 19417
rect 20810 19343 20866 19352
rect 20534 19272 20590 19281
rect 20180 19230 20484 19258
rect 20180 19174 20208 19230
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20272 18902 20300 19110
rect 20260 18896 20312 18902
rect 20260 18838 20312 18844
rect 20352 18828 20404 18834
rect 20352 18770 20404 18776
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18290 20300 18566
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 19800 17060 19852 17066
rect 19800 17002 19852 17008
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19628 15502 19656 16186
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19812 15434 19840 17002
rect 20272 16250 20300 18226
rect 20364 18222 20392 18770
rect 20456 18272 20484 19230
rect 20534 19207 20590 19216
rect 20548 19009 20576 19207
rect 20534 19000 20590 19009
rect 20534 18935 20590 18944
rect 20812 18828 20864 18834
rect 20812 18770 20864 18776
rect 20536 18760 20588 18766
rect 20536 18702 20588 18708
rect 20548 18630 20576 18702
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 20824 18329 20852 18770
rect 20810 18320 20866 18329
rect 20536 18284 20588 18290
rect 20456 18244 20536 18272
rect 20810 18255 20866 18264
rect 20536 18226 20588 18232
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20364 17338 20392 18158
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20640 17338 20668 17478
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20824 16590 20852 17614
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 20088 15706 20116 16050
rect 20824 15910 20852 16526
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 20720 15632 20772 15638
rect 20720 15574 20772 15580
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 19800 15428 19852 15434
rect 19800 15370 19852 15376
rect 20272 14618 20300 15438
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19536 13394 19564 14418
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19628 14074 19656 14214
rect 19996 14074 20024 14486
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19064 13388 19116 13394
rect 19064 13330 19116 13336
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19076 13190 19104 13330
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 18984 12974 19104 13002
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18340 12238 18368 12786
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17972 11354 18000 11698
rect 18432 11694 18460 12718
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 18616 12306 18644 12650
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18512 12164 18564 12170
rect 18512 12106 18564 12112
rect 18524 11898 18552 12106
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 18524 11200 18552 11834
rect 18616 11762 18644 12242
rect 18892 11830 18920 12582
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18696 11824 18748 11830
rect 18696 11766 18748 11772
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18708 11558 18736 11766
rect 18984 11558 19012 12174
rect 19076 11898 19104 12974
rect 19248 12436 19300 12442
rect 19536 12434 19564 13330
rect 19628 13326 19656 14010
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20272 13530 20300 13874
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20456 13326 20484 14214
rect 20732 13530 20760 15574
rect 20824 15502 20852 15846
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20824 14074 20852 14214
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20824 13326 20852 14010
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 19248 12378 19300 12384
rect 19444 12406 19564 12434
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18786 11248 18842 11257
rect 18604 11212 18656 11218
rect 18524 11172 18604 11200
rect 18786 11183 18842 11192
rect 18604 11154 18656 11160
rect 18800 11150 18828 11183
rect 18984 11150 19012 11494
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 19076 10713 19104 10950
rect 19062 10704 19118 10713
rect 19062 10639 19118 10648
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17788 9574 17908 9602
rect 17788 8430 17816 9574
rect 17972 9518 18000 9862
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17604 7206 17632 7686
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 16776 4690 16804 5170
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16960 4622 16988 5170
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16580 3528 16632 3534
rect 17592 3528 17644 3534
rect 16580 3470 16632 3476
rect 17498 3496 17554 3505
rect 16212 3460 16264 3466
rect 17592 3470 17644 3476
rect 17498 3431 17554 3440
rect 16212 3402 16264 3408
rect 16224 3194 16252 3402
rect 17512 3398 17540 3431
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 17144 3126 17172 3334
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 16040 2446 16068 3062
rect 17604 3058 17632 3470
rect 17788 3126 17816 8366
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18248 6866 18276 7890
rect 18420 7880 18472 7886
rect 18604 7880 18656 7886
rect 18420 7822 18472 7828
rect 18524 7840 18604 7868
rect 18432 7750 18460 7822
rect 18420 7744 18472 7750
rect 18340 7704 18420 7732
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18248 6322 18276 6802
rect 18340 6798 18368 7704
rect 18420 7686 18472 7692
rect 18524 7206 18552 7840
rect 18604 7822 18656 7828
rect 18708 7818 18736 8774
rect 18892 8090 18920 9590
rect 19064 8356 19116 8362
rect 19064 8298 19116 8304
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 19076 7954 19104 8298
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 18696 7812 18748 7818
rect 18748 7772 18920 7800
rect 18696 7754 18748 7760
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18524 6798 18552 7142
rect 18328 6792 18380 6798
rect 18512 6792 18564 6798
rect 18380 6752 18460 6780
rect 18328 6734 18380 6740
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18340 6118 18368 6598
rect 18328 6112 18380 6118
rect 18328 6054 18380 6060
rect 18340 5710 18368 6054
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18432 5642 18460 6752
rect 18512 6734 18564 6740
rect 18524 5914 18552 6734
rect 18696 6724 18748 6730
rect 18696 6666 18748 6672
rect 18708 6390 18736 6666
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 18892 6322 18920 7772
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 18800 5914 18828 6190
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18892 5778 18920 6258
rect 18984 5778 19012 6734
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 19076 5642 19104 6258
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 19064 5636 19116 5642
rect 19064 5578 19116 5584
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18052 3528 18104 3534
rect 18050 3496 18052 3505
rect 18104 3496 18106 3505
rect 18050 3431 18106 3440
rect 18248 3398 18276 3878
rect 18340 3466 18368 4762
rect 18616 4146 18644 5170
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18328 3460 18380 3466
rect 18328 3402 18380 3408
rect 18616 3398 18644 4082
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18708 3738 18736 4014
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 3194 18644 3334
rect 18708 3194 18736 3674
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18156 2650 18184 2994
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 2228 2304 2280 2310
rect 2228 2246 2280 2252
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2240 2038 2268 2246
rect 2228 2032 2280 2038
rect 2228 1974 2280 1980
rect 2608 800 2636 2246
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5828 800 5856 2382
rect 9048 800 9076 2382
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 11624 800 11652 2246
rect 14844 800 14872 2246
rect 18064 800 18092 2382
rect 19168 2378 19196 12106
rect 19260 11937 19288 12378
rect 19246 11928 19302 11937
rect 19246 11863 19302 11872
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 11286 19288 11698
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19248 11076 19300 11082
rect 19444 11064 19472 12406
rect 19524 12232 19576 12238
rect 19984 12232 20036 12238
rect 19524 12174 19576 12180
rect 19890 12200 19946 12209
rect 19536 11626 19564 12174
rect 19984 12174 20036 12180
rect 19890 12135 19892 12144
rect 19944 12135 19946 12144
rect 19892 12106 19944 12112
rect 19708 12096 19760 12102
rect 19708 12038 19760 12044
rect 19720 11762 19748 12038
rect 19996 11762 20024 12174
rect 20916 11801 20944 24550
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21008 22094 21036 23054
rect 21100 22778 21128 26438
rect 21180 26308 21232 26314
rect 21180 26250 21232 26256
rect 21192 24818 21220 26250
rect 21284 26246 21312 26522
rect 21836 26450 21864 32830
rect 22284 32778 22336 32784
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 22100 32768 22152 32774
rect 22100 32710 22152 32716
rect 21824 26444 21876 26450
rect 21824 26386 21876 26392
rect 21364 26376 21416 26382
rect 21364 26318 21416 26324
rect 21916 26376 21968 26382
rect 21916 26318 21968 26324
rect 21272 26240 21324 26246
rect 21272 26182 21324 26188
rect 21376 25974 21404 26318
rect 21548 26308 21600 26314
rect 21548 26250 21600 26256
rect 21364 25968 21416 25974
rect 21364 25910 21416 25916
rect 21180 24812 21232 24818
rect 21180 24754 21232 24760
rect 21560 24750 21588 26250
rect 21732 25900 21784 25906
rect 21732 25842 21784 25848
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 21548 24744 21600 24750
rect 21548 24686 21600 24692
rect 21284 24410 21312 24686
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21272 24404 21324 24410
rect 21272 24346 21324 24352
rect 21364 24336 21416 24342
rect 21364 24278 21416 24284
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 21180 22432 21232 22438
rect 21180 22374 21232 22380
rect 21192 22098 21220 22374
rect 21008 22066 21128 22094
rect 20996 21480 21048 21486
rect 20994 21448 20996 21457
rect 21048 21448 21050 21457
rect 20994 21383 21050 21392
rect 21008 21146 21036 21383
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 20994 20360 21050 20369
rect 20994 20295 21050 20304
rect 21008 19922 21036 20295
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20996 19780 21048 19786
rect 20996 19722 21048 19728
rect 21008 19446 21036 19722
rect 20996 19440 21048 19446
rect 20996 19382 21048 19388
rect 21100 19281 21128 22066
rect 21180 22092 21232 22098
rect 21180 22034 21232 22040
rect 21192 21162 21220 22034
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 21284 21690 21312 21966
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21192 21134 21312 21162
rect 21180 21072 21232 21078
rect 21180 21014 21232 21020
rect 21192 20942 21220 21014
rect 21180 20936 21232 20942
rect 21180 20878 21232 20884
rect 21180 20324 21232 20330
rect 21180 20266 21232 20272
rect 21086 19272 21142 19281
rect 21086 19207 21142 19216
rect 21192 18426 21220 20266
rect 21284 19854 21312 21134
rect 21376 20346 21404 24278
rect 21456 24268 21508 24274
rect 21456 24210 21508 24216
rect 21468 23866 21496 24210
rect 21456 23860 21508 23866
rect 21456 23802 21508 23808
rect 21560 23526 21588 24550
rect 21640 24336 21692 24342
rect 21640 24278 21692 24284
rect 21744 24290 21772 25842
rect 21928 25702 21956 26318
rect 21916 25696 21968 25702
rect 21916 25638 21968 25644
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21836 24410 21864 24754
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21652 23866 21680 24278
rect 21744 24262 21864 24290
rect 21732 24064 21784 24070
rect 21732 24006 21784 24012
rect 21744 23866 21772 24006
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 21732 23860 21784 23866
rect 21732 23802 21784 23808
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21836 23338 21864 24262
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 21560 23310 21864 23338
rect 21468 22982 21496 23258
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 21468 21010 21496 21286
rect 21456 21004 21508 21010
rect 21456 20946 21508 20952
rect 21376 20318 21496 20346
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21272 19848 21324 19854
rect 21376 19850 21404 20198
rect 21272 19790 21324 19796
rect 21364 19844 21416 19850
rect 21364 19786 21416 19792
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21284 19514 21312 19654
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21468 18970 21496 20318
rect 21560 20244 21588 23310
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 21652 21418 21680 22918
rect 22020 21554 22048 32710
rect 22112 32570 22140 32710
rect 22296 32570 22324 32778
rect 22100 32564 22152 32570
rect 22100 32506 22152 32512
rect 22284 32564 22336 32570
rect 22284 32506 22336 32512
rect 22192 30592 22244 30598
rect 22192 30534 22244 30540
rect 22204 30394 22232 30534
rect 22192 30388 22244 30394
rect 22192 30330 22244 30336
rect 22284 30320 22336 30326
rect 22284 30262 22336 30268
rect 22296 30054 22324 30262
rect 22468 30184 22520 30190
rect 22468 30126 22520 30132
rect 22284 30048 22336 30054
rect 22284 29990 22336 29996
rect 22480 29238 22508 30126
rect 22468 29232 22520 29238
rect 22468 29174 22520 29180
rect 22376 28416 22428 28422
rect 22376 28358 22428 28364
rect 22388 26586 22416 28358
rect 22376 26580 22428 26586
rect 22376 26522 22428 26528
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22112 25226 22140 25842
rect 22480 25537 22508 26250
rect 22466 25528 22522 25537
rect 22466 25463 22522 25472
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 22112 24410 22140 25162
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22204 21690 22232 21830
rect 22296 21690 22324 23462
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 21640 21412 21692 21418
rect 21640 21354 21692 21360
rect 22296 20602 22324 21626
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 21824 20528 21876 20534
rect 21824 20470 21876 20476
rect 21560 20216 21680 20244
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 21560 19514 21588 19722
rect 21548 19508 21600 19514
rect 21548 19450 21600 19456
rect 21548 19372 21600 19378
rect 21548 19314 21600 19320
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 21560 18766 21588 19314
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 21008 17338 21036 17546
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 21560 16250 21588 18702
rect 21652 18426 21680 20216
rect 21836 19718 21864 20470
rect 22284 20392 22336 20398
rect 22282 20360 22284 20369
rect 22336 20360 22338 20369
rect 22282 20295 22338 20304
rect 22008 19780 22060 19786
rect 22008 19722 22060 19728
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21744 19122 21772 19246
rect 21836 19242 21864 19654
rect 22020 19514 22048 19722
rect 22388 19530 22416 24550
rect 22468 24200 22520 24206
rect 22468 24142 22520 24148
rect 22480 23730 22508 24142
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22480 19666 22508 23666
rect 22572 22094 22600 36722
rect 22744 36644 22796 36650
rect 22744 36586 22796 36592
rect 22756 36378 22784 36586
rect 22744 36372 22796 36378
rect 22744 36314 22796 36320
rect 22848 35086 22876 36722
rect 24124 36576 24176 36582
rect 24124 36518 24176 36524
rect 22836 35080 22888 35086
rect 22836 35022 22888 35028
rect 23940 35080 23992 35086
rect 23940 35022 23992 35028
rect 22744 33516 22796 33522
rect 22744 33458 22796 33464
rect 22652 32972 22704 32978
rect 22652 32914 22704 32920
rect 22664 32026 22692 32914
rect 22756 32570 22784 33458
rect 22744 32564 22796 32570
rect 22744 32506 22796 32512
rect 22848 32366 22876 35022
rect 23952 34746 23980 35022
rect 23940 34740 23992 34746
rect 23940 34682 23992 34688
rect 23848 34604 23900 34610
rect 23848 34546 23900 34552
rect 23480 32972 23532 32978
rect 23480 32914 23532 32920
rect 23020 32904 23072 32910
rect 23020 32846 23072 32852
rect 23032 32774 23060 32846
rect 23020 32768 23072 32774
rect 23020 32710 23072 32716
rect 22836 32360 22888 32366
rect 22836 32302 22888 32308
rect 22652 32020 22704 32026
rect 22652 31962 22704 31968
rect 23492 31958 23520 32914
rect 23480 31952 23532 31958
rect 23480 31894 23532 31900
rect 23492 31482 23520 31894
rect 23860 31754 23888 34546
rect 23940 32836 23992 32842
rect 23940 32778 23992 32784
rect 23952 32026 23980 32778
rect 24032 32768 24084 32774
rect 24032 32710 24084 32716
rect 24044 32502 24072 32710
rect 24032 32496 24084 32502
rect 24032 32438 24084 32444
rect 23940 32020 23992 32026
rect 23940 31962 23992 31968
rect 23768 31726 23888 31754
rect 23480 31476 23532 31482
rect 23480 31418 23532 31424
rect 23296 31204 23348 31210
rect 23296 31146 23348 31152
rect 22652 30728 22704 30734
rect 22652 30670 22704 30676
rect 22664 29714 22692 30670
rect 22652 29708 22704 29714
rect 22652 29650 22704 29656
rect 22664 29170 22692 29650
rect 23308 29646 23336 31146
rect 23768 30258 23796 31726
rect 23848 31340 23900 31346
rect 23848 31282 23900 31288
rect 23756 30252 23808 30258
rect 23756 30194 23808 30200
rect 23388 30116 23440 30122
rect 23388 30058 23440 30064
rect 23296 29640 23348 29646
rect 23296 29582 23348 29588
rect 23308 29170 23336 29582
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22928 29164 22980 29170
rect 22928 29106 22980 29112
rect 23296 29164 23348 29170
rect 23296 29106 23348 29112
rect 22940 28762 22968 29106
rect 22928 28756 22980 28762
rect 22928 28698 22980 28704
rect 23400 28626 23428 30058
rect 23664 28960 23716 28966
rect 23664 28902 23716 28908
rect 23388 28620 23440 28626
rect 23388 28562 23440 28568
rect 23676 28490 23704 28902
rect 23664 28484 23716 28490
rect 23664 28426 23716 28432
rect 23388 28416 23440 28422
rect 23388 28358 23440 28364
rect 23400 28218 23428 28358
rect 23388 28212 23440 28218
rect 23388 28154 23440 28160
rect 23664 28008 23716 28014
rect 23664 27950 23716 27956
rect 23570 27568 23626 27577
rect 23676 27538 23704 27950
rect 23860 27946 23888 31282
rect 23952 31210 23980 31962
rect 23940 31204 23992 31210
rect 23940 31146 23992 31152
rect 24032 30252 24084 30258
rect 24032 30194 24084 30200
rect 24044 29102 24072 30194
rect 24032 29096 24084 29102
rect 24032 29038 24084 29044
rect 23848 27940 23900 27946
rect 23848 27882 23900 27888
rect 24032 27872 24084 27878
rect 24032 27814 24084 27820
rect 24044 27674 24072 27814
rect 24032 27668 24084 27674
rect 24032 27610 24084 27616
rect 23570 27503 23572 27512
rect 23624 27503 23626 27512
rect 23664 27532 23716 27538
rect 23572 27474 23624 27480
rect 23664 27474 23716 27480
rect 23664 27124 23716 27130
rect 23664 27066 23716 27072
rect 22836 27056 22888 27062
rect 22836 26998 22888 27004
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 22756 26518 22784 26930
rect 22744 26512 22796 26518
rect 22744 26454 22796 26460
rect 22756 26042 22784 26454
rect 22744 26036 22796 26042
rect 22744 25978 22796 25984
rect 22848 25974 22876 26998
rect 23480 26784 23532 26790
rect 23480 26726 23532 26732
rect 23204 26444 23256 26450
rect 23204 26386 23256 26392
rect 22928 26308 22980 26314
rect 22928 26250 22980 26256
rect 22836 25968 22888 25974
rect 22836 25910 22888 25916
rect 22940 24818 22968 26250
rect 23216 25770 23244 26386
rect 23204 25764 23256 25770
rect 23204 25706 23256 25712
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 23112 24812 23164 24818
rect 23112 24754 23164 24760
rect 22836 24608 22888 24614
rect 22836 24550 22888 24556
rect 22848 23730 22876 24550
rect 23124 24410 23152 24754
rect 23204 24744 23256 24750
rect 23204 24686 23256 24692
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 23216 24206 23244 24686
rect 23492 24206 23520 26726
rect 23572 25696 23624 25702
rect 23572 25638 23624 25644
rect 23584 24410 23612 25638
rect 23572 24404 23624 24410
rect 23572 24346 23624 24352
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23020 24064 23072 24070
rect 23020 24006 23072 24012
rect 22836 23724 22888 23730
rect 22836 23666 22888 23672
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22572 22066 22784 22094
rect 22480 19638 22600 19666
rect 22008 19508 22060 19514
rect 22388 19502 22508 19530
rect 22008 19450 22060 19456
rect 21824 19236 21876 19242
rect 21824 19178 21876 19184
rect 22008 19168 22060 19174
rect 21928 19128 22008 19156
rect 21928 19122 21956 19128
rect 21744 19094 21956 19122
rect 22008 19110 22060 19116
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21836 17202 21864 18022
rect 22112 17882 22140 18158
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22112 15178 22140 15438
rect 22020 15150 22140 15178
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21008 13258 21036 14418
rect 21376 14346 21404 14418
rect 21364 14340 21416 14346
rect 21364 14282 21416 14288
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21192 13394 21220 14214
rect 21272 14000 21324 14006
rect 21272 13942 21324 13948
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 21192 12986 21220 13330
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 21100 12345 21128 12378
rect 21086 12336 21142 12345
rect 21086 12271 21142 12280
rect 20902 11792 20958 11801
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 20444 11756 20496 11762
rect 20902 11727 20958 11736
rect 20444 11698 20496 11704
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19300 11036 19472 11064
rect 19248 11018 19300 11024
rect 19248 10532 19300 10538
rect 19248 10474 19300 10480
rect 19260 10130 19288 10474
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19260 7886 19288 10066
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19260 6254 19288 6938
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19352 5710 19380 6054
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 4078 19380 5646
rect 19444 4282 19472 11036
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19260 3482 19288 3538
rect 19432 3528 19484 3534
rect 19260 3454 19380 3482
rect 19432 3470 19484 3476
rect 19352 2990 19380 3454
rect 19444 3194 19472 3470
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19536 2650 19564 11018
rect 19812 7857 19840 11698
rect 19996 11558 20024 11698
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 19996 11150 20024 11222
rect 20456 11150 20484 11698
rect 19984 11144 20036 11150
rect 20260 11144 20312 11150
rect 19984 11086 20036 11092
rect 20258 11112 20260 11121
rect 20444 11144 20496 11150
rect 20312 11112 20314 11121
rect 20444 11086 20496 11092
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20258 11047 20314 11056
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20640 9926 20668 10610
rect 20824 10146 20852 11086
rect 21192 11082 21220 12922
rect 21284 12306 21312 13942
rect 21376 13394 21404 14282
rect 21548 14000 21600 14006
rect 22020 13954 22048 15150
rect 21600 13948 22048 13954
rect 21548 13942 22048 13948
rect 21560 13926 22048 13942
rect 22020 13870 22048 13926
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 21836 13530 21864 13806
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22006 12336 22062 12345
rect 21272 12300 21324 12306
rect 22006 12271 22062 12280
rect 21272 12242 21324 12248
rect 22020 12238 22048 12271
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21824 12164 21876 12170
rect 21824 12106 21876 12112
rect 21836 11898 21864 12106
rect 21928 11898 21956 12174
rect 22112 11898 22140 13126
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22204 11218 22232 16594
rect 22376 15428 22428 15434
rect 22376 15370 22428 15376
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22296 14618 22324 14962
rect 22388 14822 22416 15370
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22284 14000 22336 14006
rect 22284 13942 22336 13948
rect 22296 13734 22324 13942
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22480 12238 22508 19502
rect 22572 15706 22600 19638
rect 22756 18170 22784 22066
rect 22848 21486 22876 22578
rect 22836 21480 22888 21486
rect 22836 21422 22888 21428
rect 22928 21344 22980 21350
rect 22928 21286 22980 21292
rect 22940 20398 22968 21286
rect 22928 20392 22980 20398
rect 22928 20334 22980 20340
rect 22928 18284 22980 18290
rect 22928 18226 22980 18232
rect 22756 18142 22876 18170
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22756 17678 22784 18022
rect 22744 17672 22796 17678
rect 22744 17614 22796 17620
rect 22652 17604 22704 17610
rect 22652 17546 22704 17552
rect 22664 16046 22692 17546
rect 22848 16538 22876 18142
rect 22940 17338 22968 18226
rect 22928 17332 22980 17338
rect 22928 17274 22980 17280
rect 22756 16510 22876 16538
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22756 14346 22784 16510
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22848 16114 22876 16390
rect 22836 16108 22888 16114
rect 22836 16050 22888 16056
rect 23032 15094 23060 24006
rect 23216 23798 23244 24142
rect 23400 23866 23428 24142
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 23204 23792 23256 23798
rect 23676 23769 23704 27066
rect 23940 24744 23992 24750
rect 23940 24686 23992 24692
rect 23756 24676 23808 24682
rect 23756 24618 23808 24624
rect 23768 24206 23796 24618
rect 23952 24410 23980 24686
rect 23940 24404 23992 24410
rect 23940 24346 23992 24352
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23940 24200 23992 24206
rect 23940 24142 23992 24148
rect 23204 23734 23256 23740
rect 23662 23760 23718 23769
rect 23662 23695 23718 23704
rect 23388 23588 23440 23594
rect 23388 23530 23440 23536
rect 23400 23497 23428 23530
rect 23386 23488 23442 23497
rect 23386 23423 23442 23432
rect 23112 22568 23164 22574
rect 23112 22510 23164 22516
rect 23124 22098 23152 22510
rect 23112 22092 23164 22098
rect 23112 22034 23164 22040
rect 23124 21554 23152 22034
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23400 21146 23428 21490
rect 23388 21140 23440 21146
rect 23388 21082 23440 21088
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23296 20324 23348 20330
rect 23296 20266 23348 20272
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 23124 19009 23152 19654
rect 23308 19310 23336 20266
rect 23584 20058 23612 20402
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23676 19922 23704 23695
rect 23952 23662 23980 24142
rect 24032 24064 24084 24070
rect 24032 24006 24084 24012
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 24044 23594 24072 24006
rect 24032 23588 24084 23594
rect 24032 23530 24084 23536
rect 23756 22976 23808 22982
rect 23756 22918 23808 22924
rect 23768 22710 23796 22918
rect 23756 22704 23808 22710
rect 23756 22646 23808 22652
rect 24136 20346 24164 36518
rect 25148 35894 25176 37130
rect 25884 36553 25912 37198
rect 26068 37126 26096 39358
rect 28354 39358 28488 39386
rect 28354 39280 28410 39358
rect 28460 37330 28488 39358
rect 31574 39358 31708 39386
rect 31574 39280 31630 39358
rect 31680 38298 31708 39358
rect 34794 39280 34850 40080
rect 37370 39280 37426 40080
rect 31680 38270 31800 38298
rect 31772 37398 31800 38270
rect 29920 37392 29972 37398
rect 29920 37334 29972 37340
rect 31760 37392 31812 37398
rect 31760 37334 31812 37340
rect 28448 37324 28500 37330
rect 28448 37266 28500 37272
rect 28632 37256 28684 37262
rect 28632 37198 28684 37204
rect 26056 37120 26108 37126
rect 26056 37062 26108 37068
rect 25870 36544 25926 36553
rect 25870 36479 25926 36488
rect 25056 35866 25176 35894
rect 28644 35894 28672 37198
rect 29276 36236 29328 36242
rect 29276 36178 29328 36184
rect 28644 35866 28764 35894
rect 24492 35284 24544 35290
rect 24492 35226 24544 35232
rect 24308 34944 24360 34950
rect 24308 34886 24360 34892
rect 24320 34746 24348 34886
rect 24308 34740 24360 34746
rect 24308 34682 24360 34688
rect 24504 34542 24532 35226
rect 24952 35080 25004 35086
rect 24952 35022 25004 35028
rect 24860 34944 24912 34950
rect 24780 34904 24860 34932
rect 24780 34610 24808 34904
rect 24860 34886 24912 34892
rect 24964 34746 24992 35022
rect 24952 34740 25004 34746
rect 24952 34682 25004 34688
rect 24768 34604 24820 34610
rect 24768 34546 24820 34552
rect 25056 34542 25084 35866
rect 25504 35012 25556 35018
rect 25504 34954 25556 34960
rect 25412 34672 25464 34678
rect 25412 34614 25464 34620
rect 24492 34536 24544 34542
rect 24492 34478 24544 34484
rect 25044 34536 25096 34542
rect 25044 34478 25096 34484
rect 24400 33516 24452 33522
rect 24400 33458 24452 33464
rect 24308 33448 24360 33454
rect 24308 33390 24360 33396
rect 24216 33312 24268 33318
rect 24216 33254 24268 33260
rect 24228 32910 24256 33254
rect 24320 33017 24348 33390
rect 24306 33008 24362 33017
rect 24306 32943 24362 32952
rect 24216 32904 24268 32910
rect 24216 32846 24268 32852
rect 24320 31958 24348 32943
rect 24412 32774 24440 33458
rect 24768 32972 24820 32978
rect 24768 32914 24820 32920
rect 24492 32904 24544 32910
rect 24492 32846 24544 32852
rect 24400 32768 24452 32774
rect 24400 32710 24452 32716
rect 24412 32298 24440 32710
rect 24504 32570 24532 32846
rect 24492 32564 24544 32570
rect 24492 32506 24544 32512
rect 24780 32434 24808 32914
rect 24768 32428 24820 32434
rect 24768 32370 24820 32376
rect 24400 32292 24452 32298
rect 24400 32234 24452 32240
rect 24308 31952 24360 31958
rect 24308 31894 24360 31900
rect 24768 31340 24820 31346
rect 24768 31282 24820 31288
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24216 30592 24268 30598
rect 24216 30534 24268 30540
rect 24228 30258 24256 30534
rect 24596 30394 24624 30670
rect 24584 30388 24636 30394
rect 24584 30330 24636 30336
rect 24780 30326 24808 31282
rect 24952 31272 25004 31278
rect 24952 31214 25004 31220
rect 24964 30734 24992 31214
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 24768 30320 24820 30326
rect 24768 30262 24820 30268
rect 24216 30252 24268 30258
rect 24216 30194 24268 30200
rect 24400 30252 24452 30258
rect 24400 30194 24452 30200
rect 24412 28082 24440 30194
rect 24492 29232 24544 29238
rect 24492 29174 24544 29180
rect 24504 28218 24532 29174
rect 24584 28960 24636 28966
rect 24584 28902 24636 28908
rect 24492 28212 24544 28218
rect 24492 28154 24544 28160
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24216 27940 24268 27946
rect 24216 27882 24268 27888
rect 24228 20466 24256 27882
rect 24412 27334 24440 28018
rect 24504 27470 24532 28154
rect 24596 28082 24624 28902
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24780 27996 24808 30262
rect 25056 30258 25084 34478
rect 25424 32910 25452 34614
rect 25516 34542 25544 34954
rect 25596 34944 25648 34950
rect 25596 34886 25648 34892
rect 26516 34944 26568 34950
rect 26516 34886 26568 34892
rect 25608 34610 25636 34886
rect 25596 34604 25648 34610
rect 25596 34546 25648 34552
rect 26528 34542 26556 34886
rect 25504 34536 25556 34542
rect 25504 34478 25556 34484
rect 26332 34536 26384 34542
rect 26332 34478 26384 34484
rect 26516 34536 26568 34542
rect 26516 34478 26568 34484
rect 26344 33454 26372 34478
rect 26332 33448 26384 33454
rect 26332 33390 26384 33396
rect 26424 33380 26476 33386
rect 26424 33322 26476 33328
rect 25688 33108 25740 33114
rect 25688 33050 25740 33056
rect 26148 33108 26200 33114
rect 26148 33050 26200 33056
rect 25700 32910 25728 33050
rect 25412 32904 25464 32910
rect 25412 32846 25464 32852
rect 25504 32904 25556 32910
rect 25504 32846 25556 32852
rect 25688 32904 25740 32910
rect 25688 32846 25740 32852
rect 25424 32348 25452 32846
rect 25516 32774 25544 32846
rect 25504 32768 25556 32774
rect 25504 32710 25556 32716
rect 25688 32768 25740 32774
rect 25688 32710 25740 32716
rect 25516 32450 25544 32710
rect 25516 32434 25636 32450
rect 25516 32428 25648 32434
rect 25516 32422 25596 32428
rect 25596 32370 25648 32376
rect 25504 32360 25556 32366
rect 25424 32320 25504 32348
rect 25700 32314 25728 32710
rect 25504 32302 25556 32308
rect 25228 32292 25280 32298
rect 25228 32234 25280 32240
rect 25608 32286 25728 32314
rect 25780 32360 25832 32366
rect 25780 32302 25832 32308
rect 25240 31929 25268 32234
rect 25226 31920 25282 31929
rect 25226 31855 25282 31864
rect 25240 30870 25268 31855
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 25228 30864 25280 30870
rect 25228 30806 25280 30812
rect 25332 30802 25360 31282
rect 25320 30796 25372 30802
rect 25320 30738 25372 30744
rect 25136 30728 25188 30734
rect 25136 30670 25188 30676
rect 25148 30394 25176 30670
rect 25136 30388 25188 30394
rect 25136 30330 25188 30336
rect 25044 30252 25096 30258
rect 25044 30194 25096 30200
rect 24952 30184 25004 30190
rect 24952 30126 25004 30132
rect 24964 29714 24992 30126
rect 24952 29708 25004 29714
rect 24952 29650 25004 29656
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24872 29306 24900 29582
rect 25504 29504 25556 29510
rect 25504 29446 25556 29452
rect 25516 29306 25544 29446
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 25504 29300 25556 29306
rect 25504 29242 25556 29248
rect 25044 29096 25096 29102
rect 25044 29038 25096 29044
rect 24952 28212 25004 28218
rect 24952 28154 25004 28160
rect 24860 28008 24912 28014
rect 24780 27968 24860 27996
rect 24492 27464 24544 27470
rect 24492 27406 24544 27412
rect 24400 27328 24452 27334
rect 24400 27270 24452 27276
rect 24780 27130 24808 27968
rect 24964 27985 24992 28154
rect 24860 27950 24912 27956
rect 24950 27976 25006 27985
rect 24950 27911 25006 27920
rect 24860 27872 24912 27878
rect 24860 27814 24912 27820
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24584 26376 24636 26382
rect 24584 26318 24636 26324
rect 24400 26240 24452 26246
rect 24400 26182 24452 26188
rect 24412 25974 24440 26182
rect 24400 25968 24452 25974
rect 24400 25910 24452 25916
rect 24596 25498 24624 26318
rect 24584 25492 24636 25498
rect 24584 25434 24636 25440
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24688 24274 24716 25434
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24688 23730 24716 24210
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 24676 22976 24728 22982
rect 24780 22964 24808 26930
rect 24872 25906 24900 27814
rect 24964 27538 24992 27911
rect 24952 27532 25004 27538
rect 24952 27474 25004 27480
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 24872 23866 24900 24142
rect 24860 23860 24912 23866
rect 24860 23802 24912 23808
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 24728 22936 24808 22964
rect 24676 22918 24728 22924
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 24504 21350 24532 21490
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 24308 20868 24360 20874
rect 24308 20810 24360 20816
rect 24320 20505 24348 20810
rect 24306 20496 24362 20505
rect 24216 20460 24268 20466
rect 24306 20431 24308 20440
rect 24216 20402 24268 20408
rect 24360 20431 24362 20440
rect 24308 20402 24360 20408
rect 24136 20318 24348 20346
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 23664 19916 23716 19922
rect 23664 19858 23716 19864
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23400 19378 23428 19790
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23110 19000 23166 19009
rect 23110 18935 23166 18944
rect 23124 18834 23152 18935
rect 23112 18828 23164 18834
rect 23112 18770 23164 18776
rect 23204 18692 23256 18698
rect 23204 18634 23256 18640
rect 23216 18290 23244 18634
rect 23204 18284 23256 18290
rect 23204 18226 23256 18232
rect 23400 15706 23428 19314
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23584 18222 23612 18702
rect 23676 18222 23704 19110
rect 23848 18896 23900 18902
rect 23848 18838 23900 18844
rect 23572 18216 23624 18222
rect 23664 18216 23716 18222
rect 23572 18158 23624 18164
rect 23662 18184 23664 18193
rect 23756 18216 23808 18222
rect 23716 18184 23718 18193
rect 23756 18158 23808 18164
rect 23860 18170 23888 18838
rect 23940 18624 23992 18630
rect 23940 18566 23992 18572
rect 23952 18290 23980 18566
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 24032 18216 24084 18222
rect 23860 18164 24032 18170
rect 23860 18158 24084 18164
rect 23662 18119 23718 18128
rect 23664 17264 23716 17270
rect 23664 17206 23716 17212
rect 23676 16658 23704 17206
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 23664 16516 23716 16522
rect 23768 16504 23796 18158
rect 23860 18142 24072 18158
rect 23860 17882 23888 18142
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 23860 17338 23888 17818
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23716 16476 23796 16504
rect 23664 16458 23716 16464
rect 23768 16250 23796 16476
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23952 15502 23980 16594
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 24136 15162 24164 20198
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24228 18290 24256 18906
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 24124 15156 24176 15162
rect 24124 15098 24176 15104
rect 23020 15088 23072 15094
rect 23020 15030 23072 15036
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 22744 14340 22796 14346
rect 22744 14282 22796 14288
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22664 14074 22692 14214
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22664 13326 22692 14010
rect 22756 13326 22784 14282
rect 22928 13388 22980 13394
rect 22928 13330 22980 13336
rect 22652 13320 22704 13326
rect 22652 13262 22704 13268
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22756 13190 22784 13262
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22756 12238 22784 12582
rect 22940 12442 22968 13330
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22282 11792 22338 11801
rect 22664 11762 22692 12038
rect 22652 11756 22704 11762
rect 22338 11736 22416 11744
rect 22282 11727 22284 11736
rect 22336 11716 22416 11736
rect 22284 11698 22336 11704
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 21272 10736 21324 10742
rect 21324 10696 21404 10724
rect 21272 10678 21324 10684
rect 21376 10606 21404 10696
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21284 10169 21312 10474
rect 20732 10118 20852 10146
rect 21270 10160 21326 10169
rect 20628 9920 20680 9926
rect 19982 9888 20038 9897
rect 20628 9862 20680 9868
rect 19982 9823 20038 9832
rect 19798 7848 19854 7857
rect 19798 7783 19854 7792
rect 19996 7546 20024 9823
rect 20076 8560 20128 8566
rect 20076 8502 20128 8508
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 20088 7410 20116 8502
rect 20732 8294 20760 10118
rect 21270 10095 21326 10104
rect 21376 10062 21404 10542
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21836 10130 21864 10406
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 20824 9518 20852 9998
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21732 9988 21784 9994
rect 21732 9930 21784 9936
rect 21560 9761 21588 9930
rect 21744 9897 21772 9930
rect 21836 9926 21864 10066
rect 21824 9920 21876 9926
rect 21730 9888 21786 9897
rect 21824 9862 21876 9868
rect 21730 9823 21786 9832
rect 21546 9752 21602 9761
rect 21546 9687 21548 9696
rect 21600 9687 21602 9696
rect 21548 9658 21600 9664
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20916 8974 20944 9522
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 21008 8498 21036 9046
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20812 7880 20864 7886
rect 20864 7840 20944 7868
rect 20812 7822 20864 7828
rect 20444 7472 20496 7478
rect 20444 7414 20496 7420
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 19720 5302 19748 5646
rect 19904 5370 19932 7346
rect 20456 6866 20484 7414
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19996 5710 20024 6394
rect 20168 5840 20220 5846
rect 20168 5782 20220 5788
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19708 5296 19760 5302
rect 19708 5238 19760 5244
rect 19996 5234 20024 5646
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 20088 5098 20116 5646
rect 20180 5302 20208 5782
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20272 5370 20300 5646
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20168 5296 20220 5302
rect 20168 5238 20220 5244
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 20456 5030 20484 5170
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19628 3058 19656 3878
rect 19996 3534 20024 4218
rect 20548 3534 20576 7346
rect 20916 7002 20944 7840
rect 21008 7546 21036 8434
rect 21100 8362 21128 9318
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21284 8498 21312 8910
rect 21744 8498 21772 9522
rect 21928 9042 21956 10610
rect 22112 10198 22140 11018
rect 22296 10674 22324 11290
rect 22388 11098 22416 11716
rect 22652 11698 22704 11704
rect 22756 11354 22784 12174
rect 23032 11762 23060 14418
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24136 13938 24164 14214
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24216 13932 24268 13938
rect 24320 13920 24348 20318
rect 24504 18766 24532 21286
rect 24596 20942 24624 21286
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 24688 17270 24716 22918
rect 24872 22778 24900 23054
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24872 20466 24900 20810
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24964 20346 24992 27474
rect 25056 26790 25084 29038
rect 25504 28960 25556 28966
rect 25504 28902 25556 28908
rect 25412 28416 25464 28422
rect 25412 28358 25464 28364
rect 25424 28014 25452 28358
rect 25412 28008 25464 28014
rect 25412 27950 25464 27956
rect 25136 27872 25188 27878
rect 25136 27814 25188 27820
rect 25044 26784 25096 26790
rect 25044 26726 25096 26732
rect 25056 25158 25084 26726
rect 25044 25152 25096 25158
rect 25044 25094 25096 25100
rect 24780 20318 24992 20346
rect 24780 19446 24808 20318
rect 25056 19514 25084 25094
rect 25148 24954 25176 27814
rect 25516 27538 25544 28902
rect 25504 27532 25556 27538
rect 25504 27474 25556 27480
rect 25320 27464 25372 27470
rect 25240 27424 25320 27452
rect 25240 27334 25268 27424
rect 25320 27406 25372 27412
rect 25228 27328 25280 27334
rect 25228 27270 25280 27276
rect 25608 26450 25636 32286
rect 25792 31890 25820 32302
rect 25780 31884 25832 31890
rect 25780 31826 25832 31832
rect 25792 31754 25820 31826
rect 26160 31770 26188 33050
rect 25792 31726 25912 31754
rect 26160 31742 26280 31770
rect 25884 30802 25912 31726
rect 26252 31634 26280 31742
rect 26160 31606 26280 31634
rect 26160 31346 26188 31606
rect 26148 31340 26200 31346
rect 26148 31282 26200 31288
rect 26056 31272 26108 31278
rect 26108 31220 26188 31226
rect 26056 31214 26188 31220
rect 26068 31198 26188 31214
rect 26056 31136 26108 31142
rect 26056 31078 26108 31084
rect 26068 30938 26096 31078
rect 26056 30932 26108 30938
rect 26056 30874 26108 30880
rect 25780 30796 25832 30802
rect 25780 30738 25832 30744
rect 25872 30796 25924 30802
rect 25872 30738 25924 30744
rect 25792 30598 25820 30738
rect 25780 30592 25832 30598
rect 25780 30534 25832 30540
rect 25884 28762 25912 30738
rect 26068 30734 26096 30874
rect 26160 30734 26188 31198
rect 26056 30728 26108 30734
rect 26056 30670 26108 30676
rect 26148 30728 26200 30734
rect 26148 30670 26200 30676
rect 26240 30592 26292 30598
rect 26240 30534 26292 30540
rect 26148 30320 26200 30326
rect 26148 30262 26200 30268
rect 26160 28762 26188 30262
rect 25872 28756 25924 28762
rect 25872 28698 25924 28704
rect 26148 28756 26200 28762
rect 26148 28698 26200 28704
rect 25780 28552 25832 28558
rect 25780 28494 25832 28500
rect 25792 27538 25820 28494
rect 26056 28484 26108 28490
rect 26056 28426 26108 28432
rect 25964 28076 26016 28082
rect 25964 28018 26016 28024
rect 25780 27532 25832 27538
rect 25780 27474 25832 27480
rect 25596 26444 25648 26450
rect 25596 26386 25648 26392
rect 25504 25696 25556 25702
rect 25504 25638 25556 25644
rect 25516 25294 25544 25638
rect 25504 25288 25556 25294
rect 25504 25230 25556 25236
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 25228 24880 25280 24886
rect 25228 24822 25280 24828
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25148 21078 25176 23462
rect 25136 21072 25188 21078
rect 25136 21014 25188 21020
rect 25240 20890 25268 24822
rect 25412 24608 25464 24614
rect 25412 24550 25464 24556
rect 25424 24342 25452 24550
rect 25320 24336 25372 24342
rect 25318 24304 25320 24313
rect 25412 24336 25464 24342
rect 25372 24304 25374 24313
rect 25412 24278 25464 24284
rect 25318 24239 25374 24248
rect 25516 24188 25544 25230
rect 25596 24200 25648 24206
rect 25516 24160 25596 24188
rect 25596 24142 25648 24148
rect 25688 24200 25740 24206
rect 25688 24142 25740 24148
rect 25608 23730 25636 24142
rect 25700 23730 25728 24142
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 25318 23624 25374 23633
rect 25318 23559 25320 23568
rect 25372 23559 25374 23568
rect 25320 23530 25372 23536
rect 25332 23050 25360 23530
rect 25700 23118 25728 23666
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25504 22976 25556 22982
rect 25504 22918 25556 22924
rect 25516 22030 25544 22918
rect 25596 22432 25648 22438
rect 25596 22374 25648 22380
rect 25608 22098 25636 22374
rect 25596 22092 25648 22098
rect 25596 22034 25648 22040
rect 25504 22024 25556 22030
rect 25504 21966 25556 21972
rect 25320 21616 25372 21622
rect 25320 21558 25372 21564
rect 25148 20862 25268 20890
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24860 19372 24912 19378
rect 24860 19314 24912 19320
rect 24872 18850 24900 19314
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 24780 18822 24900 18850
rect 24780 18766 24808 18822
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24872 17610 24900 18158
rect 24964 17678 24992 19110
rect 25042 18864 25098 18873
rect 25042 18799 25044 18808
rect 25096 18799 25098 18808
rect 25044 18770 25096 18776
rect 25148 18426 25176 20862
rect 25332 20806 25360 21558
rect 25228 20800 25280 20806
rect 25228 20742 25280 20748
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25240 20262 25268 20742
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25792 19394 25820 27474
rect 25872 27328 25924 27334
rect 25872 27270 25924 27276
rect 25884 20602 25912 27270
rect 25976 27130 26004 28018
rect 25964 27124 26016 27130
rect 25964 27066 26016 27072
rect 25964 25900 26016 25906
rect 25964 25842 26016 25848
rect 25976 25294 26004 25842
rect 25964 25288 26016 25294
rect 25964 25230 26016 25236
rect 26068 24750 26096 28426
rect 26252 28218 26280 30534
rect 26436 28626 26464 33322
rect 26528 32570 26556 34478
rect 26608 34468 26660 34474
rect 26608 34410 26660 34416
rect 28632 34468 28684 34474
rect 28632 34410 28684 34416
rect 26620 34202 26648 34410
rect 26608 34196 26660 34202
rect 26608 34138 26660 34144
rect 26700 33516 26752 33522
rect 26700 33458 26752 33464
rect 26712 33114 26740 33458
rect 26884 33380 26936 33386
rect 26884 33322 26936 33328
rect 26700 33108 26752 33114
rect 26700 33050 26752 33056
rect 26896 32978 26924 33322
rect 28356 33312 28408 33318
rect 28356 33254 28408 33260
rect 26884 32972 26936 32978
rect 26884 32914 26936 32920
rect 27620 32972 27672 32978
rect 27620 32914 27672 32920
rect 28172 32972 28224 32978
rect 28172 32914 28224 32920
rect 26516 32564 26568 32570
rect 26516 32506 26568 32512
rect 26884 32360 26936 32366
rect 26884 32302 26936 32308
rect 26896 31822 26924 32302
rect 27632 32298 27660 32914
rect 27620 32292 27672 32298
rect 27620 32234 27672 32240
rect 27252 32224 27304 32230
rect 27252 32166 27304 32172
rect 26884 31816 26936 31822
rect 26884 31758 26936 31764
rect 26516 31136 26568 31142
rect 26516 31078 26568 31084
rect 26424 28620 26476 28626
rect 26424 28562 26476 28568
rect 26240 28212 26292 28218
rect 26240 28154 26292 28160
rect 26332 27328 26384 27334
rect 26332 27270 26384 27276
rect 26344 27130 26372 27270
rect 26436 27130 26464 28562
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 26424 27124 26476 27130
rect 26424 27066 26476 27072
rect 26436 25838 26464 27066
rect 26528 26042 26556 31078
rect 26608 30592 26660 30598
rect 26608 30534 26660 30540
rect 26516 26036 26568 26042
rect 26516 25978 26568 25984
rect 26424 25832 26476 25838
rect 26424 25774 26476 25780
rect 26240 25696 26292 25702
rect 26240 25638 26292 25644
rect 26252 25294 26280 25638
rect 26240 25288 26292 25294
rect 26240 25230 26292 25236
rect 26056 24744 26108 24750
rect 26056 24686 26108 24692
rect 26068 23746 26096 24686
rect 26238 24304 26294 24313
rect 26238 24239 26240 24248
rect 26292 24239 26294 24248
rect 26240 24210 26292 24216
rect 26148 23860 26200 23866
rect 26200 23820 26280 23848
rect 26148 23802 26200 23808
rect 25976 23718 26096 23746
rect 25976 22642 26004 23718
rect 26056 23656 26108 23662
rect 26056 23598 26108 23604
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 25962 21040 26018 21049
rect 25962 20975 25964 20984
rect 26016 20975 26018 20984
rect 25964 20946 26016 20952
rect 25872 20596 25924 20602
rect 25872 20538 25924 20544
rect 26068 19514 26096 23598
rect 26252 22982 26280 23820
rect 26436 23186 26464 25774
rect 26424 23180 26476 23186
rect 26424 23122 26476 23128
rect 26516 23180 26568 23186
rect 26516 23122 26568 23128
rect 26240 22976 26292 22982
rect 26240 22918 26292 22924
rect 26252 22234 26280 22918
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 26436 22094 26464 23122
rect 26528 22642 26556 23122
rect 26516 22636 26568 22642
rect 26516 22578 26568 22584
rect 26344 22066 26464 22094
rect 26344 21690 26372 22066
rect 26332 21684 26384 21690
rect 26332 21626 26384 21632
rect 26620 21010 26648 30534
rect 26896 29714 26924 31758
rect 27160 30048 27212 30054
rect 27160 29990 27212 29996
rect 26884 29708 26936 29714
rect 26884 29650 26936 29656
rect 27172 29646 27200 29990
rect 27160 29640 27212 29646
rect 27160 29582 27212 29588
rect 27264 28994 27292 32166
rect 28080 31816 28132 31822
rect 28080 31758 28132 31764
rect 27344 31748 27396 31754
rect 27344 31690 27396 31696
rect 27356 31482 27384 31690
rect 27896 31680 27948 31686
rect 27896 31622 27948 31628
rect 27908 31482 27936 31622
rect 27344 31476 27396 31482
rect 27344 31418 27396 31424
rect 27896 31476 27948 31482
rect 27896 31418 27948 31424
rect 28092 31414 28120 31758
rect 28080 31408 28132 31414
rect 28080 31350 28132 31356
rect 28092 30258 28120 31350
rect 28184 31278 28212 32914
rect 28368 32910 28396 33254
rect 28356 32904 28408 32910
rect 28356 32846 28408 32852
rect 28540 32428 28592 32434
rect 28540 32370 28592 32376
rect 28552 32026 28580 32370
rect 28540 32020 28592 32026
rect 28540 31962 28592 31968
rect 28644 31890 28672 34410
rect 28632 31884 28684 31890
rect 28632 31826 28684 31832
rect 28172 31272 28224 31278
rect 28172 31214 28224 31220
rect 28540 31272 28592 31278
rect 28540 31214 28592 31220
rect 27804 30252 27856 30258
rect 27804 30194 27856 30200
rect 28080 30252 28132 30258
rect 28080 30194 28132 30200
rect 27816 29850 27844 30194
rect 27988 30184 28040 30190
rect 27988 30126 28040 30132
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 27436 29300 27488 29306
rect 27436 29242 27488 29248
rect 27172 28966 27292 28994
rect 26792 27872 26844 27878
rect 26792 27814 26844 27820
rect 26804 27470 26832 27814
rect 26882 27568 26938 27577
rect 26882 27503 26884 27512
rect 26936 27503 26938 27512
rect 26884 27474 26936 27480
rect 26792 27464 26844 27470
rect 26792 27406 26844 27412
rect 26792 27328 26844 27334
rect 26792 27270 26844 27276
rect 26804 26994 26832 27270
rect 26896 27130 26924 27474
rect 26884 27124 26936 27130
rect 26884 27066 26936 27072
rect 26792 26988 26844 26994
rect 26792 26930 26844 26936
rect 26792 24200 26844 24206
rect 26792 24142 26844 24148
rect 26804 23798 26832 24142
rect 26976 24064 27028 24070
rect 26976 24006 27028 24012
rect 26792 23792 26844 23798
rect 26792 23734 26844 23740
rect 26988 23730 27016 24006
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 26608 21004 26660 21010
rect 26608 20946 26660 20952
rect 26332 20936 26384 20942
rect 26332 20878 26384 20884
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26148 20800 26200 20806
rect 26148 20742 26200 20748
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 25870 19408 25926 19417
rect 25412 19372 25464 19378
rect 25792 19366 25870 19394
rect 25870 19343 25872 19352
rect 25412 19314 25464 19320
rect 25924 19343 25926 19352
rect 25872 19314 25924 19320
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 25332 18630 25360 18702
rect 25320 18624 25372 18630
rect 25320 18566 25372 18572
rect 25424 18426 25452 19314
rect 25688 19304 25740 19310
rect 25688 19246 25740 19252
rect 25596 19168 25648 19174
rect 25596 19110 25648 19116
rect 25608 18834 25636 19110
rect 25596 18828 25648 18834
rect 25596 18770 25648 18776
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 25056 17882 25084 18226
rect 25700 18086 25728 19246
rect 25884 18737 25912 19314
rect 26068 19281 26096 19450
rect 26054 19272 26110 19281
rect 26054 19207 26110 19216
rect 26160 19156 26188 20742
rect 26344 20534 26372 20878
rect 26516 20800 26568 20806
rect 26516 20742 26568 20748
rect 26240 20528 26292 20534
rect 26240 20470 26292 20476
rect 26332 20528 26384 20534
rect 26332 20470 26384 20476
rect 26068 19128 26188 19156
rect 25870 18728 25926 18737
rect 25870 18663 25926 18672
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25688 18080 25740 18086
rect 25688 18022 25740 18028
rect 25044 17876 25096 17882
rect 25044 17818 25096 17824
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 25148 17134 25176 17818
rect 25976 17762 26004 18226
rect 25884 17734 26004 17762
rect 25884 17678 25912 17734
rect 25872 17672 25924 17678
rect 25872 17614 25924 17620
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24872 16250 24900 16526
rect 25884 16250 25912 17614
rect 26068 16454 26096 19128
rect 26252 18970 26280 20470
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 26344 19446 26372 19654
rect 26332 19440 26384 19446
rect 26332 19382 26384 19388
rect 26424 19168 26476 19174
rect 26422 19136 26424 19145
rect 26476 19136 26478 19145
rect 26422 19071 26478 19080
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 26146 18864 26202 18873
rect 26146 18799 26202 18808
rect 26160 18698 26188 18799
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 26424 17604 26476 17610
rect 26424 17546 26476 17552
rect 26252 17338 26280 17546
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 26436 17202 26464 17546
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26332 16516 26384 16522
rect 26332 16458 26384 16464
rect 26056 16448 26108 16454
rect 26056 16390 26108 16396
rect 26344 16250 26372 16458
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 25872 16244 25924 16250
rect 25872 16186 25924 16192
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26148 16176 26200 16182
rect 26148 16118 26200 16124
rect 25872 16108 25924 16114
rect 25872 16050 25924 16056
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 24400 15360 24452 15366
rect 24400 15302 24452 15308
rect 24268 13892 24348 13920
rect 24216 13874 24268 13880
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 23860 13462 23888 13670
rect 24044 13530 24072 13874
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 23400 12434 23428 13126
rect 24044 12434 24072 13330
rect 23400 12406 23520 12434
rect 23112 12232 23164 12238
rect 23112 12174 23164 12180
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 22836 11688 22888 11694
rect 22836 11630 22888 11636
rect 22928 11688 22980 11694
rect 23124 11642 23152 12174
rect 22928 11630 22980 11636
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 22388 11070 22508 11098
rect 22848 11082 22876 11630
rect 22940 11150 22968 11630
rect 23032 11626 23152 11642
rect 23020 11620 23152 11626
rect 23072 11614 23152 11620
rect 23020 11562 23072 11568
rect 23032 11218 23060 11562
rect 23020 11212 23072 11218
rect 23020 11154 23072 11160
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22388 10266 22416 10950
rect 22376 10260 22428 10266
rect 22376 10202 22428 10208
rect 22100 10192 22152 10198
rect 22100 10134 22152 10140
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 22020 9674 22048 10066
rect 22480 9926 22508 11070
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 22560 10192 22612 10198
rect 22560 10134 22612 10140
rect 22468 9920 22520 9926
rect 22468 9862 22520 9868
rect 22020 9646 22140 9674
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 22020 9110 22048 9386
rect 22112 9178 22140 9646
rect 22572 9518 22600 10134
rect 23032 10010 23060 11154
rect 23296 10464 23348 10470
rect 23296 10406 23348 10412
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 23216 10062 23244 10202
rect 22940 9982 23060 10010
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 22652 9920 22704 9926
rect 22652 9862 22704 9868
rect 22664 9722 22692 9862
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22940 9450 22968 9982
rect 23124 9926 23152 9998
rect 23308 9994 23336 10406
rect 23296 9988 23348 9994
rect 23296 9930 23348 9936
rect 23020 9920 23072 9926
rect 23020 9862 23072 9868
rect 23112 9920 23164 9926
rect 23112 9862 23164 9868
rect 23032 9654 23060 9862
rect 23020 9648 23072 9654
rect 23020 9590 23072 9596
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22008 9104 22060 9110
rect 22008 9046 22060 9052
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21088 8356 21140 8362
rect 21088 8298 21140 8304
rect 21100 7818 21128 8298
rect 21272 7948 21324 7954
rect 21272 7890 21324 7896
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21284 7546 21312 7890
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21284 7410 21312 7482
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20720 6316 20772 6322
rect 20824 6304 20852 6734
rect 20772 6276 20852 6304
rect 20720 6258 20772 6264
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20640 5710 20668 6054
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20640 5302 20668 5646
rect 20628 5296 20680 5302
rect 20628 5238 20680 5244
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 20088 3058 20116 3334
rect 20548 3074 20576 3470
rect 20824 3398 20852 6276
rect 20916 5642 20944 6938
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21192 5710 21220 6054
rect 21376 5914 21404 7822
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21468 7410 21496 7686
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21652 7206 21680 7822
rect 21640 7200 21692 7206
rect 21640 7142 21692 7148
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 21560 5234 21588 5646
rect 21744 5642 21772 8434
rect 21928 8022 21956 8978
rect 22112 8498 22140 9114
rect 22940 9042 22968 9386
rect 23216 9110 23244 9454
rect 23204 9104 23256 9110
rect 23204 9046 23256 9052
rect 22928 9036 22980 9042
rect 22928 8978 22980 8984
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22572 8634 22600 8910
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22100 8492 22152 8498
rect 22020 8452 22100 8480
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21836 6662 21864 7822
rect 22020 7478 22048 8452
rect 22100 8434 22152 8440
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 22848 7886 22876 8434
rect 23492 7886 23520 12406
rect 23952 12406 24072 12434
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 23768 11898 23796 12106
rect 23756 11892 23808 11898
rect 23756 11834 23808 11840
rect 23768 11762 23796 11834
rect 23756 11756 23808 11762
rect 23756 11698 23808 11704
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23768 11354 23796 11698
rect 23756 11348 23808 11354
rect 23756 11290 23808 11296
rect 23860 10470 23888 11698
rect 23952 10674 23980 12406
rect 24136 12374 24164 13874
rect 24412 13512 24440 15302
rect 24504 14346 24532 15438
rect 25136 15428 25188 15434
rect 25136 15370 25188 15376
rect 25148 15162 25176 15370
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25424 15026 25452 15846
rect 25884 15366 25912 16050
rect 26160 15502 26188 16118
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25688 15088 25740 15094
rect 25688 15030 25740 15036
rect 25412 15020 25464 15026
rect 25412 14962 25464 14968
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 24492 14340 24544 14346
rect 24492 14282 24544 14288
rect 24228 13484 24440 13512
rect 24228 12646 24256 13484
rect 24308 13252 24360 13258
rect 24308 13194 24360 13200
rect 24320 12850 24348 13194
rect 24768 13184 24820 13190
rect 24768 13126 24820 13132
rect 24780 12986 24808 13126
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 24032 12368 24084 12374
rect 24032 12310 24084 12316
rect 24124 12368 24176 12374
rect 24124 12310 24176 12316
rect 24044 11762 24072 12310
rect 24228 12238 24256 12582
rect 24596 12434 24624 12922
rect 24504 12406 24624 12434
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 24136 11801 24164 12174
rect 24400 12164 24452 12170
rect 24400 12106 24452 12112
rect 24412 11830 24440 12106
rect 24400 11824 24452 11830
rect 24122 11792 24178 11801
rect 24032 11756 24084 11762
rect 24400 11766 24452 11772
rect 24122 11727 24178 11736
rect 24032 11698 24084 11704
rect 24136 11694 24164 11727
rect 24124 11688 24176 11694
rect 24124 11630 24176 11636
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23676 9722 23704 9998
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23584 9178 23612 9522
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 23676 9058 23704 9658
rect 23584 9030 23704 9058
rect 23584 8974 23612 9030
rect 23952 8974 23980 9862
rect 24032 9512 24084 9518
rect 24032 9454 24084 9460
rect 24044 9178 24072 9454
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 23584 8430 23612 8910
rect 23952 8634 23980 8910
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 23572 8424 23624 8430
rect 23572 8366 23624 8372
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 22376 7812 22428 7818
rect 22376 7754 22428 7760
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22008 7472 22060 7478
rect 22008 7414 22060 7420
rect 22204 7410 22232 7686
rect 22388 7410 22416 7754
rect 22756 7546 22784 7822
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 21928 6798 21956 7142
rect 22020 7002 22048 7142
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 22112 6866 22140 7346
rect 22376 7268 22428 7274
rect 22376 7210 22428 7216
rect 22388 6866 22416 7210
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21836 6322 21864 6598
rect 21928 6322 21956 6734
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 22020 6458 22048 6666
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22112 6458 22140 6598
rect 22008 6452 22060 6458
rect 22008 6394 22060 6400
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 22112 6322 22140 6394
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21916 6316 21968 6322
rect 21916 6258 21968 6264
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 21732 5636 21784 5642
rect 21732 5578 21784 5584
rect 21836 5370 21864 5646
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21088 5092 21140 5098
rect 21088 5034 21140 5040
rect 21100 3602 21128 5034
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21376 4282 21404 4558
rect 21928 4434 21956 6258
rect 22008 5636 22060 5642
rect 22008 5578 22060 5584
rect 22020 5250 22048 5578
rect 22112 5370 22140 6258
rect 22480 5914 22508 6734
rect 22560 6724 22612 6730
rect 22560 6666 22612 6672
rect 22572 6322 22600 6666
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22572 5914 22600 6258
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22204 5574 22232 5646
rect 22284 5636 22336 5642
rect 22284 5578 22336 5584
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 22296 5250 22324 5578
rect 22020 5222 22324 5250
rect 22008 5160 22060 5166
rect 22008 5102 22060 5108
rect 22020 4622 22048 5102
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 21928 4406 22048 4434
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 21088 3596 21140 3602
rect 21088 3538 21140 3544
rect 20916 3398 20944 3538
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20824 3194 20852 3334
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20364 3058 20576 3074
rect 19616 3052 19668 3058
rect 19616 2994 19668 3000
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 20352 3052 20576 3058
rect 20404 3046 20576 3052
rect 20352 2994 20404 3000
rect 21100 2990 21128 3538
rect 21560 3534 21588 3878
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 21836 3194 21864 4082
rect 22020 3738 22048 4406
rect 22008 3732 22060 3738
rect 22008 3674 22060 3680
rect 22020 3194 22048 3674
rect 22112 3602 22140 5222
rect 22480 4078 22508 5850
rect 22664 5166 22692 6258
rect 22848 5642 22876 7822
rect 23492 7546 23520 7822
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 23572 7336 23624 7342
rect 23572 7278 23624 7284
rect 23584 7002 23612 7278
rect 23572 6996 23624 7002
rect 23572 6938 23624 6944
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23676 5710 23704 6054
rect 23860 5710 23888 7414
rect 23952 7206 23980 8570
rect 24136 8242 24164 11290
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24228 9586 24256 10610
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 24228 8362 24256 9522
rect 24216 8356 24268 8362
rect 24216 8298 24268 8304
rect 24136 8214 24256 8242
rect 24124 7812 24176 7818
rect 24124 7754 24176 7760
rect 24136 7546 24164 7754
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24228 7342 24256 8214
rect 24320 7410 24348 10950
rect 24400 10056 24452 10062
rect 24400 9998 24452 10004
rect 24412 9761 24440 9998
rect 24398 9752 24454 9761
rect 24398 9687 24454 9696
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 24228 6458 24256 7278
rect 24216 6452 24268 6458
rect 24136 6412 24216 6440
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 23664 5704 23716 5710
rect 23664 5646 23716 5652
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 22836 5636 22888 5642
rect 22836 5578 22888 5584
rect 22652 5160 22704 5166
rect 23860 5148 23888 5646
rect 23952 5370 23980 6258
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 24136 5166 24164 6412
rect 24216 6394 24268 6400
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 24228 5914 24256 6190
rect 24216 5908 24268 5914
rect 24216 5850 24268 5856
rect 24228 5302 24256 5850
rect 24216 5296 24268 5302
rect 24216 5238 24268 5244
rect 23940 5160 23992 5166
rect 23860 5120 23940 5148
rect 22652 5102 22704 5108
rect 23940 5102 23992 5108
rect 24124 5160 24176 5166
rect 24124 5102 24176 5108
rect 23848 4548 23900 4554
rect 23848 4490 23900 4496
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 22664 3194 22692 3470
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22848 3058 22876 3878
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 22940 2922 22968 4218
rect 23480 4208 23532 4214
rect 23480 4150 23532 4156
rect 23492 3738 23520 4150
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 23400 3126 23428 3334
rect 23388 3120 23440 3126
rect 23388 3062 23440 3068
rect 22928 2916 22980 2922
rect 22928 2858 22980 2864
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 23860 2446 23888 4490
rect 23952 4146 23980 5102
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 24504 3738 24532 12406
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24596 11218 24624 11698
rect 24584 11212 24636 11218
rect 24584 11154 24636 11160
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 24688 9586 24716 10406
rect 24780 10169 24808 10474
rect 24766 10160 24822 10169
rect 24766 10095 24768 10104
rect 24820 10095 24822 10104
rect 24768 10066 24820 10072
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 24872 9450 24900 14894
rect 25424 14550 25452 14962
rect 25412 14544 25464 14550
rect 25412 14486 25464 14492
rect 25412 14408 25464 14414
rect 25412 14350 25464 14356
rect 25424 14074 25452 14350
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25502 13832 25558 13841
rect 25502 13767 25504 13776
rect 25556 13767 25558 13776
rect 25504 13738 25556 13744
rect 25516 13394 25544 13738
rect 25504 13388 25556 13394
rect 25504 13330 25556 13336
rect 25596 13184 25648 13190
rect 25410 13152 25466 13161
rect 25596 13126 25648 13132
rect 25410 13087 25466 13096
rect 25424 12782 25452 13087
rect 25608 12850 25636 13126
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25412 12776 25464 12782
rect 25412 12718 25464 12724
rect 25700 11286 25728 15030
rect 25884 13938 25912 15302
rect 26160 14482 26188 15438
rect 26148 14476 26200 14482
rect 26148 14418 26200 14424
rect 26424 14408 26476 14414
rect 26528 14396 26556 20742
rect 26804 20505 26832 20878
rect 26790 20496 26846 20505
rect 26790 20431 26846 20440
rect 26988 19378 27016 21490
rect 27068 21140 27120 21146
rect 27068 21082 27120 21088
rect 27080 20856 27108 21082
rect 27172 21078 27200 28966
rect 27448 28626 27476 29242
rect 27528 29096 27580 29102
rect 27580 29044 27660 29050
rect 27528 29038 27660 29044
rect 27540 29022 27660 29038
rect 27436 28620 27488 28626
rect 27436 28562 27488 28568
rect 27528 28620 27580 28626
rect 27528 28562 27580 28568
rect 27540 28150 27568 28562
rect 27632 28558 27660 29022
rect 28000 28694 28028 30126
rect 27988 28688 28040 28694
rect 27988 28630 28040 28636
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27632 28150 27660 28494
rect 27528 28144 27580 28150
rect 27528 28086 27580 28092
rect 27620 28144 27672 28150
rect 27620 28086 27672 28092
rect 27896 27872 27948 27878
rect 27896 27814 27948 27820
rect 27908 27470 27936 27814
rect 28000 27606 28028 28630
rect 27988 27600 28040 27606
rect 27988 27542 28040 27548
rect 27896 27464 27948 27470
rect 27896 27406 27948 27412
rect 27988 27464 28040 27470
rect 27988 27406 28040 27412
rect 27344 25900 27396 25906
rect 27344 25842 27396 25848
rect 27356 25498 27384 25842
rect 27528 25832 27580 25838
rect 27528 25774 27580 25780
rect 27344 25492 27396 25498
rect 27344 25434 27396 25440
rect 27540 24818 27568 25774
rect 27896 25696 27948 25702
rect 27896 25638 27948 25644
rect 27908 25294 27936 25638
rect 28000 25498 28028 27406
rect 28092 26790 28120 30194
rect 28448 30048 28500 30054
rect 28448 29990 28500 29996
rect 28264 29844 28316 29850
rect 28264 29786 28316 29792
rect 28276 29170 28304 29786
rect 28460 29170 28488 29990
rect 28172 29164 28224 29170
rect 28172 29106 28224 29112
rect 28264 29164 28316 29170
rect 28264 29106 28316 29112
rect 28448 29164 28500 29170
rect 28448 29106 28500 29112
rect 28184 28966 28212 29106
rect 28172 28960 28224 28966
rect 28172 28902 28224 28908
rect 28184 28626 28212 28902
rect 28172 28620 28224 28626
rect 28276 28608 28304 29106
rect 28448 28620 28500 28626
rect 28276 28580 28448 28608
rect 28172 28562 28224 28568
rect 28448 28562 28500 28568
rect 28080 26784 28132 26790
rect 28080 26726 28132 26732
rect 28448 26784 28500 26790
rect 28448 26726 28500 26732
rect 28080 25900 28132 25906
rect 28080 25842 28132 25848
rect 27988 25492 28040 25498
rect 27988 25434 28040 25440
rect 27896 25288 27948 25294
rect 27896 25230 27948 25236
rect 28092 24954 28120 25842
rect 28264 25152 28316 25158
rect 28264 25094 28316 25100
rect 28276 24954 28304 25094
rect 28080 24948 28132 24954
rect 28080 24890 28132 24896
rect 28264 24948 28316 24954
rect 28264 24890 28316 24896
rect 27528 24812 27580 24818
rect 27528 24754 27580 24760
rect 28172 24744 28224 24750
rect 28172 24686 28224 24692
rect 27528 24676 27580 24682
rect 27528 24618 27580 24624
rect 27540 24274 27568 24618
rect 27804 24608 27856 24614
rect 27804 24550 27856 24556
rect 27528 24268 27580 24274
rect 27528 24210 27580 24216
rect 27540 23746 27568 24210
rect 27816 24206 27844 24550
rect 28184 24274 28212 24686
rect 27988 24268 28040 24274
rect 27988 24210 28040 24216
rect 28172 24268 28224 24274
rect 28172 24210 28224 24216
rect 27804 24200 27856 24206
rect 27804 24142 27856 24148
rect 28000 23866 28028 24210
rect 28276 24070 28304 24890
rect 28356 24744 28408 24750
rect 28460 24698 28488 26726
rect 28552 26382 28580 31214
rect 28632 28552 28684 28558
rect 28632 28494 28684 28500
rect 28644 28422 28672 28494
rect 28632 28416 28684 28422
rect 28632 28358 28684 28364
rect 28632 27940 28684 27946
rect 28632 27882 28684 27888
rect 28644 27130 28672 27882
rect 28632 27124 28684 27130
rect 28632 27066 28684 27072
rect 28540 26376 28592 26382
rect 28540 26318 28592 26324
rect 28408 24692 28488 24698
rect 28356 24686 28488 24692
rect 28368 24670 28488 24686
rect 28264 24064 28316 24070
rect 28264 24006 28316 24012
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 27540 23730 27936 23746
rect 28000 23730 28028 23802
rect 27540 23724 27948 23730
rect 27540 23718 27896 23724
rect 27896 23666 27948 23672
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 27528 23656 27580 23662
rect 27528 23598 27580 23604
rect 27618 23624 27674 23633
rect 27540 23474 27568 23598
rect 27618 23559 27620 23568
rect 27672 23559 27674 23568
rect 27620 23530 27672 23536
rect 27988 23520 28040 23526
rect 27540 23446 27752 23474
rect 27988 23462 28040 23468
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27632 22778 27660 23054
rect 27620 22772 27672 22778
rect 27620 22714 27672 22720
rect 27724 22710 27752 23446
rect 27804 23112 27856 23118
rect 27804 23054 27856 23060
rect 27712 22704 27764 22710
rect 27712 22646 27764 22652
rect 27160 21072 27212 21078
rect 27160 21014 27212 21020
rect 27816 21010 27844 23054
rect 28000 21146 28028 23462
rect 28356 22976 28408 22982
rect 28356 22918 28408 22924
rect 28368 22710 28396 22918
rect 28356 22704 28408 22710
rect 28356 22646 28408 22652
rect 28460 22574 28488 24670
rect 28448 22568 28500 22574
rect 28448 22510 28500 22516
rect 28460 21690 28488 22510
rect 28448 21684 28500 21690
rect 28448 21626 28500 21632
rect 28632 21548 28684 21554
rect 28632 21490 28684 21496
rect 28644 21146 28672 21490
rect 27988 21140 28040 21146
rect 27988 21082 28040 21088
rect 28632 21140 28684 21146
rect 28632 21082 28684 21088
rect 27804 21004 27856 21010
rect 27804 20946 27856 20952
rect 27160 20868 27212 20874
rect 27080 20828 27160 20856
rect 27160 20810 27212 20816
rect 27172 20602 27200 20810
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 28092 20602 28120 20742
rect 27160 20596 27212 20602
rect 27160 20538 27212 20544
rect 28080 20596 28132 20602
rect 28080 20538 28132 20544
rect 28632 19848 28684 19854
rect 28632 19790 28684 19796
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27068 19304 27120 19310
rect 27066 19272 27068 19281
rect 27120 19272 27122 19281
rect 27066 19207 27122 19216
rect 27356 18766 27384 19314
rect 27528 19304 27580 19310
rect 27528 19246 27580 19252
rect 28080 19304 28132 19310
rect 28540 19304 28592 19310
rect 28080 19246 28132 19252
rect 28354 19272 28410 19281
rect 27540 18766 27568 19246
rect 28092 18834 28120 19246
rect 28540 19246 28592 19252
rect 28354 19207 28410 19216
rect 28368 19174 28396 19207
rect 28264 19168 28316 19174
rect 28264 19110 28316 19116
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 27896 18828 27948 18834
rect 27896 18770 27948 18776
rect 28080 18828 28132 18834
rect 28080 18770 28132 18776
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 27344 18760 27396 18766
rect 27344 18702 27396 18708
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 26988 18465 27016 18702
rect 26974 18456 27030 18465
rect 26974 18391 27030 18400
rect 26884 18216 26936 18222
rect 26884 18158 26936 18164
rect 26476 14368 26556 14396
rect 26424 14350 26476 14356
rect 26424 14272 26476 14278
rect 26424 14214 26476 14220
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 26332 13388 26384 13394
rect 26332 13330 26384 13336
rect 26148 13184 26200 13190
rect 26146 13152 26148 13161
rect 26240 13184 26292 13190
rect 26200 13152 26202 13161
rect 26240 13126 26292 13132
rect 26146 13087 26202 13096
rect 26160 12850 26188 13087
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26252 12102 26280 13126
rect 26240 12096 26292 12102
rect 26240 12038 26292 12044
rect 25044 11280 25096 11286
rect 25044 11222 25096 11228
rect 25688 11280 25740 11286
rect 25688 11222 25740 11228
rect 25056 10674 25084 11222
rect 25412 11076 25464 11082
rect 25412 11018 25464 11024
rect 25044 10668 25096 10674
rect 24964 10628 25044 10656
rect 24964 9926 24992 10628
rect 25044 10610 25096 10616
rect 25424 10606 25452 11018
rect 26344 11014 26372 13330
rect 26332 11008 26384 11014
rect 26332 10950 26384 10956
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 25044 10532 25096 10538
rect 25044 10474 25096 10480
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24964 9654 24992 9862
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 24860 9444 24912 9450
rect 24860 9386 24912 9392
rect 25056 7886 25084 10474
rect 25148 9586 25176 10542
rect 25964 10124 26016 10130
rect 25964 10066 26016 10072
rect 25976 9586 26004 10066
rect 26056 9988 26108 9994
rect 26056 9930 26108 9936
rect 26068 9722 26096 9930
rect 26056 9716 26108 9722
rect 26056 9658 26108 9664
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25148 8974 25176 9522
rect 26436 9382 26464 14214
rect 26896 11150 26924 18158
rect 27908 18154 27936 18770
rect 28276 18766 28304 19110
rect 28552 19009 28580 19246
rect 28538 19000 28594 19009
rect 28538 18935 28594 18944
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28356 18760 28408 18766
rect 28356 18702 28408 18708
rect 28446 18728 28502 18737
rect 27896 18148 27948 18154
rect 27896 18090 27948 18096
rect 28172 17536 28224 17542
rect 28172 17478 28224 17484
rect 27712 17264 27764 17270
rect 27712 17206 27764 17212
rect 27724 16794 27752 17206
rect 27712 16788 27764 16794
rect 27712 16730 27764 16736
rect 28184 16658 28212 17478
rect 28276 17338 28304 18702
rect 28368 17678 28396 18702
rect 28446 18663 28502 18672
rect 28460 18426 28488 18663
rect 28538 18456 28594 18465
rect 28448 18420 28500 18426
rect 28538 18391 28594 18400
rect 28448 18362 28500 18368
rect 28552 18358 28580 18391
rect 28540 18352 28592 18358
rect 28540 18294 28592 18300
rect 28644 18222 28672 19790
rect 28632 18216 28684 18222
rect 28632 18158 28684 18164
rect 28644 18086 28672 18158
rect 28632 18080 28684 18086
rect 28632 18022 28684 18028
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 28264 17332 28316 17338
rect 28264 17274 28316 17280
rect 27804 16652 27856 16658
rect 27804 16594 27856 16600
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 26988 15706 27016 16050
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 27252 15564 27304 15570
rect 27252 15506 27304 15512
rect 27264 15162 27292 15506
rect 27436 15496 27488 15502
rect 27436 15438 27488 15444
rect 27252 15156 27304 15162
rect 27252 15098 27304 15104
rect 27448 15026 27476 15438
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27436 15020 27488 15026
rect 27436 14962 27488 14968
rect 27160 14816 27212 14822
rect 27160 14758 27212 14764
rect 26976 14340 27028 14346
rect 26976 14282 27028 14288
rect 26988 14074 27016 14282
rect 26976 14068 27028 14074
rect 26976 14010 27028 14016
rect 27172 13938 27200 14758
rect 27448 14618 27476 14962
rect 27540 14958 27568 15302
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27540 14804 27568 14894
rect 27540 14776 27660 14804
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 27160 13320 27212 13326
rect 27160 13262 27212 13268
rect 27172 12442 27200 13262
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27264 12850 27292 13126
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27632 12646 27660 14776
rect 27620 12640 27672 12646
rect 27620 12582 27672 12588
rect 27160 12436 27212 12442
rect 27160 12378 27212 12384
rect 27816 12170 27844 16594
rect 28276 16590 28304 17274
rect 28264 16584 28316 16590
rect 28264 16526 28316 16532
rect 28448 15904 28500 15910
rect 28448 15846 28500 15852
rect 28460 15570 28488 15846
rect 28448 15564 28500 15570
rect 28448 15506 28500 15512
rect 28632 15496 28684 15502
rect 28632 15438 28684 15444
rect 28264 15360 28316 15366
rect 28264 15302 28316 15308
rect 27988 14884 28040 14890
rect 27988 14826 28040 14832
rect 28000 14618 28028 14826
rect 27988 14612 28040 14618
rect 27988 14554 28040 14560
rect 28172 14476 28224 14482
rect 28172 14418 28224 14424
rect 28184 14006 28212 14418
rect 28172 14000 28224 14006
rect 28172 13942 28224 13948
rect 28184 13870 28212 13942
rect 28172 13864 28224 13870
rect 28172 13806 28224 13812
rect 27988 13728 28040 13734
rect 27988 13670 28040 13676
rect 28000 13190 28028 13670
rect 27988 13184 28040 13190
rect 27988 13126 28040 13132
rect 28184 12918 28212 13806
rect 28276 12986 28304 15302
rect 28644 15094 28672 15438
rect 28632 15088 28684 15094
rect 28632 15030 28684 15036
rect 28448 13932 28500 13938
rect 28448 13874 28500 13880
rect 28460 13530 28488 13874
rect 28540 13728 28592 13734
rect 28540 13670 28592 13676
rect 28448 13524 28500 13530
rect 28448 13466 28500 13472
rect 28552 13190 28580 13670
rect 28448 13184 28500 13190
rect 28448 13126 28500 13132
rect 28540 13184 28592 13190
rect 28540 13126 28592 13132
rect 28460 12986 28488 13126
rect 28264 12980 28316 12986
rect 28264 12922 28316 12928
rect 28448 12980 28500 12986
rect 28448 12922 28500 12928
rect 28172 12912 28224 12918
rect 28172 12854 28224 12860
rect 27988 12640 28040 12646
rect 27988 12582 28040 12588
rect 28000 12238 28028 12582
rect 27988 12232 28040 12238
rect 27988 12174 28040 12180
rect 27804 12164 27856 12170
rect 27804 12106 27856 12112
rect 27988 12096 28040 12102
rect 27988 12038 28040 12044
rect 28000 11150 28028 12038
rect 28736 11257 28764 35866
rect 29288 35698 29316 36178
rect 29932 36174 29960 37334
rect 34808 37262 34836 39280
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 36176 37256 36228 37262
rect 36176 37198 36228 37204
rect 31484 37188 31536 37194
rect 31484 37130 31536 37136
rect 30104 37120 30156 37126
rect 30104 37062 30156 37068
rect 30116 36854 30144 37062
rect 30104 36848 30156 36854
rect 30104 36790 30156 36796
rect 30840 36644 30892 36650
rect 30840 36586 30892 36592
rect 30288 36372 30340 36378
rect 30288 36314 30340 36320
rect 29920 36168 29972 36174
rect 29920 36110 29972 36116
rect 30196 35828 30248 35834
rect 30196 35770 30248 35776
rect 29276 35692 29328 35698
rect 29276 35634 29328 35640
rect 29736 35692 29788 35698
rect 29736 35634 29788 35640
rect 29288 34678 29316 35634
rect 29748 35290 29776 35634
rect 29736 35284 29788 35290
rect 29736 35226 29788 35232
rect 30208 35154 30236 35770
rect 30300 35154 30328 36314
rect 30852 36174 30880 36586
rect 30840 36168 30892 36174
rect 30838 36136 30840 36145
rect 30892 36136 30894 36145
rect 30838 36071 30894 36080
rect 30564 35488 30616 35494
rect 30564 35430 30616 35436
rect 30196 35148 30248 35154
rect 30196 35090 30248 35096
rect 30288 35148 30340 35154
rect 30288 35090 30340 35096
rect 30104 34944 30156 34950
rect 30104 34886 30156 34892
rect 29276 34672 29328 34678
rect 29276 34614 29328 34620
rect 29276 32224 29328 32230
rect 29276 32166 29328 32172
rect 29368 32224 29420 32230
rect 29368 32166 29420 32172
rect 29288 31346 29316 32166
rect 29380 31754 29408 32166
rect 29828 31816 29880 31822
rect 29828 31758 29880 31764
rect 29368 31748 29420 31754
rect 29368 31690 29420 31696
rect 29276 31340 29328 31346
rect 29276 31282 29328 31288
rect 29380 31142 29408 31690
rect 29644 31680 29696 31686
rect 29644 31622 29696 31628
rect 29656 31414 29684 31622
rect 29644 31408 29696 31414
rect 29644 31350 29696 31356
rect 29368 31136 29420 31142
rect 29368 31078 29420 31084
rect 29840 30938 29868 31758
rect 30012 31680 30064 31686
rect 30012 31622 30064 31628
rect 29828 30932 29880 30938
rect 29828 30874 29880 30880
rect 30024 30598 30052 31622
rect 29828 30592 29880 30598
rect 29828 30534 29880 30540
rect 30012 30592 30064 30598
rect 30012 30534 30064 30540
rect 29368 29640 29420 29646
rect 29368 29582 29420 29588
rect 29380 29306 29408 29582
rect 29368 29300 29420 29306
rect 29368 29242 29420 29248
rect 29840 29102 29868 30534
rect 29920 29504 29972 29510
rect 29920 29446 29972 29452
rect 29932 29306 29960 29446
rect 29920 29300 29972 29306
rect 29920 29242 29972 29248
rect 29828 29096 29880 29102
rect 29828 29038 29880 29044
rect 29092 29028 29144 29034
rect 29092 28970 29144 28976
rect 28816 28960 28868 28966
rect 28816 28902 28868 28908
rect 28828 28626 28856 28902
rect 28816 28620 28868 28626
rect 28816 28562 28868 28568
rect 28908 28144 28960 28150
rect 28908 28086 28960 28092
rect 28816 28008 28868 28014
rect 28816 27950 28868 27956
rect 28828 26994 28856 27950
rect 28920 27674 28948 28086
rect 28908 27668 28960 27674
rect 28908 27610 28960 27616
rect 28816 26988 28868 26994
rect 28816 26930 28868 26936
rect 29104 26858 29132 28970
rect 29840 28422 29868 29038
rect 29276 28416 29328 28422
rect 29276 28358 29328 28364
rect 29828 28416 29880 28422
rect 29828 28358 29880 28364
rect 29092 26852 29144 26858
rect 29092 26794 29144 26800
rect 29092 25220 29144 25226
rect 29092 25162 29144 25168
rect 29104 24614 29132 25162
rect 29092 24608 29144 24614
rect 29092 24550 29144 24556
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 29184 23724 29236 23730
rect 29184 23666 29236 23672
rect 28814 23488 28870 23497
rect 28814 23423 28870 23432
rect 28828 19310 28856 23423
rect 28920 23118 28948 23666
rect 29196 23322 29224 23666
rect 29184 23316 29236 23322
rect 29184 23258 29236 23264
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 29288 20602 29316 28358
rect 29840 26858 29868 28358
rect 29828 26852 29880 26858
rect 29828 26794 29880 26800
rect 29368 25288 29420 25294
rect 29368 25230 29420 25236
rect 29380 24954 29408 25230
rect 29840 24954 29868 26794
rect 30012 25832 30064 25838
rect 30012 25774 30064 25780
rect 29368 24948 29420 24954
rect 29368 24890 29420 24896
rect 29828 24948 29880 24954
rect 29828 24890 29880 24896
rect 29736 21344 29788 21350
rect 29736 21286 29788 21292
rect 29748 20942 29776 21286
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29276 20596 29328 20602
rect 29276 20538 29328 20544
rect 29184 20528 29236 20534
rect 29184 20470 29236 20476
rect 28816 19304 28868 19310
rect 28816 19246 28868 19252
rect 29196 18970 29224 20470
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29748 19446 29776 19654
rect 29736 19440 29788 19446
rect 29736 19382 29788 19388
rect 29552 19372 29604 19378
rect 29552 19314 29604 19320
rect 29184 18964 29236 18970
rect 29184 18906 29236 18912
rect 29564 17746 29592 19314
rect 29840 18766 29868 24890
rect 30024 24750 30052 25774
rect 30012 24744 30064 24750
rect 30012 24686 30064 24692
rect 29920 23860 29972 23866
rect 29920 23802 29972 23808
rect 29932 23118 29960 23802
rect 29920 23112 29972 23118
rect 29920 23054 29972 23060
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 29932 18970 29960 19790
rect 29920 18964 29972 18970
rect 29920 18906 29972 18912
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29184 17740 29236 17746
rect 29184 17682 29236 17688
rect 29552 17740 29604 17746
rect 29552 17682 29604 17688
rect 29196 16998 29224 17682
rect 29460 17604 29512 17610
rect 29460 17546 29512 17552
rect 29472 17338 29500 17546
rect 29460 17332 29512 17338
rect 29460 17274 29512 17280
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 29196 16046 29224 16934
rect 29656 16794 29684 17138
rect 29644 16788 29696 16794
rect 29644 16730 29696 16736
rect 30116 16726 30144 34886
rect 30288 34196 30340 34202
rect 30288 34138 30340 34144
rect 30196 31340 30248 31346
rect 30196 31282 30248 31288
rect 30208 30682 30236 31282
rect 30300 30802 30328 34138
rect 30576 31278 30604 35430
rect 31208 31816 31260 31822
rect 31208 31758 31260 31764
rect 30564 31272 30616 31278
rect 30564 31214 30616 31220
rect 30288 30796 30340 30802
rect 30288 30738 30340 30744
rect 30380 30728 30432 30734
rect 30208 30676 30380 30682
rect 30208 30670 30432 30676
rect 30208 30654 30420 30670
rect 30208 29646 30236 30654
rect 30196 29640 30248 29646
rect 30196 29582 30248 29588
rect 30576 29170 30604 31214
rect 30748 31136 30800 31142
rect 30748 31078 30800 31084
rect 30760 30870 30788 31078
rect 30748 30864 30800 30870
rect 30748 30806 30800 30812
rect 31220 30598 31248 31758
rect 31208 30592 31260 30598
rect 31208 30534 31260 30540
rect 31220 30394 31248 30534
rect 31208 30388 31260 30394
rect 31208 30330 31260 30336
rect 31208 29640 31260 29646
rect 31208 29582 31260 29588
rect 31024 29504 31076 29510
rect 31024 29446 31076 29452
rect 31036 29238 31064 29446
rect 31024 29232 31076 29238
rect 31024 29174 31076 29180
rect 30564 29164 30616 29170
rect 30564 29106 30616 29112
rect 30472 29096 30524 29102
rect 30472 29038 30524 29044
rect 30196 26988 30248 26994
rect 30196 26930 30248 26936
rect 30208 22982 30236 26930
rect 30484 25498 30512 29038
rect 31220 28762 31248 29582
rect 31208 28756 31260 28762
rect 31208 28698 31260 28704
rect 30932 27532 30984 27538
rect 30932 27474 30984 27480
rect 30656 27328 30708 27334
rect 30656 27270 30708 27276
rect 30748 27328 30800 27334
rect 30748 27270 30800 27276
rect 30668 26450 30696 27270
rect 30760 27010 30788 27270
rect 30760 26994 30880 27010
rect 30760 26988 30892 26994
rect 30760 26982 30840 26988
rect 30840 26930 30892 26936
rect 30748 26920 30800 26926
rect 30748 26862 30800 26868
rect 30656 26444 30708 26450
rect 30656 26386 30708 26392
rect 30472 25492 30524 25498
rect 30472 25434 30524 25440
rect 30760 25294 30788 26862
rect 30852 26314 30880 26930
rect 30944 26926 30972 27474
rect 31116 27396 31168 27402
rect 31116 27338 31168 27344
rect 31128 27130 31156 27338
rect 31116 27124 31168 27130
rect 31116 27066 31168 27072
rect 30932 26920 30984 26926
rect 30932 26862 30984 26868
rect 30840 26308 30892 26314
rect 30840 26250 30892 26256
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30748 25288 30800 25294
rect 30748 25230 30800 25236
rect 30392 24614 30420 25230
rect 30760 24750 30788 25230
rect 30656 24744 30708 24750
rect 30656 24686 30708 24692
rect 30748 24744 30800 24750
rect 30748 24686 30800 24692
rect 30380 24608 30432 24614
rect 30380 24550 30432 24556
rect 30668 23118 30696 24686
rect 30656 23112 30708 23118
rect 30656 23054 30708 23060
rect 30196 22976 30248 22982
rect 30196 22918 30248 22924
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30656 22976 30708 22982
rect 30656 22918 30708 22924
rect 30208 17542 30236 22918
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30484 22030 30512 22714
rect 30576 22574 30604 22918
rect 30564 22568 30616 22574
rect 30564 22510 30616 22516
rect 30472 22024 30524 22030
rect 30472 21966 30524 21972
rect 30668 21962 30696 22918
rect 30760 22522 30788 24686
rect 30852 22964 30880 26250
rect 31128 25770 31156 27066
rect 31300 26988 31352 26994
rect 31300 26930 31352 26936
rect 31208 26444 31260 26450
rect 31208 26386 31260 26392
rect 31116 25764 31168 25770
rect 31116 25706 31168 25712
rect 31128 25362 31156 25706
rect 31220 25702 31248 26386
rect 31312 26314 31340 26930
rect 31300 26308 31352 26314
rect 31300 26250 31352 26256
rect 31312 25906 31340 26250
rect 31300 25900 31352 25906
rect 31300 25842 31352 25848
rect 31208 25696 31260 25702
rect 31208 25638 31260 25644
rect 31116 25356 31168 25362
rect 31116 25298 31168 25304
rect 30932 25152 30984 25158
rect 30932 25094 30984 25100
rect 30944 24818 30972 25094
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30932 22976 30984 22982
rect 30852 22936 30932 22964
rect 30932 22918 30984 22924
rect 30944 22778 30972 22918
rect 30932 22772 30984 22778
rect 30932 22714 30984 22720
rect 30840 22636 30892 22642
rect 30840 22578 30892 22584
rect 30852 22522 30880 22578
rect 30760 22494 30880 22522
rect 30932 22568 30984 22574
rect 30932 22510 30984 22516
rect 30760 22098 30788 22494
rect 30748 22092 30800 22098
rect 30748 22034 30800 22040
rect 30656 21956 30708 21962
rect 30656 21898 30708 21904
rect 30748 21956 30800 21962
rect 30748 21898 30800 21904
rect 30564 21888 30616 21894
rect 30564 21830 30616 21836
rect 30576 20942 30604 21830
rect 30564 20936 30616 20942
rect 30564 20878 30616 20884
rect 30380 20800 30432 20806
rect 30380 20742 30432 20748
rect 30392 19174 30420 20742
rect 30576 20534 30604 20878
rect 30668 20602 30696 21898
rect 30760 21010 30788 21898
rect 30840 21888 30892 21894
rect 30840 21830 30892 21836
rect 30852 21486 30880 21830
rect 30840 21480 30892 21486
rect 30840 21422 30892 21428
rect 30944 21010 30972 22510
rect 31220 22094 31248 25638
rect 31312 24750 31340 25842
rect 31392 25220 31444 25226
rect 31392 25162 31444 25168
rect 31404 24750 31432 25162
rect 31300 24744 31352 24750
rect 31300 24686 31352 24692
rect 31392 24744 31444 24750
rect 31392 24686 31444 24692
rect 31312 22794 31340 24686
rect 31404 22982 31432 24686
rect 31392 22976 31444 22982
rect 31392 22918 31444 22924
rect 31312 22766 31432 22794
rect 31404 22234 31432 22766
rect 31392 22228 31444 22234
rect 31392 22170 31444 22176
rect 31220 22066 31340 22094
rect 31024 21344 31076 21350
rect 31024 21286 31076 21292
rect 31036 21078 31064 21286
rect 31208 21140 31260 21146
rect 31208 21082 31260 21088
rect 31024 21072 31076 21078
rect 31024 21014 31076 21020
rect 30748 21004 30800 21010
rect 30748 20946 30800 20952
rect 30932 21004 30984 21010
rect 30932 20946 30984 20952
rect 30656 20596 30708 20602
rect 30656 20538 30708 20544
rect 30564 20528 30616 20534
rect 30564 20470 30616 20476
rect 30472 20460 30524 20466
rect 30472 20402 30524 20408
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 30392 18834 30420 19110
rect 30484 18970 30512 20402
rect 30760 20398 30788 20946
rect 30838 20632 30894 20641
rect 30838 20567 30894 20576
rect 30748 20392 30800 20398
rect 30748 20334 30800 20340
rect 30656 20256 30708 20262
rect 30656 20198 30708 20204
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30380 18828 30432 18834
rect 30380 18770 30432 18776
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 30392 18170 30420 18226
rect 30564 18216 30616 18222
rect 30392 18142 30512 18170
rect 30564 18158 30616 18164
rect 30484 17882 30512 18142
rect 30472 17876 30524 17882
rect 30472 17818 30524 17824
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30288 17060 30340 17066
rect 30288 17002 30340 17008
rect 30104 16720 30156 16726
rect 30104 16662 30156 16668
rect 29552 16584 29604 16590
rect 30116 16538 30144 16662
rect 30300 16658 30328 17002
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 29552 16526 29604 16532
rect 29184 16040 29236 16046
rect 29184 15982 29236 15988
rect 29564 15706 29592 16526
rect 30024 16510 30144 16538
rect 30196 16516 30248 16522
rect 29736 16108 29788 16114
rect 29736 16050 29788 16056
rect 29748 15706 29776 16050
rect 29552 15700 29604 15706
rect 29552 15642 29604 15648
rect 29736 15700 29788 15706
rect 29736 15642 29788 15648
rect 29368 14408 29420 14414
rect 29368 14350 29420 14356
rect 29276 14272 29328 14278
rect 29276 14214 29328 14220
rect 29288 13938 29316 14214
rect 29380 14074 29408 14350
rect 30024 14278 30052 16510
rect 30196 16458 30248 16464
rect 30104 16448 30156 16454
rect 30104 16390 30156 16396
rect 30116 16250 30144 16390
rect 30104 16244 30156 16250
rect 30104 16186 30156 16192
rect 30116 15502 30144 16186
rect 30208 15570 30236 16458
rect 30576 16454 30604 18158
rect 30668 17678 30696 20198
rect 30852 19990 30880 20567
rect 30944 20466 30972 20946
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 30840 19984 30892 19990
rect 30840 19926 30892 19932
rect 30932 19916 30984 19922
rect 30932 19858 30984 19864
rect 30840 19168 30892 19174
rect 30840 19110 30892 19116
rect 30852 18766 30880 19110
rect 30840 18760 30892 18766
rect 30840 18702 30892 18708
rect 30944 18222 30972 19858
rect 31036 18630 31064 21014
rect 31220 20942 31248 21082
rect 31208 20936 31260 20942
rect 31208 20878 31260 20884
rect 31312 20806 31340 22066
rect 31404 21350 31432 22170
rect 31392 21344 31444 21350
rect 31392 21286 31444 21292
rect 31300 20800 31352 20806
rect 31300 20742 31352 20748
rect 31208 18692 31260 18698
rect 31208 18634 31260 18640
rect 31024 18624 31076 18630
rect 31024 18566 31076 18572
rect 31220 18426 31248 18634
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31312 18358 31340 20742
rect 31300 18352 31352 18358
rect 31300 18294 31352 18300
rect 31392 18284 31444 18290
rect 31392 18226 31444 18232
rect 30932 18216 30984 18222
rect 30932 18158 30984 18164
rect 30656 17672 30708 17678
rect 30656 17614 30708 17620
rect 30564 16448 30616 16454
rect 30564 16390 30616 16396
rect 30196 15564 30248 15570
rect 30196 15506 30248 15512
rect 30104 15496 30156 15502
rect 30104 15438 30156 15444
rect 30208 14550 30236 15506
rect 30748 15020 30800 15026
rect 30748 14962 30800 14968
rect 30288 14884 30340 14890
rect 30288 14826 30340 14832
rect 30196 14544 30248 14550
rect 30196 14486 30248 14492
rect 30012 14272 30064 14278
rect 30012 14214 30064 14220
rect 30208 14074 30236 14486
rect 30300 14482 30328 14826
rect 30760 14550 30788 14962
rect 30748 14544 30800 14550
rect 30748 14486 30800 14492
rect 30288 14476 30340 14482
rect 30288 14418 30340 14424
rect 29368 14068 29420 14074
rect 29368 14010 29420 14016
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29092 13456 29144 13462
rect 29092 13398 29144 13404
rect 29104 13326 29132 13398
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 29092 13320 29144 13326
rect 29092 13262 29144 13268
rect 29012 13190 29040 13262
rect 29000 13184 29052 13190
rect 29000 13126 29052 13132
rect 29288 12986 29316 13874
rect 30300 13870 30328 14418
rect 30748 13932 30800 13938
rect 30748 13874 30800 13880
rect 30288 13864 30340 13870
rect 30288 13806 30340 13812
rect 29920 13796 29972 13802
rect 29920 13738 29972 13744
rect 29276 12980 29328 12986
rect 29276 12922 29328 12928
rect 29644 12980 29696 12986
rect 29644 12922 29696 12928
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 29196 12442 29224 12786
rect 29184 12436 29236 12442
rect 29184 12378 29236 12384
rect 29276 12436 29328 12442
rect 29656 12434 29684 12922
rect 29932 12442 29960 13738
rect 30656 13728 30708 13734
rect 30656 13670 30708 13676
rect 30104 13184 30156 13190
rect 30104 13126 30156 13132
rect 29276 12378 29328 12384
rect 29564 12406 29684 12434
rect 29920 12436 29972 12442
rect 29288 12306 29316 12378
rect 29564 12306 29592 12406
rect 29920 12378 29972 12384
rect 30012 12436 30064 12442
rect 30012 12378 30064 12384
rect 30024 12322 30052 12378
rect 29276 12300 29328 12306
rect 29276 12242 29328 12248
rect 29552 12300 29604 12306
rect 29552 12242 29604 12248
rect 29932 12294 30052 12322
rect 30116 12306 30144 13126
rect 30668 12374 30696 13670
rect 30760 13530 30788 13874
rect 30748 13524 30800 13530
rect 30748 13466 30800 13472
rect 30656 12368 30708 12374
rect 30656 12310 30708 12316
rect 30104 12300 30156 12306
rect 29288 11354 29316 12242
rect 29276 11348 29328 11354
rect 29276 11290 29328 11296
rect 28722 11248 28778 11257
rect 28722 11183 28778 11192
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 28172 11144 28224 11150
rect 28172 11086 28224 11092
rect 28724 11144 28776 11150
rect 28724 11086 28776 11092
rect 27896 10804 27948 10810
rect 27896 10746 27948 10752
rect 27712 10600 27764 10606
rect 27712 10542 27764 10548
rect 27620 10532 27672 10538
rect 27620 10474 27672 10480
rect 27160 10464 27212 10470
rect 27160 10406 27212 10412
rect 27172 10062 27200 10406
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 27252 10056 27304 10062
rect 27252 9998 27304 10004
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 26436 9178 26464 9318
rect 26424 9172 26476 9178
rect 26424 9114 26476 9120
rect 26792 9036 26844 9042
rect 26792 8978 26844 8984
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 26804 8634 26832 8978
rect 26792 8628 26844 8634
rect 26792 8570 26844 8576
rect 26516 8492 26568 8498
rect 26516 8434 26568 8440
rect 26332 8288 26384 8294
rect 26332 8230 26384 8236
rect 26344 8090 26372 8230
rect 26528 8090 26556 8434
rect 26332 8084 26384 8090
rect 26332 8026 26384 8032
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 26608 7948 26660 7954
rect 26608 7890 26660 7896
rect 25044 7880 25096 7886
rect 24964 7840 25044 7868
rect 24964 7342 24992 7840
rect 25044 7822 25096 7828
rect 25964 7812 26016 7818
rect 25964 7754 26016 7760
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 25976 7206 26004 7754
rect 26620 7342 26648 7890
rect 26804 7886 26832 8570
rect 27264 8294 27292 9998
rect 27344 9104 27396 9110
rect 27344 9046 27396 9052
rect 27356 8498 27384 9046
rect 27632 8566 27660 10474
rect 27724 10266 27752 10542
rect 27804 10464 27856 10470
rect 27804 10406 27856 10412
rect 27712 10260 27764 10266
rect 27712 10202 27764 10208
rect 27724 9450 27752 10202
rect 27712 9444 27764 9450
rect 27712 9386 27764 9392
rect 27816 8974 27844 10406
rect 27908 8974 27936 10746
rect 28000 10606 28028 11086
rect 28184 10674 28212 11086
rect 28540 11008 28592 11014
rect 28540 10950 28592 10956
rect 28632 11008 28684 11014
rect 28632 10950 28684 10956
rect 28172 10668 28224 10674
rect 28172 10610 28224 10616
rect 28552 10606 28580 10950
rect 28644 10674 28672 10950
rect 28632 10668 28684 10674
rect 28632 10610 28684 10616
rect 27988 10600 28040 10606
rect 27988 10542 28040 10548
rect 28540 10600 28592 10606
rect 28540 10542 28592 10548
rect 27804 8968 27856 8974
rect 27804 8910 27856 8916
rect 27896 8968 27948 8974
rect 27896 8910 27948 8916
rect 27908 8838 27936 8910
rect 27896 8832 27948 8838
rect 27896 8774 27948 8780
rect 27620 8560 27672 8566
rect 27620 8502 27672 8508
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27436 8356 27488 8362
rect 27436 8298 27488 8304
rect 27252 8288 27304 8294
rect 27252 8230 27304 8236
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 26608 7336 26660 7342
rect 26608 7278 26660 7284
rect 25964 7200 26016 7206
rect 25964 7142 26016 7148
rect 25976 6934 26004 7142
rect 25964 6928 26016 6934
rect 25964 6870 26016 6876
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 25688 6316 25740 6322
rect 25688 6258 25740 6264
rect 24860 6180 24912 6186
rect 24860 6122 24912 6128
rect 24872 5710 24900 6122
rect 25056 5846 25084 6258
rect 25044 5840 25096 5846
rect 25044 5782 25096 5788
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24872 5234 24900 5646
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 25056 4826 25084 5782
rect 25700 5098 25728 6258
rect 25872 6112 25924 6118
rect 25872 6054 25924 6060
rect 25884 5846 25912 6054
rect 25872 5840 25924 5846
rect 25872 5782 25924 5788
rect 25884 5710 25912 5782
rect 26620 5778 26648 7278
rect 26700 7268 26752 7274
rect 26700 7210 26752 7216
rect 26712 6730 26740 7210
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26712 6186 26740 6666
rect 26700 6180 26752 6186
rect 26700 6122 26752 6128
rect 26608 5772 26660 5778
rect 26608 5714 26660 5720
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 25964 5704 26016 5710
rect 25964 5646 26016 5652
rect 25976 5370 26004 5646
rect 26712 5642 26740 6122
rect 27252 5704 27304 5710
rect 27252 5646 27304 5652
rect 26700 5636 26752 5642
rect 26700 5578 26752 5584
rect 25964 5364 26016 5370
rect 25964 5306 26016 5312
rect 27264 5302 27292 5646
rect 27448 5642 27476 8298
rect 27540 7886 27568 8366
rect 27632 7954 27660 8502
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27724 8022 27752 8434
rect 27712 8016 27764 8022
rect 27712 7958 27764 7964
rect 27908 7954 27936 8774
rect 27620 7948 27672 7954
rect 27620 7890 27672 7896
rect 27896 7948 27948 7954
rect 27896 7890 27948 7896
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27540 7546 27568 7822
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27540 5778 27568 6258
rect 27620 6112 27672 6118
rect 27620 6054 27672 6060
rect 27712 6112 27764 6118
rect 27712 6054 27764 6060
rect 27528 5772 27580 5778
rect 27528 5714 27580 5720
rect 27436 5636 27488 5642
rect 27436 5578 27488 5584
rect 27448 5370 27476 5578
rect 27436 5364 27488 5370
rect 27436 5306 27488 5312
rect 27252 5296 27304 5302
rect 27252 5238 27304 5244
rect 25688 5092 25740 5098
rect 25688 5034 25740 5040
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 25700 4758 25728 5034
rect 26240 5024 26292 5030
rect 26240 4966 26292 4972
rect 25688 4752 25740 4758
rect 25688 4694 25740 4700
rect 25700 4622 25728 4694
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25688 4616 25740 4622
rect 25688 4558 25740 4564
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 25056 4146 25084 4422
rect 25240 4146 25268 4558
rect 25700 4146 25728 4558
rect 26252 4146 26280 4966
rect 26700 4684 26752 4690
rect 26700 4626 26752 4632
rect 26516 4480 26568 4486
rect 26516 4422 26568 4428
rect 26528 4146 26556 4422
rect 26712 4146 26740 4626
rect 27264 4622 27292 5238
rect 27252 4616 27304 4622
rect 27252 4558 27304 4564
rect 27448 4554 27476 5306
rect 27632 4826 27660 6054
rect 27724 5710 27752 6054
rect 27712 5704 27764 5710
rect 27712 5646 27764 5652
rect 27804 5568 27856 5574
rect 27804 5510 27856 5516
rect 27816 5234 27844 5510
rect 27804 5228 27856 5234
rect 27804 5170 27856 5176
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 27816 4690 27844 5170
rect 27804 4684 27856 4690
rect 27804 4626 27856 4632
rect 27436 4548 27488 4554
rect 27436 4490 27488 4496
rect 27896 4548 27948 4554
rect 27896 4490 27948 4496
rect 27908 4214 27936 4490
rect 27896 4208 27948 4214
rect 27896 4150 27948 4156
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 25228 4140 25280 4146
rect 25228 4082 25280 4088
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26700 4140 26752 4146
rect 26700 4082 26752 4088
rect 24492 3732 24544 3738
rect 24492 3674 24544 3680
rect 25056 3194 25084 4082
rect 26148 3936 26200 3942
rect 26148 3878 26200 3884
rect 26160 3602 26188 3878
rect 26252 3602 26280 4082
rect 26608 4072 26660 4078
rect 26608 4014 26660 4020
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 26240 3596 26292 3602
rect 26240 3538 26292 3544
rect 26620 3534 26648 4014
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26608 3528 26660 3534
rect 26608 3470 26660 3476
rect 25136 3392 25188 3398
rect 25136 3334 25188 3340
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 23952 2961 23980 2994
rect 25148 2990 25176 3334
rect 25700 3194 25728 3470
rect 25688 3188 25740 3194
rect 25688 3130 25740 3136
rect 24308 2984 24360 2990
rect 23938 2952 23994 2961
rect 24308 2926 24360 2932
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 23938 2887 23994 2896
rect 24320 2854 24348 2926
rect 25320 2916 25372 2922
rect 25320 2858 25372 2864
rect 24308 2848 24360 2854
rect 24308 2790 24360 2796
rect 24320 2514 24348 2790
rect 24308 2508 24360 2514
rect 24308 2450 24360 2456
rect 25332 2446 25360 2858
rect 25976 2650 26004 3470
rect 26528 3380 26556 3470
rect 26712 3380 26740 4082
rect 28000 4010 28028 10542
rect 28552 10062 28580 10542
rect 28644 10266 28672 10610
rect 28736 10282 28764 11086
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 28816 10804 28868 10810
rect 28816 10746 28868 10752
rect 28828 10674 28856 10746
rect 29012 10742 29040 10950
rect 29000 10736 29052 10742
rect 29000 10678 29052 10684
rect 29368 10736 29420 10742
rect 29368 10678 29420 10684
rect 28816 10668 28868 10674
rect 28816 10610 28868 10616
rect 28828 10470 28856 10610
rect 28908 10532 28960 10538
rect 28908 10474 28960 10480
rect 28816 10464 28868 10470
rect 28816 10406 28868 10412
rect 28736 10266 28856 10282
rect 28632 10260 28684 10266
rect 28736 10260 28868 10266
rect 28736 10254 28816 10260
rect 28632 10202 28684 10208
rect 28816 10202 28868 10208
rect 28920 10130 28948 10474
rect 29092 10464 29144 10470
rect 29092 10406 29144 10412
rect 29104 10130 29132 10406
rect 29380 10198 29408 10678
rect 29368 10192 29420 10198
rect 29368 10134 29420 10140
rect 28908 10124 28960 10130
rect 28908 10066 28960 10072
rect 29092 10124 29144 10130
rect 29092 10066 29144 10072
rect 28540 10056 28592 10062
rect 28540 9998 28592 10004
rect 29276 9512 29328 9518
rect 29276 9454 29328 9460
rect 28908 9444 28960 9450
rect 28908 9386 28960 9392
rect 28264 8900 28316 8906
rect 28264 8842 28316 8848
rect 28172 7744 28224 7750
rect 28276 7732 28304 8842
rect 28448 8628 28500 8634
rect 28448 8570 28500 8576
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28368 8090 28396 8434
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 28460 7750 28488 8570
rect 28224 7704 28304 7732
rect 28448 7744 28500 7750
rect 28172 7686 28224 7692
rect 28448 7686 28500 7692
rect 28184 6458 28212 7686
rect 28172 6452 28224 6458
rect 28172 6394 28224 6400
rect 28460 6322 28488 7686
rect 28920 6798 28948 9386
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 29196 8566 29224 8774
rect 29184 8560 29236 8566
rect 29184 8502 29236 8508
rect 29184 8288 29236 8294
rect 29288 8276 29316 9454
rect 29236 8248 29316 8276
rect 29368 8288 29420 8294
rect 29184 8230 29236 8236
rect 29368 8230 29420 8236
rect 29196 7818 29224 8230
rect 29184 7812 29236 7818
rect 29184 7754 29236 7760
rect 29092 7744 29144 7750
rect 29092 7686 29144 7692
rect 29104 7410 29132 7686
rect 29092 7404 29144 7410
rect 29092 7346 29144 7352
rect 29104 6798 29132 7346
rect 29380 6934 29408 8230
rect 29460 7200 29512 7206
rect 29460 7142 29512 7148
rect 29368 6928 29420 6934
rect 29368 6870 29420 6876
rect 28908 6792 28960 6798
rect 28908 6734 28960 6740
rect 29092 6792 29144 6798
rect 29092 6734 29144 6740
rect 28920 6322 28948 6734
rect 29000 6656 29052 6662
rect 29000 6598 29052 6604
rect 28448 6316 28500 6322
rect 28448 6258 28500 6264
rect 28908 6316 28960 6322
rect 28908 6258 28960 6264
rect 28540 5704 28592 5710
rect 28540 5646 28592 5652
rect 28264 4752 28316 4758
rect 28264 4694 28316 4700
rect 28276 4622 28304 4694
rect 28356 4684 28408 4690
rect 28356 4626 28408 4632
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28264 4616 28316 4622
rect 28264 4558 28316 4564
rect 28184 4468 28212 4558
rect 28368 4468 28396 4626
rect 28448 4616 28500 4622
rect 28448 4558 28500 4564
rect 28184 4440 28396 4468
rect 28460 4214 28488 4558
rect 28448 4208 28500 4214
rect 28448 4150 28500 4156
rect 27988 4004 28040 4010
rect 27988 3946 28040 3952
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 27068 3528 27120 3534
rect 27068 3470 27120 3476
rect 26528 3352 26740 3380
rect 27080 3194 27108 3470
rect 27540 3194 27568 3538
rect 26148 3188 26200 3194
rect 26148 3130 26200 3136
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 26056 3052 26108 3058
rect 26056 2994 26108 3000
rect 25964 2644 26016 2650
rect 25964 2586 26016 2592
rect 26068 2530 26096 2994
rect 25976 2514 26096 2530
rect 26160 2514 26188 3130
rect 28552 3058 28580 5646
rect 29012 4554 29040 6598
rect 29104 6390 29132 6734
rect 29380 6662 29408 6870
rect 29368 6656 29420 6662
rect 29368 6598 29420 6604
rect 29092 6384 29144 6390
rect 29092 6326 29144 6332
rect 29472 6322 29500 7142
rect 29460 6316 29512 6322
rect 29460 6258 29512 6264
rect 29460 5704 29512 5710
rect 29458 5672 29460 5681
rect 29512 5672 29514 5681
rect 29458 5607 29514 5616
rect 29564 5522 29592 12242
rect 29644 12232 29696 12238
rect 29644 12174 29696 12180
rect 29656 10674 29684 12174
rect 29932 12102 29960 12294
rect 30104 12242 30156 12248
rect 29920 12096 29972 12102
rect 29920 12038 29972 12044
rect 30288 12096 30340 12102
rect 30288 12038 30340 12044
rect 29932 11558 29960 12038
rect 30300 11762 30328 12038
rect 30668 11762 30696 12310
rect 30944 12306 30972 18158
rect 31404 18154 31432 18226
rect 31392 18148 31444 18154
rect 31392 18090 31444 18096
rect 31496 17218 31524 37130
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 32772 36236 32824 36242
rect 32772 36178 32824 36184
rect 31852 32020 31904 32026
rect 31852 31962 31904 31968
rect 31760 31136 31812 31142
rect 31760 31078 31812 31084
rect 31772 30734 31800 31078
rect 31760 30728 31812 30734
rect 31760 30670 31812 30676
rect 31864 27606 31892 31962
rect 31944 31952 31996 31958
rect 31944 31894 31996 31900
rect 31956 31346 31984 31894
rect 32588 31884 32640 31890
rect 32588 31826 32640 31832
rect 31944 31340 31996 31346
rect 31944 31282 31996 31288
rect 32404 30660 32456 30666
rect 32404 30602 32456 30608
rect 31944 28960 31996 28966
rect 31944 28902 31996 28908
rect 31956 28558 31984 28902
rect 32036 28620 32088 28626
rect 32036 28562 32088 28568
rect 31944 28552 31996 28558
rect 31944 28494 31996 28500
rect 31852 27600 31904 27606
rect 31852 27542 31904 27548
rect 31576 27328 31628 27334
rect 31628 27276 31708 27282
rect 31576 27270 31708 27276
rect 31588 27254 31708 27270
rect 31680 26994 31708 27254
rect 31668 26988 31720 26994
rect 31668 26930 31720 26936
rect 31680 26450 31708 26930
rect 31852 26920 31904 26926
rect 31852 26862 31904 26868
rect 31668 26444 31720 26450
rect 31668 26386 31720 26392
rect 31864 26382 31892 26862
rect 31944 26512 31996 26518
rect 31944 26454 31996 26460
rect 31576 26376 31628 26382
rect 31576 26318 31628 26324
rect 31852 26376 31904 26382
rect 31852 26318 31904 26324
rect 31588 25158 31616 26318
rect 31956 26234 31984 26454
rect 31772 26206 31984 26234
rect 31576 25152 31628 25158
rect 31576 25094 31628 25100
rect 31588 24954 31616 25094
rect 31576 24948 31628 24954
rect 31576 24890 31628 24896
rect 31772 23338 31800 26206
rect 32048 25158 32076 28562
rect 32416 26586 32444 30602
rect 32600 27062 32628 31826
rect 32588 27056 32640 27062
rect 32588 26998 32640 27004
rect 32404 26580 32456 26586
rect 32404 26522 32456 26528
rect 32404 25832 32456 25838
rect 32324 25780 32404 25786
rect 32324 25774 32456 25780
rect 32324 25758 32444 25774
rect 32324 25498 32352 25758
rect 32312 25492 32364 25498
rect 32312 25434 32364 25440
rect 32036 25152 32088 25158
rect 32036 25094 32088 25100
rect 32036 24948 32088 24954
rect 32036 24890 32088 24896
rect 31680 23310 31800 23338
rect 31680 23254 31708 23310
rect 31668 23248 31720 23254
rect 31668 23190 31720 23196
rect 31668 22432 31720 22438
rect 31668 22374 31720 22380
rect 31680 21146 31708 22374
rect 31668 21140 31720 21146
rect 31668 21082 31720 21088
rect 31772 21078 31800 23310
rect 31852 23044 31904 23050
rect 31852 22986 31904 22992
rect 31864 22506 31892 22986
rect 31852 22500 31904 22506
rect 31852 22442 31904 22448
rect 32048 21146 32076 24890
rect 32220 24812 32272 24818
rect 32220 24754 32272 24760
rect 32232 24342 32260 24754
rect 32220 24336 32272 24342
rect 32220 24278 32272 24284
rect 32128 24200 32180 24206
rect 32128 24142 32180 24148
rect 32140 21894 32168 24142
rect 32220 22976 32272 22982
rect 32220 22918 32272 22924
rect 32232 22642 32260 22918
rect 32324 22778 32352 25434
rect 32404 25424 32456 25430
rect 32404 25366 32456 25372
rect 32416 23186 32444 25366
rect 32784 25362 32812 36178
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 36188 35834 36216 37198
rect 37384 37194 37412 39280
rect 37372 37188 37424 37194
rect 37372 37130 37424 37136
rect 36360 37120 36412 37126
rect 36360 37062 36412 37068
rect 36372 36825 36400 37062
rect 36358 36816 36414 36825
rect 36358 36751 36414 36760
rect 36176 35828 36228 35834
rect 36176 35770 36228 35776
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 35992 33516 36044 33522
rect 35992 33458 36044 33464
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35440 27464 35492 27470
rect 35440 27406 35492 27412
rect 33324 27396 33376 27402
rect 33324 27338 33376 27344
rect 33336 26994 33364 27338
rect 33324 26988 33376 26994
rect 33324 26930 33376 26936
rect 32864 26920 32916 26926
rect 32864 26862 32916 26868
rect 32876 26518 32904 26862
rect 32864 26512 32916 26518
rect 32864 26454 32916 26460
rect 32876 26382 32904 26454
rect 33336 26450 33364 26930
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 33324 26444 33376 26450
rect 33324 26386 33376 26392
rect 32864 26376 32916 26382
rect 32864 26318 32916 26324
rect 33336 26042 33364 26386
rect 33324 26036 33376 26042
rect 33324 25978 33376 25984
rect 33140 25900 33192 25906
rect 33140 25842 33192 25848
rect 32956 25832 33008 25838
rect 32956 25774 33008 25780
rect 32968 25362 32996 25774
rect 32772 25356 32824 25362
rect 32772 25298 32824 25304
rect 32956 25356 33008 25362
rect 32956 25298 33008 25304
rect 33048 25288 33100 25294
rect 33048 25230 33100 25236
rect 33060 24886 33088 25230
rect 33152 25226 33180 25842
rect 33876 25764 33928 25770
rect 33876 25706 33928 25712
rect 33888 25294 33916 25706
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 33876 25288 33928 25294
rect 33876 25230 33928 25236
rect 33140 25220 33192 25226
rect 33140 25162 33192 25168
rect 33048 24880 33100 24886
rect 33048 24822 33100 24828
rect 32588 24812 32640 24818
rect 32588 24754 32640 24760
rect 32600 24410 32628 24754
rect 32588 24404 32640 24410
rect 32588 24346 32640 24352
rect 33060 23798 33088 24822
rect 33048 23792 33100 23798
rect 33048 23734 33100 23740
rect 32864 23248 32916 23254
rect 32864 23190 32916 23196
rect 32404 23180 32456 23186
rect 32404 23122 32456 23128
rect 32416 22778 32444 23122
rect 32312 22772 32364 22778
rect 32312 22714 32364 22720
rect 32404 22772 32456 22778
rect 32404 22714 32456 22720
rect 32220 22636 32272 22642
rect 32220 22578 32272 22584
rect 32312 22636 32364 22642
rect 32312 22578 32364 22584
rect 32128 21888 32180 21894
rect 32128 21830 32180 21836
rect 32036 21140 32088 21146
rect 32036 21082 32088 21088
rect 31760 21072 31812 21078
rect 31760 21014 31812 21020
rect 32048 20874 32076 21082
rect 32128 20936 32180 20942
rect 32232 20924 32260 22578
rect 32324 22234 32352 22578
rect 32312 22228 32364 22234
rect 32312 22170 32364 22176
rect 32416 22030 32444 22714
rect 32876 22642 32904 23190
rect 32496 22636 32548 22642
rect 32496 22578 32548 22584
rect 32864 22636 32916 22642
rect 32864 22578 32916 22584
rect 32508 22506 32536 22578
rect 33152 22574 33180 25162
rect 33888 24954 33916 25230
rect 33876 24948 33928 24954
rect 33876 24890 33928 24896
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 33232 23860 33284 23866
rect 33232 23802 33284 23808
rect 33244 23118 33272 23802
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 33232 23112 33284 23118
rect 33232 23054 33284 23060
rect 33244 22794 33272 23054
rect 33784 23044 33836 23050
rect 33784 22986 33836 22992
rect 33244 22766 33364 22794
rect 33796 22778 33824 22986
rect 33232 22636 33284 22642
rect 33232 22578 33284 22584
rect 33140 22568 33192 22574
rect 33140 22510 33192 22516
rect 32496 22500 32548 22506
rect 32496 22442 32548 22448
rect 32680 22160 32732 22166
rect 32680 22102 32732 22108
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 32588 21888 32640 21894
rect 32588 21830 32640 21836
rect 32180 20896 32260 20924
rect 32128 20878 32180 20884
rect 32036 20868 32088 20874
rect 32036 20810 32088 20816
rect 31944 20800 31996 20806
rect 31944 20742 31996 20748
rect 31668 20460 31720 20466
rect 31668 20402 31720 20408
rect 31852 20460 31904 20466
rect 31852 20402 31904 20408
rect 31680 19922 31708 20402
rect 31864 20262 31892 20402
rect 31852 20256 31904 20262
rect 31852 20198 31904 20204
rect 31668 19916 31720 19922
rect 31668 19858 31720 19864
rect 31576 18760 31628 18766
rect 31576 18702 31628 18708
rect 31312 17190 31524 17218
rect 31116 16652 31168 16658
rect 31116 16594 31168 16600
rect 31128 15910 31156 16594
rect 31116 15904 31168 15910
rect 31116 15846 31168 15852
rect 31208 14272 31260 14278
rect 31128 14232 31208 14260
rect 31128 13190 31156 14232
rect 31208 14214 31260 14220
rect 31116 13184 31168 13190
rect 31116 13126 31168 13132
rect 30932 12300 30984 12306
rect 30932 12242 30984 12248
rect 31128 12238 31156 13126
rect 31312 12322 31340 17190
rect 31588 16658 31616 18702
rect 31956 16794 31984 20742
rect 32048 20466 32076 20810
rect 32140 20602 32168 20878
rect 32128 20596 32180 20602
rect 32128 20538 32180 20544
rect 32036 20460 32088 20466
rect 32036 20402 32088 20408
rect 32140 20330 32168 20538
rect 32128 20324 32180 20330
rect 32128 20266 32180 20272
rect 32404 19304 32456 19310
rect 32404 19246 32456 19252
rect 32416 18834 32444 19246
rect 32404 18828 32456 18834
rect 32404 18770 32456 18776
rect 32220 18692 32272 18698
rect 32220 18634 32272 18640
rect 32232 18426 32260 18634
rect 32416 18426 32444 18770
rect 32220 18420 32272 18426
rect 32220 18362 32272 18368
rect 32404 18420 32456 18426
rect 32404 18362 32456 18368
rect 32404 18284 32456 18290
rect 32404 18226 32456 18232
rect 32416 17338 32444 18226
rect 32404 17332 32456 17338
rect 32404 17274 32456 17280
rect 32496 17196 32548 17202
rect 32496 17138 32548 17144
rect 32508 16794 32536 17138
rect 31944 16788 31996 16794
rect 31944 16730 31996 16736
rect 32496 16788 32548 16794
rect 32496 16730 32548 16736
rect 31576 16652 31628 16658
rect 31576 16594 31628 16600
rect 31852 16516 31904 16522
rect 31852 16458 31904 16464
rect 31864 16250 31892 16458
rect 32508 16250 32536 16730
rect 32600 16250 32628 21830
rect 32692 19922 32720 22102
rect 33152 22030 33180 22510
rect 33140 22024 33192 22030
rect 33140 21966 33192 21972
rect 33244 21894 33272 22578
rect 33232 21888 33284 21894
rect 33232 21830 33284 21836
rect 33336 21706 33364 22766
rect 33784 22772 33836 22778
rect 33784 22714 33836 22720
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 33416 21888 33468 21894
rect 33416 21830 33468 21836
rect 33152 21678 33364 21706
rect 33048 21072 33100 21078
rect 33048 21014 33100 21020
rect 32680 19916 32732 19922
rect 32680 19858 32732 19864
rect 33060 19854 33088 21014
rect 33152 21010 33180 21678
rect 33324 21548 33376 21554
rect 33324 21490 33376 21496
rect 33232 21344 33284 21350
rect 33232 21286 33284 21292
rect 33140 21004 33192 21010
rect 33140 20946 33192 20952
rect 33152 20466 33180 20946
rect 33244 20942 33272 21286
rect 33232 20936 33284 20942
rect 33232 20878 33284 20884
rect 33140 20460 33192 20466
rect 33140 20402 33192 20408
rect 33336 20058 33364 21490
rect 33324 20052 33376 20058
rect 33324 19994 33376 20000
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 33140 19712 33192 19718
rect 33140 19654 33192 19660
rect 32680 17128 32732 17134
rect 32680 17070 32732 17076
rect 31852 16244 31904 16250
rect 31852 16186 31904 16192
rect 32496 16244 32548 16250
rect 32496 16186 32548 16192
rect 32588 16244 32640 16250
rect 32588 16186 32640 16192
rect 32692 16130 32720 17070
rect 32600 16102 32720 16130
rect 32600 16046 32628 16102
rect 32588 16040 32640 16046
rect 32588 15982 32640 15988
rect 32680 16040 32732 16046
rect 32680 15982 32732 15988
rect 31852 14816 31904 14822
rect 31852 14758 31904 14764
rect 31864 14414 31892 14758
rect 31852 14408 31904 14414
rect 31852 14350 31904 14356
rect 32600 14278 32628 15982
rect 32692 15570 32720 15982
rect 32680 15564 32732 15570
rect 32680 15506 32732 15512
rect 32864 14476 32916 14482
rect 32864 14418 32916 14424
rect 32876 14346 32904 14418
rect 32864 14340 32916 14346
rect 32864 14282 32916 14288
rect 32588 14272 32640 14278
rect 32588 14214 32640 14220
rect 31944 13932 31996 13938
rect 31944 13874 31996 13880
rect 31956 13258 31984 13874
rect 32036 13388 32088 13394
rect 32036 13330 32088 13336
rect 31944 13252 31996 13258
rect 31944 13194 31996 13200
rect 32048 12442 32076 13330
rect 32876 13326 32904 14282
rect 33152 14074 33180 19654
rect 33324 18284 33376 18290
rect 33324 18226 33376 18232
rect 33336 17882 33364 18226
rect 33324 17876 33376 17882
rect 33324 17818 33376 17824
rect 33428 15638 33456 21830
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 20256 34848 20262
rect 34796 20198 34848 20204
rect 34704 19780 34756 19786
rect 34704 19722 34756 19728
rect 34612 19712 34664 19718
rect 34612 19654 34664 19660
rect 34624 19446 34652 19654
rect 34612 19440 34664 19446
rect 34612 19382 34664 19388
rect 34152 19372 34204 19378
rect 34152 19314 34204 19320
rect 34164 18834 34192 19314
rect 34152 18828 34204 18834
rect 34152 18770 34204 18776
rect 33600 17672 33652 17678
rect 33600 17614 33652 17620
rect 33612 17338 33640 17614
rect 33600 17332 33652 17338
rect 33600 17274 33652 17280
rect 34060 17128 34112 17134
rect 34060 17070 34112 17076
rect 33784 16584 33836 16590
rect 33784 16526 33836 16532
rect 33796 16250 33824 16526
rect 33784 16244 33836 16250
rect 33784 16186 33836 16192
rect 34072 16182 34100 17070
rect 34164 16794 34192 18770
rect 34624 18766 34652 19382
rect 34612 18760 34664 18766
rect 34612 18702 34664 18708
rect 34520 18216 34572 18222
rect 34520 18158 34572 18164
rect 34428 17196 34480 17202
rect 34428 17138 34480 17144
rect 34336 17128 34388 17134
rect 34336 17070 34388 17076
rect 34152 16788 34204 16794
rect 34152 16730 34204 16736
rect 33508 16176 33560 16182
rect 33508 16118 33560 16124
rect 34060 16176 34112 16182
rect 34060 16118 34112 16124
rect 33416 15632 33468 15638
rect 33416 15574 33468 15580
rect 33416 14952 33468 14958
rect 33416 14894 33468 14900
rect 33232 14816 33284 14822
rect 33232 14758 33284 14764
rect 33324 14816 33376 14822
rect 33324 14758 33376 14764
rect 33244 14414 33272 14758
rect 33336 14482 33364 14758
rect 33324 14476 33376 14482
rect 33324 14418 33376 14424
rect 33232 14408 33284 14414
rect 33232 14350 33284 14356
rect 33140 14068 33192 14074
rect 33140 14010 33192 14016
rect 32956 13728 33008 13734
rect 32956 13670 33008 13676
rect 32968 13394 32996 13670
rect 32956 13388 33008 13394
rect 32956 13330 33008 13336
rect 32864 13320 32916 13326
rect 32864 13262 32916 13268
rect 32968 13274 32996 13330
rect 32968 13246 33088 13274
rect 33060 12850 33088 13246
rect 33324 12980 33376 12986
rect 33324 12922 33376 12928
rect 32956 12844 33008 12850
rect 32956 12786 33008 12792
rect 33048 12844 33100 12850
rect 33048 12786 33100 12792
rect 32968 12442 32996 12786
rect 32036 12436 32088 12442
rect 32036 12378 32088 12384
rect 32956 12436 33008 12442
rect 32956 12378 33008 12384
rect 31576 12368 31628 12374
rect 31312 12294 31432 12322
rect 31628 12316 31708 12322
rect 31576 12310 31708 12316
rect 31588 12294 31708 12310
rect 33336 12306 33364 12922
rect 33428 12306 33456 14894
rect 33520 13938 33548 16118
rect 33692 16040 33744 16046
rect 33692 15982 33744 15988
rect 33508 13932 33560 13938
rect 33508 13874 33560 13880
rect 33704 13870 33732 15982
rect 34072 15162 34100 16118
rect 34348 16046 34376 17070
rect 34440 16794 34468 17138
rect 34428 16788 34480 16794
rect 34428 16730 34480 16736
rect 34440 16250 34468 16730
rect 34428 16244 34480 16250
rect 34428 16186 34480 16192
rect 34336 16040 34388 16046
rect 34336 15982 34388 15988
rect 34060 15156 34112 15162
rect 34060 15098 34112 15104
rect 34072 14550 34100 15098
rect 34244 15020 34296 15026
rect 34244 14962 34296 14968
rect 34060 14544 34112 14550
rect 34060 14486 34112 14492
rect 34072 14074 34100 14486
rect 34060 14068 34112 14074
rect 34060 14010 34112 14016
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33692 13864 33744 13870
rect 33692 13806 33744 13812
rect 33612 12986 33640 13806
rect 33600 12980 33652 12986
rect 33600 12922 33652 12928
rect 31116 12232 31168 12238
rect 31114 12200 31116 12209
rect 31300 12232 31352 12238
rect 31168 12200 31170 12209
rect 31114 12135 31170 12144
rect 31220 12192 31300 12220
rect 30288 11756 30340 11762
rect 30288 11698 30340 11704
rect 30656 11756 30708 11762
rect 30656 11698 30708 11704
rect 30380 11620 30432 11626
rect 30380 11562 30432 11568
rect 29920 11552 29972 11558
rect 29920 11494 29972 11500
rect 30392 10962 30420 11562
rect 31024 11552 31076 11558
rect 31024 11494 31076 11500
rect 30300 10934 30420 10962
rect 29644 10668 29696 10674
rect 29644 10610 29696 10616
rect 30300 10538 30328 10934
rect 31036 10606 31064 11494
rect 31024 10600 31076 10606
rect 31024 10542 31076 10548
rect 30288 10532 30340 10538
rect 30288 10474 30340 10480
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 30116 10062 30144 10406
rect 30196 10192 30248 10198
rect 30196 10134 30248 10140
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 29828 9988 29880 9994
rect 29828 9930 29880 9936
rect 29840 9586 29868 9930
rect 29920 9920 29972 9926
rect 29920 9862 29972 9868
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 29932 9178 29960 9862
rect 30024 9722 30052 9862
rect 30012 9716 30064 9722
rect 30012 9658 30064 9664
rect 30116 9654 30144 9998
rect 30104 9648 30156 9654
rect 30104 9590 30156 9596
rect 29920 9172 29972 9178
rect 29920 9114 29972 9120
rect 29736 7744 29788 7750
rect 29736 7686 29788 7692
rect 29748 7478 29776 7686
rect 29736 7472 29788 7478
rect 29736 7414 29788 7420
rect 29932 7342 29960 9114
rect 30012 8288 30064 8294
rect 30012 8230 30064 8236
rect 30024 7886 30052 8230
rect 30208 7954 30236 10134
rect 30300 10062 30328 10474
rect 30656 10260 30708 10266
rect 30656 10202 30708 10208
rect 30288 10056 30340 10062
rect 30288 9998 30340 10004
rect 30300 9926 30328 9998
rect 30288 9920 30340 9926
rect 30288 9862 30340 9868
rect 30196 7948 30248 7954
rect 30196 7890 30248 7896
rect 30012 7880 30064 7886
rect 30012 7822 30064 7828
rect 30300 7698 30328 9862
rect 30472 9376 30524 9382
rect 30472 9318 30524 9324
rect 30484 7954 30512 9318
rect 30564 8832 30616 8838
rect 30564 8774 30616 8780
rect 30576 8090 30604 8774
rect 30564 8084 30616 8090
rect 30564 8026 30616 8032
rect 30472 7948 30524 7954
rect 30472 7890 30524 7896
rect 30472 7812 30524 7818
rect 30472 7754 30524 7760
rect 30116 7670 30328 7698
rect 29920 7336 29972 7342
rect 29920 7278 29972 7284
rect 29644 6112 29696 6118
rect 29644 6054 29696 6060
rect 29656 5710 29684 6054
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 29564 5494 29684 5522
rect 29000 4548 29052 4554
rect 29000 4490 29052 4496
rect 29012 3466 29040 4490
rect 29000 3460 29052 3466
rect 29000 3402 29052 3408
rect 29552 3392 29604 3398
rect 29552 3334 29604 3340
rect 29564 3126 29592 3334
rect 29552 3120 29604 3126
rect 29552 3062 29604 3068
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 28540 3052 28592 3058
rect 28540 2994 28592 3000
rect 25964 2508 26096 2514
rect 26016 2502 26096 2508
rect 26148 2508 26200 2514
rect 25964 2450 26016 2456
rect 26148 2450 26200 2456
rect 26252 2446 26280 2994
rect 29656 2446 29684 5494
rect 29736 4480 29788 4486
rect 29736 4422 29788 4428
rect 29748 3398 29776 4422
rect 29828 3528 29880 3534
rect 29828 3470 29880 3476
rect 29736 3392 29788 3398
rect 29840 3369 29868 3470
rect 29736 3334 29788 3340
rect 29826 3360 29882 3369
rect 29826 3295 29882 3304
rect 30116 2774 30144 7670
rect 30484 7546 30512 7754
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30380 7404 30432 7410
rect 30380 7346 30432 7352
rect 30564 7404 30616 7410
rect 30564 7346 30616 7352
rect 30392 6730 30420 7346
rect 30576 7290 30604 7346
rect 30484 7262 30604 7290
rect 30380 6724 30432 6730
rect 30380 6666 30432 6672
rect 30196 5296 30248 5302
rect 30196 5238 30248 5244
rect 30208 3534 30236 5238
rect 30288 4140 30340 4146
rect 30484 4128 30512 7262
rect 30564 7200 30616 7206
rect 30564 7142 30616 7148
rect 30576 6866 30604 7142
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30668 5574 30696 10202
rect 31220 10062 31248 12192
rect 31300 12174 31352 12180
rect 31300 11824 31352 11830
rect 31300 11766 31352 11772
rect 31312 11354 31340 11766
rect 31404 11694 31432 12294
rect 31576 12232 31628 12238
rect 31576 12174 31628 12180
rect 31588 11778 31616 12174
rect 31680 11914 31708 12294
rect 33324 12300 33376 12306
rect 33324 12242 33376 12248
rect 33416 12300 33468 12306
rect 33416 12242 33468 12248
rect 32128 12232 32180 12238
rect 32126 12200 32128 12209
rect 32180 12200 32182 12209
rect 32126 12135 32182 12144
rect 31944 12096 31996 12102
rect 31944 12038 31996 12044
rect 32036 12096 32088 12102
rect 32036 12038 32088 12044
rect 31680 11886 31800 11914
rect 31772 11830 31800 11886
rect 31760 11824 31812 11830
rect 31588 11762 31708 11778
rect 31760 11766 31812 11772
rect 31588 11756 31720 11762
rect 31588 11750 31668 11756
rect 31668 11698 31720 11704
rect 31392 11688 31444 11694
rect 31392 11630 31444 11636
rect 31760 11688 31812 11694
rect 31760 11630 31812 11636
rect 31404 11354 31432 11630
rect 31576 11620 31628 11626
rect 31576 11562 31628 11568
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 31392 11348 31444 11354
rect 31392 11290 31444 11296
rect 31484 11212 31536 11218
rect 31484 11154 31536 11160
rect 31392 11144 31444 11150
rect 31392 11086 31444 11092
rect 31300 11076 31352 11082
rect 31300 11018 31352 11024
rect 31312 10674 31340 11018
rect 31404 10674 31432 11086
rect 31496 10810 31524 11154
rect 31484 10804 31536 10810
rect 31484 10746 31536 10752
rect 31300 10668 31352 10674
rect 31300 10610 31352 10616
rect 31392 10668 31444 10674
rect 31392 10610 31444 10616
rect 31024 10056 31076 10062
rect 31024 9998 31076 10004
rect 31208 10056 31260 10062
rect 31208 9998 31260 10004
rect 30748 9988 30800 9994
rect 30748 9930 30800 9936
rect 30760 9586 30788 9930
rect 30748 9580 30800 9586
rect 30748 9522 30800 9528
rect 30932 9376 30984 9382
rect 30932 9318 30984 9324
rect 30944 8974 30972 9318
rect 30932 8968 30984 8974
rect 30932 8910 30984 8916
rect 30748 7880 30800 7886
rect 30748 7822 30800 7828
rect 30840 7880 30892 7886
rect 30840 7822 30892 7828
rect 30760 7546 30788 7822
rect 30748 7540 30800 7546
rect 30748 7482 30800 7488
rect 30852 7410 30880 7822
rect 30840 7404 30892 7410
rect 30840 7346 30892 7352
rect 30748 7336 30800 7342
rect 30746 7304 30748 7313
rect 30800 7304 30802 7313
rect 30746 7239 30802 7248
rect 31036 7002 31064 9998
rect 31404 9926 31432 10610
rect 31392 9920 31444 9926
rect 31392 9862 31444 9868
rect 31588 9722 31616 11562
rect 31772 11506 31800 11630
rect 31956 11626 31984 12038
rect 31944 11620 31996 11626
rect 31944 11562 31996 11568
rect 31680 11478 31800 11506
rect 31680 11218 31708 11478
rect 31668 11212 31720 11218
rect 31668 11154 31720 11160
rect 31956 11150 31984 11562
rect 32048 11150 32076 12038
rect 32140 11778 32168 12135
rect 32140 11750 32260 11778
rect 32128 11688 32180 11694
rect 32128 11630 32180 11636
rect 31944 11144 31996 11150
rect 31944 11086 31996 11092
rect 32036 11144 32088 11150
rect 32036 11086 32088 11092
rect 31956 10690 31984 11086
rect 32140 11082 32168 11630
rect 32232 11558 32260 11750
rect 33140 11756 33192 11762
rect 33140 11698 33192 11704
rect 33152 11665 33180 11698
rect 33138 11656 33194 11665
rect 33138 11591 33194 11600
rect 32220 11552 32272 11558
rect 32220 11494 32272 11500
rect 33152 11354 33180 11591
rect 33140 11348 33192 11354
rect 33140 11290 33192 11296
rect 32220 11144 32272 11150
rect 32220 11086 32272 11092
rect 32128 11076 32180 11082
rect 32128 11018 32180 11024
rect 31668 10668 31720 10674
rect 31956 10662 32076 10690
rect 32232 10674 32260 11086
rect 33232 10736 33284 10742
rect 33232 10678 33284 10684
rect 31668 10610 31720 10616
rect 31680 10130 31708 10610
rect 32048 10606 32076 10662
rect 32220 10668 32272 10674
rect 32220 10610 32272 10616
rect 32864 10668 32916 10674
rect 32864 10610 32916 10616
rect 31944 10600 31996 10606
rect 31944 10542 31996 10548
rect 32036 10600 32088 10606
rect 32036 10542 32088 10548
rect 31852 10464 31904 10470
rect 31852 10406 31904 10412
rect 31668 10124 31720 10130
rect 31668 10066 31720 10072
rect 31760 9920 31812 9926
rect 31760 9862 31812 9868
rect 31576 9716 31628 9722
rect 31576 9658 31628 9664
rect 31772 9586 31800 9862
rect 31760 9580 31812 9586
rect 31760 9522 31812 9528
rect 31864 8906 31892 10406
rect 31956 9926 31984 10542
rect 32036 10192 32088 10198
rect 32036 10134 32088 10140
rect 31944 9920 31996 9926
rect 31944 9862 31996 9868
rect 31956 9722 31984 9862
rect 31944 9716 31996 9722
rect 31944 9658 31996 9664
rect 31852 8900 31904 8906
rect 31852 8842 31904 8848
rect 32048 8634 32076 10134
rect 32232 10062 32260 10610
rect 32680 10464 32732 10470
rect 32680 10406 32732 10412
rect 32692 10062 32720 10406
rect 32876 10062 32904 10610
rect 33244 10606 33272 10678
rect 33428 10674 33456 12242
rect 33508 11688 33560 11694
rect 33506 11656 33508 11665
rect 33560 11656 33562 11665
rect 33506 11591 33562 11600
rect 33600 11552 33652 11558
rect 33600 11494 33652 11500
rect 33612 10674 33640 11494
rect 34256 10810 34284 14962
rect 34532 11014 34560 18158
rect 34624 12646 34652 18702
rect 34716 18358 34744 19722
rect 34704 18352 34756 18358
rect 34704 18294 34756 18300
rect 34716 18086 34744 18294
rect 34808 18222 34836 20198
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35452 19514 35480 27406
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 35440 19508 35492 19514
rect 35440 19450 35492 19456
rect 35348 19372 35400 19378
rect 35348 19314 35400 19320
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18426 35388 19314
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 35452 18290 35480 19450
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35440 18284 35492 18290
rect 35440 18226 35492 18232
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 34704 18080 34756 18086
rect 34704 18022 34756 18028
rect 34704 12844 34756 12850
rect 34704 12786 34756 12792
rect 34612 12640 34664 12646
rect 34612 12582 34664 12588
rect 34624 11762 34652 12582
rect 34716 12442 34744 12786
rect 34704 12436 34756 12442
rect 34704 12378 34756 12384
rect 34808 12102 34836 18158
rect 35348 18080 35400 18086
rect 35348 18022 35400 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34888 12232 34940 12238
rect 34888 12174 34940 12180
rect 34796 12096 34848 12102
rect 34796 12038 34848 12044
rect 34612 11756 34664 11762
rect 34612 11698 34664 11704
rect 34808 11286 34836 12038
rect 34900 11898 34928 12174
rect 34888 11892 34940 11898
rect 34888 11834 34940 11840
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11280 34848 11286
rect 34796 11222 34848 11228
rect 35360 11150 35388 18022
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 36004 12986 36032 33458
rect 36358 33416 36414 33425
rect 36358 33351 36360 33360
rect 36412 33351 36414 33360
rect 36360 33322 36412 33328
rect 36544 30252 36596 30258
rect 36544 30194 36596 30200
rect 36360 30048 36412 30054
rect 36358 30016 36360 30025
rect 36412 30016 36414 30025
rect 36358 29951 36414 29960
rect 36360 27328 36412 27334
rect 36358 27296 36360 27305
rect 36412 27296 36414 27305
rect 36358 27231 36414 27240
rect 36084 24200 36136 24206
rect 36084 24142 36136 24148
rect 35992 12980 36044 12986
rect 35992 12922 36044 12928
rect 36004 12238 36032 12922
rect 35992 12232 36044 12238
rect 35992 12174 36044 12180
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 35348 11144 35400 11150
rect 35348 11086 35400 11092
rect 34520 11008 34572 11014
rect 34520 10950 34572 10956
rect 34704 11008 34756 11014
rect 34704 10950 34756 10956
rect 34244 10804 34296 10810
rect 34244 10746 34296 10752
rect 33968 10736 34020 10742
rect 33968 10678 34020 10684
rect 33416 10668 33468 10674
rect 33416 10610 33468 10616
rect 33600 10668 33652 10674
rect 33600 10610 33652 10616
rect 33784 10668 33836 10674
rect 33784 10610 33836 10616
rect 32956 10600 33008 10606
rect 33232 10600 33284 10606
rect 33008 10560 33088 10588
rect 32956 10542 33008 10548
rect 32220 10056 32272 10062
rect 32220 9998 32272 10004
rect 32680 10056 32732 10062
rect 32680 9998 32732 10004
rect 32864 10056 32916 10062
rect 32864 9998 32916 10004
rect 32956 10056 33008 10062
rect 32956 9998 33008 10004
rect 32312 9376 32364 9382
rect 32312 9318 32364 9324
rect 32128 8832 32180 8838
rect 32128 8774 32180 8780
rect 32036 8628 32088 8634
rect 32036 8570 32088 8576
rect 31852 8492 31904 8498
rect 31852 8434 31904 8440
rect 31668 8356 31720 8362
rect 31668 8298 31720 8304
rect 31116 7880 31168 7886
rect 31116 7822 31168 7828
rect 31208 7880 31260 7886
rect 31208 7822 31260 7828
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 31024 6996 31076 7002
rect 31024 6938 31076 6944
rect 31128 6322 31156 7822
rect 31220 7562 31248 7822
rect 31392 7812 31444 7818
rect 31392 7754 31444 7760
rect 31220 7534 31340 7562
rect 31208 7404 31260 7410
rect 31208 7346 31260 7352
rect 31220 6798 31248 7346
rect 31312 7206 31340 7534
rect 31404 7410 31432 7754
rect 31484 7744 31536 7750
rect 31484 7686 31536 7692
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 31496 6798 31524 7686
rect 31208 6792 31260 6798
rect 31208 6734 31260 6740
rect 31484 6792 31536 6798
rect 31484 6734 31536 6740
rect 31116 6316 31168 6322
rect 31116 6258 31168 6264
rect 30840 6180 30892 6186
rect 30840 6122 30892 6128
rect 30656 5568 30708 5574
rect 30656 5510 30708 5516
rect 30668 5234 30696 5510
rect 30656 5228 30708 5234
rect 30656 5170 30708 5176
rect 30564 4208 30616 4214
rect 30564 4150 30616 4156
rect 30340 4100 30512 4128
rect 30288 4082 30340 4088
rect 30300 3890 30328 4082
rect 30380 4004 30432 4010
rect 30432 3964 30512 3992
rect 30380 3946 30432 3952
rect 30300 3862 30420 3890
rect 30392 3738 30420 3862
rect 30288 3732 30340 3738
rect 30288 3674 30340 3680
rect 30380 3732 30432 3738
rect 30380 3674 30432 3680
rect 30196 3528 30248 3534
rect 30196 3470 30248 3476
rect 30300 2854 30328 3674
rect 30392 3058 30420 3674
rect 30484 3602 30512 3964
rect 30472 3596 30524 3602
rect 30472 3538 30524 3544
rect 30484 3194 30512 3538
rect 30576 3194 30604 4150
rect 30668 3482 30696 5170
rect 30852 4128 30880 6122
rect 31024 6112 31076 6118
rect 31024 6054 31076 6060
rect 31036 5778 31064 6054
rect 31024 5772 31076 5778
rect 31024 5714 31076 5720
rect 31220 5574 31248 6734
rect 31392 6656 31444 6662
rect 31392 6598 31444 6604
rect 31404 6322 31432 6598
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 31392 6316 31444 6322
rect 31392 6258 31444 6264
rect 31312 6202 31340 6258
rect 31312 6174 31432 6202
rect 31300 6112 31352 6118
rect 31300 6054 31352 6060
rect 31312 5914 31340 6054
rect 31300 5908 31352 5914
rect 31300 5850 31352 5856
rect 31116 5568 31168 5574
rect 31116 5510 31168 5516
rect 31208 5568 31260 5574
rect 31208 5510 31260 5516
rect 31128 5166 31156 5510
rect 31116 5160 31168 5166
rect 31116 5102 31168 5108
rect 31116 4752 31168 4758
rect 31116 4694 31168 4700
rect 31128 4214 31156 4694
rect 31116 4208 31168 4214
rect 31116 4150 31168 4156
rect 30932 4140 30984 4146
rect 30852 4100 30932 4128
rect 30932 4082 30984 4088
rect 30748 3936 30800 3942
rect 30748 3878 30800 3884
rect 30760 3602 30788 3878
rect 30748 3596 30800 3602
rect 30748 3538 30800 3544
rect 30944 3534 30972 4082
rect 30840 3528 30892 3534
rect 30838 3496 30840 3505
rect 30932 3528 30984 3534
rect 30892 3496 30894 3505
rect 30668 3454 30788 3482
rect 30656 3392 30708 3398
rect 30656 3334 30708 3340
rect 30668 3194 30696 3334
rect 30472 3188 30524 3194
rect 30472 3130 30524 3136
rect 30564 3188 30616 3194
rect 30564 3130 30616 3136
rect 30656 3188 30708 3194
rect 30656 3130 30708 3136
rect 30380 3052 30432 3058
rect 30380 2994 30432 3000
rect 30196 2848 30248 2854
rect 30196 2790 30248 2796
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 29932 2746 30144 2774
rect 29932 2582 29960 2746
rect 29920 2576 29972 2582
rect 29920 2518 29972 2524
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 25320 2440 25372 2446
rect 25320 2382 25372 2388
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 19156 2372 19208 2378
rect 19156 2314 19208 2320
rect 21284 800 21312 2382
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 23860 800 23888 2246
rect 27080 800 27108 2382
rect 30208 2378 30236 2790
rect 30484 2582 30512 3130
rect 30472 2576 30524 2582
rect 30472 2518 30524 2524
rect 30196 2372 30248 2378
rect 30196 2314 30248 2320
rect 30380 2304 30432 2310
rect 30380 2246 30432 2252
rect 30392 1442 30420 2246
rect 30760 2038 30788 3454
rect 30932 3470 30984 3476
rect 30838 3431 30894 3440
rect 30944 3058 30972 3470
rect 31128 3398 31156 4150
rect 31220 4078 31248 5510
rect 31312 5302 31340 5850
rect 31300 5296 31352 5302
rect 31300 5238 31352 5244
rect 31300 5024 31352 5030
rect 31300 4966 31352 4972
rect 31312 4622 31340 4966
rect 31300 4616 31352 4622
rect 31300 4558 31352 4564
rect 31208 4072 31260 4078
rect 31208 4014 31260 4020
rect 31300 3732 31352 3738
rect 31300 3674 31352 3680
rect 31312 3534 31340 3674
rect 31404 3534 31432 6174
rect 31496 5370 31524 6734
rect 31588 6322 31616 7822
rect 31680 7342 31708 8298
rect 31760 8084 31812 8090
rect 31760 8026 31812 8032
rect 31772 7392 31800 8026
rect 31864 7886 31892 8434
rect 31944 8288 31996 8294
rect 31944 8230 31996 8236
rect 31852 7880 31904 7886
rect 31852 7822 31904 7828
rect 31956 7750 31984 8230
rect 32048 7886 32076 8570
rect 32140 8566 32168 8774
rect 32128 8560 32180 8566
rect 32128 8502 32180 8508
rect 32036 7880 32088 7886
rect 32036 7822 32088 7828
rect 32140 7834 32168 8502
rect 32048 7750 32076 7822
rect 32140 7818 32260 7834
rect 32140 7812 32272 7818
rect 32140 7806 32220 7812
rect 32220 7754 32272 7760
rect 31944 7744 31996 7750
rect 31944 7686 31996 7692
rect 32036 7744 32088 7750
rect 32036 7686 32088 7692
rect 31944 7404 31996 7410
rect 31772 7364 31944 7392
rect 32324 7392 32352 9318
rect 32968 8634 32996 9998
rect 33060 9586 33088 10560
rect 33232 10542 33284 10548
rect 33140 10532 33192 10538
rect 33140 10474 33192 10480
rect 33152 10130 33180 10474
rect 33140 10124 33192 10130
rect 33192 10084 33272 10112
rect 33140 10066 33192 10072
rect 33140 9920 33192 9926
rect 33140 9862 33192 9868
rect 33152 9654 33180 9862
rect 33140 9648 33192 9654
rect 33140 9590 33192 9596
rect 33048 9580 33100 9586
rect 33048 9522 33100 9528
rect 33060 8838 33088 9522
rect 33244 9518 33272 10084
rect 33232 9512 33284 9518
rect 33232 9454 33284 9460
rect 33428 9382 33456 10610
rect 33612 10554 33640 10610
rect 33520 10538 33640 10554
rect 33508 10532 33640 10538
rect 33560 10526 33640 10532
rect 33508 10474 33560 10480
rect 33796 10470 33824 10610
rect 33876 10600 33928 10606
rect 33876 10542 33928 10548
rect 33600 10464 33652 10470
rect 33600 10406 33652 10412
rect 33784 10464 33836 10470
rect 33784 10406 33836 10412
rect 33612 9654 33640 10406
rect 33784 10124 33836 10130
rect 33784 10066 33836 10072
rect 33692 10056 33744 10062
rect 33692 9998 33744 10004
rect 33704 9722 33732 9998
rect 33692 9716 33744 9722
rect 33692 9658 33744 9664
rect 33600 9648 33652 9654
rect 33600 9590 33652 9596
rect 33140 9376 33192 9382
rect 33140 9318 33192 9324
rect 33416 9376 33468 9382
rect 33416 9318 33468 9324
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 32956 8628 33008 8634
rect 32956 8570 33008 8576
rect 33060 8566 33088 8774
rect 33048 8560 33100 8566
rect 33048 8502 33100 8508
rect 32864 8492 32916 8498
rect 32864 8434 32916 8440
rect 32404 8424 32456 8430
rect 32404 8366 32456 8372
rect 32416 8294 32444 8366
rect 32404 8288 32456 8294
rect 32404 8230 32456 8236
rect 32496 8288 32548 8294
rect 32496 8230 32548 8236
rect 32404 7404 32456 7410
rect 32324 7364 32404 7392
rect 31944 7346 31996 7352
rect 32404 7346 32456 7352
rect 31668 7336 31720 7342
rect 31668 7278 31720 7284
rect 31760 7268 31812 7274
rect 31760 7210 31812 7216
rect 31772 6866 31800 7210
rect 31760 6860 31812 6866
rect 31760 6802 31812 6808
rect 31668 6792 31720 6798
rect 31668 6734 31720 6740
rect 31576 6316 31628 6322
rect 31576 6258 31628 6264
rect 31484 5364 31536 5370
rect 31484 5306 31536 5312
rect 31588 3618 31616 6258
rect 31680 5846 31708 6734
rect 31772 5846 31800 6802
rect 31852 6180 31904 6186
rect 31852 6122 31904 6128
rect 31864 5914 31892 6122
rect 31956 6118 31984 7346
rect 32508 7274 32536 8230
rect 32680 7812 32732 7818
rect 32680 7754 32732 7760
rect 32692 7410 32720 7754
rect 32876 7750 32904 8434
rect 32956 8016 33008 8022
rect 32956 7958 33008 7964
rect 32968 7818 32996 7958
rect 32956 7812 33008 7818
rect 32956 7754 33008 7760
rect 32864 7744 32916 7750
rect 32864 7686 32916 7692
rect 32680 7404 32732 7410
rect 32680 7346 32732 7352
rect 32496 7268 32548 7274
rect 32496 7210 32548 7216
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 31944 6112 31996 6118
rect 31944 6054 31996 6060
rect 31852 5908 31904 5914
rect 31852 5850 31904 5856
rect 31668 5840 31720 5846
rect 31668 5782 31720 5788
rect 31760 5840 31812 5846
rect 31760 5782 31812 5788
rect 31680 5624 31708 5782
rect 32324 5710 32352 7142
rect 33152 6458 33180 9318
rect 33598 8256 33654 8265
rect 33598 8191 33654 8200
rect 33612 8022 33640 8191
rect 33600 8016 33652 8022
rect 33600 7958 33652 7964
rect 33324 7880 33376 7886
rect 33324 7822 33376 7828
rect 33336 7546 33364 7822
rect 33692 7812 33744 7818
rect 33692 7754 33744 7760
rect 33704 7546 33732 7754
rect 33324 7540 33376 7546
rect 33324 7482 33376 7488
rect 33692 7540 33744 7546
rect 33692 7482 33744 7488
rect 33796 7410 33824 10066
rect 33888 9602 33916 10542
rect 33980 10470 34008 10678
rect 34152 10668 34204 10674
rect 34152 10610 34204 10616
rect 33968 10464 34020 10470
rect 33968 10406 34020 10412
rect 33980 10130 34008 10406
rect 33968 10124 34020 10130
rect 33968 10066 34020 10072
rect 33888 9574 34008 9602
rect 33876 9376 33928 9382
rect 33876 9318 33928 9324
rect 33888 7478 33916 9318
rect 33876 7472 33928 7478
rect 33876 7414 33928 7420
rect 33784 7404 33836 7410
rect 33784 7346 33836 7352
rect 33600 6996 33652 7002
rect 33600 6938 33652 6944
rect 33140 6452 33192 6458
rect 33140 6394 33192 6400
rect 33612 5914 33640 6938
rect 33796 6934 33824 7346
rect 33980 7342 34008 9574
rect 34060 8016 34112 8022
rect 34060 7958 34112 7964
rect 34072 7818 34100 7958
rect 34060 7812 34112 7818
rect 34060 7754 34112 7760
rect 33968 7336 34020 7342
rect 33874 7304 33930 7313
rect 33968 7278 34020 7284
rect 33874 7239 33930 7248
rect 33784 6928 33836 6934
rect 33784 6870 33836 6876
rect 33888 6798 33916 7239
rect 33876 6792 33928 6798
rect 33876 6734 33928 6740
rect 33968 6656 34020 6662
rect 33968 6598 34020 6604
rect 33980 6458 34008 6598
rect 33968 6452 34020 6458
rect 33968 6394 34020 6400
rect 33600 5908 33652 5914
rect 33600 5850 33652 5856
rect 31944 5704 31996 5710
rect 32220 5704 32272 5710
rect 31944 5646 31996 5652
rect 32218 5672 32220 5681
rect 32312 5704 32364 5710
rect 32272 5672 32274 5681
rect 31852 5636 31904 5642
rect 31680 5596 31852 5624
rect 31680 4758 31708 5596
rect 31852 5578 31904 5584
rect 31956 5370 31984 5646
rect 32312 5646 32364 5652
rect 32218 5607 32274 5616
rect 31944 5364 31996 5370
rect 31944 5306 31996 5312
rect 32232 5234 32260 5607
rect 32220 5228 32272 5234
rect 32220 5170 32272 5176
rect 32772 5228 32824 5234
rect 32772 5170 32824 5176
rect 31668 4752 31720 4758
rect 31668 4694 31720 4700
rect 31852 3732 31904 3738
rect 31852 3674 31904 3680
rect 31588 3602 31708 3618
rect 31588 3596 31720 3602
rect 31588 3590 31668 3596
rect 31668 3538 31720 3544
rect 31300 3528 31352 3534
rect 31300 3470 31352 3476
rect 31392 3528 31444 3534
rect 31392 3470 31444 3476
rect 31484 3528 31536 3534
rect 31484 3470 31536 3476
rect 31116 3392 31168 3398
rect 31116 3334 31168 3340
rect 31208 3392 31260 3398
rect 31300 3392 31352 3398
rect 31208 3334 31260 3340
rect 31298 3360 31300 3369
rect 31352 3360 31354 3369
rect 30932 3052 30984 3058
rect 30932 2994 30984 3000
rect 31220 2582 31248 3334
rect 31298 3295 31354 3304
rect 31404 3058 31432 3470
rect 31496 3126 31524 3470
rect 31576 3460 31628 3466
rect 31576 3402 31628 3408
rect 31588 3194 31616 3402
rect 31680 3380 31708 3538
rect 31864 3534 31892 3674
rect 32220 3664 32272 3670
rect 32220 3606 32272 3612
rect 31852 3528 31904 3534
rect 31850 3496 31852 3505
rect 31904 3496 31906 3505
rect 32232 3466 32260 3606
rect 32784 3534 32812 5170
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 32772 3528 32824 3534
rect 32772 3470 32824 3476
rect 31850 3431 31906 3440
rect 32220 3460 32272 3466
rect 32220 3402 32272 3408
rect 31760 3392 31812 3398
rect 31680 3352 31760 3380
rect 31576 3188 31628 3194
rect 31576 3130 31628 3136
rect 31484 3120 31536 3126
rect 31484 3062 31536 3068
rect 31680 3058 31708 3352
rect 31760 3334 31812 3340
rect 32416 3126 32444 3470
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 32784 3058 32812 3470
rect 34164 3194 34192 10610
rect 34716 10606 34744 10950
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 35900 10804 35952 10810
rect 35900 10746 35952 10752
rect 34796 10668 34848 10674
rect 34796 10610 34848 10616
rect 34704 10600 34756 10606
rect 34704 10542 34756 10548
rect 34336 10056 34388 10062
rect 34336 9998 34388 10004
rect 34348 9518 34376 9998
rect 34244 9512 34296 9518
rect 34244 9454 34296 9460
rect 34336 9512 34388 9518
rect 34336 9454 34388 9460
rect 34256 9178 34284 9454
rect 34244 9172 34296 9178
rect 34244 9114 34296 9120
rect 34256 8566 34284 9114
rect 34348 8634 34376 9454
rect 34336 8628 34388 8634
rect 34336 8570 34388 8576
rect 34244 8560 34296 8566
rect 34244 8502 34296 8508
rect 34348 7410 34376 8570
rect 34612 8356 34664 8362
rect 34612 8298 34664 8304
rect 34520 7880 34572 7886
rect 34520 7822 34572 7828
rect 34532 7750 34560 7822
rect 34520 7744 34572 7750
rect 34520 7686 34572 7692
rect 34532 7410 34560 7686
rect 34624 7546 34652 8298
rect 34716 7886 34744 10542
rect 34808 10266 34836 10610
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 10260 34848 10266
rect 34796 10202 34848 10208
rect 35912 10062 35940 10746
rect 35900 10056 35952 10062
rect 35900 9998 35952 10004
rect 34888 9920 34940 9926
rect 34888 9862 34940 9868
rect 34900 9722 34928 9862
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 34888 9716 34940 9722
rect 34888 9658 34940 9664
rect 34900 9466 34928 9658
rect 34808 9438 34928 9466
rect 34704 7880 34756 7886
rect 34704 7822 34756 7828
rect 34612 7540 34664 7546
rect 34612 7482 34664 7488
rect 34336 7404 34388 7410
rect 34336 7346 34388 7352
rect 34520 7404 34572 7410
rect 34520 7346 34572 7352
rect 34716 5778 34744 7822
rect 34808 7546 34836 9438
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 34796 7540 34848 7546
rect 34796 7482 34848 7488
rect 34796 7336 34848 7342
rect 34796 7278 34848 7284
rect 34808 6798 34836 7278
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34796 6792 34848 6798
rect 34796 6734 34848 6740
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34704 5772 34756 5778
rect 34704 5714 34756 5720
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 36096 3738 36124 24142
rect 36360 24064 36412 24070
rect 36360 24006 36412 24012
rect 36372 23905 36400 24006
rect 36358 23896 36414 23905
rect 36358 23831 36414 23840
rect 36268 20868 36320 20874
rect 36268 20810 36320 20816
rect 36176 16992 36228 16998
rect 36176 16934 36228 16940
rect 36188 15026 36216 16934
rect 36176 15020 36228 15026
rect 36176 14962 36228 14968
rect 36280 12434 36308 20810
rect 36360 20800 36412 20806
rect 36360 20742 36412 20748
rect 36372 20505 36400 20742
rect 36358 20496 36414 20505
rect 36358 20431 36414 20440
rect 36452 17196 36504 17202
rect 36452 17138 36504 17144
rect 36464 17105 36492 17138
rect 36450 17096 36506 17105
rect 36450 17031 36506 17040
rect 36358 14376 36414 14385
rect 36358 14311 36414 14320
rect 36372 14278 36400 14311
rect 36360 14272 36412 14278
rect 36360 14214 36412 14220
rect 36280 12406 36400 12434
rect 36268 11756 36320 11762
rect 36268 11698 36320 11704
rect 36280 11354 36308 11698
rect 36268 11348 36320 11354
rect 36268 11290 36320 11296
rect 36372 10810 36400 12406
rect 36452 11144 36504 11150
rect 36452 11086 36504 11092
rect 36464 10985 36492 11086
rect 36450 10976 36506 10985
rect 36450 10911 36506 10920
rect 36360 10804 36412 10810
rect 36360 10746 36412 10752
rect 36176 9036 36228 9042
rect 36176 8978 36228 8984
rect 36188 5234 36216 8978
rect 36452 7880 36504 7886
rect 36266 7848 36322 7857
rect 36452 7822 36504 7828
rect 36266 7783 36322 7792
rect 36280 7750 36308 7783
rect 36268 7744 36320 7750
rect 36268 7686 36320 7692
rect 36464 7585 36492 7822
rect 36450 7576 36506 7585
rect 36450 7511 36506 7520
rect 36556 5370 36584 30194
rect 36544 5364 36596 5370
rect 36544 5306 36596 5312
rect 36176 5228 36228 5234
rect 36176 5170 36228 5176
rect 36360 5024 36412 5030
rect 36360 4966 36412 4972
rect 36372 4865 36400 4966
rect 36358 4856 36414 4865
rect 36358 4791 36414 4800
rect 36084 3732 36136 3738
rect 36084 3674 36136 3680
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 34152 3188 34204 3194
rect 34152 3130 34204 3136
rect 31392 3052 31444 3058
rect 31392 2994 31444 3000
rect 31668 3052 31720 3058
rect 31668 2994 31720 3000
rect 32772 3052 32824 3058
rect 32772 2994 32824 3000
rect 33048 3052 33100 3058
rect 33048 2994 33100 3000
rect 33060 2650 33088 2994
rect 35440 2916 35492 2922
rect 35440 2858 35492 2864
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 33048 2644 33100 2650
rect 33048 2586 33100 2592
rect 31208 2576 31260 2582
rect 31208 2518 31260 2524
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 30748 2032 30800 2038
rect 30748 1974 30800 1980
rect 30300 1414 30420 1442
rect 30300 800 30328 1414
rect 32876 800 32904 2382
rect 35452 1465 35480 2858
rect 35898 2544 35954 2553
rect 35898 2479 35954 2488
rect 36084 2508 36136 2514
rect 35912 2446 35940 2479
rect 36084 2450 36136 2456
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 35438 1456 35494 1465
rect 35438 1391 35494 1400
rect 36096 800 36124 2450
rect 18 0 74 800
rect 2594 0 2650 800
rect 5814 0 5870 800
rect 9034 0 9090 800
rect 11610 0 11666 800
rect 14830 0 14886 800
rect 18050 0 18106 800
rect 21270 0 21326 800
rect 23846 0 23902 800
rect 27066 0 27122 800
rect 30286 0 30342 800
rect 32862 0 32918 800
rect 36082 0 36138 800
<< via2 >>
rect 938 38120 994 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 938 34720 994 34776
rect 938 32000 994 32056
rect 1582 28600 1638 28656
rect 1398 25200 1454 25256
rect 938 22500 994 22536
rect 938 22480 940 22500
rect 940 22480 992 22500
rect 992 22480 994 22500
rect 938 19116 940 19136
rect 940 19116 992 19136
rect 992 19116 994 19136
rect 938 19080 994 19116
rect 938 15680 994 15736
rect 1582 12280 1638 12336
rect 1582 9560 1638 9616
rect 1766 12144 1822 12200
rect 1306 6160 1362 6216
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 6918 32292 6974 32328
rect 6918 32272 6920 32292
rect 6920 32272 6972 32292
rect 6972 32272 6974 32292
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 7102 30368 7158 30424
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 5354 18264 5410 18320
rect 5538 18264 5594 18320
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4158 11756 4214 11792
rect 4158 11736 4160 11756
rect 4160 11736 4212 11756
rect 4212 11736 4214 11756
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 6642 18128 6698 18184
rect 7010 19216 7066 19272
rect 8114 31728 8170 31784
rect 7194 21800 7250 21856
rect 7562 18128 7618 18184
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 5722 12008 5778 12064
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 8390 23740 8392 23760
rect 8392 23740 8444 23760
rect 8444 23740 8446 23760
rect 8390 23704 8446 23740
rect 9126 23724 9182 23760
rect 9126 23704 9128 23724
rect 9128 23704 9180 23724
rect 9180 23704 9182 23724
rect 8850 18300 8852 18320
rect 8852 18300 8904 18320
rect 8904 18300 8906 18320
rect 8850 18264 8906 18300
rect 9678 32272 9734 32328
rect 10230 19216 10286 19272
rect 10138 18148 10194 18184
rect 10138 18128 10140 18148
rect 10140 18128 10192 18148
rect 10192 18128 10194 18148
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 6090 5752 6146 5808
rect 8390 12008 8446 12064
rect 10690 18284 10746 18320
rect 10690 18264 10692 18284
rect 10692 18264 10744 18284
rect 10744 18264 10746 18284
rect 11610 23724 11666 23760
rect 11610 23704 11612 23724
rect 11612 23704 11664 23724
rect 11664 23704 11666 23724
rect 11702 18264 11758 18320
rect 9218 5772 9274 5808
rect 9218 5752 9220 5772
rect 9220 5752 9272 5772
rect 9272 5752 9274 5772
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4250 2916 4306 2952
rect 4250 2896 4252 2916
rect 4252 2896 4304 2916
rect 4304 2896 4306 2916
rect 938 2760 994 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 11518 13812 11520 13832
rect 11520 13812 11572 13832
rect 11572 13812 11574 13832
rect 11518 13776 11574 13812
rect 11794 12300 11850 12336
rect 11794 12280 11796 12300
rect 11796 12280 11848 12300
rect 11848 12280 11850 12300
rect 11702 11892 11758 11928
rect 11702 11872 11704 11892
rect 11704 11872 11756 11892
rect 11756 11872 11758 11892
rect 10322 10668 10378 10704
rect 10322 10648 10324 10668
rect 10324 10648 10376 10668
rect 10376 10648 10378 10668
rect 10506 9580 10562 9616
rect 10506 9560 10508 9580
rect 10508 9560 10560 9580
rect 10560 9560 10562 9580
rect 11610 8916 11612 8936
rect 11612 8916 11664 8936
rect 11664 8916 11666 8936
rect 11610 8880 11666 8916
rect 14186 33108 14242 33144
rect 14186 33088 14188 33108
rect 14188 33088 14240 33108
rect 14240 33088 14242 33108
rect 13818 31864 13874 31920
rect 14738 31884 14794 31920
rect 14738 31864 14740 31884
rect 14740 31864 14792 31884
rect 14792 31864 14794 31884
rect 15290 31764 15292 31784
rect 15292 31764 15344 31784
rect 15344 31764 15346 31784
rect 15290 31728 15346 31764
rect 14922 25780 14924 25800
rect 14924 25780 14976 25800
rect 14976 25780 14978 25800
rect 14922 25744 14978 25780
rect 13174 21664 13230 21720
rect 13450 19252 13452 19272
rect 13452 19252 13504 19272
rect 13504 19252 13506 19272
rect 13450 19216 13506 19252
rect 13726 22208 13782 22264
rect 13726 20848 13782 20904
rect 13634 17992 13690 18048
rect 16118 21120 16174 21176
rect 16026 20984 16082 21040
rect 14278 18944 14334 19000
rect 14462 18264 14518 18320
rect 14554 18028 14556 18048
rect 14556 18028 14608 18048
rect 14608 18028 14610 18048
rect 14554 17992 14610 18028
rect 13174 13948 13176 13968
rect 13176 13948 13228 13968
rect 13228 13948 13230 13968
rect 13174 13912 13230 13948
rect 14186 13948 14188 13968
rect 14188 13948 14240 13968
rect 14240 13948 14242 13968
rect 14186 13912 14242 13948
rect 13266 13776 13322 13832
rect 14002 12280 14058 12336
rect 12622 8492 12678 8528
rect 12622 8472 12624 8492
rect 12624 8472 12676 8492
rect 12676 8472 12678 8492
rect 12898 8880 12954 8936
rect 16210 9560 16266 9616
rect 16854 21800 16910 21856
rect 17774 31900 17776 31920
rect 17776 31900 17828 31920
rect 17828 31900 17830 31920
rect 17774 31864 17830 31900
rect 18234 31764 18236 31784
rect 18236 31764 18288 31784
rect 18288 31764 18290 31784
rect 18234 31728 18290 31764
rect 17222 22092 17278 22128
rect 17222 22072 17224 22092
rect 17224 22072 17276 22092
rect 17276 22072 17278 22092
rect 16946 21664 17002 21720
rect 16762 20984 16818 21040
rect 16946 20984 17002 21040
rect 17130 20324 17186 20360
rect 17130 20304 17132 20324
rect 17132 20304 17184 20324
rect 17184 20304 17186 20324
rect 17038 18828 17094 18864
rect 17038 18808 17040 18828
rect 17040 18808 17092 18828
rect 17092 18808 17094 18828
rect 17406 20460 17462 20496
rect 17406 20440 17408 20460
rect 17408 20440 17460 20460
rect 17460 20440 17462 20460
rect 17682 25492 17738 25528
rect 17682 25472 17684 25492
rect 17684 25472 17736 25492
rect 17736 25472 17738 25492
rect 17590 22208 17646 22264
rect 17590 21120 17646 21176
rect 18326 25780 18328 25800
rect 18328 25780 18380 25800
rect 18380 25780 18382 25800
rect 18326 25744 18382 25780
rect 17866 20848 17922 20904
rect 17866 20304 17922 20360
rect 17866 18284 17922 18320
rect 17866 18264 17868 18284
rect 17868 18264 17920 18284
rect 17920 18264 17922 18284
rect 16486 8472 16542 8528
rect 18418 20440 18474 20496
rect 19338 21392 19394 21448
rect 19430 18264 19486 18320
rect 19982 32972 20038 33008
rect 19982 32952 19984 32972
rect 19984 32952 20036 32972
rect 20036 32952 20038 32972
rect 20994 33088 21050 33144
rect 20350 27920 20406 27976
rect 21362 33088 21418 33144
rect 19706 20984 19762 21040
rect 19982 21664 20038 21720
rect 20258 19352 20314 19408
rect 20810 19388 20812 19408
rect 20812 19388 20864 19408
rect 20864 19388 20866 19408
rect 20810 19352 20866 19388
rect 20534 19216 20590 19272
rect 20534 18944 20590 19000
rect 20810 18264 20866 18320
rect 18786 11192 18842 11248
rect 19062 10648 19118 10704
rect 17498 3440 17554 3496
rect 18050 3476 18052 3496
rect 18052 3476 18104 3496
rect 18104 3476 18106 3496
rect 18050 3440 18106 3476
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 19246 11872 19302 11928
rect 19890 12164 19946 12200
rect 19890 12144 19892 12164
rect 19892 12144 19944 12164
rect 19944 12144 19946 12164
rect 20994 21428 20996 21448
rect 20996 21428 21048 21448
rect 21048 21428 21050 21448
rect 20994 21392 21050 21428
rect 20994 20304 21050 20360
rect 21086 19216 21142 19272
rect 22466 25472 22522 25528
rect 22282 20340 22284 20360
rect 22284 20340 22336 20360
rect 22336 20340 22338 20360
rect 22282 20304 22338 20340
rect 23570 27532 23626 27568
rect 23570 27512 23572 27532
rect 23572 27512 23624 27532
rect 23624 27512 23626 27532
rect 21086 12280 21142 12336
rect 20902 11736 20958 11792
rect 20258 11092 20260 11112
rect 20260 11092 20312 11112
rect 20312 11092 20314 11112
rect 20258 11056 20314 11092
rect 22006 12280 22062 12336
rect 23662 23704 23718 23760
rect 23386 23432 23442 23488
rect 25870 36488 25926 36544
rect 24306 32952 24362 33008
rect 25226 31864 25282 31920
rect 24950 27920 25006 27976
rect 24306 20460 24362 20496
rect 24306 20440 24308 20460
rect 24308 20440 24360 20460
rect 24360 20440 24362 20460
rect 23110 18944 23166 19000
rect 23662 18164 23664 18184
rect 23664 18164 23716 18184
rect 23716 18164 23718 18184
rect 23662 18128 23718 18164
rect 22282 11756 22338 11792
rect 22282 11736 22284 11756
rect 22284 11736 22336 11756
rect 22336 11736 22338 11756
rect 19982 9832 20038 9888
rect 19798 7792 19854 7848
rect 21270 10104 21326 10160
rect 21730 9832 21786 9888
rect 21546 9716 21602 9752
rect 21546 9696 21548 9716
rect 21548 9696 21600 9716
rect 21600 9696 21602 9716
rect 25318 24284 25320 24304
rect 25320 24284 25372 24304
rect 25372 24284 25374 24304
rect 25318 24248 25374 24284
rect 25318 23588 25374 23624
rect 25318 23568 25320 23588
rect 25320 23568 25372 23588
rect 25372 23568 25374 23588
rect 25042 18828 25098 18864
rect 25042 18808 25044 18828
rect 25044 18808 25096 18828
rect 25096 18808 25098 18828
rect 26238 24268 26294 24304
rect 26238 24248 26240 24268
rect 26240 24248 26292 24268
rect 26292 24248 26294 24268
rect 25962 21004 26018 21040
rect 25962 20984 25964 21004
rect 25964 20984 26016 21004
rect 26016 20984 26018 21004
rect 26882 27532 26938 27568
rect 26882 27512 26884 27532
rect 26884 27512 26936 27532
rect 26936 27512 26938 27532
rect 25870 19372 25926 19408
rect 25870 19352 25872 19372
rect 25872 19352 25924 19372
rect 25924 19352 25926 19372
rect 26054 19216 26110 19272
rect 25870 18672 25926 18728
rect 26422 19116 26424 19136
rect 26424 19116 26476 19136
rect 26476 19116 26478 19136
rect 26422 19080 26478 19116
rect 26146 18808 26202 18864
rect 24122 11736 24178 11792
rect 24398 9696 24454 9752
rect 24766 10124 24822 10160
rect 24766 10104 24768 10124
rect 24768 10104 24820 10124
rect 24820 10104 24822 10124
rect 25502 13796 25558 13832
rect 25502 13776 25504 13796
rect 25504 13776 25556 13796
rect 25556 13776 25558 13796
rect 25410 13096 25466 13152
rect 26790 20440 26846 20496
rect 27618 23588 27674 23624
rect 27618 23568 27620 23588
rect 27620 23568 27672 23588
rect 27672 23568 27674 23588
rect 27066 19252 27068 19272
rect 27068 19252 27120 19272
rect 27120 19252 27122 19272
rect 27066 19216 27122 19252
rect 28354 19216 28410 19272
rect 26974 18400 27030 18456
rect 26146 13132 26148 13152
rect 26148 13132 26200 13152
rect 26200 13132 26202 13152
rect 26146 13096 26202 13132
rect 28538 18944 28594 19000
rect 28446 18672 28502 18728
rect 28538 18400 28594 18456
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 30838 36116 30840 36136
rect 30840 36116 30892 36136
rect 30892 36116 30894 36136
rect 30838 36080 30894 36116
rect 28814 23432 28870 23488
rect 30838 20576 30894 20632
rect 28722 11192 28778 11248
rect 23938 2896 23994 2952
rect 29458 5652 29460 5672
rect 29460 5652 29512 5672
rect 29512 5652 29514 5672
rect 29458 5616 29514 5652
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 36358 36760 36414 36816
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 31114 12180 31116 12200
rect 31116 12180 31168 12200
rect 31168 12180 31170 12200
rect 31114 12144 31170 12180
rect 29826 3304 29882 3360
rect 32126 12180 32128 12200
rect 32128 12180 32180 12200
rect 32180 12180 32182 12200
rect 32126 12144 32182 12180
rect 30746 7284 30748 7304
rect 30748 7284 30800 7304
rect 30800 7284 30802 7304
rect 30746 7248 30802 7284
rect 33138 11600 33194 11656
rect 33506 11636 33508 11656
rect 33508 11636 33560 11656
rect 33560 11636 33562 11656
rect 33506 11600 33562 11636
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 36358 33380 36414 33416
rect 36358 33360 36360 33380
rect 36360 33360 36412 33380
rect 36412 33360 36414 33380
rect 36358 29996 36360 30016
rect 36360 29996 36412 30016
rect 36412 29996 36414 30016
rect 36358 29960 36414 29996
rect 36358 27276 36360 27296
rect 36360 27276 36412 27296
rect 36412 27276 36414 27296
rect 36358 27240 36414 27276
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 30838 3476 30840 3496
rect 30840 3476 30892 3496
rect 30892 3476 30894 3496
rect 30838 3440 30894 3476
rect 33598 8200 33654 8256
rect 33874 7248 33930 7304
rect 32218 5652 32220 5672
rect 32220 5652 32272 5672
rect 32272 5652 32274 5672
rect 32218 5616 32274 5652
rect 31298 3340 31300 3360
rect 31300 3340 31352 3360
rect 31352 3340 31354 3360
rect 31298 3304 31354 3340
rect 31850 3476 31852 3496
rect 31852 3476 31904 3496
rect 31904 3476 31906 3496
rect 31850 3440 31906 3476
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 36358 23840 36414 23896
rect 36358 20440 36414 20496
rect 36450 17040 36506 17096
rect 36358 14320 36414 14376
rect 36450 10920 36506 10976
rect 36266 7792 36322 7848
rect 36450 7520 36506 7576
rect 36358 4800 36414 4856
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35898 2488 35954 2544
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 35438 1400 35494 1456
<< metal3 >>
rect 0 38178 800 38208
rect 933 38178 999 38181
rect 0 38176 999 38178
rect 0 38120 938 38176
rect 994 38120 999 38176
rect 0 38118 999 38120
rect 0 38088 800 38118
rect 933 38115 999 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 36353 36818 36419 36821
rect 37136 36818 37936 36848
rect 36353 36816 37936 36818
rect 36353 36760 36358 36816
rect 36414 36760 37936 36816
rect 36353 36758 37936 36760
rect 36353 36755 36419 36758
rect 37136 36728 37936 36758
rect 25630 36484 25636 36548
rect 25700 36546 25706 36548
rect 25865 36546 25931 36549
rect 25700 36544 25931 36546
rect 25700 36488 25870 36544
rect 25926 36488 25931 36544
rect 25700 36486 25931 36488
rect 25700 36484 25706 36486
rect 25865 36483 25931 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 30833 36138 30899 36141
rect 30966 36138 30972 36140
rect 30833 36136 30972 36138
rect 30833 36080 30838 36136
rect 30894 36080 30972 36136
rect 30833 36078 30972 36080
rect 30833 36075 30899 36078
rect 30966 36076 30972 36078
rect 31036 36076 31042 36140
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 4870 34848 5186 34849
rect 0 34778 800 34808
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 933 34778 999 34781
rect 0 34776 999 34778
rect 0 34720 938 34776
rect 994 34720 999 34776
rect 0 34718 999 34720
rect 0 34688 800 34718
rect 933 34715 999 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 36353 33418 36419 33421
rect 37136 33418 37936 33448
rect 36353 33416 37936 33418
rect 36353 33360 36358 33416
rect 36414 33360 37936 33416
rect 36353 33358 37936 33360
rect 36353 33355 36419 33358
rect 37136 33328 37936 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 14181 33146 14247 33149
rect 20989 33146 21055 33149
rect 21357 33146 21423 33149
rect 14181 33144 21423 33146
rect 14181 33088 14186 33144
rect 14242 33088 20994 33144
rect 21050 33088 21362 33144
rect 21418 33088 21423 33144
rect 14181 33086 21423 33088
rect 14181 33083 14247 33086
rect 20989 33083 21055 33086
rect 21357 33083 21423 33086
rect 19977 33010 20043 33013
rect 24301 33010 24367 33013
rect 19977 33008 24367 33010
rect 19977 32952 19982 33008
rect 20038 32952 24306 33008
rect 24362 32952 24367 33008
rect 19977 32950 24367 32952
rect 19977 32947 20043 32950
rect 24301 32947 24367 32950
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 6913 32330 6979 32333
rect 9673 32330 9739 32333
rect 6913 32328 9739 32330
rect 6913 32272 6918 32328
rect 6974 32272 9678 32328
rect 9734 32272 9739 32328
rect 6913 32270 9739 32272
rect 6913 32267 6979 32270
rect 9673 32267 9739 32270
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 933 32058 999 32061
rect 0 32056 999 32058
rect 0 32000 938 32056
rect 994 32000 999 32056
rect 0 31998 999 32000
rect 0 31968 800 31998
rect 933 31995 999 31998
rect 13813 31922 13879 31925
rect 14733 31922 14799 31925
rect 17769 31922 17835 31925
rect 25221 31922 25287 31925
rect 13813 31920 25287 31922
rect 13813 31864 13818 31920
rect 13874 31864 14738 31920
rect 14794 31864 17774 31920
rect 17830 31864 25226 31920
rect 25282 31864 25287 31920
rect 13813 31862 25287 31864
rect 13813 31859 13879 31862
rect 14733 31859 14799 31862
rect 17769 31859 17835 31862
rect 25221 31859 25287 31862
rect 8109 31786 8175 31789
rect 15285 31786 15351 31789
rect 18229 31786 18295 31789
rect 8109 31784 18295 31786
rect 8109 31728 8114 31784
rect 8170 31728 15290 31784
rect 15346 31728 18234 31784
rect 18290 31728 18295 31784
rect 8109 31726 18295 31728
rect 8109 31723 8175 31726
rect 15285 31723 15351 31726
rect 18229 31723 18295 31726
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 7097 30426 7163 30429
rect 7230 30426 7236 30428
rect 7097 30424 7236 30426
rect 7097 30368 7102 30424
rect 7158 30368 7236 30424
rect 7097 30366 7236 30368
rect 7097 30363 7163 30366
rect 7230 30364 7236 30366
rect 7300 30364 7306 30428
rect 36353 30018 36419 30021
rect 37136 30018 37936 30048
rect 36353 30016 37936 30018
rect 36353 29960 36358 30016
rect 36414 29960 37936 30016
rect 36353 29958 37936 29960
rect 36353 29955 36419 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 37136 29928 37936 29958
rect 34930 29887 35246 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 0 28658 800 28688
rect 1577 28658 1643 28661
rect 0 28656 1643 28658
rect 0 28600 1582 28656
rect 1638 28600 1643 28656
rect 0 28598 1643 28600
rect 0 28568 800 28598
rect 1577 28595 1643 28598
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 20345 27978 20411 27981
rect 24945 27978 25011 27981
rect 20345 27976 25011 27978
rect 20345 27920 20350 27976
rect 20406 27920 24950 27976
rect 25006 27920 25011 27976
rect 20345 27918 25011 27920
rect 20345 27915 20411 27918
rect 24945 27915 25011 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 23565 27570 23631 27573
rect 26877 27570 26943 27573
rect 23565 27568 26943 27570
rect 23565 27512 23570 27568
rect 23626 27512 26882 27568
rect 26938 27512 26943 27568
rect 23565 27510 26943 27512
rect 23565 27507 23631 27510
rect 26877 27507 26943 27510
rect 36353 27298 36419 27301
rect 37136 27298 37936 27328
rect 36353 27296 37936 27298
rect 36353 27240 36358 27296
rect 36414 27240 37936 27296
rect 36353 27238 37936 27240
rect 36353 27235 36419 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 37136 27208 37936 27238
rect 35590 27167 35906 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 14917 25802 14983 25805
rect 18321 25802 18387 25805
rect 14917 25800 18387 25802
rect 14917 25744 14922 25800
rect 14978 25744 18326 25800
rect 18382 25744 18387 25800
rect 14917 25742 18387 25744
rect 14917 25739 14983 25742
rect 18321 25739 18387 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 17677 25530 17743 25533
rect 22461 25530 22527 25533
rect 17677 25528 22527 25530
rect 17677 25472 17682 25528
rect 17738 25472 22466 25528
rect 22522 25472 22527 25528
rect 17677 25470 22527 25472
rect 17677 25467 17743 25470
rect 22461 25467 22527 25470
rect 0 25258 800 25288
rect 1393 25258 1459 25261
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25168 800 25198
rect 1393 25195 1459 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 25313 24306 25379 24309
rect 26233 24306 26299 24309
rect 25313 24304 26299 24306
rect 25313 24248 25318 24304
rect 25374 24248 26238 24304
rect 26294 24248 26299 24304
rect 25313 24246 26299 24248
rect 25313 24243 25379 24246
rect 26233 24243 26299 24246
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 36353 23898 36419 23901
rect 37136 23898 37936 23928
rect 36353 23896 37936 23898
rect 36353 23840 36358 23896
rect 36414 23840 37936 23896
rect 36353 23838 37936 23840
rect 36353 23835 36419 23838
rect 37136 23808 37936 23838
rect 8385 23762 8451 23765
rect 9121 23762 9187 23765
rect 8385 23760 9187 23762
rect 8385 23704 8390 23760
rect 8446 23704 9126 23760
rect 9182 23704 9187 23760
rect 8385 23702 9187 23704
rect 8385 23699 8451 23702
rect 9121 23699 9187 23702
rect 11605 23762 11671 23765
rect 23657 23762 23723 23765
rect 11605 23760 23723 23762
rect 11605 23704 11610 23760
rect 11666 23704 23662 23760
rect 23718 23704 23723 23760
rect 11605 23702 23723 23704
rect 11605 23699 11671 23702
rect 23657 23699 23723 23702
rect 25313 23626 25379 23629
rect 27613 23626 27679 23629
rect 25313 23624 27679 23626
rect 25313 23568 25318 23624
rect 25374 23568 27618 23624
rect 27674 23568 27679 23624
rect 25313 23566 27679 23568
rect 25313 23563 25379 23566
rect 27613 23563 27679 23566
rect 23381 23490 23447 23493
rect 28809 23490 28875 23493
rect 23381 23488 28875 23490
rect 23381 23432 23386 23488
rect 23442 23432 28814 23488
rect 28870 23432 28875 23488
rect 23381 23430 28875 23432
rect 23381 23427 23447 23430
rect 28809 23427 28875 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 0 22538 800 22568
rect 933 22538 999 22541
rect 0 22536 999 22538
rect 0 22480 938 22536
rect 994 22480 999 22536
rect 0 22478 999 22480
rect 0 22448 800 22478
rect 933 22475 999 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 13721 22266 13787 22269
rect 17585 22266 17651 22269
rect 13721 22264 17651 22266
rect 13721 22208 13726 22264
rect 13782 22208 17590 22264
rect 17646 22208 17651 22264
rect 13721 22206 17651 22208
rect 13721 22203 13787 22206
rect 17585 22203 17651 22206
rect 17217 22130 17283 22133
rect 17174 22128 17283 22130
rect 17174 22072 17222 22128
rect 17278 22072 17283 22128
rect 17174 22067 17283 22072
rect 7189 21860 7255 21861
rect 7189 21856 7236 21860
rect 7300 21858 7306 21860
rect 16849 21858 16915 21861
rect 17174 21858 17234 22067
rect 7189 21800 7194 21856
rect 7189 21796 7236 21800
rect 7300 21798 7346 21858
rect 16849 21856 17234 21858
rect 16849 21800 16854 21856
rect 16910 21800 17234 21856
rect 16849 21798 17234 21800
rect 7300 21796 7306 21798
rect 7189 21795 7255 21796
rect 16849 21795 16915 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 13169 21722 13235 21725
rect 16941 21722 17007 21725
rect 19977 21722 20043 21725
rect 13169 21720 20043 21722
rect 13169 21664 13174 21720
rect 13230 21664 16946 21720
rect 17002 21664 19982 21720
rect 20038 21664 20043 21720
rect 13169 21662 20043 21664
rect 13169 21659 13235 21662
rect 16941 21659 17007 21662
rect 19977 21659 20043 21662
rect 19333 21450 19399 21453
rect 20989 21450 21055 21453
rect 19333 21448 21055 21450
rect 19333 21392 19338 21448
rect 19394 21392 20994 21448
rect 21050 21392 21055 21448
rect 19333 21390 21055 21392
rect 19333 21387 19399 21390
rect 20989 21387 21055 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 16113 21178 16179 21181
rect 17585 21178 17651 21181
rect 16113 21176 17651 21178
rect 16113 21120 16118 21176
rect 16174 21120 17590 21176
rect 17646 21120 17651 21176
rect 16113 21118 17651 21120
rect 16113 21115 16179 21118
rect 17585 21115 17651 21118
rect 16021 21042 16087 21045
rect 16757 21042 16823 21045
rect 16941 21042 17007 21045
rect 16021 21040 17007 21042
rect 16021 20984 16026 21040
rect 16082 20984 16762 21040
rect 16818 20984 16946 21040
rect 17002 20984 17007 21040
rect 16021 20982 17007 20984
rect 16021 20979 16087 20982
rect 16757 20979 16823 20982
rect 16941 20979 17007 20982
rect 19701 21042 19767 21045
rect 25957 21042 26023 21045
rect 19701 21040 26023 21042
rect 19701 20984 19706 21040
rect 19762 20984 25962 21040
rect 26018 20984 26023 21040
rect 19701 20982 26023 20984
rect 19701 20979 19767 20982
rect 25957 20979 26023 20982
rect 13721 20906 13787 20909
rect 17861 20906 17927 20909
rect 13721 20904 17927 20906
rect 13721 20848 13726 20904
rect 13782 20848 17866 20904
rect 17922 20848 17927 20904
rect 13721 20846 17927 20848
rect 13721 20843 13787 20846
rect 17861 20843 17927 20846
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 30833 20634 30899 20637
rect 30966 20634 30972 20636
rect 30833 20632 30972 20634
rect 30833 20576 30838 20632
rect 30894 20576 30972 20632
rect 30833 20574 30972 20576
rect 30833 20571 30899 20574
rect 30966 20572 30972 20574
rect 31036 20572 31042 20636
rect 17401 20498 17467 20501
rect 18413 20498 18479 20501
rect 17401 20496 18479 20498
rect 17401 20440 17406 20496
rect 17462 20440 18418 20496
rect 18474 20440 18479 20496
rect 17401 20438 18479 20440
rect 17401 20435 17467 20438
rect 18413 20435 18479 20438
rect 24301 20498 24367 20501
rect 26785 20498 26851 20501
rect 24301 20496 26851 20498
rect 24301 20440 24306 20496
rect 24362 20440 26790 20496
rect 26846 20440 26851 20496
rect 24301 20438 26851 20440
rect 24301 20435 24367 20438
rect 26785 20435 26851 20438
rect 36353 20498 36419 20501
rect 37136 20498 37936 20528
rect 36353 20496 37936 20498
rect 36353 20440 36358 20496
rect 36414 20440 37936 20496
rect 36353 20438 37936 20440
rect 36353 20435 36419 20438
rect 37136 20408 37936 20438
rect 17125 20362 17191 20365
rect 17861 20362 17927 20365
rect 17125 20360 17927 20362
rect 17125 20304 17130 20360
rect 17186 20304 17866 20360
rect 17922 20304 17927 20360
rect 17125 20302 17927 20304
rect 17125 20299 17191 20302
rect 17861 20299 17927 20302
rect 20989 20362 21055 20365
rect 22277 20362 22343 20365
rect 20989 20360 22343 20362
rect 20989 20304 20994 20360
rect 21050 20304 22282 20360
rect 22338 20304 22343 20360
rect 20989 20302 22343 20304
rect 20989 20299 21055 20302
rect 22277 20299 22343 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 20253 19410 20319 19413
rect 20805 19410 20871 19413
rect 25865 19410 25931 19413
rect 20253 19408 20362 19410
rect 20253 19352 20258 19408
rect 20314 19352 20362 19408
rect 20253 19347 20362 19352
rect 20805 19408 25931 19410
rect 20805 19352 20810 19408
rect 20866 19352 25870 19408
rect 25926 19352 25931 19408
rect 20805 19350 25931 19352
rect 20805 19347 20871 19350
rect 25865 19347 25931 19350
rect 7005 19274 7071 19277
rect 10225 19274 10291 19277
rect 13445 19274 13511 19277
rect 20302 19274 20362 19347
rect 7005 19272 20362 19274
rect 7005 19216 7010 19272
rect 7066 19216 10230 19272
rect 10286 19216 13450 19272
rect 13506 19216 20362 19272
rect 7005 19214 20362 19216
rect 7005 19211 7071 19214
rect 10225 19211 10291 19214
rect 13445 19211 13511 19214
rect 0 19138 800 19168
rect 933 19138 999 19141
rect 0 19136 999 19138
rect 0 19080 938 19136
rect 994 19080 999 19136
rect 0 19078 999 19080
rect 20302 19138 20362 19214
rect 20529 19274 20595 19277
rect 21081 19274 21147 19277
rect 26049 19274 26115 19277
rect 20529 19272 26115 19274
rect 20529 19216 20534 19272
rect 20590 19216 21086 19272
rect 21142 19216 26054 19272
rect 26110 19216 26115 19272
rect 20529 19214 26115 19216
rect 20529 19211 20595 19214
rect 21081 19211 21147 19214
rect 26049 19211 26115 19214
rect 27061 19274 27127 19277
rect 28349 19274 28415 19277
rect 27061 19272 28415 19274
rect 27061 19216 27066 19272
rect 27122 19216 28354 19272
rect 28410 19216 28415 19272
rect 27061 19214 28415 19216
rect 27061 19211 27127 19214
rect 28349 19211 28415 19214
rect 26417 19138 26483 19141
rect 20302 19136 26483 19138
rect 20302 19080 26422 19136
rect 26478 19080 26483 19136
rect 20302 19078 26483 19080
rect 0 19048 800 19078
rect 933 19075 999 19078
rect 26417 19075 26483 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 14273 19002 14339 19005
rect 20529 19002 20595 19005
rect 14273 19000 20595 19002
rect 14273 18944 14278 19000
rect 14334 18944 20534 19000
rect 20590 18944 20595 19000
rect 14273 18942 20595 18944
rect 14273 18939 14339 18942
rect 20529 18939 20595 18942
rect 23105 19002 23171 19005
rect 28533 19002 28599 19005
rect 23105 19000 28599 19002
rect 23105 18944 23110 19000
rect 23166 18944 28538 19000
rect 28594 18944 28599 19000
rect 23105 18942 28599 18944
rect 23105 18939 23171 18942
rect 28533 18939 28599 18942
rect 17033 18866 17099 18869
rect 25037 18866 25103 18869
rect 26141 18866 26207 18869
rect 17033 18864 26207 18866
rect 17033 18808 17038 18864
rect 17094 18808 25042 18864
rect 25098 18808 26146 18864
rect 26202 18808 26207 18864
rect 17033 18806 26207 18808
rect 17033 18803 17099 18806
rect 25037 18803 25103 18806
rect 26141 18803 26207 18806
rect 25865 18730 25931 18733
rect 28441 18730 28507 18733
rect 25865 18728 28507 18730
rect 25865 18672 25870 18728
rect 25926 18672 28446 18728
rect 28502 18672 28507 18728
rect 25865 18670 28507 18672
rect 25865 18667 25931 18670
rect 28441 18667 28507 18670
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 26969 18458 27035 18461
rect 28533 18458 28599 18461
rect 26969 18456 28599 18458
rect 26969 18400 26974 18456
rect 27030 18400 28538 18456
rect 28594 18400 28599 18456
rect 26969 18398 28599 18400
rect 26969 18395 27035 18398
rect 28533 18395 28599 18398
rect 5349 18322 5415 18325
rect 5533 18322 5599 18325
rect 5349 18320 5599 18322
rect 5349 18264 5354 18320
rect 5410 18264 5538 18320
rect 5594 18264 5599 18320
rect 5349 18262 5599 18264
rect 5349 18259 5415 18262
rect 5533 18259 5599 18262
rect 8845 18322 8911 18325
rect 10685 18322 10751 18325
rect 11697 18322 11763 18325
rect 8845 18320 11763 18322
rect 8845 18264 8850 18320
rect 8906 18264 10690 18320
rect 10746 18264 11702 18320
rect 11758 18264 11763 18320
rect 8845 18262 11763 18264
rect 8845 18259 8911 18262
rect 10685 18259 10751 18262
rect 11697 18259 11763 18262
rect 14457 18322 14523 18325
rect 17861 18322 17927 18325
rect 14457 18320 17927 18322
rect 14457 18264 14462 18320
rect 14518 18264 17866 18320
rect 17922 18264 17927 18320
rect 14457 18262 17927 18264
rect 14457 18259 14523 18262
rect 17861 18259 17927 18262
rect 19425 18322 19491 18325
rect 20805 18322 20871 18325
rect 19425 18320 20871 18322
rect 19425 18264 19430 18320
rect 19486 18264 20810 18320
rect 20866 18264 20871 18320
rect 19425 18262 20871 18264
rect 19425 18259 19491 18262
rect 20805 18259 20871 18262
rect 6637 18186 6703 18189
rect 7557 18186 7623 18189
rect 10133 18186 10199 18189
rect 23657 18186 23723 18189
rect 6637 18184 23723 18186
rect 6637 18128 6642 18184
rect 6698 18128 7562 18184
rect 7618 18128 10138 18184
rect 10194 18128 23662 18184
rect 23718 18128 23723 18184
rect 6637 18126 23723 18128
rect 6637 18123 6703 18126
rect 7557 18123 7623 18126
rect 10133 18123 10199 18126
rect 23657 18123 23723 18126
rect 13629 18050 13695 18053
rect 14549 18050 14615 18053
rect 13629 18048 14615 18050
rect 13629 17992 13634 18048
rect 13690 17992 14554 18048
rect 14610 17992 14615 18048
rect 13629 17990 14615 17992
rect 13629 17987 13695 17990
rect 14549 17987 14615 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 36445 17098 36511 17101
rect 37136 17098 37936 17128
rect 36445 17096 37936 17098
rect 36445 17040 36450 17096
rect 36506 17040 37936 17096
rect 36445 17038 37936 17040
rect 36445 17035 36511 17038
rect 37136 17008 37936 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 933 15738 999 15741
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 36353 14378 36419 14381
rect 37136 14378 37936 14408
rect 36353 14376 37936 14378
rect 36353 14320 36358 14376
rect 36414 14320 37936 14376
rect 36353 14318 37936 14320
rect 36353 14315 36419 14318
rect 37136 14288 37936 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 13169 13970 13235 13973
rect 14181 13970 14247 13973
rect 13169 13968 14247 13970
rect 13169 13912 13174 13968
rect 13230 13912 14186 13968
rect 14242 13912 14247 13968
rect 13169 13910 14247 13912
rect 13169 13907 13235 13910
rect 14181 13907 14247 13910
rect 11513 13834 11579 13837
rect 13261 13834 13327 13837
rect 11513 13832 13327 13834
rect 11513 13776 11518 13832
rect 11574 13776 13266 13832
rect 13322 13776 13327 13832
rect 11513 13774 13327 13776
rect 11513 13771 11579 13774
rect 13261 13771 13327 13774
rect 25497 13834 25563 13837
rect 25630 13834 25636 13836
rect 25497 13832 25636 13834
rect 25497 13776 25502 13832
rect 25558 13776 25636 13832
rect 25497 13774 25636 13776
rect 25497 13771 25563 13774
rect 25630 13772 25636 13774
rect 25700 13772 25706 13836
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 25405 13154 25471 13157
rect 26141 13154 26207 13157
rect 25405 13152 26207 13154
rect 25405 13096 25410 13152
rect 25466 13096 26146 13152
rect 26202 13096 26207 13152
rect 25405 13094 26207 13096
rect 25405 13091 25471 13094
rect 26141 13091 26207 13094
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12338 800 12368
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 800 12278
rect 1577 12275 1643 12278
rect 11789 12338 11855 12341
rect 13997 12338 14063 12341
rect 11789 12336 14063 12338
rect 11789 12280 11794 12336
rect 11850 12280 14002 12336
rect 14058 12280 14063 12336
rect 11789 12278 14063 12280
rect 11789 12275 11855 12278
rect 13997 12275 14063 12278
rect 21081 12338 21147 12341
rect 22001 12338 22067 12341
rect 21081 12336 22067 12338
rect 21081 12280 21086 12336
rect 21142 12280 22006 12336
rect 22062 12280 22067 12336
rect 21081 12278 22067 12280
rect 21081 12275 21147 12278
rect 22001 12275 22067 12278
rect 1761 12202 1827 12205
rect 19885 12202 19951 12205
rect 1761 12200 19951 12202
rect 1761 12144 1766 12200
rect 1822 12144 19890 12200
rect 19946 12144 19951 12200
rect 1761 12142 19951 12144
rect 1761 12139 1827 12142
rect 19885 12139 19951 12142
rect 31109 12202 31175 12205
rect 32121 12202 32187 12205
rect 31109 12200 32187 12202
rect 31109 12144 31114 12200
rect 31170 12144 32126 12200
rect 32182 12144 32187 12200
rect 31109 12142 32187 12144
rect 31109 12139 31175 12142
rect 32121 12139 32187 12142
rect 5717 12066 5783 12069
rect 8385 12066 8451 12069
rect 5717 12064 8451 12066
rect 5717 12008 5722 12064
rect 5778 12008 8390 12064
rect 8446 12008 8451 12064
rect 5717 12006 8451 12008
rect 5717 12003 5783 12006
rect 8385 12003 8451 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 11697 11930 11763 11933
rect 19241 11930 19307 11933
rect 11697 11928 19307 11930
rect 11697 11872 11702 11928
rect 11758 11872 19246 11928
rect 19302 11872 19307 11928
rect 11697 11870 19307 11872
rect 11697 11867 11763 11870
rect 19241 11867 19307 11870
rect 4153 11794 4219 11797
rect 20897 11794 20963 11797
rect 4153 11792 20963 11794
rect 4153 11736 4158 11792
rect 4214 11736 20902 11792
rect 20958 11736 20963 11792
rect 4153 11734 20963 11736
rect 4153 11731 4219 11734
rect 20897 11731 20963 11734
rect 22277 11794 22343 11797
rect 24117 11794 24183 11797
rect 22277 11792 24183 11794
rect 22277 11736 22282 11792
rect 22338 11736 24122 11792
rect 24178 11736 24183 11792
rect 22277 11734 24183 11736
rect 22277 11731 22343 11734
rect 24117 11731 24183 11734
rect 33133 11658 33199 11661
rect 33501 11660 33567 11661
rect 33501 11658 33548 11660
rect 33133 11656 33548 11658
rect 33133 11600 33138 11656
rect 33194 11600 33506 11656
rect 33133 11598 33548 11600
rect 33133 11595 33199 11598
rect 33501 11596 33548 11598
rect 33612 11596 33618 11660
rect 33501 11595 33567 11596
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 18781 11250 18847 11253
rect 28717 11250 28783 11253
rect 18781 11248 28783 11250
rect 18781 11192 18786 11248
rect 18842 11192 28722 11248
rect 28778 11192 28783 11248
rect 18781 11190 28783 11192
rect 18781 11187 18847 11190
rect 28717 11187 28783 11190
rect 20253 11116 20319 11117
rect 20253 11112 20300 11116
rect 20364 11114 20370 11116
rect 20253 11056 20258 11112
rect 20253 11052 20300 11056
rect 20364 11054 20410 11114
rect 20364 11052 20370 11054
rect 20253 11051 20319 11052
rect 36445 10978 36511 10981
rect 37136 10978 37936 11008
rect 36445 10976 37936 10978
rect 36445 10920 36450 10976
rect 36506 10920 37936 10976
rect 36445 10918 37936 10920
rect 36445 10915 36511 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 37136 10888 37936 10918
rect 35590 10847 35906 10848
rect 10317 10706 10383 10709
rect 19057 10706 19123 10709
rect 10317 10704 19123 10706
rect 10317 10648 10322 10704
rect 10378 10648 19062 10704
rect 19118 10648 19123 10704
rect 10317 10646 19123 10648
rect 10317 10643 10383 10646
rect 19057 10643 19123 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 21265 10162 21331 10165
rect 24761 10162 24827 10165
rect 21265 10160 24827 10162
rect 21265 10104 21270 10160
rect 21326 10104 24766 10160
rect 24822 10104 24827 10160
rect 21265 10102 24827 10104
rect 21265 10099 21331 10102
rect 24761 10099 24827 10102
rect 19977 9890 20043 9893
rect 21725 9890 21791 9893
rect 19977 9888 21791 9890
rect 19977 9832 19982 9888
rect 20038 9832 21730 9888
rect 21786 9832 21791 9888
rect 19977 9830 21791 9832
rect 19977 9827 20043 9830
rect 21725 9827 21791 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 21541 9754 21607 9757
rect 24393 9754 24459 9757
rect 21541 9752 24459 9754
rect 21541 9696 21546 9752
rect 21602 9696 24398 9752
rect 24454 9696 24459 9752
rect 21541 9694 24459 9696
rect 21541 9691 21607 9694
rect 24393 9691 24459 9694
rect 0 9618 800 9648
rect 1577 9618 1643 9621
rect 0 9616 1643 9618
rect 0 9560 1582 9616
rect 1638 9560 1643 9616
rect 0 9558 1643 9560
rect 0 9528 800 9558
rect 1577 9555 1643 9558
rect 10501 9618 10567 9621
rect 16205 9618 16271 9621
rect 10501 9616 16271 9618
rect 10501 9560 10506 9616
rect 10562 9560 16210 9616
rect 16266 9560 16271 9616
rect 10501 9558 16271 9560
rect 10501 9555 10567 9558
rect 16205 9555 16271 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 11605 8938 11671 8941
rect 12893 8938 12959 8941
rect 11605 8936 12959 8938
rect 11605 8880 11610 8936
rect 11666 8880 12898 8936
rect 12954 8880 12959 8936
rect 11605 8878 12959 8880
rect 11605 8875 11671 8878
rect 12893 8875 12959 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 12617 8530 12683 8533
rect 16481 8530 16547 8533
rect 12617 8528 16547 8530
rect 12617 8472 12622 8528
rect 12678 8472 16486 8528
rect 16542 8472 16547 8528
rect 12617 8470 16547 8472
rect 12617 8467 12683 8470
rect 16481 8467 16547 8470
rect 33593 8260 33659 8261
rect 33542 8258 33548 8260
rect 33502 8198 33548 8258
rect 33612 8256 33659 8260
rect 33654 8200 33659 8256
rect 33542 8196 33548 8198
rect 33612 8196 33659 8200
rect 33593 8195 33659 8196
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19793 7850 19859 7853
rect 36261 7850 36327 7853
rect 19793 7848 36327 7850
rect 19793 7792 19798 7848
rect 19854 7792 36266 7848
rect 36322 7792 36327 7848
rect 19793 7790 36327 7792
rect 19793 7787 19859 7790
rect 36261 7787 36327 7790
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 36445 7578 36511 7581
rect 37136 7578 37936 7608
rect 36445 7576 37936 7578
rect 36445 7520 36450 7576
rect 36506 7520 37936 7576
rect 36445 7518 37936 7520
rect 36445 7515 36511 7518
rect 37136 7488 37936 7518
rect 30741 7306 30807 7309
rect 33869 7306 33935 7309
rect 30741 7304 33935 7306
rect 30741 7248 30746 7304
rect 30802 7248 33874 7304
rect 33930 7248 33935 7304
rect 30741 7246 33935 7248
rect 30741 7243 30807 7246
rect 33869 7243 33935 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 0 6218 800 6248
rect 1301 6218 1367 6221
rect 0 6216 1367 6218
rect 0 6160 1306 6216
rect 1362 6160 1367 6216
rect 0 6158 1367 6160
rect 0 6128 800 6158
rect 1301 6155 1367 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 6085 5810 6151 5813
rect 9213 5810 9279 5813
rect 6085 5808 9279 5810
rect 6085 5752 6090 5808
rect 6146 5752 9218 5808
rect 9274 5752 9279 5808
rect 6085 5750 9279 5752
rect 6085 5747 6151 5750
rect 9213 5747 9279 5750
rect 29453 5674 29519 5677
rect 32213 5674 32279 5677
rect 29453 5672 32279 5674
rect 29453 5616 29458 5672
rect 29514 5616 32218 5672
rect 32274 5616 32279 5672
rect 29453 5614 32279 5616
rect 29453 5611 29519 5614
rect 32213 5611 32279 5614
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 36353 4858 36419 4861
rect 37136 4858 37936 4888
rect 36353 4856 37936 4858
rect 36353 4800 36358 4856
rect 36414 4800 37936 4856
rect 36353 4798 37936 4800
rect 36353 4795 36419 4798
rect 37136 4768 37936 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 17493 3498 17559 3501
rect 18045 3498 18111 3501
rect 17493 3496 18111 3498
rect 17493 3440 17498 3496
rect 17554 3440 18050 3496
rect 18106 3440 18111 3496
rect 17493 3438 18111 3440
rect 17493 3435 17559 3438
rect 18045 3435 18111 3438
rect 30833 3498 30899 3501
rect 31845 3498 31911 3501
rect 30833 3496 31911 3498
rect 30833 3440 30838 3496
rect 30894 3440 31850 3496
rect 31906 3440 31911 3496
rect 30833 3438 31911 3440
rect 30833 3435 30899 3438
rect 31845 3435 31911 3438
rect 29821 3362 29887 3365
rect 31293 3362 31359 3365
rect 29821 3360 31359 3362
rect 29821 3304 29826 3360
rect 29882 3304 31298 3360
rect 31354 3304 31359 3360
rect 29821 3302 31359 3304
rect 29821 3299 29887 3302
rect 31293 3299 31359 3302
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4245 2954 4311 2957
rect 23933 2954 23999 2957
rect 4245 2952 23999 2954
rect 4245 2896 4250 2952
rect 4306 2896 23938 2952
rect 23994 2896 23999 2952
rect 4245 2894 23999 2896
rect 4245 2891 4311 2894
rect 23933 2891 23999 2894
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 20294 2484 20300 2548
rect 20364 2546 20370 2548
rect 35893 2546 35959 2549
rect 20364 2544 35959 2546
rect 20364 2488 35898 2544
rect 35954 2488 35959 2544
rect 20364 2486 35959 2488
rect 20364 2484 20370 2486
rect 35893 2483 35959 2486
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 35433 1458 35499 1461
rect 37136 1458 37936 1488
rect 35433 1456 37936 1458
rect 35433 1400 35438 1456
rect 35494 1400 37936 1456
rect 35433 1398 37936 1400
rect 35433 1395 35499 1398
rect 37136 1368 37936 1398
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 25636 36484 25700 36548
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 30972 36076 31036 36140
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 7236 30364 7300 30428
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 7236 21856 7300 21860
rect 7236 21800 7250 21856
rect 7250 21800 7300 21856
rect 7236 21796 7300 21800
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 30972 20572 31036 20636
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 25636 13772 25700 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 33548 11656 33612 11660
rect 33548 11600 33562 11656
rect 33562 11600 33612 11656
rect 33548 11596 33612 11600
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 20300 11112 20364 11116
rect 20300 11056 20314 11112
rect 20314 11056 20364 11112
rect 20300 11052 20364 11056
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 33548 8256 33612 8260
rect 33548 8200 33598 8256
rect 33598 8200 33612 8256
rect 33548 8196 33612 8200
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 20300 2484 20364 2548
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 37024 5188 37584
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 25635 36548 25701 36549
rect 25635 36484 25636 36548
rect 25700 36484 25701 36548
rect 25635 36483 25701 36484
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 7235 30428 7301 30429
rect 7235 30364 7236 30428
rect 7300 30364 7301 30428
rect 7235 30363 7301 30364
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 7238 21861 7298 30363
rect 7235 21860 7301 21861
rect 7235 21796 7236 21860
rect 7300 21796 7301 21860
rect 7235 21795 7301 21796
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 25638 13837 25698 36483
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36260 35248 36416
rect 30971 36140 31037 36141
rect 30971 36076 30972 36140
rect 31036 36076 31037 36140
rect 30971 36075 31037 36076
rect 30974 20637 31034 36075
rect 34928 36024 34970 36260
rect 35206 36024 35248 36260
rect 34928 35392 35248 36024
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 30971 20636 31037 20637
rect 30971 20572 30972 20636
rect 31036 20572 31037 20636
rect 30971 20571 31037 20572
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 25635 13836 25701 13837
rect 25635 13772 25636 13836
rect 25700 13772 25701 13836
rect 25635 13771 25701 13772
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 33547 11660 33613 11661
rect 33547 11596 33548 11660
rect 33612 11596 33613 11660
rect 33547 11595 33613 11596
rect 20299 11116 20365 11117
rect 20299 11052 20300 11116
rect 20364 11052 20365 11116
rect 20299 11051 20365 11052
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 20302 2549 20362 11051
rect 33550 8261 33610 11595
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 33547 8260 33613 8261
rect 33547 8196 33548 8260
rect 33612 8196 33613 8260
rect 33547 8195 33613 8196
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 20299 2548 20365 2549
rect 20299 2484 20300 2548
rect 20364 2484 20365 2548
rect 20299 2483 20365 2484
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 2128 35248 2688
rect 35588 37024 35908 37584
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 36920 35908 36960
rect 35588 36684 35630 36920
rect 35866 36684 35908 36920
rect 35588 35936 35908 36684
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
<< via4 >>
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 36684 5146 36920
rect 34970 36024 35206 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 36684 35866 36920
rect 35630 6048 35866 6284
<< metal5 >>
rect 1056 36920 36848 36962
rect 1056 36684 4910 36920
rect 5146 36684 35630 36920
rect 35866 36684 36848 36920
rect 1056 36642 36848 36684
rect 1056 36260 36848 36302
rect 1056 36024 4250 36260
rect 4486 36024 34970 36260
rect 35206 36024 36848 36260
rect 1056 35982 36848 36024
rect 1056 6284 36848 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 36848 6284
rect 1056 6006 36848 6048
rect 1056 5624 36848 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 36848 5624
rect 1056 5346 36848 5388
use sky130_fd_sc_hd__dlymetal6s2s_1  _0889_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14076 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0890_
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0891_
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0892_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0893_
timestamp 1679235063
transform 1 0 12144 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0894_
timestamp 1679235063
transform 1 0 12328 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0895_
timestamp 1679235063
transform 1 0 11500 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _0896_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9936 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0897_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0898_
timestamp 1679235063
transform 1 0 10028 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0899_
timestamp 1679235063
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0900_
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1679235063
transform 1 0 12512 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0902_
timestamp 1679235063
transform 1 0 10948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0903_
timestamp 1679235063
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0904_
timestamp 1679235063
transform 1 0 9936 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0905_
timestamp 1679235063
transform 1 0 10028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0906_
timestamp 1679235063
transform 1 0 10948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0907_
timestamp 1679235063
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0908_
timestamp 1679235063
transform 1 0 12880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0909_
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0910_
timestamp 1679235063
transform 1 0 14352 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 1679235063
transform 1 0 15088 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0912_
timestamp 1679235063
transform 1 0 17572 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17020 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0914_
timestamp 1679235063
transform 1 0 22448 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0915_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0916_
timestamp 1679235063
transform 1 0 17296 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0917_
timestamp 1679235063
transform 1 0 17204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0918_
timestamp 1679235063
transform 1 0 16652 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_2  _0919_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0920_
timestamp 1679235063
transform 1 0 17940 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor4b_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15916 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0922_
timestamp 1679235063
transform 1 0 20424 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_1  _0923_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19780 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0924_
timestamp 1679235063
transform 1 0 19872 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0925_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 21988 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _0926_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18308 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17204 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_1  _0928_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16284 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0929_
timestamp 1679235063
transform 1 0 9200 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0930_
timestamp 1679235063
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0931_
timestamp 1679235063
transform 1 0 10212 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_1  _0932_
timestamp 1679235063
transform 1 0 11684 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0933_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _0934_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18124 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_1  _0935_
timestamp 1679235063
transform 1 0 18492 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0936_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0937_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0938_
timestamp 1679235063
transform 1 0 21068 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0939_
timestamp 1679235063
transform 1 0 23736 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0940_
timestamp 1679235063
transform 1 0 19136 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_2  _0941_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0943_
timestamp 1679235063
transform 1 0 20976 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _0944_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20700 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0945_
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0946_
timestamp 1679235063
transform 1 0 22908 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0947_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 21436 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0948_
timestamp 1679235063
transform 1 0 21620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0949_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0950_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22448 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0951_
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0952_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13064 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0953_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14536 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1679235063
transform 1 0 14996 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0955_
timestamp 1679235063
transform 1 0 22264 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0956_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23368 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0957_
timestamp 1679235063
transform 1 0 11868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0958_
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0959_
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _0960_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 12604 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _0961_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14812 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0962_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23000 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0963_
timestamp 1679235063
transform 1 0 23184 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _0964_
timestamp 1679235063
transform 1 0 13708 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _0965_
timestamp 1679235063
transform 1 0 21896 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0966_
timestamp 1679235063
transform 1 0 22540 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0967_
timestamp 1679235063
transform 1 0 22448 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _0968_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14352 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0969_
timestamp 1679235063
transform 1 0 22172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0970_
timestamp 1679235063
transform 1 0 23000 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0971_
timestamp 1679235063
transform 1 0 22908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _0972_
timestamp 1679235063
transform 1 0 12880 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _0973_
timestamp 1679235063
transform 1 0 13616 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0974_
timestamp 1679235063
transform 1 0 14076 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _0975_
timestamp 1679235063
transform 1 0 7820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0976_
timestamp 1679235063
transform 1 0 14628 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0977_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14168 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0978_
timestamp 1679235063
transform 1 0 23736 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0979_
timestamp 1679235063
transform 1 0 24288 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _0980_
timestamp 1679235063
transform 1 0 6440 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _0981_
timestamp 1679235063
transform 1 0 8188 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _0982_
timestamp 1679235063
transform 1 0 7452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _0983_
timestamp 1679235063
transform 1 0 4324 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _0984_
timestamp 1679235063
transform 1 0 6532 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0985_
timestamp 1679235063
transform 1 0 23276 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0986_
timestamp 1679235063
transform 1 0 21804 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _0987_
timestamp 1679235063
transform 1 0 5980 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0988_
timestamp 1679235063
transform 1 0 6624 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0989_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7176 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _0990_
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _0991_
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _0992_
timestamp 1679235063
transform 1 0 17572 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0993_
timestamp 1679235063
transform 1 0 17020 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _0994_
timestamp 1679235063
transform 1 0 17848 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _0995_
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _0996_
timestamp 1679235063
transform 1 0 18124 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0997_
timestamp 1679235063
transform 1 0 16836 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _0998_
timestamp 1679235063
transform 1 0 18584 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0999_
timestamp 1679235063
transform 1 0 17388 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1000_
timestamp 1679235063
transform 1 0 5428 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1001_
timestamp 1679235063
transform 1 0 7084 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1002_
timestamp 1679235063
transform 1 0 4784 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1003_
timestamp 1679235063
transform 1 0 7084 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1004_
timestamp 1679235063
transform 1 0 4324 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1005_
timestamp 1679235063
transform 1 0 4968 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1006_
timestamp 1679235063
transform 1 0 6348 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1007_
timestamp 1679235063
transform 1 0 6348 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1008_
timestamp 1679235063
transform 1 0 26588 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1009_
timestamp 1679235063
transform 1 0 23000 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1010_
timestamp 1679235063
transform 1 0 24932 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1011_
timestamp 1679235063
transform 1 0 22908 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1012_
timestamp 1679235063
transform 1 0 26956 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1013_
timestamp 1679235063
transform 1 0 23092 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1014_
timestamp 1679235063
transform 1 0 27232 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1015_
timestamp 1679235063
transform 1 0 22724 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1016_
timestamp 1679235063
transform 1 0 23184 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1017_
timestamp 1679235063
transform 1 0 24472 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1018_
timestamp 1679235063
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1019_
timestamp 1679235063
transform 1 0 24656 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1020_
timestamp 1679235063
transform 1 0 23644 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1021_
timestamp 1679235063
transform 1 0 23000 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1022_
timestamp 1679235063
transform 1 0 23460 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1023_
timestamp 1679235063
transform 1 0 23644 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1024_
timestamp 1679235063
transform 1 0 22356 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1025_
timestamp 1679235063
transform 1 0 19780 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1026_
timestamp 1679235063
transform 1 0 21344 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1027_
timestamp 1679235063
transform 1 0 22080 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1028_
timestamp 1679235063
transform 1 0 21436 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1029_
timestamp 1679235063
transform 1 0 19596 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1030_
timestamp 1679235063
transform 1 0 20792 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1031_
timestamp 1679235063
transform 1 0 20516 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1032_
timestamp 1679235063
transform 1 0 20884 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1033_
timestamp 1679235063
transform 1 0 20884 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1034_
timestamp 1679235063
transform 1 0 10028 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1035_
timestamp 1679235063
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1036_
timestamp 1679235063
transform 1 0 9844 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1037_
timestamp 1679235063
transform 1 0 11040 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1038_
timestamp 1679235063
transform 1 0 9476 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1039_
timestamp 1679235063
transform 1 0 10212 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1040_
timestamp 1679235063
transform 1 0 10764 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1041_
timestamp 1679235063
transform 1 0 10120 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1042_
timestamp 1679235063
transform 1 0 27968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1043_
timestamp 1679235063
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1044_
timestamp 1679235063
transform 1 0 28428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1045_
timestamp 1679235063
transform 1 0 25208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1046_
timestamp 1679235063
transform 1 0 14076 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _1047_
timestamp 1679235063
transform 1 0 28888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1048_
timestamp 1679235063
transform 1 0 26036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1049_
timestamp 1679235063
transform 1 0 9660 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1050_
timestamp 1679235063
transform 1 0 14168 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1051_
timestamp 1679235063
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1052_
timestamp 1679235063
transform 1 0 19872 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1053_
timestamp 1679235063
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1054_
timestamp 1679235063
transform 1 0 12512 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1055_
timestamp 1679235063
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1056_
timestamp 1679235063
transform 1 0 9292 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1057_
timestamp 1679235063
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1058_
timestamp 1679235063
transform 1 0 25852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1059_
timestamp 1679235063
transform 1 0 12880 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_4  _1060_
timestamp 1679235063
transform 1 0 27876 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1061_
timestamp 1679235063
transform 1 0 26956 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1062_
timestamp 1679235063
transform 1 0 13340 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _1063_
timestamp 1679235063
transform 1 0 27508 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1064_
timestamp 1679235063
transform 1 0 13984 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1065_
timestamp 1679235063
transform 1 0 13340 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1066_
timestamp 1679235063
transform 1 0 6624 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1067_
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1068_
timestamp 1679235063
transform 1 0 4600 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1069_
timestamp 1679235063
transform 1 0 7360 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1070_
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1071_
timestamp 1679235063
transform 1 0 6900 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1072_
timestamp 1679235063
transform 1 0 8280 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1073_
timestamp 1679235063
transform 1 0 8004 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1074_
timestamp 1679235063
transform 1 0 17020 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1075_
timestamp 1679235063
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1076_
timestamp 1679235063
transform 1 0 16192 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1077_
timestamp 1679235063
transform 1 0 16744 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1078_
timestamp 1679235063
transform 1 0 16376 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1079_
timestamp 1679235063
transform 1 0 16928 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1080_
timestamp 1679235063
transform 1 0 17848 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1081_
timestamp 1679235063
transform 1 0 17204 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1082_
timestamp 1679235063
transform 1 0 20240 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1083_
timestamp 1679235063
transform 1 0 20792 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1084_
timestamp 1679235063
transform 1 0 5152 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1085_
timestamp 1679235063
transform 1 0 7544 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1086_
timestamp 1679235063
transform 1 0 4324 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1087_
timestamp 1679235063
transform 1 0 6348 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1088_
timestamp 1679235063
transform 1 0 5244 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _1089_
timestamp 1679235063
transform 1 0 19504 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1090_
timestamp 1679235063
transform 1 0 6808 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1091_
timestamp 1679235063
transform 1 0 4876 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1092_
timestamp 1679235063
transform 1 0 6624 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1093_
timestamp 1679235063
transform 1 0 6716 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1094_
timestamp 1679235063
transform 1 0 25116 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1095_
timestamp 1679235063
transform 1 0 26036 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1096_
timestamp 1679235063
transform 1 0 26956 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1097_
timestamp 1679235063
transform 1 0 27416 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1098_
timestamp 1679235063
transform 1 0 27324 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1099_
timestamp 1679235063
transform 1 0 27416 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1100_
timestamp 1679235063
transform 1 0 28060 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1101_
timestamp 1679235063
transform 1 0 26772 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1102_
timestamp 1679235063
transform 1 0 24564 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1103_
timestamp 1679235063
transform 1 0 25300 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1104_
timestamp 1679235063
transform 1 0 24656 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1105_
timestamp 1679235063
transform 1 0 24748 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1106_
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1107_
timestamp 1679235063
transform 1 0 24380 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1108_
timestamp 1679235063
transform 1 0 24748 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1109_
timestamp 1679235063
transform 1 0 24104 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1110_
timestamp 1679235063
transform 1 0 19780 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1111_
timestamp 1679235063
transform 1 0 20976 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1112_
timestamp 1679235063
transform 1 0 20148 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1113_
timestamp 1679235063
transform 1 0 20240 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1114_
timestamp 1679235063
transform 1 0 19320 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1115_
timestamp 1679235063
transform 1 0 20148 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1116_
timestamp 1679235063
transform 1 0 19780 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1117_
timestamp 1679235063
transform 1 0 20516 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1118_
timestamp 1679235063
transform 1 0 19872 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1119_
timestamp 1679235063
transform 1 0 9476 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1120_
timestamp 1679235063
transform 1 0 10488 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1121_
timestamp 1679235063
transform 1 0 10028 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _1122_
timestamp 1679235063
transform 1 0 11040 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1123_
timestamp 1679235063
transform 1 0 9384 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1124_
timestamp 1679235063
transform 1 0 10488 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1125_
timestamp 1679235063
transform 1 0 10028 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1126_
timestamp 1679235063
transform 1 0 11776 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1127_
timestamp 1679235063
transform 1 0 10672 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1128_
timestamp 1679235063
transform 1 0 22356 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _1129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22080 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1130_
timestamp 1679235063
transform 1 0 22724 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1131_
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1132_
timestamp 1679235063
transform 1 0 22264 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1133_
timestamp 1679235063
transform 1 0 22356 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1134_
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1135_
timestamp 1679235063
transform 1 0 20056 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1136_
timestamp 1679235063
transform 1 0 20700 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1137_
timestamp 1679235063
transform 1 0 20424 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1138_
timestamp 1679235063
transform 1 0 16744 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1139_
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _1140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20148 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_4  _1141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__nor3_2  _1142_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22264 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1143_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23000 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o32ai_4  _1144_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23460 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1145_
timestamp 1679235063
transform 1 0 28612 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1146_
timestamp 1679235063
transform 1 0 33580 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1147_
timestamp 1679235063
transform 1 0 33488 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1148_
timestamp 1679235063
transform 1 0 29716 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1149_
timestamp 1679235063
transform 1 0 29440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1150_
timestamp 1679235063
transform 1 0 32108 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1151_
timestamp 1679235063
transform 1 0 32200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1152_
timestamp 1679235063
transform 1 0 26956 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1153_
timestamp 1679235063
transform 1 0 26312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1154_
timestamp 1679235063
transform 1 0 34408 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1155_
timestamp 1679235063
transform 1 0 23368 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1156_
timestamp 1679235063
transform 1 0 32936 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1157_
timestamp 1679235063
transform 1 0 32752 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1158_
timestamp 1679235063
transform 1 0 28060 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1159_
timestamp 1679235063
transform 1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1160_
timestamp 1679235063
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1161_
timestamp 1679235063
transform 1 0 30912 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1162_
timestamp 1679235063
transform 1 0 30544 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1163_
timestamp 1679235063
transform 1 0 25760 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1164_
timestamp 1679235063
transform 1 0 25392 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1165_
timestamp 1679235063
transform 1 0 23092 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1166_
timestamp 1679235063
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1167_
timestamp 1679235063
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1168_
timestamp 1679235063
transform 1 0 19596 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1169_
timestamp 1679235063
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1170_
timestamp 1679235063
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1171_
timestamp 1679235063
transform 1 0 22356 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1172_
timestamp 1679235063
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1173_
timestamp 1679235063
transform 1 0 18216 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1174_
timestamp 1679235063
transform 1 0 17480 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1175_
timestamp 1679235063
transform 1 0 23368 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1176_
timestamp 1679235063
transform 1 0 33212 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1177_
timestamp 1679235063
transform 1 0 33028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1178_
timestamp 1679235063
transform 1 0 29532 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1179_
timestamp 1679235063
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1180_
timestamp 1679235063
transform 1 0 30728 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1679235063
transform 1 0 31648 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1182_
timestamp 1679235063
transform 1 0 27048 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1183_
timestamp 1679235063
transform 1 0 26956 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1184_
timestamp 1679235063
transform 1 0 23460 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1185_
timestamp 1679235063
transform 1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1186_
timestamp 1679235063
transform 1 0 21988 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1187_
timestamp 1679235063
transform 1 0 21620 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1188_
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1189_
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1190_
timestamp 1679235063
transform 1 0 20424 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1191_
timestamp 1679235063
transform 1 0 19872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1192_
timestamp 1679235063
transform 1 0 15088 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1193_
timestamp 1679235063
transform 1 0 14720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1194_
timestamp 1679235063
transform 1 0 16744 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1195_
timestamp 1679235063
transform 1 0 15088 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1196_
timestamp 1679235063
transform 1 0 14720 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1197_
timestamp 1679235063
transform 1 0 15824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15088 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1199_
timestamp 1679235063
transform 1 0 11408 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1200_
timestamp 1679235063
transform 1 0 10120 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1201_
timestamp 1679235063
transform 1 0 9752 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1202_
timestamp 1679235063
transform 1 0 10488 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 11408 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1204_
timestamp 1679235063
transform 1 0 10672 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1206_
timestamp 1679235063
transform 1 0 9108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1207_
timestamp 1679235063
transform 1 0 9384 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9752 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1209_
timestamp 1679235063
transform 1 0 10212 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1210_
timestamp 1679235063
transform 1 0 7360 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1211_
timestamp 1679235063
transform 1 0 7084 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 1679235063
transform 1 0 7728 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1213_
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1214_
timestamp 1679235063
transform 1 0 9292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1215_
timestamp 1679235063
transform 1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1216_
timestamp 1679235063
transform 1 0 8740 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1217_
timestamp 1679235063
transform 1 0 7728 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1218_
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1219_
timestamp 1679235063
transform 1 0 7820 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1220_
timestamp 1679235063
transform 1 0 8280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1221_
timestamp 1679235063
transform 1 0 8648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 8188 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1223_
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1224_
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1225_
timestamp 1679235063
transform 1 0 7268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1226_
timestamp 1679235063
transform 1 0 5704 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1227_
timestamp 1679235063
transform 1 0 5888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1228_
timestamp 1679235063
transform 1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1229_
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1230_
timestamp 1679235063
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1231_
timestamp 1679235063
transform 1 0 7820 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1232_
timestamp 1679235063
transform 1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1233_
timestamp 1679235063
transform 1 0 4048 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1234_
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1235_
timestamp 1679235063
transform 1 0 4508 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1236_
timestamp 1679235063
transform 1 0 4968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1237_
timestamp 1679235063
transform 1 0 5336 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1238_
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5520 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1240_
timestamp 1679235063
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _1241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4508 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _1242_
timestamp 1679235063
transform 1 0 4416 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1243_
timestamp 1679235063
transform 1 0 5244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1244_
timestamp 1679235063
transform 1 0 4692 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1245_
timestamp 1679235063
transform 1 0 4416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1246_
timestamp 1679235063
transform 1 0 18216 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1247_
timestamp 1679235063
transform 1 0 17848 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1248_
timestamp 1679235063
transform 1 0 18216 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1249_
timestamp 1679235063
transform 1 0 18768 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1250_
timestamp 1679235063
transform 1 0 13432 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _1251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13892 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1252_
timestamp 1679235063
transform 1 0 14444 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1253_
timestamp 1679235063
transform 1 0 13708 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1254_
timestamp 1679235063
transform 1 0 14996 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1256_
timestamp 1679235063
transform 1 0 19412 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1257_
timestamp 1679235063
transform 1 0 13340 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1258_
timestamp 1679235063
transform 1 0 31096 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1259_
timestamp 1679235063
transform 1 0 32108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1260_
timestamp 1679235063
transform 1 0 32844 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1261_
timestamp 1679235063
transform 1 0 33488 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1262_
timestamp 1679235063
transform 1 0 30728 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_2  _1263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 31004 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1264_
timestamp 1679235063
transform 1 0 18676 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1265_
timestamp 1679235063
transform 1 0 14076 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1266_
timestamp 1679235063
transform 1 0 14076 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1267_
timestamp 1679235063
transform 1 0 12512 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1268_
timestamp 1679235063
transform 1 0 13340 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1269_
timestamp 1679235063
transform 1 0 13340 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _1270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13984 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13800 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13800 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1273_
timestamp 1679235063
transform 1 0 14904 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _1274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13156 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1275_
timestamp 1679235063
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1276_
timestamp 1679235063
transform 1 0 6992 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1277_
timestamp 1679235063
transform 1 0 7820 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1278_
timestamp 1679235063
transform 1 0 12144 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1279_
timestamp 1679235063
transform 1 0 11960 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_2  _1280_
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1281_
timestamp 1679235063
transform 1 0 11500 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1282_
timestamp 1679235063
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 12144 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _1284_
timestamp 1679235063
transform 1 0 18216 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1285_
timestamp 1679235063
transform 1 0 16836 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1286_
timestamp 1679235063
transform 1 0 17388 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1287_
timestamp 1679235063
transform 1 0 16928 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1288_
timestamp 1679235063
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1289_
timestamp 1679235063
transform 1 0 9384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1290_
timestamp 1679235063
transform 1 0 9752 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1291_
timestamp 1679235063
transform 1 0 10396 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1293_
timestamp 1679235063
transform 1 0 12328 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1294_
timestamp 1679235063
transform 1 0 15548 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _1295_
timestamp 1679235063
transform 1 0 11684 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1296_
timestamp 1679235063
transform 1 0 4600 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1297_
timestamp 1679235063
transform 1 0 5244 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1298_
timestamp 1679235063
transform 1 0 4968 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1299_
timestamp 1679235063
transform 1 0 8372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _1300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 8556 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1301_
timestamp 1679235063
transform 1 0 8096 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1302_
timestamp 1679235063
transform 1 0 6808 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1303_
timestamp 1679235063
transform 1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7268 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1305_
timestamp 1679235063
transform 1 0 8004 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1306_
timestamp 1679235063
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1307_
timestamp 1679235063
transform 1 0 7084 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _1308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 12604 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1309_
timestamp 1679235063
transform 1 0 15732 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1310_
timestamp 1679235063
transform 1 0 15272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_2  _1311_
timestamp 1679235063
transform 1 0 19504 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1312_
timestamp 1679235063
transform 1 0 29532 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1313_
timestamp 1679235063
transform 1 0 29532 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1314_
timestamp 1679235063
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1315_
timestamp 1679235063
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6900 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7636 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1318_
timestamp 1679235063
transform 1 0 8096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1319_
timestamp 1679235063
transform 1 0 13248 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1320_
timestamp 1679235063
transform 1 0 12328 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1321_
timestamp 1679235063
transform 1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _1322_
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1323_
timestamp 1679235063
transform 1 0 20700 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1324_
timestamp 1679235063
transform 1 0 24932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1325_
timestamp 1679235063
transform 1 0 25116 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1326_
timestamp 1679235063
transform 1 0 24656 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _1327_
timestamp 1679235063
transform 1 0 7084 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1328_
timestamp 1679235063
transform 1 0 6808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1329_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6164 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1330_
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1331_
timestamp 1679235063
transform 1 0 5888 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1332_
timestamp 1679235063
transform 1 0 10488 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7176 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _1334_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19780 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_4  _1335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17020 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _1336_
timestamp 1679235063
transform 1 0 20884 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1337_
timestamp 1679235063
transform 1 0 21804 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1338_
timestamp 1679235063
transform 1 0 20976 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1340_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4876 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1341_
timestamp 1679235063
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1342_
timestamp 1679235063
transform 1 0 5060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1343_
timestamp 1679235063
transform 1 0 5520 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1344_
timestamp 1679235063
transform 1 0 10856 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1345_
timestamp 1679235063
transform 1 0 10948 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1346_
timestamp 1679235063
transform 1 0 18492 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _1347_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10120 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _1348_
timestamp 1679235063
transform 1 0 9292 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1349_
timestamp 1679235063
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1350_
timestamp 1679235063
transform 1 0 10304 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1351_
timestamp 1679235063
transform 1 0 13432 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1352_
timestamp 1679235063
transform 1 0 31280 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1353_
timestamp 1679235063
transform 1 0 31004 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_2  _1354_
timestamp 1679235063
transform 1 0 30360 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1355_
timestamp 1679235063
transform 1 0 19504 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1356_
timestamp 1679235063
transform 1 0 12512 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1357_
timestamp 1679235063
transform 1 0 12328 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1358_
timestamp 1679235063
transform 1 0 4232 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1359_
timestamp 1679235063
transform 1 0 2852 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1360_
timestamp 1679235063
transform 1 0 1748 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1361_
timestamp 1679235063
transform 1 0 17204 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1362_
timestamp 1679235063
transform 1 0 15732 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1679235063
transform 1 0 15456 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1364_
timestamp 1679235063
transform 1 0 3864 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1365_
timestamp 1679235063
transform 1 0 2392 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1366_
timestamp 1679235063
transform 1 0 2024 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1367_
timestamp 1679235063
transform 1 0 28244 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1368_
timestamp 1679235063
transform 1 0 27416 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1369_
timestamp 1679235063
transform 1 0 27140 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1370_
timestamp 1679235063
transform 1 0 26220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1371_
timestamp 1679235063
transform 1 0 23276 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1372_
timestamp 1679235063
transform 1 0 23000 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1373_
timestamp 1679235063
transform 1 0 20424 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1374_
timestamp 1679235063
transform 1 0 19504 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1375_
timestamp 1679235063
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1376_
timestamp 1679235063
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1377_
timestamp 1679235063
transform 1 0 9292 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1378_
timestamp 1679235063
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1379_
timestamp 1679235063
transform 1 0 32108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1380_
timestamp 1679235063
transform 1 0 33672 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_2  _1381_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 31832 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1382_
timestamp 1679235063
transform 1 0 19504 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1383_
timestamp 1679235063
transform 1 0 12604 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1384_
timestamp 1679235063
transform 1 0 12328 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1385_
timestamp 1679235063
transform 1 0 6716 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1386_
timestamp 1679235063
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1387_
timestamp 1679235063
transform 1 0 16100 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1388_
timestamp 1679235063
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1389_
timestamp 1679235063
transform 1 0 4232 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1390_
timestamp 1679235063
transform 1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1391_
timestamp 1679235063
transform 1 0 30728 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1392_
timestamp 1679235063
transform 1 0 31004 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1393_
timestamp 1679235063
transform 1 0 23736 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1394_
timestamp 1679235063
transform 1 0 24380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1395_
timestamp 1679235063
transform 1 0 19872 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1396_
timestamp 1679235063
transform 1 0 19688 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1397_
timestamp 1679235063
transform 1 0 9568 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1398_
timestamp 1679235063
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1399_
timestamp 1679235063
transform 1 0 32660 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1400_
timestamp 1679235063
transform 1 0 32384 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_2  _1401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 30360 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1402_
timestamp 1679235063
transform 1 0 18124 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1403_
timestamp 1679235063
transform 1 0 14168 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1404_
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1405_
timestamp 1679235063
transform 1 0 2208 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1406_
timestamp 1679235063
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1407_
timestamp 1679235063
transform 1 0 17296 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1408_
timestamp 1679235063
transform 1 0 16744 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1409_
timestamp 1679235063
transform 1 0 2116 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1410_
timestamp 1679235063
transform 1 0 1748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1411_
timestamp 1679235063
transform 1 0 27968 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1412_
timestamp 1679235063
transform 1 0 27416 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1413_
timestamp 1679235063
transform 1 0 25852 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1414_
timestamp 1679235063
transform 1 0 25300 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1415_
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1416_
timestamp 1679235063
transform 1 0 21068 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1417_
timestamp 1679235063
transform 1 0 10672 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1418_
timestamp 1679235063
transform 1 0 9292 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _1419_
timestamp 1679235063
transform 1 0 30268 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1420_
timestamp 1679235063
transform 1 0 18032 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1421_
timestamp 1679235063
transform 1 0 12604 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1422_
timestamp 1679235063
transform 1 0 12328 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1423_
timestamp 1679235063
transform 1 0 2208 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1424_
timestamp 1679235063
transform 1 0 1932 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1425_
timestamp 1679235063
transform 1 0 15916 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1426_
timestamp 1679235063
transform 1 0 15640 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1427_
timestamp 1679235063
transform 1 0 2208 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1428_
timestamp 1679235063
transform 1 0 1840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1429_
timestamp 1679235063
transform 1 0 27876 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1430_
timestamp 1679235063
transform 1 0 27876 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1431_
timestamp 1679235063
transform 1 0 26956 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1432_
timestamp 1679235063
transform 1 0 26128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1433_
timestamp 1679235063
transform 1 0 19596 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1434_
timestamp 1679235063
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1435_
timestamp 1679235063
transform 1 0 9016 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1436_
timestamp 1679235063
transform 1 0 8372 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1437_
timestamp 1679235063
transform 1 0 31648 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _1438_
timestamp 1679235063
transform 1 0 30176 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1439_
timestamp 1679235063
transform 1 0 16744 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1440_
timestamp 1679235063
transform 1 0 12052 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1679235063
transform 1 0 11868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1442_
timestamp 1679235063
transform 1 0 2300 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1679235063
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1444_
timestamp 1679235063
transform 1 0 15916 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1679235063
transform 1 0 15180 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1446_
timestamp 1679235063
transform 1 0 2484 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1447_
timestamp 1679235063
transform 1 0 2208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1448_
timestamp 1679235063
transform 1 0 28244 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1449_
timestamp 1679235063
transform 1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1450_
timestamp 1679235063
transform 1 0 24564 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1451_
timestamp 1679235063
transform 1 0 23368 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1452_
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1453_
timestamp 1679235063
transform 1 0 21160 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1454_
timestamp 1679235063
transform 1 0 8924 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1455_
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _1456_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 32936 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _1457_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 31188 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1458_
timestamp 1679235063
transform 1 0 19780 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1459_
timestamp 1679235063
transform 1 0 12512 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1460_
timestamp 1679235063
transform 1 0 12236 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1461_
timestamp 1679235063
transform 1 0 6164 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1462_
timestamp 1679235063
transform 1 0 6348 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1463_
timestamp 1679235063
transform 1 0 16192 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1464_
timestamp 1679235063
transform 1 0 16652 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1465_
timestamp 1679235063
transform 1 0 5244 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1466_
timestamp 1679235063
transform 1 0 4232 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 1679235063
transform 1 0 29716 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1468_
timestamp 1679235063
transform 1 0 29624 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1469_
timestamp 1679235063
transform 1 0 23828 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1470_
timestamp 1679235063
transform 1 0 24380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1471_
timestamp 1679235063
transform 1 0 19964 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1472_
timestamp 1679235063
transform 1 0 19688 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1473_
timestamp 1679235063
transform 1 0 9568 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1474_
timestamp 1679235063
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _1475_
timestamp 1679235063
transform 1 0 31188 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1476_
timestamp 1679235063
transform 1 0 19596 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1477_
timestamp 1679235063
transform 1 0 12420 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1478_
timestamp 1679235063
transform 1 0 12236 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1479_
timestamp 1679235063
transform 1 0 3864 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1480_
timestamp 1679235063
transform 1 0 3404 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1481_
timestamp 1679235063
transform 1 0 15732 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1482_
timestamp 1679235063
transform 1 0 16008 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1483_
timestamp 1679235063
transform 1 0 3864 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1484_
timestamp 1679235063
transform 1 0 3220 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1485_
timestamp 1679235063
transform 1 0 28520 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1486_
timestamp 1679235063
transform 1 0 27692 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1487_
timestamp 1679235063
transform 1 0 23644 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1488_
timestamp 1679235063
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1489_
timestamp 1679235063
transform 1 0 19320 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1490_
timestamp 1679235063
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1491_
timestamp 1679235063
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1492_
timestamp 1679235063
transform 1 0 8372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_4  _1493_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 32108 0 -1 27200
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1494_
timestamp 1679235063
transform 1 0 19044 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1495_
timestamp 1679235063
transform 1 0 14076 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1679235063
transform 1 0 13616 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1497_
timestamp 1679235063
transform 1 0 7084 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 1679235063
transform 1 0 6624 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1499_
timestamp 1679235063
transform 1 0 18216 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1679235063
transform 1 0 17020 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1501_
timestamp 1679235063
transform 1 0 6256 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1502_
timestamp 1679235063
transform 1 0 5152 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1503_
timestamp 1679235063
transform 1 0 30728 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1504_
timestamp 1679235063
transform 1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1505_
timestamp 1679235063
transform 1 0 26036 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1506_
timestamp 1679235063
transform 1 0 24748 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1507_
timestamp 1679235063
transform 1 0 21804 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1508_
timestamp 1679235063
transform 1 0 20884 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1509_
timestamp 1679235063
transform 1 0 11500 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1510_
timestamp 1679235063
transform 1 0 10212 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_2  _1511_
timestamp 1679235063
transform 1 0 30268 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1512_
timestamp 1679235063
transform 1 0 19228 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1513_
timestamp 1679235063
transform 1 0 14260 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1514_
timestamp 1679235063
transform 1 0 14260 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1515_
timestamp 1679235063
transform 1 0 2300 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1516_
timestamp 1679235063
transform 1 0 1932 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1517_
timestamp 1679235063
transform 1 0 17480 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1518_
timestamp 1679235063
transform 1 0 17112 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1519_
timestamp 1679235063
transform 1 0 2300 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1520_
timestamp 1679235063
transform 1 0 1932 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 1679235063
transform 1 0 27508 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1522_
timestamp 1679235063
transform 1 0 27232 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1523_
timestamp 1679235063
transform 1 0 26404 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1524_
timestamp 1679235063
transform 1 0 26496 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1525_
timestamp 1679235063
transform 1 0 21988 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1526_
timestamp 1679235063
transform 1 0 22816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1527_
timestamp 1679235063
transform 1 0 9752 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1528_
timestamp 1679235063
transform 1 0 9292 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1529_
timestamp 1679235063
transform 1 0 27600 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1530_
timestamp 1679235063
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1531_
timestamp 1679235063
transform 1 0 28796 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1532_
timestamp 1679235063
transform 1 0 34684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1533_
timestamp 1679235063
transform 1 0 33948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1534_
timestamp 1679235063
transform 1 0 33856 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1535_
timestamp 1679235063
transform 1 0 33764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _1536_
timestamp 1679235063
transform 1 0 26864 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1537_
timestamp 1679235063
transform 1 0 33764 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1538_
timestamp 1679235063
transform 1 0 33212 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1539_
timestamp 1679235063
transform 1 0 33672 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1540_
timestamp 1679235063
transform 1 0 30544 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1541_
timestamp 1679235063
transform 1 0 30268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1542_
timestamp 1679235063
transform 1 0 33488 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1543_
timestamp 1679235063
transform 1 0 33028 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 33212 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_2  _1545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 33488 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1546_
timestamp 1679235063
transform 1 0 34592 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1547_
timestamp 1679235063
transform 1 0 34224 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1548_
timestamp 1679235063
transform 1 0 34316 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1549_
timestamp 1679235063
transform 1 0 33488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1550_
timestamp 1679235063
transform 1 0 33120 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1551_
timestamp 1679235063
transform 1 0 30176 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1552_
timestamp 1679235063
transform 1 0 29072 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1553_
timestamp 1679235063
transform 1 0 32568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1554_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 32108 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _1555_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 31464 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1556_
timestamp 1679235063
transform 1 0 31188 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1557_
timestamp 1679235063
transform 1 0 31924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1558_
timestamp 1679235063
transform 1 0 31740 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 32384 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1560_
timestamp 1679235063
transform 1 0 30912 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_4  _1561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 30544 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__a21boi_1  _1562_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 31464 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a2111oi_1  _1563_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 32108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1564_
timestamp 1679235063
transform 1 0 32108 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1565_
timestamp 1679235063
transform 1 0 30636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1566_
timestamp 1679235063
transform 1 0 30452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1567_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 32200 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_2  _1568_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 32200 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1569_
timestamp 1679235063
transform 1 0 28060 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1570_
timestamp 1679235063
transform 1 0 28520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1571_
timestamp 1679235063
transform 1 0 27600 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _1572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 29256 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1573_
timestamp 1679235063
transform 1 0 28612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1574_
timestamp 1679235063
transform 1 0 29808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1575_
timestamp 1679235063
transform 1 0 29808 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _1576_
timestamp 1679235063
transform 1 0 30360 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1577_
timestamp 1679235063
transform 1 0 29532 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1578_
timestamp 1679235063
transform 1 0 29256 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1579_
timestamp 1679235063
transform 1 0 25852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1580_
timestamp 1679235063
transform 1 0 30728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1581_
timestamp 1679235063
transform 1 0 31004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1582_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 31464 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1583_
timestamp 1679235063
transform 1 0 30820 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1584_
timestamp 1679235063
transform 1 0 26128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1585_
timestamp 1679235063
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1586_
timestamp 1679235063
transform 1 0 27508 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1587_
timestamp 1679235063
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1588_
timestamp 1679235063
transform 1 0 31188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1589_
timestamp 1679235063
transform 1 0 30268 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1590_
timestamp 1679235063
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1591_
timestamp 1679235063
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1592_
timestamp 1679235063
transform 1 0 28612 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 27876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1594_
timestamp 1679235063
transform 1 0 27232 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1595_
timestamp 1679235063
transform 1 0 28060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1596_
timestamp 1679235063
transform 1 0 29164 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1597_
timestamp 1679235063
transform 1 0 29716 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1598_
timestamp 1679235063
transform 1 0 31096 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1599_
timestamp 1679235063
transform 1 0 31096 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1600_
timestamp 1679235063
transform 1 0 31740 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1601_
timestamp 1679235063
transform 1 0 31004 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1602_
timestamp 1679235063
transform 1 0 25300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1603_
timestamp 1679235063
transform 1 0 25024 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1604_
timestamp 1679235063
transform 1 0 26312 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1605_
timestamp 1679235063
transform 1 0 25668 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1606_
timestamp 1679235063
transform 1 0 26772 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1607_
timestamp 1679235063
transform 1 0 27968 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1608_
timestamp 1679235063
transform 1 0 27508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _1609_
timestamp 1679235063
transform 1 0 27140 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__a311o_1  _1610_
timestamp 1679235063
transform 1 0 27968 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1611_
timestamp 1679235063
transform 1 0 27600 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1612_
timestamp 1679235063
transform 1 0 31096 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1613_
timestamp 1679235063
transform 1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1614_
timestamp 1679235063
transform 1 0 30084 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1615_
timestamp 1679235063
transform 1 0 30360 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _1616_
timestamp 1679235063
transform 1 0 31372 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1617_
timestamp 1679235063
transform 1 0 27600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1618_
timestamp 1679235063
transform 1 0 24196 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24840 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1620_
timestamp 1679235063
transform 1 0 25484 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1621_
timestamp 1679235063
transform 1 0 28244 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1622_
timestamp 1679235063
transform 1 0 27508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1623_
timestamp 1679235063
transform 1 0 28796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1625_
timestamp 1679235063
transform 1 0 31832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1626_
timestamp 1679235063
transform 1 0 24840 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1627_
timestamp 1679235063
transform 1 0 25668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1628_
timestamp 1679235063
transform 1 0 25760 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1629_
timestamp 1679235063
transform 1 0 26496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1630_
timestamp 1679235063
transform 1 0 27232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1631_
timestamp 1679235063
transform 1 0 24840 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _1632_
timestamp 1679235063
transform 1 0 25944 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1633_
timestamp 1679235063
transform 1 0 25852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1634_
timestamp 1679235063
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 27508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _1636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 26496 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1637_
timestamp 1679235063
transform 1 0 28152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1638_
timestamp 1679235063
transform 1 0 32108 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1639_
timestamp 1679235063
transform 1 0 30636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1640_
timestamp 1679235063
transform 1 0 31280 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_1  _1641_
timestamp 1679235063
transform 1 0 32108 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_2  _1642_
timestamp 1679235063
transform 1 0 30452 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1643_
timestamp 1679235063
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1644_
timestamp 1679235063
transform 1 0 14076 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1645_
timestamp 1679235063
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1646_
timestamp 1679235063
transform 1 0 4140 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1647_
timestamp 1679235063
transform 1 0 2760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1648_
timestamp 1679235063
transform 1 0 18216 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1649_
timestamp 1679235063
transform 1 0 17572 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1650_
timestamp 1679235063
transform 1 0 4140 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1651_
timestamp 1679235063
transform 1 0 3864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1652_
timestamp 1679235063
transform 1 0 28336 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1653_
timestamp 1679235063
transform 1 0 27692 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1654_
timestamp 1679235063
transform 1 0 26312 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1655_
timestamp 1679235063
transform 1 0 25944 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1656_
timestamp 1679235063
transform 1 0 21160 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1657_
timestamp 1679235063
transform 1 0 21344 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1658_
timestamp 1679235063
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1659_
timestamp 1679235063
transform 1 0 10120 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1661_
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1662_
timestamp 1679235063
transform 1 0 24840 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _1663_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 31372 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1664_
timestamp 1679235063
transform 1 0 17572 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 1679235063
transform 1 0 12880 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1666_
timestamp 1679235063
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1667_
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1668_
timestamp 1679235063
transform 1 0 5336 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1669_
timestamp 1679235063
transform 1 0 16100 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1670_
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1671_
timestamp 1679235063
transform 1 0 4048 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1672_
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1673_
timestamp 1679235063
transform 1 0 27692 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1674_
timestamp 1679235063
transform 1 0 27048 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1675_
timestamp 1679235063
transform 1 0 23276 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1676_
timestamp 1679235063
transform 1 0 22632 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1677_
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1678_
timestamp 1679235063
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1679_
timestamp 1679235063
transform 1 0 10304 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1680_
timestamp 1679235063
transform 1 0 9016 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _1681_
timestamp 1679235063
transform 1 0 31280 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1682_
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1683_
timestamp 1679235063
transform 1 0 12880 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1684_
timestamp 1679235063
transform 1 0 11776 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1685_
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1686_
timestamp 1679235063
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1687_
timestamp 1679235063
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1688_
timestamp 1679235063
transform 1 0 15272 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 1679235063
transform 1 0 2852 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1690_
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1691_
timestamp 1679235063
transform 1 0 29532 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1692_
timestamp 1679235063
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1693_
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1694_
timestamp 1679235063
transform 1 0 23736 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1695_
timestamp 1679235063
transform 1 0 18952 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1696_
timestamp 1679235063
transform 1 0 18768 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1697_
timestamp 1679235063
transform 1 0 9016 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1698_
timestamp 1679235063
transform 1 0 7912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _1699_
timestamp 1679235063
transform 1 0 30360 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1700_
timestamp 1679235063
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1701_
timestamp 1679235063
transform 1 0 12052 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1702_
timestamp 1679235063
transform 1 0 11776 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1703_
timestamp 1679235063
transform 1 0 4784 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1704_
timestamp 1679235063
transform 1 0 4600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1705_
timestamp 1679235063
transform 1 0 16376 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1706_
timestamp 1679235063
transform 1 0 15272 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1707_
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1708_
timestamp 1679235063
transform 1 0 2852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1709_
timestamp 1679235063
transform 1 0 27416 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1710_
timestamp 1679235063
transform 1 0 26220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1711_
timestamp 1679235063
transform 1 0 22816 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1679235063
transform 1 0 22724 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1713_
timestamp 1679235063
transform 1 0 18860 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1714_
timestamp 1679235063
transform 1 0 18768 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1715_
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1716_
timestamp 1679235063
transform 1 0 8004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_4  _1717_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 30268 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1718_
timestamp 1679235063
transform 1 0 18584 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1719_
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1720_
timestamp 1679235063
transform 1 0 13248 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1721_
timestamp 1679235063
transform 1 0 6440 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1722_
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1723_
timestamp 1679235063
transform 1 0 17020 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1724_
timestamp 1679235063
transform 1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1725_
timestamp 1679235063
transform 1 0 4416 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1726_
timestamp 1679235063
transform 1 0 3956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1727_
timestamp 1679235063
transform 1 0 29808 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1728_
timestamp 1679235063
transform 1 0 29716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1729_
timestamp 1679235063
transform 1 0 24932 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1730_
timestamp 1679235063
transform 1 0 24932 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1731_
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1732_
timestamp 1679235063
transform 1 0 20976 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1733_
timestamp 1679235063
transform 1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1734_
timestamp 1679235063
transform 1 0 9568 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1735_
timestamp 1679235063
transform 1 0 23092 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1736_
timestamp 1679235063
transform 1 0 24288 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1737_
timestamp 1679235063
transform 1 0 21528 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _1738_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23736 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1739_
timestamp 1679235063
transform 1 0 22540 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1740_
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1741_
timestamp 1679235063
transform 1 0 23644 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1742_
timestamp 1679235063
transform 1 0 25484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a2111oi_1  _1743_
timestamp 1679235063
transform 1 0 23920 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_4  _1744_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 32108 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1745_
timestamp 1679235063
transform 1 0 17480 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1746_
timestamp 1679235063
transform 1 0 12420 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1747_
timestamp 1679235063
transform 1 0 12236 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1748_
timestamp 1679235063
transform 1 0 5060 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1749_
timestamp 1679235063
transform 1 0 4600 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1750_
timestamp 1679235063
transform 1 0 16652 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1751_
timestamp 1679235063
transform 1 0 15916 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1752_
timestamp 1679235063
transform 1 0 4048 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1753_
timestamp 1679235063
transform 1 0 3772 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1754_
timestamp 1679235063
transform 1 0 29440 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1755_
timestamp 1679235063
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1756_
timestamp 1679235063
transform 1 0 24472 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1757_
timestamp 1679235063
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1758_
timestamp 1679235063
transform 1 0 19872 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1759_
timestamp 1679235063
transform 1 0 19688 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1760_
timestamp 1679235063
transform 1 0 10304 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1761_
timestamp 1679235063
transform 1 0 9108 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1762_
timestamp 1679235063
transform 1 0 18032 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1763_
timestamp 1679235063
transform 1 0 29532 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1764_
timestamp 1679235063
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1765_
timestamp 1679235063
transform 1 0 29716 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1766_
timestamp 1679235063
transform 1 0 29348 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1767_
timestamp 1679235063
transform 1 0 17940 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1768_
timestamp 1679235063
transform 1 0 17112 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1769_
timestamp 1679235063
transform 1 0 16652 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1770_
timestamp 1679235063
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1771_
timestamp 1679235063
transform 1 0 21804 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1772_
timestamp 1679235063
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1773_
timestamp 1679235063
transform 1 0 19504 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1774_
timestamp 1679235063
transform 1 0 18952 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1775_
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1776_
timestamp 1679235063
transform 1 0 23828 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1777_
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1778_
timestamp 1679235063
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1779_
timestamp 1679235063
transform 1 0 34684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1780_
timestamp 1679235063
transform 1 0 24380 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1781_
timestamp 1679235063
transform 1 0 34684 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1782_
timestamp 1679235063
transform 1 0 15456 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1783_
timestamp 1679235063
transform 1 0 15088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1784_
timestamp 1679235063
transform 1 0 14536 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1785_
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1786_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20700 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1787_
timestamp 1679235063
transform 1 0 25116 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _1788_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23552 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1789_
timestamp 1679235063
transform 1 0 31464 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1790_
timestamp 1679235063
transform 1 0 22264 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1791_
timestamp 1679235063
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1792_
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1793_
timestamp 1679235063
transform 1 0 18308 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1794_
timestamp 1679235063
transform 1 0 20424 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1795_
timestamp 1679235063
transform 1 0 20240 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1796_
timestamp 1679235063
transform 1 0 16744 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1797_
timestamp 1679235063
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1798_
timestamp 1679235063
transform 1 0 33764 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1799_
timestamp 1679235063
transform 1 0 34684 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1800_
timestamp 1679235063
transform 1 0 29716 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1801_
timestamp 1679235063
transform 1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1802_
timestamp 1679235063
transform 1 0 32108 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1803_
timestamp 1679235063
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1804_
timestamp 1679235063
transform 1 0 27048 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1805_
timestamp 1679235063
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1806_
timestamp 1679235063
transform 1 0 33120 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1807_
timestamp 1679235063
transform 1 0 32660 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1808_
timestamp 1679235063
transform 1 0 33120 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1809_
timestamp 1679235063
transform 1 0 30544 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1810_
timestamp 1679235063
transform 1 0 30360 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1811_
timestamp 1679235063
transform 1 0 31188 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1812_
timestamp 1679235063
transform 1 0 32936 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1813_
timestamp 1679235063
transform 1 0 32108 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1814_
timestamp 1679235063
transform 1 0 32384 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1815_
timestamp 1679235063
transform 1 0 27784 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1816_
timestamp 1679235063
transform 1 0 32936 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1817_
timestamp 1679235063
transform 1 0 33764 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1818_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13616 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1679235063
transform 1 0 7176 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1679235063
transform 1 0 17204 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1679235063
transform 1 0 4600 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1679235063
transform 1 0 29532 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1679235063
transform 1 0 24932 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1679235063
transform 1 0 21252 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1679235063
transform 1 0 9936 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtp_1  _1826_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13800 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1827_
timestamp 1679235063
transform 1 0 6900 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1828_
timestamp 1679235063
transform 1 0 15364 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1829_
timestamp 1679235063
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1830_
timestamp 1679235063
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1831_
timestamp 1679235063
transform -1 0 6072 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1832_
timestamp 1679235063
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1833_
timestamp 1679235063
transform 1 0 4416 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1834_
timestamp 1679235063
transform 1 0 12696 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1835_
timestamp 1679235063
transform 1 0 7820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1836_
timestamp 1679235063
transform 1 0 17296 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1837_
timestamp 1679235063
transform 1 0 7084 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1838_
timestamp 1679235063
transform 1 0 25392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1839_
timestamp 1679235063
transform 1 0 15456 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1840_
timestamp 1679235063
transform 1 0 18216 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1841_
timestamp 1679235063
transform 1 0 10488 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1679235063
transform 1 0 12144 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1679235063
transform 1 0 1380 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1679235063
transform 1 0 15180 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1679235063
transform 1 0 1748 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1679235063
transform 1 0 26864 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1679235063
transform 1 0 22632 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1679235063
transform 1 0 18308 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1679235063
transform 1 0 8372 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1679235063
transform 1 0 11960 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1679235063
transform 1 0 6440 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1679235063
transform 1 0 15088 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1679235063
transform 1 0 3772 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1679235063
transform 1 0 30544 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1679235063
transform 1 0 22816 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1679235063
transform 1 0 19412 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1679235063
transform 1 0 8464 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1679235063
transform 1 0 14444 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1679235063
transform 1 0 1472 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1679235063
transform 1 0 17020 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1679235063
transform 1 0 27692 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1679235063
transform 1 0 25576 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1679235063
transform 1 0 21344 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1679235063
transform 1 0 9200 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1679235063
transform 1 0 33028 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1679235063
transform 1 0 29532 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1679235063
transform 1 0 32384 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1869_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24840 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1679235063
transform 1 0 12052 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1679235063
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1679235063
transform 1 0 15088 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1679235063
transform 1 0 1472 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1679235063
transform 1 0 27600 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1679235063
transform 1 0 25944 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1679235063
transform 1 0 19228 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1679235063
transform 1 0 11500 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1679235063
transform 1 0 14812 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1679235063
transform 1 0 1840 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1679235063
transform 1 0 27968 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1679235063
transform 1 0 23092 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1679235063
transform 1 0 21436 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1679235063
transform 1 0 8004 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1679235063
transform 1 0 11868 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1679235063
transform 1 0 5796 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1679235063
transform 1 0 15088 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1679235063
transform 1 0 3772 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1679235063
transform 1 0 29348 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1679235063
transform 1 0 22816 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1679235063
transform 1 0 19412 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1679235063
transform 1 0 8464 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1679235063
transform 1 0 11868 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1679235063
transform 1 0 3772 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1679235063
transform 1 0 15456 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1679235063
transform 1 0 3496 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1679235063
transform 1 0 27968 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1679235063
transform 1 0 23092 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1679235063
transform 1 0 19136 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1679235063
transform 1 0 8372 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1679235063
transform 1 0 13432 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1679235063
transform 1 0 6900 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1679235063
transform 1 0 17204 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1679235063
transform 1 0 4784 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1679235063
transform 1 0 30728 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1679235063
transform 1 0 25024 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1679235063
transform 1 0 21160 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1679235063
transform 1 0 9936 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1679235063
transform 1 0 14076 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1679235063
transform 1 0 1656 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1679235063
transform 1 0 17388 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1679235063
transform 1 0 1564 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1679235063
transform 1 0 27048 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1679235063
transform 1 0 26956 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1679235063
transform 1 0 21896 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1679235063
transform 1 0 9292 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1679235063
transform 1 0 34960 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1919_
timestamp 1679235063
transform 1 0 34684 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1679235063
transform 1 0 32200 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1921_
timestamp 1679235063
transform 1 0 29532 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1679235063
transform 1 0 24932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1679235063
transform 1 0 32752 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1924_
timestamp 1679235063
transform 1 0 28520 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1925_
timestamp 1679235063
transform 1 0 32752 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1679235063
transform 1 0 13616 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1679235063
transform 1 0 3036 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1679235063
transform 1 0 17296 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1679235063
transform 1 0 3588 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1679235063
transform 1 0 27968 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1679235063
transform 1 0 25392 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1679235063
transform 1 0 21804 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1679235063
transform 1 0 9936 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1679235063
transform 1 0 32752 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1935_
timestamp 1679235063
transform 1 0 22724 0 -1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1679235063
transform 1 0 34960 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1937_
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1938_
timestamp 1679235063
transform 1 0 9292 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1679235063
transform 1 0 2852 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1679235063
transform 1 0 17572 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1679235063
transform 1 0 25392 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1679235063
transform 1 0 22264 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1944_
timestamp 1679235063
transform 1 0 20148 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1945_
timestamp 1679235063
transform 1 0 20700 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1946_
timestamp 1679235063
transform 1 0 16468 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1679235063
transform 1 0 12512 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1679235063
transform 1 0 5060 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1679235063
transform 1 0 15088 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1950_
timestamp 1679235063
transform 1 0 3128 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1951_
timestamp 1679235063
transform 1 0 27324 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1952_
timestamp 1679235063
transform 1 0 22908 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1679235063
transform 1 0 18400 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1954_
timestamp 1679235063
transform 1 0 8832 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1679235063
transform 1 0 11408 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1679235063
transform 1 0 3036 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1679235063
transform 1 0 14904 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1958_
timestamp 1679235063
transform 1 0 2944 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1679235063
transform 1 0 28888 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1679235063
transform 1 0 23368 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1961_
timestamp 1679235063
transform 1 0 18492 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1962_
timestamp 1679235063
transform 1 0 7544 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1964_
timestamp 1679235063
transform 1 0 4324 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1965_
timestamp 1679235063
transform 1 0 14904 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1966_
timestamp 1679235063
transform 1 0 2392 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1967_
timestamp 1679235063
transform 1 0 25944 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1968_
timestamp 1679235063
transform 1 0 22448 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1970_
timestamp 1679235063
transform 1 0 7360 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1971_
timestamp 1679235063
transform 1 0 13524 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1972_
timestamp 1679235063
transform 1 0 5888 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1973_
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1974_
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1975_
timestamp 1679235063
transform 1 0 29440 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1976_
timestamp 1679235063
transform 1 0 24932 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1977_
timestamp 1679235063
transform 1 0 20700 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1978_
timestamp 1679235063
transform 1 0 9660 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1979_
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1980_
timestamp 1679235063
transform 1 0 21252 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1981_
timestamp 1679235063
transform 1 0 17296 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1982_
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1983_
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1984_
timestamp 1679235063
transform 1 0 17940 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1985_
timestamp 1679235063
transform 1 0 24748 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1986_
timestamp 1679235063
transform 1 0 24472 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1987_
timestamp 1679235063
transform 1 0 11868 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1988_
timestamp 1679235063
transform 1 0 4048 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1989_
timestamp 1679235063
transform 1 0 15088 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1990_
timestamp 1679235063
transform 1 0 3312 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1991_
timestamp 1679235063
transform 1 0 29532 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1992_
timestamp 1679235063
transform 1 0 24104 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1993_
timestamp 1679235063
transform 1 0 19320 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1994_
timestamp 1679235063
transform 1 0 8832 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _1995_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 33028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _1996_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 28152 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _1997_
timestamp 1679235063
transform 1 0 30820 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _1998_
timestamp 1679235063
transform 1 0 25668 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _1999_
timestamp 1679235063
transform 1 0 22816 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _2000_
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _2001_
timestamp 1679235063
transform 1 0 22448 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2002_
timestamp 1679235063
transform 1 0 17756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2003_
timestamp 1679235063
transform 1 0 28888 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2004_
timestamp 1679235063
transform 1 0 29624 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2005_
timestamp 1679235063
transform 1 0 17388 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2006_
timestamp 1679235063
transform 1 0 15824 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2007_
timestamp 1679235063
transform 1 0 21252 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2008_
timestamp 1679235063
transform 1 0 19228 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2009_
timestamp 1679235063
transform 1 0 24104 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2010_
timestamp 1679235063
transform 1 0 15732 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2011_
timestamp 1679235063
transform 1 0 34592 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2012_
timestamp 1679235063
transform 1 0 34132 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _2013_
timestamp 1679235063
transform 1 0 33304 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2014_
timestamp 1679235063
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2015_
timestamp 1679235063
transform 1 0 31556 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2016_
timestamp 1679235063
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2017_
timestamp 1679235063
transform 1 0 23184 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2018_
timestamp 1679235063
transform 1 0 21896 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2019_
timestamp 1679235063
transform 1 0 21252 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2020_
timestamp 1679235063
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2021_
timestamp 1679235063
transform 1 0 14536 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2022_
timestamp 1679235063
transform 1 0 13156 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2023_
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2024_
timestamp 1679235063
transform 1 0 24564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2025_
timestamp 1679235063
transform 1 0 32108 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2026_
timestamp 1679235063
transform 1 0 21988 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2027_
timestamp 1679235063
transform 1 0 17940 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2028_
timestamp 1679235063
transform 1 0 19964 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2029_
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2030_
timestamp 1679235063
transform 1 0 33120 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2031_
timestamp 1679235063
transform 1 0 29164 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2032_
timestamp 1679235063
transform 1 0 31556 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2033_
timestamp 1679235063
transform 1 0 26496 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2034_
timestamp 1679235063
transform 1 0 33120 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2035_
timestamp 1679235063
transform 1 0 30912 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2036_
timestamp 1679235063
transform 1 0 32476 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2037_
timestamp 1679235063
transform 1 0 33120 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _2039_
timestamp 1679235063
transform 1 0 6808 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2040_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14720 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2041_
timestamp 1679235063
transform 1 0 13064 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2042_
timestamp 1679235063
transform 1 0 11592 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2043_
timestamp 1679235063
transform 1 0 9752 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2044_
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2045_
timestamp 1679235063
transform 1 0 11500 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2046_
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2047_
timestamp 1679235063
transform 1 0 9844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 30544 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform -1 0 4784 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 35604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1679235063
transform -1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1679235063
transform -1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1679235063
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout51
timestamp 1679235063
transform 1 0 7636 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 1679235063
transform 1 0 25944 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout53
timestamp 1679235063
transform 1 0 25668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout54
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout55
timestamp 1679235063
transform 1 0 21344 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout56
timestamp 1679235063
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout57
timestamp 1679235063
transform 1 0 31096 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout58
timestamp 1679235063
transform 1 0 21344 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout59
timestamp 1679235063
transform 1 0 24104 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout60
timestamp 1679235063
transform 1 0 23184 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout61
timestamp 1679235063
transform 1 0 33028 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout62
timestamp 1679235063
transform 1 0 34040 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout63
timestamp 1679235063
transform 1 0 18032 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout64
timestamp 1679235063
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout65
timestamp 1679235063
transform 1 0 7912 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout66
timestamp 1679235063
transform 1 0 9292 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout67
timestamp 1679235063
transform 1 0 9936 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout68
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout69
timestamp 1679235063
transform 1 0 14996 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout70
timestamp 1679235063
transform 1 0 14996 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout71
timestamp 1679235063
transform 1 0 33672 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout72
timestamp 1679235063
transform 1 0 26220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout73
timestamp 1679235063
transform 1 0 35052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout74
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout75
timestamp 1679235063
transform 1 0 25576 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout76
timestamp 1679235063
transform 1 0 25668 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout77
timestamp 1679235063
transform 1 0 26956 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout78
timestamp 1679235063
transform 1 0 33120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout79
timestamp 1679235063
transform 1 0 34684 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout80
timestamp 1679235063
transform 1 0 34684 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout81
timestamp 1679235063
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout82
timestamp 1679235063
transform 1 0 4692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout83
timestamp 1679235063
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout84
timestamp 1679235063
transform 1 0 8924 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout85
timestamp 1679235063
transform 1 0 17296 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout86
timestamp 1679235063
transform 1 0 18768 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout87
timestamp 1679235063
transform 1 0 19136 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout88
timestamp 1679235063
transform 1 0 6900 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout89
timestamp 1679235063
transform 1 0 9844 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout90
timestamp 1679235063
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout91
timestamp 1679235063
transform 1 0 7084 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout92
timestamp 1679235063
transform 1 0 17204 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout93
timestamp 1679235063
transform 1 0 17296 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout94
timestamp 1679235063
transform 1 0 17480 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout95
timestamp 1679235063
transform 1 0 17664 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout96
timestamp 1679235063
transform 1 0 19228 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout97
timestamp 1679235063
transform 1 0 25576 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout98
timestamp 1679235063
transform 1 0 25760 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout99
timestamp 1679235063
transform 1 0 33212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout100
timestamp 1679235063
transform 1 0 32200 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout101
timestamp 1679235063
transform 1 0 32752 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout102
timestamp 1679235063
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout103
timestamp 1679235063
transform 1 0 25116 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout104
timestamp 1679235063
transform 1 0 25024 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout105
timestamp 1679235063
transform 1 0 30820 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout106
timestamp 1679235063
transform 1 0 29072 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout107
timestamp 1679235063
transform 1 0 29900 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout108
timestamp 1679235063
transform 1 0 30820 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout109
timestamp 1679235063
transform 1 0 29992 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13
timestamp 1679235063
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21
timestamp 1679235063
transform 1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49
timestamp 1679235063
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1679235063
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1679235063
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90
timestamp 1679235063
transform 1 0 9384 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102
timestamp 1679235063
transform 1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1679235063
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119
timestamp 1679235063
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1679235063
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1679235063
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1679235063
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154
timestamp 1679235063
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1679235063
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1679235063
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_209
timestamp 1679235063
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_217
timestamp 1679235063
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1679235063
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_237
timestamp 1679235063
transform 1 0 22908 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_245
timestamp 1679235063
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_265
timestamp 1679235063
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1679235063
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_286
timestamp 1679235063
transform 1 0 27416 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_298
timestamp 1679235063
transform 1 0 28520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1679235063
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309
timestamp 1679235063
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_325
timestamp 1679235063
transform 1 0 31004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1679235063
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1679235063
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1679235063
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1679235063
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1679235063
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1679235063
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_373
timestamp 1679235063
transform 1 0 35420 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6
timestamp 1679235063
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_18
timestamp 1679235063
transform 1 0 2760 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_35
timestamp 1679235063
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1679235063
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1679235063
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1679235063
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1679235063
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1679235063
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1679235063
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1679235063
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1679235063
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1679235063
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1679235063
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_161
timestamp 1679235063
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1679235063
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_178
timestamp 1679235063
transform 1 0 17480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1679235063
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_202
timestamp 1679235063
transform 1 0 19688 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1679235063
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1679235063
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_237
timestamp 1679235063
transform 1 0 22908 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_245
timestamp 1679235063
transform 1 0 23644 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_265
timestamp 1679235063
transform 1 0 25484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_275
timestamp 1679235063
transform 1 0 26404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1679235063
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_291
timestamp 1679235063
transform 1 0 27876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_297
timestamp 1679235063
transform 1 0 28428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_315
timestamp 1679235063
transform 1 0 30084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_323
timestamp 1679235063
transform 1 0 30820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_327
timestamp 1679235063
transform 1 0 31188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1679235063
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_342
timestamp 1679235063
transform 1 0 32568 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_360
timestamp 1679235063
transform 1 0 34224 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_372
timestamp 1679235063
transform 1 0 35328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_377
timestamp 1679235063
transform 1 0 35788 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1679235063
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1679235063
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1679235063
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1679235063
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1679235063
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1679235063
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1679235063
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1679235063
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1679235063
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1679235063
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1679235063
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1679235063
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_153
timestamp 1679235063
transform 1 0 15180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_175
timestamp 1679235063
transform 1 0 17204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 1679235063
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_231
timestamp 1679235063
transform 1 0 22356 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp 1679235063
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp 1679235063
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_273
timestamp 1679235063
transform 1 0 26220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_283
timestamp 1679235063
transform 1 0 27140 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_291
timestamp 1679235063
transform 1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_298
timestamp 1679235063
transform 1 0 28520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1679235063
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_317
timestamp 1679235063
transform 1 0 30268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_343
timestamp 1679235063
transform 1 0 32660 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_361
timestamp 1679235063
transform 1 0 34316 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1679235063
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_377
timestamp 1679235063
transform 1 0 35788 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1679235063
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1679235063
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1679235063
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1679235063
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1679235063
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_74
timestamp 1679235063
transform 1 0 7912 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_86
timestamp 1679235063
transform 1 0 9016 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1679235063
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1679235063
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1679235063
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1679235063
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1679235063
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1679235063
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_185
timestamp 1679235063
transform 1 0 18124 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_195
timestamp 1679235063
transform 1 0 19044 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_210
timestamp 1679235063
transform 1 0 20424 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1679235063
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_228
timestamp 1679235063
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_240
timestamp 1679235063
transform 1 0 23184 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_252
timestamp 1679235063
transform 1 0 24288 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_264
timestamp 1679235063
transform 1 0 25392 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1679235063
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1679235063
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1679235063
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_305
timestamp 1679235063
transform 1 0 29164 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_313
timestamp 1679235063
transform 1 0 29900 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_326
timestamp 1679235063
transform 1 0 31096 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1679235063
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1679235063
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1679235063
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1679235063
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1679235063
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1679235063
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1679235063
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1679235063
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1679235063
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1679235063
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1679235063
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1679235063
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1679235063
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1679235063
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1679235063
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1679235063
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_165
timestamp 1679235063
transform 1 0 16284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_169
timestamp 1679235063
transform 1 0 16652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_176
timestamp 1679235063
transform 1 0 17296 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_188
timestamp 1679235063
transform 1 0 18400 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1679235063
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1679235063
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1679235063
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1679235063
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1679235063
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_257
timestamp 1679235063
transform 1 0 24748 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_270
timestamp 1679235063
transform 1 0 25944 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_282
timestamp 1679235063
transform 1 0 27048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_286
timestamp 1679235063
transform 1 0 27416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1679235063
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1679235063
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1679235063
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_325
timestamp 1679235063
transform 1 0 31004 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_330
timestamp 1679235063
transform 1 0 31464 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_342
timestamp 1679235063
transform 1 0 32568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_354
timestamp 1679235063
transform 1 0 33672 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1679235063
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1679235063
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_377
timestamp 1679235063
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1679235063
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1679235063
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1679235063
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1679235063
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_73
timestamp 1679235063
transform 1 0 7820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_85
timestamp 1679235063
transform 1 0 8924 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_91
timestamp 1679235063
transform 1 0 9476 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_96
timestamp 1679235063
transform 1 0 9936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1679235063
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_119
timestamp 1679235063
transform 1 0 12052 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_127
timestamp 1679235063
transform 1 0 12788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_139
timestamp 1679235063
transform 1 0 13892 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_147
timestamp 1679235063
transform 1 0 14628 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_160
timestamp 1679235063
transform 1 0 15824 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_180
timestamp 1679235063
transform 1 0 17664 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_192
timestamp 1679235063
transform 1 0 18768 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_200
timestamp 1679235063
transform 1 0 19504 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_214
timestamp 1679235063
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1679235063
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_236
timestamp 1679235063
transform 1 0 22816 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_242
timestamp 1679235063
transform 1 0 23368 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_252
timestamp 1679235063
transform 1 0 24288 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_265
timestamp 1679235063
transform 1 0 25484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 1679235063
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp 1679235063
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_288
timestamp 1679235063
transform 1 0 27600 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_300
timestamp 1679235063
transform 1 0 28704 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_312
timestamp 1679235063
transform 1 0 29808 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_320
timestamp 1679235063
transform 1 0 30544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_325
timestamp 1679235063
transform 1 0 31004 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_331
timestamp 1679235063
transform 1 0 31556 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_337
timestamp 1679235063
transform 1 0 32108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_343
timestamp 1679235063
transform 1 0 32660 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_360
timestamp 1679235063
transform 1 0 34224 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_372
timestamp 1679235063
transform 1 0 35328 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_380
timestamp 1679235063
transform 1 0 36064 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7
timestamp 1679235063
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1679235063
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1679235063
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1679235063
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1679235063
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_90
timestamp 1679235063
transform 1 0 9384 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_105
timestamp 1679235063
transform 1 0 10764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_129
timestamp 1679235063
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 1679235063
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_147
timestamp 1679235063
transform 1 0 14628 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_163
timestamp 1679235063
transform 1 0 16100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_187
timestamp 1679235063
transform 1 0 18308 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1679235063
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_238
timestamp 1679235063
transform 1 0 23000 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_259
timestamp 1679235063
transform 1 0 24932 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_284
timestamp 1679235063
transform 1 0 27232 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_295
timestamp 1679235063
transform 1 0 28244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1679235063
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1679235063
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_377
timestamp 1679235063
transform 1 0 35788 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_19
timestamp 1679235063
transform 1 0 2852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_31
timestamp 1679235063
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_43
timestamp 1679235063
transform 1 0 5060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1679235063
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_60
timestamp 1679235063
transform 1 0 6624 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_68
timestamp 1679235063
transform 1 0 7360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_86
timestamp 1679235063
transform 1 0 9016 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_94
timestamp 1679235063
transform 1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_102
timestamp 1679235063
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1679235063
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_123
timestamp 1679235063
transform 1 0 12420 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_147
timestamp 1679235063
transform 1 0 14628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_151
timestamp 1679235063
transform 1 0 14996 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_159
timestamp 1679235063
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1679235063
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_178
timestamp 1679235063
transform 1 0 17480 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_200
timestamp 1679235063
transform 1 0 19504 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1679235063
transform 1 0 20884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1679235063
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_236
timestamp 1679235063
transform 1 0 22816 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1679235063
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_261
timestamp 1679235063
transform 1 0 25116 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_266
timestamp 1679235063
transform 1 0 25576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1679235063
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_281
timestamp 1679235063
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_287
timestamp 1679235063
transform 1 0 27508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_300
timestamp 1679235063
transform 1 0 28704 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_309
timestamp 1679235063
transform 1 0 29532 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_321
timestamp 1679235063
transform 1 0 30636 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1679235063
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1679235063
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1679235063
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1679235063
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1679235063
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1679235063
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1679235063
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1679235063
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_45
timestamp 1679235063
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_52
timestamp 1679235063
transform 1 0 5888 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_64
timestamp 1679235063
transform 1 0 6992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1679235063
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1679235063
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_102
timestamp 1679235063
transform 1 0 10488 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_106
timestamp 1679235063
transform 1 0 10856 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_123
timestamp 1679235063
transform 1 0 12420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1679235063
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1679235063
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1679235063
transform 1 0 14352 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_155
timestamp 1679235063
transform 1 0 15364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_167
timestamp 1679235063
transform 1 0 16468 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_179
timestamp 1679235063
transform 1 0 17572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1679235063
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1679235063
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_232
timestamp 1679235063
transform 1 0 22448 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_240
timestamp 1679235063
transform 1 0 23184 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1679235063
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_265
timestamp 1679235063
transform 1 0 25484 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_273
timestamp 1679235063
transform 1 0 26220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_285
timestamp 1679235063
transform 1 0 27324 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_297
timestamp 1679235063
transform 1 0 28428 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1679235063
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1679235063
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_321
timestamp 1679235063
transform 1 0 30636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_325
timestamp 1679235063
transform 1 0 31004 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1679235063
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_345
timestamp 1679235063
transform 1 0 32844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_353
timestamp 1679235063
transform 1 0 33580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 1679235063
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1679235063
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1679235063
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_377
timestamp 1679235063
transform 1 0 35788 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1679235063
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1679235063
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1679235063
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_51
timestamp 1679235063
transform 1 0 5796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_70
timestamp 1679235063
transform 1 0 7544 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_75
timestamp 1679235063
transform 1 0 8004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_87
timestamp 1679235063
transform 1 0 9108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_95
timestamp 1679235063
transform 1 0 9844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1679235063
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1679235063
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp 1679235063
transform 1 0 12052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_138
timestamp 1679235063
transform 1 0 13800 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_151
timestamp 1679235063
transform 1 0 14996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1679235063
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1679235063
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_185
timestamp 1679235063
transform 1 0 18124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_197
timestamp 1679235063
transform 1 0 19228 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_203
timestamp 1679235063
transform 1 0 19780 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_207
timestamp 1679235063
transform 1 0 20148 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_215
timestamp 1679235063
transform 1 0 20884 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_233
timestamp 1679235063
transform 1 0 22540 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_256
timestamp 1679235063
transform 1 0 24656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1679235063
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1679235063
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_287
timestamp 1679235063
transform 1 0 27508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_299
timestamp 1679235063
transform 1 0 28612 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_303
timestamp 1679235063
transform 1 0 28980 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_307
timestamp 1679235063
transform 1 0 29348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_318
timestamp 1679235063
transform 1 0 30360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_323
timestamp 1679235063
transform 1 0 30820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_328
timestamp 1679235063
transform 1 0 31280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_344
timestamp 1679235063
transform 1 0 32752 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_368
timestamp 1679235063
transform 1 0 34960 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_380
timestamp 1679235063
transform 1 0 36064 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_384
timestamp 1679235063
transform 1 0 36432 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1679235063
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_35
timestamp 1679235063
transform 1 0 4324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1679235063
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1679235063
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1679235063
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_103
timestamp 1679235063
transform 1 0 10580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_112
timestamp 1679235063
transform 1 0 11408 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_116
timestamp 1679235063
transform 1 0 11776 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_130
timestamp 1679235063
transform 1 0 13064 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_151
timestamp 1679235063
transform 1 0 14996 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_155
timestamp 1679235063
transform 1 0 15364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_167
timestamp 1679235063
transform 1 0 16468 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_183
timestamp 1679235063
transform 1 0 17940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_226
timestamp 1679235063
transform 1 0 21896 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_232
timestamp 1679235063
transform 1 0 22448 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp 1679235063
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_270
timestamp 1679235063
transform 1 0 25944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_278
timestamp 1679235063
transform 1 0 26680 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_292
timestamp 1679235063
transform 1 0 27968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_299
timestamp 1679235063
transform 1 0 28612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_303
timestamp 1679235063
transform 1 0 28980 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1679235063
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_345
timestamp 1679235063
transform 1 0 32844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_358
timestamp 1679235063
transform 1 0 34040 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1679235063
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1679235063
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1679235063
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_68
timestamp 1679235063
transform 1 0 7360 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_80
timestamp 1679235063
transform 1 0 8464 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1679235063
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_102
timestamp 1679235063
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1679235063
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1679235063
transform 1 0 12236 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_130
timestamp 1679235063
transform 1 0 13064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1679235063
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_176
timestamp 1679235063
transform 1 0 17296 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_188
timestamp 1679235063
transform 1 0 18400 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_200
timestamp 1679235063
transform 1 0 19504 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_212
timestamp 1679235063
transform 1 0 20608 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_216
timestamp 1679235063
transform 1 0 20976 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1679235063
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_239
timestamp 1679235063
transform 1 0 23092 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_245
timestamp 1679235063
transform 1 0 23644 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_260
timestamp 1679235063
transform 1 0 25024 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_272
timestamp 1679235063
transform 1 0 26128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1679235063
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_310
timestamp 1679235063
transform 1 0 29624 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_322
timestamp 1679235063
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1679235063
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_346
timestamp 1679235063
transform 1 0 32936 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_354
timestamp 1679235063
transform 1 0 33672 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_365
timestamp 1679235063
transform 1 0 34684 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_377
timestamp 1679235063
transform 1 0 35788 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1679235063
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1679235063
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_35
timestamp 1679235063
transform 1 0 4324 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_42
timestamp 1679235063
transform 1 0 4968 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_54
timestamp 1679235063
transform 1 0 6072 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_66
timestamp 1679235063
transform 1 0 7176 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_78
timestamp 1679235063
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_97
timestamp 1679235063
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_104
timestamp 1679235063
transform 1 0 10672 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_115
timestamp 1679235063
transform 1 0 11684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_127
timestamp 1679235063
transform 1 0 12788 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1679235063
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_150
timestamp 1679235063
transform 1 0 14904 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_174
timestamp 1679235063
transform 1 0 17112 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1679235063
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_209
timestamp 1679235063
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_217
timestamp 1679235063
transform 1 0 21068 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1679235063
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1679235063
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_277
timestamp 1679235063
transform 1 0 26588 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_285
timestamp 1679235063
transform 1 0 27324 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_299
timestamp 1679235063
transform 1 0 28612 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1679235063
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_309
timestamp 1679235063
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1679235063
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1679235063
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1679235063
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1679235063
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1679235063
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1679235063
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_377
timestamp 1679235063
transform 1 0 35788 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1679235063
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1679235063
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_39
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1679235063
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1679235063
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_62
timestamp 1679235063
transform 1 0 6808 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_74
timestamp 1679235063
transform 1 0 7912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_82
timestamp 1679235063
transform 1 0 8648 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_98
timestamp 1679235063
transform 1 0 10120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1679235063
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_119
timestamp 1679235063
transform 1 0 12052 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_131
timestamp 1679235063
transform 1 0 13156 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_143
timestamp 1679235063
transform 1 0 14260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_151
timestamp 1679235063
transform 1 0 14996 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_155
timestamp 1679235063
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1679235063
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_173
timestamp 1679235063
transform 1 0 17020 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1679235063
transform 1 0 17756 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_199
timestamp 1679235063
transform 1 0 19412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_211
timestamp 1679235063
transform 1 0 20516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1679235063
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_241
timestamp 1679235063
transform 1 0 23276 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1679235063
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1679235063
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1679235063
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1679235063
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_305
timestamp 1679235063
transform 1 0 29164 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_311
timestamp 1679235063
transform 1 0 29716 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_325
timestamp 1679235063
transform 1 0 31004 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_333
timestamp 1679235063
transform 1 0 31740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_345
timestamp 1679235063
transform 1 0 32844 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_364
timestamp 1679235063
transform 1 0 34592 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_376
timestamp 1679235063
transform 1 0 35696 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_384
timestamp 1679235063
transform 1 0 36432 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_9
timestamp 1679235063
transform 1 0 1932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1679235063
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1679235063
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_46
timestamp 1679235063
transform 1 0 5336 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1679235063
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1679235063
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_95
timestamp 1679235063
transform 1 0 9844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_107
timestamp 1679235063
transform 1 0 10948 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_127
timestamp 1679235063
transform 1 0 12788 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_133
timestamp 1679235063
transform 1 0 13340 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1679235063
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_144
timestamp 1679235063
transform 1 0 14352 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_156
timestamp 1679235063
transform 1 0 15456 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_168
timestamp 1679235063
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_179
timestamp 1679235063
transform 1 0 17572 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_188
timestamp 1679235063
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_221
timestamp 1679235063
transform 1 0 21436 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_230
timestamp 1679235063
transform 1 0 22264 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1679235063
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_273
timestamp 1679235063
transform 1 0 26220 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_279
timestamp 1679235063
transform 1 0 26772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_292
timestamp 1679235063
transform 1 0 27968 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_298
timestamp 1679235063
transform 1 0 28520 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1679235063
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1679235063
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_309
timestamp 1679235063
transform 1 0 29532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_336
timestamp 1679235063
transform 1 0 32016 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1679235063
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_369
timestamp 1679235063
transform 1 0 35052 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_381
timestamp 1679235063
transform 1 0 36156 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1679235063
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1679235063
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_39
timestamp 1679235063
transform 1 0 4692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_47
timestamp 1679235063
transform 1 0 5428 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1679235063
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_65
timestamp 1679235063
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_70
timestamp 1679235063
transform 1 0 7544 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_82
timestamp 1679235063
transform 1 0 8648 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_94
timestamp 1679235063
transform 1 0 9752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1679235063
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1679235063
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_142
timestamp 1679235063
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_154
timestamp 1679235063
transform 1 0 15272 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_162
timestamp 1679235063
transform 1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_185
timestamp 1679235063
transform 1 0 18124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_197
timestamp 1679235063
transform 1 0 19228 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_209
timestamp 1679235063
transform 1 0 20332 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_217
timestamp 1679235063
transform 1 0 21068 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1679235063
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_229
timestamp 1679235063
transform 1 0 22172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_241
timestamp 1679235063
transform 1 0 23276 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1679235063
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_287
timestamp 1679235063
transform 1 0 27508 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_311
timestamp 1679235063
transform 1 0 29716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_323
timestamp 1679235063
transform 1 0 30820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_337
timestamp 1679235063
transform 1 0 32108 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_350
timestamp 1679235063
transform 1 0 33304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_366
timestamp 1679235063
transform 1 0 34776 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_384
timestamp 1679235063
transform 1 0 36432 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1679235063
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1679235063
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1679235063
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1679235063
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_71
timestamp 1679235063
transform 1 0 7636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1679235063
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp 1679235063
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_94
timestamp 1679235063
transform 1 0 9752 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_106
timestamp 1679235063
transform 1 0 10856 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_122
timestamp 1679235063
transform 1 0 12328 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_134
timestamp 1679235063
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_154
timestamp 1679235063
transform 1 0 15272 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1679235063
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_179
timestamp 1679235063
transform 1 0 17572 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_187
timestamp 1679235063
transform 1 0 18308 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_218
timestamp 1679235063
transform 1 0 21160 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_226
timestamp 1679235063
transform 1 0 21896 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_234
timestamp 1679235063
transform 1 0 22632 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_238
timestamp 1679235063
transform 1 0 23000 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1679235063
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_265
timestamp 1679235063
transform 1 0 25484 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1679235063
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_289
timestamp 1679235063
transform 1 0 27692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_302
timestamp 1679235063
transform 1 0 28888 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1679235063
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_321
timestamp 1679235063
transform 1 0 30636 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_329
timestamp 1679235063
transform 1 0 31372 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_339
timestamp 1679235063
transform 1 0 32292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_351
timestamp 1679235063
transform 1 0 33396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1679235063
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_365
timestamp 1679235063
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_372
timestamp 1679235063
transform 1 0 35328 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_380
timestamp 1679235063
transform 1 0 36064 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1679235063
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_27
timestamp 1679235063
transform 1 0 3588 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_42
timestamp 1679235063
transform 1 0 4968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1679235063
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 1679235063
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_82
timestamp 1679235063
transform 1 0 8648 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1679235063
transform 1 0 9200 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_95
timestamp 1679235063
transform 1 0 9844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1679235063
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_127
timestamp 1679235063
transform 1 0 12788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_145
timestamp 1679235063
transform 1 0 14444 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_153
timestamp 1679235063
transform 1 0 15180 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1679235063
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_196
timestamp 1679235063
transform 1 0 19136 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_208
timestamp 1679235063
transform 1 0 20240 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1679235063
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_240
timestamp 1679235063
transform 1 0 23184 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_256
timestamp 1679235063
transform 1 0 24656 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_268
timestamp 1679235063
transform 1 0 25760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1679235063
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1679235063
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1679235063
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_341
timestamp 1679235063
transform 1 0 32476 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_357
timestamp 1679235063
transform 1 0 33948 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_365
timestamp 1679235063
transform 1 0 34684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_384
timestamp 1679235063
transform 1 0 36432 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1679235063
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1679235063
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_37
timestamp 1679235063
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_40
timestamp 1679235063
transform 1 0 4784 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_54
timestamp 1679235063
transform 1 0 6072 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_62
timestamp 1679235063
transform 1 0 6808 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_70
timestamp 1679235063
transform 1 0 7544 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1679235063
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1679235063
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_117
timestamp 1679235063
transform 1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_126
timestamp 1679235063
transform 1 0 12696 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1679235063
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_156
timestamp 1679235063
transform 1 0 15456 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_164
timestamp 1679235063
transform 1 0 16192 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_176
timestamp 1679235063
transform 1 0 17296 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1679235063
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_209
timestamp 1679235063
transform 1 0 20332 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_217
timestamp 1679235063
transform 1 0 21068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_239
timestamp 1679235063
transform 1 0 23092 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_243
timestamp 1679235063
transform 1 0 23460 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_269
timestamp 1679235063
transform 1 0 25852 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_281
timestamp 1679235063
transform 1 0 26956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_291
timestamp 1679235063
transform 1 0 27876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_303
timestamp 1679235063
transform 1 0 28980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_318
timestamp 1679235063
transform 1 0 30360 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_326
timestamp 1679235063
transform 1 0 31096 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_331
timestamp 1679235063
transform 1 0 31556 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_338
timestamp 1679235063
transform 1 0 32200 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_355
timestamp 1679235063
transform 1 0 33764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1679235063
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_371
timestamp 1679235063
transform 1 0 35236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_383
timestamp 1679235063
transform 1 0 36340 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1679235063
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_21
timestamp 1679235063
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_33
timestamp 1679235063
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1679235063
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_67
timestamp 1679235063
transform 1 0 7268 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_86
timestamp 1679235063
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_95
timestamp 1679235063
transform 1 0 9844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1679235063
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1679235063
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_125
timestamp 1679235063
transform 1 0 12604 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1679235063
transform 1 0 14444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_149
timestamp 1679235063
transform 1 0 14812 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1679235063
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_172
timestamp 1679235063
transform 1 0 16928 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1679235063
transform 1 0 18032 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_192
timestamp 1679235063
transform 1 0 18768 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_204
timestamp 1679235063
transform 1 0 19872 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_216
timestamp 1679235063
transform 1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1679235063
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1679235063
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_261
timestamp 1679235063
transform 1 0 25116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_293
timestamp 1679235063
transform 1 0 28060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_301
timestamp 1679235063
transform 1 0 28796 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_318
timestamp 1679235063
transform 1 0 30360 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_330
timestamp 1679235063
transform 1 0 31464 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_337
timestamp 1679235063
transform 1 0 32108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_343
timestamp 1679235063
transform 1 0 32660 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_359
timestamp 1679235063
transform 1 0 34132 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_363
timestamp 1679235063
transform 1 0 34500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_380
timestamp 1679235063
transform 1 0 36064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_384
timestamp 1679235063
transform 1 0 36432 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1679235063
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1679235063
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_35
timestamp 1679235063
transform 1 0 4324 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_48
timestamp 1679235063
transform 1 0 5520 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_52
timestamp 1679235063
transform 1 0 5888 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_65
timestamp 1679235063
transform 1 0 7084 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_73
timestamp 1679235063
transform 1 0 7820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1679235063
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1679235063
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_103
timestamp 1679235063
transform 1 0 10580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_111
timestamp 1679235063
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_119
timestamp 1679235063
transform 1 0 12052 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_131
timestamp 1679235063
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1679235063
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_153
timestamp 1679235063
transform 1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1679235063
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1679235063
transform 1 0 20056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_211
timestamp 1679235063
transform 1 0 20516 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_222
timestamp 1679235063
transform 1 0 21528 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_239
timestamp 1679235063
transform 1 0 23092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1679235063
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_262
timestamp 1679235063
transform 1 0 25208 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_277
timestamp 1679235063
transform 1 0 26588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_284
timestamp 1679235063
transform 1 0 27232 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_292
timestamp 1679235063
transform 1 0 27968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_305
timestamp 1679235063
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1679235063
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_317
timestamp 1679235063
transform 1 0 30268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_322
timestamp 1679235063
transform 1 0 30728 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1679235063
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_345
timestamp 1679235063
transform 1 0 32844 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1679235063
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1679235063
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1679235063
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_377
timestamp 1679235063
transform 1 0 35788 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_15
timestamp 1679235063
transform 1 0 2484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_21
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_38
timestamp 1679235063
transform 1 0 4600 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1679235063
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_75
timestamp 1679235063
transform 1 0 8004 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_82
timestamp 1679235063
transform 1 0 8648 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_92
timestamp 1679235063
transform 1 0 9568 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1679235063
transform 1 0 12420 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_151
timestamp 1679235063
transform 1 0 14996 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1679235063
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1679235063
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1679235063
transform 1 0 17756 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_199
timestamp 1679235063
transform 1 0 19412 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_243
timestamp 1679235063
transform 1 0 23460 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_266
timestamp 1679235063
transform 1 0 25576 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_270
timestamp 1679235063
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1679235063
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_284
timestamp 1679235063
transform 1 0 27232 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_292
timestamp 1679235063
transform 1 0 27968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_307
timestamp 1679235063
transform 1 0 29348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_318
timestamp 1679235063
transform 1 0 30360 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1679235063
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_345
timestamp 1679235063
transform 1 0 32844 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_357
timestamp 1679235063
transform 1 0 33948 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_369
timestamp 1679235063
transform 1 0 35052 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_381
timestamp 1679235063
transform 1 0 36156 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1679235063
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1679235063
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_32
timestamp 1679235063
transform 1 0 4048 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_40
timestamp 1679235063
transform 1 0 4784 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_59
timestamp 1679235063
transform 1 0 6532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1679235063
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1679235063
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_93
timestamp 1679235063
transform 1 0 9660 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_100
timestamp 1679235063
transform 1 0 10304 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_105
timestamp 1679235063
transform 1 0 10764 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 1679235063
transform 1 0 11316 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_123
timestamp 1679235063
transform 1 0 12420 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1679235063
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_146
timestamp 1679235063
transform 1 0 14536 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1679235063
transform 1 0 15272 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_168
timestamp 1679235063
transform 1 0 16560 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_180
timestamp 1679235063
transform 1 0 17664 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_186
timestamp 1679235063
transform 1 0 18216 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1679235063
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_206
timestamp 1679235063
transform 1 0 20056 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_219
timestamp 1679235063
transform 1 0 21252 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_227
timestamp 1679235063
transform 1 0 21988 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_239
timestamp 1679235063
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1679235063
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_257
timestamp 1679235063
transform 1 0 24748 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_263
timestamp 1679235063
transform 1 0 25300 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_292
timestamp 1679235063
transform 1 0 27968 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_304
timestamp 1679235063
transform 1 0 29072 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_321
timestamp 1679235063
transform 1 0 30636 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_343
timestamp 1679235063
transform 1 0 32660 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1679235063
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1679235063
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_377
timestamp 1679235063
transform 1 0 35788 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1679235063
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1679235063
transform 1 0 3588 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_31
timestamp 1679235063
transform 1 0 3956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_41
timestamp 1679235063
transform 1 0 4876 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_45
timestamp 1679235063
transform 1 0 5244 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_49
timestamp 1679235063
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1679235063
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_66
timestamp 1679235063
transform 1 0 7176 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_72
timestamp 1679235063
transform 1 0 7728 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_85
timestamp 1679235063
transform 1 0 8924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_97
timestamp 1679235063
transform 1 0 10028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1679235063
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1679235063
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_137
timestamp 1679235063
transform 1 0 13708 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_150
timestamp 1679235063
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_172
timestamp 1679235063
transform 1 0 16928 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_188
timestamp 1679235063
transform 1 0 18400 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_200
timestamp 1679235063
transform 1 0 19504 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_212
timestamp 1679235063
transform 1 0 20608 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_234
timestamp 1679235063
transform 1 0 22632 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_246
timestamp 1679235063
transform 1 0 23736 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_258
timestamp 1679235063
transform 1 0 24840 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_267
timestamp 1679235063
transform 1 0 25668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1679235063
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_281
timestamp 1679235063
transform 1 0 26956 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_291
timestamp 1679235063
transform 1 0 27876 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_303
timestamp 1679235063
transform 1 0 28980 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_315
timestamp 1679235063
transform 1 0 30084 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_327
timestamp 1679235063
transform 1 0 31188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_331
timestamp 1679235063
transform 1 0 31556 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1679235063
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1679235063
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1679235063
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1679235063
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_15
timestamp 1679235063
transform 1 0 2484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_22
timestamp 1679235063
transform 1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_37
timestamp 1679235063
transform 1 0 4508 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_49
timestamp 1679235063
transform 1 0 5612 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_61
timestamp 1679235063
transform 1 0 6716 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_73
timestamp 1679235063
transform 1 0 7820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1679235063
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_90
timestamp 1679235063
transform 1 0 9384 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_114
timestamp 1679235063
transform 1 0 11592 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_126
timestamp 1679235063
transform 1 0 12696 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1679235063
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_153
timestamp 1679235063
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_161
timestamp 1679235063
transform 1 0 15916 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_172
timestamp 1679235063
transform 1 0 16928 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_184
timestamp 1679235063
transform 1 0 18032 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_190
timestamp 1679235063
transform 1 0 18584 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_209
timestamp 1679235063
transform 1 0 20332 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_229
timestamp 1679235063
transform 1 0 22172 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1679235063
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_271
timestamp 1679235063
transform 1 0 26036 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_279
timestamp 1679235063
transform 1 0 26772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_303
timestamp 1679235063
transform 1 0 28980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1679235063
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1679235063
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_320
timestamp 1679235063
transform 1 0 30544 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_332
timestamp 1679235063
transform 1 0 31648 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_344
timestamp 1679235063
transform 1 0 32752 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_356
timestamp 1679235063
transform 1 0 33856 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1679235063
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_377
timestamp 1679235063
transform 1 0 35788 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_7
timestamp 1679235063
transform 1 0 1748 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_13
timestamp 1679235063
transform 1 0 2300 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 1679235063
transform 1 0 3864 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_34
timestamp 1679235063
transform 1 0 4232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1679235063
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1679235063
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_60
timestamp 1679235063
transform 1 0 6624 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_72
timestamp 1679235063
transform 1 0 7728 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_79
timestamp 1679235063
transform 1 0 8372 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_83
timestamp 1679235063
transform 1 0 8740 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_103
timestamp 1679235063
transform 1 0 10580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1679235063
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_140
timestamp 1679235063
transform 1 0 13984 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_152
timestamp 1679235063
transform 1 0 15088 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_157
timestamp 1679235063
transform 1 0 15548 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1679235063
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_169
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_177
timestamp 1679235063
transform 1 0 17388 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_183
timestamp 1679235063
transform 1 0 17940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_187
timestamp 1679235063
transform 1 0 18308 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_204
timestamp 1679235063
transform 1 0 19872 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1679235063
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_233
timestamp 1679235063
transform 1 0 22540 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_253
timestamp 1679235063
transform 1 0 24380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_265
timestamp 1679235063
transform 1 0 25484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1679235063
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1679235063
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_293
timestamp 1679235063
transform 1 0 28060 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_301
timestamp 1679235063
transform 1 0 28796 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_321
timestamp 1679235063
transform 1 0 30636 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_364
timestamp 1679235063
transform 1 0 34592 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_376
timestamp 1679235063
transform 1 0 35696 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_384
timestamp 1679235063
transform 1 0 36432 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1679235063
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1679235063
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 1679235063
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_49
timestamp 1679235063
transform 1 0 5612 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_88
timestamp 1679235063
transform 1 0 9200 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_100
timestamp 1679235063
transform 1 0 10304 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1679235063
transform 1 0 11408 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_128
timestamp 1679235063
transform 1 0 12880 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_149
timestamp 1679235063
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_178
timestamp 1679235063
transform 1 0 17480 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1679235063
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1679235063
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1679235063
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_233
timestamp 1679235063
transform 1 0 22540 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 1679235063
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_275
timestamp 1679235063
transform 1 0 26404 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_287
timestamp 1679235063
transform 1 0 27508 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_298
timestamp 1679235063
transform 1 0 28520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1679235063
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1679235063
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_329
timestamp 1679235063
transform 1 0 31372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_347
timestamp 1679235063
transform 1 0 33028 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_368
timestamp 1679235063
transform 1 0 34960 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_380
timestamp 1679235063
transform 1 0 36064 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_384
timestamp 1679235063
transform 1 0 36432 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1679235063
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_11
timestamp 1679235063
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_23
timestamp 1679235063
transform 1 0 3220 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_34
timestamp 1679235063
transform 1 0 4232 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_45
timestamp 1679235063
transform 1 0 5244 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_51
timestamp 1679235063
transform 1 0 5796 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_67
timestamp 1679235063
transform 1 0 7268 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_79
timestamp 1679235063
transform 1 0 8372 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1679235063
transform 1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1679235063
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_129
timestamp 1679235063
transform 1 0 12972 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_151
timestamp 1679235063
transform 1 0 14996 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_163
timestamp 1679235063
transform 1 0 16100 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_185
timestamp 1679235063
transform 1 0 18124 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_202
timestamp 1679235063
transform 1 0 19688 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_214
timestamp 1679235063
transform 1 0 20792 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1679235063
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1679235063
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_233
timestamp 1679235063
transform 1 0 22540 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_245
timestamp 1679235063
transform 1 0 23644 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_257
timestamp 1679235063
transform 1 0 24748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_269
timestamp 1679235063
transform 1 0 25852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1679235063
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_281
timestamp 1679235063
transform 1 0 26956 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_301
timestamp 1679235063
transform 1 0 28796 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_307
timestamp 1679235063
transform 1 0 29348 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_311
timestamp 1679235063
transform 1 0 29716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_323
timestamp 1679235063
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1679235063
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_346
timestamp 1679235063
transform 1 0 32936 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_352
timestamp 1679235063
transform 1 0 33488 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_362
timestamp 1679235063
transform 1 0 34408 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_374
timestamp 1679235063
transform 1 0 35512 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1679235063
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1679235063
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_45
timestamp 1679235063
transform 1 0 5244 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_74
timestamp 1679235063
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1679235063
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1679235063
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1679235063
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1679235063
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_150
timestamp 1679235063
transform 1 0 14904 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_162
timestamp 1679235063
transform 1 0 16008 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_170
timestamp 1679235063
transform 1 0 16744 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_182
timestamp 1679235063
transform 1 0 17848 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1679235063
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1679235063
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_229
timestamp 1679235063
transform 1 0 22172 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1679235063
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_262
timestamp 1679235063
transform 1 0 25208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_266
timestamp 1679235063
transform 1 0 25576 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_295
timestamp 1679235063
transform 1 0 28244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1679235063
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_325
timestamp 1679235063
transform 1 0 31004 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_337
timestamp 1679235063
transform 1 0 32108 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_349
timestamp 1679235063
transform 1 0 33212 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_355
timestamp 1679235063
transform 1 0 33764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1679235063
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1679235063
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_377
timestamp 1679235063
transform 1 0 35788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1679235063
transform 1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_22
timestamp 1679235063
transform 1 0 3128 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_34
timestamp 1679235063
transform 1 0 4232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_78
timestamp 1679235063
transform 1 0 8280 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_84
timestamp 1679235063
transform 1 0 8832 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_88
timestamp 1679235063
transform 1 0 9200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_120
timestamp 1679235063
transform 1 0 12144 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1679235063
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_156
timestamp 1679235063
transform 1 0 15456 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_194
timestamp 1679235063
transform 1 0 18952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1679235063
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1679235063
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_234
timestamp 1679235063
transform 1 0 22632 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_275
timestamp 1679235063
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1679235063
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_301
timestamp 1679235063
transform 1 0 28796 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1679235063
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_317
timestamp 1679235063
transform 1 0 30268 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_330
timestamp 1679235063
transform 1 0 31464 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_337
timestamp 1679235063
transform 1 0 32108 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_341
timestamp 1679235063
transform 1 0 32476 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_363
timestamp 1679235063
transform 1 0 34500 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1679235063
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1679235063
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1679235063
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_56
timestamp 1679235063
transform 1 0 6256 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_68
timestamp 1679235063
transform 1 0 7360 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1679235063
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_89
timestamp 1679235063
transform 1 0 9292 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_111
timestamp 1679235063
transform 1 0 11316 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_129
timestamp 1679235063
transform 1 0 12972 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1679235063
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp 1679235063
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1679235063
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1679235063
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_222
timestamp 1679235063
transform 1 0 21528 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_229
timestamp 1679235063
transform 1 0 22172 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_241
timestamp 1679235063
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1679235063
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_274
timestamp 1679235063
transform 1 0 26312 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_280
timestamp 1679235063
transform 1 0 26864 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1679235063
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_309
timestamp 1679235063
transform 1 0 29532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_321
timestamp 1679235063
transform 1 0 30636 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 1679235063
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_375
timestamp 1679235063
transform 1 0 35604 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_383
timestamp 1679235063
transform 1 0 36340 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_9
timestamp 1679235063
transform 1 0 1932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_24
timestamp 1679235063
transform 1 0 3312 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_42
timestamp 1679235063
transform 1 0 4968 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1679235063
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_69
timestamp 1679235063
transform 1 0 7452 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_91
timestamp 1679235063
transform 1 0 9476 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_103
timestamp 1679235063
transform 1 0 10580 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1679235063
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_149
timestamp 1679235063
transform 1 0 14812 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1679235063
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1679235063
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_179
timestamp 1679235063
transform 1 0 17572 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_185
timestamp 1679235063
transform 1 0 18124 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_198
timestamp 1679235063
transform 1 0 19320 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_204
timestamp 1679235063
transform 1 0 19872 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_209
timestamp 1679235063
transform 1 0 20332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1679235063
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_229
timestamp 1679235063
transform 1 0 22172 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_247
timestamp 1679235063
transform 1 0 23828 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_268
timestamp 1679235063
transform 1 0 25760 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1679235063
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_302
timestamp 1679235063
transform 1 0 28888 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_324
timestamp 1679235063
transform 1 0 30912 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_337
timestamp 1679235063
transform 1 0 32108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_345
timestamp 1679235063
transform 1 0 32844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_352
timestamp 1679235063
transform 1 0 33488 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_358
timestamp 1679235063
transform 1 0 34040 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_375
timestamp 1679235063
transform 1 0 35604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_383
timestamp 1679235063
transform 1 0 36340 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1679235063
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_11
timestamp 1679235063
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1679235063
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1679235063
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1679235063
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_53
timestamp 1679235063
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_63
timestamp 1679235063
transform 1 0 6900 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1679235063
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1679235063
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_101
timestamp 1679235063
transform 1 0 10396 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_108
timestamp 1679235063
transform 1 0 11040 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_120
timestamp 1679235063
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_132
timestamp 1679235063
transform 1 0 13248 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1679235063
transform 1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_174
timestamp 1679235063
transform 1 0 17112 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_186
timestamp 1679235063
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_203
timestamp 1679235063
transform 1 0 19780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_210
timestamp 1679235063
transform 1 0 20424 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_241
timestamp 1679235063
transform 1 0 23276 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1679235063
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1679235063
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1679235063
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_289
timestamp 1679235063
transform 1 0 27692 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_296
timestamp 1679235063
transform 1 0 28336 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1679235063
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_314
timestamp 1679235063
transform 1 0 29992 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_326
timestamp 1679235063
transform 1 0 31096 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_338
timestamp 1679235063
transform 1 0 32200 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_342
timestamp 1679235063
transform 1 0 32568 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_352
timestamp 1679235063
transform 1 0 33488 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_369
timestamp 1679235063
transform 1 0 35052 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_381
timestamp 1679235063
transform 1 0 36156 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_20
timestamp 1679235063
transform 1 0 2944 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_37
timestamp 1679235063
transform 1 0 4508 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1679235063
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1679235063
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_77
timestamp 1679235063
transform 1 0 8188 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_87
timestamp 1679235063
transform 1 0 9108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_93
timestamp 1679235063
transform 1 0 9660 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_101
timestamp 1679235063
transform 1 0 10396 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1679235063
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1679235063
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_138
timestamp 1679235063
transform 1 0 13800 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_149
timestamp 1679235063
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_153
timestamp 1679235063
transform 1 0 15180 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_157
timestamp 1679235063
transform 1 0 15548 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1679235063
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_191
timestamp 1679235063
transform 1 0 18676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_201
timestamp 1679235063
transform 1 0 19596 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_213
timestamp 1679235063
transform 1 0 20700 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1679235063
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_234
timestamp 1679235063
transform 1 0 22632 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_244
timestamp 1679235063
transform 1 0 23552 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_266
timestamp 1679235063
transform 1 0 25576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_270
timestamp 1679235063
transform 1 0 25944 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1679235063
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1679235063
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_281
timestamp 1679235063
transform 1 0 26956 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_291
timestamp 1679235063
transform 1 0 27876 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_306
timestamp 1679235063
transform 1 0 29256 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_327
timestamp 1679235063
transform 1 0 31188 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_353
timestamp 1679235063
transform 1 0 33580 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_365
timestamp 1679235063
transform 1 0 34684 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_377
timestamp 1679235063
transform 1 0 35788 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_11
timestamp 1679235063
transform 1 0 2116 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_21
timestamp 1679235063
transform 1 0 3036 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_59
timestamp 1679235063
transform 1 0 6532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_74
timestamp 1679235063
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1679235063
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_101
timestamp 1679235063
transform 1 0 10396 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_122
timestamp 1679235063
transform 1 0 12328 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_166
timestamp 1679235063
transform 1 0 16376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1679235063
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_217
timestamp 1679235063
transform 1 0 21068 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_229
timestamp 1679235063
transform 1 0 22172 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_241
timestamp 1679235063
transform 1 0 23276 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1679235063
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1679235063
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_312
timestamp 1679235063
transform 1 0 29808 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_316
timestamp 1679235063
transform 1 0 30176 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_341
timestamp 1679235063
transform 1 0 32476 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_347
timestamp 1679235063
transform 1 0 33028 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1679235063
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_377
timestamp 1679235063
transform 1 0 35788 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1679235063
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_33
timestamp 1679235063
transform 1 0 4140 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_61
timestamp 1679235063
transform 1 0 6716 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_76
timestamp 1679235063
transform 1 0 8096 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_88
timestamp 1679235063
transform 1 0 9200 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1679235063
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1679235063
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1679235063
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_119
timestamp 1679235063
transform 1 0 12052 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_131
timestamp 1679235063
transform 1 0 13156 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_143
timestamp 1679235063
transform 1 0 14260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_155
timestamp 1679235063
transform 1 0 15364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_169
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_189
timestamp 1679235063
transform 1 0 18492 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_201
timestamp 1679235063
transform 1 0 19596 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_207
timestamp 1679235063
transform 1 0 20148 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1679235063
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_234
timestamp 1679235063
transform 1 0 22632 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_238
timestamp 1679235063
transform 1 0 23000 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_264
timestamp 1679235063
transform 1 0 25392 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1679235063
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1679235063
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_293
timestamp 1679235063
transform 1 0 28060 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_304
timestamp 1679235063
transform 1 0 29072 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_316
timestamp 1679235063
transform 1 0 30176 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_328
timestamp 1679235063
transform 1 0 31280 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_337
timestamp 1679235063
transform 1 0 32108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_345
timestamp 1679235063
transform 1 0 32844 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_351
timestamp 1679235063
transform 1 0 33396 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_363
timestamp 1679235063
transform 1 0 34500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_375
timestamp 1679235063
transform 1 0 35604 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_383
timestamp 1679235063
transform 1 0 36340 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1679235063
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1679235063
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_37
timestamp 1679235063
transform 1 0 4508 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1679235063
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_53
timestamp 1679235063
transform 1 0 5980 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_59
timestamp 1679235063
transform 1 0 6532 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_66
timestamp 1679235063
transform 1 0 7176 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_78
timestamp 1679235063
transform 1 0 8280 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_36_85
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_107
timestamp 1679235063
transform 1 0 10948 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_111
timestamp 1679235063
transform 1 0 11316 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1679235063
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_141
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_151
timestamp 1679235063
transform 1 0 14996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_163
timestamp 1679235063
transform 1 0 16100 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_185
timestamp 1679235063
transform 1 0 18124 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1679235063
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_209
timestamp 1679235063
transform 1 0 20332 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_236
timestamp 1679235063
transform 1 0 22816 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1679235063
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_261
timestamp 1679235063
transform 1 0 25116 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_282
timestamp 1679235063
transform 1 0 27048 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_294
timestamp 1679235063
transform 1 0 28152 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1679235063
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_309
timestamp 1679235063
transform 1 0 29532 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_315
timestamp 1679235063
transform 1 0 30084 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_335
timestamp 1679235063
transform 1 0 31924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_355
timestamp 1679235063
transform 1 0 33764 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1679235063
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1679235063
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_377
timestamp 1679235063
transform 1 0 35788 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_7
timestamp 1679235063
transform 1 0 1748 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_19
timestamp 1679235063
transform 1 0 2852 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_31
timestamp 1679235063
transform 1 0 3956 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 1679235063
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_69
timestamp 1679235063
transform 1 0 7452 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_89
timestamp 1679235063
transform 1 0 9292 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_101
timestamp 1679235063
transform 1 0 10396 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_109
timestamp 1679235063
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_121
timestamp 1679235063
transform 1 0 12236 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1679235063
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1679235063
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_181
timestamp 1679235063
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1679235063
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1679235063
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1679235063
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1679235063
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_241
timestamp 1679235063
transform 1 0 23276 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_258
timestamp 1679235063
transform 1 0 24840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1679235063
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1679235063
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_281
timestamp 1679235063
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_289
timestamp 1679235063
transform 1 0 27692 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_301
timestamp 1679235063
transform 1 0 28796 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_313
timestamp 1679235063
transform 1 0 29900 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_321
timestamp 1679235063
transform 1 0 30636 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1679235063
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_341
timestamp 1679235063
transform 1 0 32476 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_358
timestamp 1679235063
transform 1 0 34040 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_370
timestamp 1679235063
transform 1 0 35144 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_382
timestamp 1679235063
transform 1 0 36248 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_15
timestamp 1679235063
transform 1 0 2484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_32
timestamp 1679235063
transform 1 0 4048 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_38
timestamp 1679235063
transform 1 0 4600 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_52
timestamp 1679235063
transform 1 0 5888 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_64
timestamp 1679235063
transform 1 0 6992 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_76
timestamp 1679235063
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1679235063
transform 1 0 9660 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_116
timestamp 1679235063
transform 1 0 11776 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_128
timestamp 1679235063
transform 1 0 12880 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_146
timestamp 1679235063
transform 1 0 14536 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_170
timestamp 1679235063
transform 1 0 16744 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_182
timestamp 1679235063
transform 1 0 17848 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_190
timestamp 1679235063
transform 1 0 18584 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1679235063
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_201
timestamp 1679235063
transform 1 0 19596 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_224
timestamp 1679235063
transform 1 0 21712 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_236
timestamp 1679235063
transform 1 0 22816 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_244
timestamp 1679235063
transform 1 0 23552 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 1679235063
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_262
timestamp 1679235063
transform 1 0 25208 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_268
timestamp 1679235063
transform 1 0 25760 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_278
timestamp 1679235063
transform 1 0 26680 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_337
timestamp 1679235063
transform 1 0 32108 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_346
timestamp 1679235063
transform 1 0 32936 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1679235063
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_377
timestamp 1679235063
transform 1 0 35788 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_10
timestamp 1679235063
transform 1 0 2024 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_36
timestamp 1679235063
transform 1 0 4416 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_48
timestamp 1679235063
transform 1 0 5520 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_71
timestamp 1679235063
transform 1 0 7636 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_83
timestamp 1679235063
transform 1 0 8740 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_89
timestamp 1679235063
transform 1 0 9292 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_121
timestamp 1679235063
transform 1 0 12236 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_146
timestamp 1679235063
transform 1 0 14536 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_190
timestamp 1679235063
transform 1 0 18584 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_233
timestamp 1679235063
transform 1 0 22540 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_251
timestamp 1679235063
transform 1 0 24196 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_255
timestamp 1679235063
transform 1 0 24564 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1679235063
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_318
timestamp 1679235063
transform 1 0 30360 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_330
timestamp 1679235063
transform 1 0 31464 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1679235063
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_353
timestamp 1679235063
transform 1 0 33580 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_365
timestamp 1679235063
transform 1 0 34684 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_377
timestamp 1679235063
transform 1 0 35788 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_19
timestamp 1679235063
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1679235063
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_37
timestamp 1679235063
transform 1 0 4508 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_61
timestamp 1679235063
transform 1 0 6716 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_69
timestamp 1679235063
transform 1 0 7452 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_77
timestamp 1679235063
transform 1 0 8188 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_101
timestamp 1679235063
transform 1 0 10396 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_107
timestamp 1679235063
transform 1 0 10948 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_114
timestamp 1679235063
transform 1 0 11592 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1679235063
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1679235063
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1679235063
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_177
timestamp 1679235063
transform 1 0 17388 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1679235063
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1679235063
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1679235063
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1679235063
transform 1 0 20700 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1679235063
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1679235063
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_298
timestamp 1679235063
transform 1 0 28520 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1679235063
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1679235063
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1679235063
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_333
timestamp 1679235063
transform 1 0 31740 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_339
timestamp 1679235063
transform 1 0 32292 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_343
timestamp 1679235063
transform 1 0 32660 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_355
timestamp 1679235063
transform 1 0 33764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1679235063
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1679235063
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_377
timestamp 1679235063
transform 1 0 35788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_13
timestamp 1679235063
transform 1 0 2300 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_21
timestamp 1679235063
transform 1 0 3036 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_40
timestamp 1679235063
transform 1 0 4784 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1679235063
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_64
timestamp 1679235063
transform 1 0 6992 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_75
timestamp 1679235063
transform 1 0 8004 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_87
timestamp 1679235063
transform 1 0 9108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_99
timestamp 1679235063
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1679235063
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_113
timestamp 1679235063
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_135
timestamp 1679235063
transform 1 0 13524 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_155
timestamp 1679235063
transform 1 0 15364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1679235063
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1679235063
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_188
timestamp 1679235063
transform 1 0 18400 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_200
timestamp 1679235063
transform 1 0 19504 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_210
timestamp 1679235063
transform 1 0 20424 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_214
timestamp 1679235063
transform 1 0 20792 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1679235063
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_225
timestamp 1679235063
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_244
timestamp 1679235063
transform 1 0 23552 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_254
timestamp 1679235063
transform 1 0 24472 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_266
timestamp 1679235063
transform 1 0 25576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1679235063
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_281
timestamp 1679235063
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_289
timestamp 1679235063
transform 1 0 27692 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_300
timestamp 1679235063
transform 1 0 28704 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_337
timestamp 1679235063
transform 1 0 32108 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_357
timestamp 1679235063
transform 1 0 33948 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_369
timestamp 1679235063
transform 1 0 35052 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_381
timestamp 1679235063
transform 1 0 36156 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_3
timestamp 1679235063
transform 1 0 1380 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1679235063
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_62
timestamp 1679235063
transform 1 0 6808 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1679235063
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1679235063
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1679235063
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_91
timestamp 1679235063
transform 1 0 9476 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_97
timestamp 1679235063
transform 1 0 10028 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_114
timestamp 1679235063
transform 1 0 11592 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_126
timestamp 1679235063
transform 1 0 12696 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1679235063
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1679235063
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_153
timestamp 1679235063
transform 1 0 15180 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_164
timestamp 1679235063
transform 1 0 16192 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_176
timestamp 1679235063
transform 1 0 17296 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_188
timestamp 1679235063
transform 1 0 18400 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_192
timestamp 1679235063
transform 1 0 18768 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_213
timestamp 1679235063
transform 1 0 20700 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_225
timestamp 1679235063
transform 1 0 21804 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_237
timestamp 1679235063
transform 1 0 22908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1679235063
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_253
timestamp 1679235063
transform 1 0 24380 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_263
timestamp 1679235063
transform 1 0 25300 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_269
timestamp 1679235063
transform 1 0 25852 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_286
timestamp 1679235063
transform 1 0 27416 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_304
timestamp 1679235063
transform 1 0 29072 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_341
timestamp 1679235063
transform 1 0 32476 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1679235063
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_377
timestamp 1679235063
transform 1 0 35788 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1679235063
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1679235063
transform 1 0 1748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_11
timestamp 1679235063
transform 1 0 2116 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_21
timestamp 1679235063
transform 1 0 3036 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_33
timestamp 1679235063
transform 1 0 4140 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_45
timestamp 1679235063
transform 1 0 5244 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1679235063
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_66
timestamp 1679235063
transform 1 0 7176 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_81
timestamp 1679235063
transform 1 0 8556 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_103
timestamp 1679235063
transform 1 0 10580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1679235063
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_121
timestamp 1679235063
transform 1 0 12236 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_132
timestamp 1679235063
transform 1 0 13248 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_137
timestamp 1679235063
transform 1 0 13708 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_143
timestamp 1679235063
transform 1 0 14260 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_196
timestamp 1679235063
transform 1 0 19136 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_213
timestamp 1679235063
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1679235063
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1679235063
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_245
timestamp 1679235063
transform 1 0 23644 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_249
timestamp 1679235063
transform 1 0 24012 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_266
timestamp 1679235063
transform 1 0 25576 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1679235063
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1679235063
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_290
timestamp 1679235063
transform 1 0 27784 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_294
timestamp 1679235063
transform 1 0 28152 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_306
timestamp 1679235063
transform 1 0 29256 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_318
timestamp 1679235063
transform 1 0 30360 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_326
timestamp 1679235063
transform 1 0 31096 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1679235063
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_358
timestamp 1679235063
transform 1 0 34040 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_370
timestamp 1679235063
transform 1 0 35144 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_382
timestamp 1679235063
transform 1 0 36248 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1679235063
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1679235063
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1679235063
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_29
timestamp 1679235063
transform 1 0 3772 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_42
timestamp 1679235063
transform 1 0 4968 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_54
timestamp 1679235063
transform 1 0 6072 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_66
timestamp 1679235063
transform 1 0 7176 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_78
timestamp 1679235063
transform 1 0 8280 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_95
timestamp 1679235063
transform 1 0 9844 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_102
timestamp 1679235063
transform 1 0 10488 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_114
timestamp 1679235063
transform 1 0 11592 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_133
timestamp 1679235063
transform 1 0 13340 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1679235063
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_150
timestamp 1679235063
transform 1 0 14904 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_162
timestamp 1679235063
transform 1 0 16008 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_170
timestamp 1679235063
transform 1 0 16744 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_182
timestamp 1679235063
transform 1 0 17848 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1679235063
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_197
timestamp 1679235063
transform 1 0 19228 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_214
timestamp 1679235063
transform 1 0 20792 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_229
timestamp 1679235063
transform 1 0 22172 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_236
timestamp 1679235063
transform 1 0 22816 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1679235063
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_256
timestamp 1679235063
transform 1 0 24656 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_268
timestamp 1679235063
transform 1 0 25760 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_280
timestamp 1679235063
transform 1 0 26864 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_292
timestamp 1679235063
transform 1 0 27968 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1679235063
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_309
timestamp 1679235063
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_344
timestamp 1679235063
transform 1 0 32752 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_356
timestamp 1679235063
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1679235063
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_377
timestamp 1679235063
transform 1 0 35788 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1679235063
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_10
timestamp 1679235063
transform 1 0 2024 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_37
timestamp 1679235063
transform 1 0 4508 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_49
timestamp 1679235063
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1679235063
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_57
timestamp 1679235063
transform 1 0 6348 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_81
timestamp 1679235063
transform 1 0 8556 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_93
timestamp 1679235063
transform 1 0 9660 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_116
timestamp 1679235063
transform 1 0 11776 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_120
timestamp 1679235063
transform 1 0 12144 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_124
timestamp 1679235063
transform 1 0 12512 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_152
timestamp 1679235063
transform 1 0 15088 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1679235063
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1679235063
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_175
timestamp 1679235063
transform 1 0 17204 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_195
timestamp 1679235063
transform 1 0 19044 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_201
timestamp 1679235063
transform 1 0 19596 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1679235063
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_209
timestamp 1679235063
transform 1 0 20332 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_214
timestamp 1679235063
transform 1 0 20792 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1679235063
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1679235063
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 1679235063
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_233
timestamp 1679235063
transform 1 0 22540 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_241
timestamp 1679235063
transform 1 0 23276 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_253
timestamp 1679235063
transform 1 0 24380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_263
timestamp 1679235063
transform 1 0 25300 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_269
timestamp 1679235063
transform 1 0 25852 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1679235063
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1679235063
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_293
timestamp 1679235063
transform 1 0 28060 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_299
timestamp 1679235063
transform 1 0 28612 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_307
timestamp 1679235063
transform 1 0 29348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_313
timestamp 1679235063
transform 1 0 29900 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1679235063
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1679235063
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_356
timestamp 1679235063
transform 1 0 33856 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_368
timestamp 1679235063
transform 1 0 34960 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_380
timestamp 1679235063
transform 1 0 36064 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_384
timestamp 1679235063
transform 1 0 36432 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_29
timestamp 1679235063
transform 1 0 3772 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1679235063
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_118
timestamp 1679235063
transform 1 0 11960 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_130
timestamp 1679235063
transform 1 0 13064 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1679235063
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_144
timestamp 1679235063
transform 1 0 14352 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_152
timestamp 1679235063
transform 1 0 15088 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_169
timestamp 1679235063
transform 1 0 16652 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_175
timestamp 1679235063
transform 1 0 17204 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1679235063
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_201
timestamp 1679235063
transform 1 0 19596 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_213
timestamp 1679235063
transform 1 0 20700 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_217
timestamp 1679235063
transform 1 0 21068 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_227
timestamp 1679235063
transform 1 0 21988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_239
timestamp 1679235063
transform 1 0 23092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1679235063
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_283
timestamp 1679235063
transform 1 0 27140 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_309
timestamp 1679235063
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_317
timestamp 1679235063
transform 1 0 30268 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_336
timestamp 1679235063
transform 1 0 32016 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_348
timestamp 1679235063
transform 1 0 33120 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1679235063
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1679235063
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_377
timestamp 1679235063
transform 1 0 35788 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1679235063
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1679235063
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_43
timestamp 1679235063
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1679235063
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1679235063
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_69
timestamp 1679235063
transform 1 0 7452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_77
timestamp 1679235063
transform 1 0 8188 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_95
timestamp 1679235063
transform 1 0 9844 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_107
timestamp 1679235063
transform 1 0 10948 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1679235063
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_113
timestamp 1679235063
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_121
timestamp 1679235063
transform 1 0 12236 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_154
timestamp 1679235063
transform 1 0 15272 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1679235063
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_199
timestamp 1679235063
transform 1 0 19412 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_204
timestamp 1679235063
transform 1 0 19872 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_218
timestamp 1679235063
transform 1 0 21160 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1679235063
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_241
timestamp 1679235063
transform 1 0 23276 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_287
timestamp 1679235063
transform 1 0 27508 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_295
timestamp 1679235063
transform 1 0 28244 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1679235063
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1679235063
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1679235063
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1679235063
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1679235063
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1679235063
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1679235063
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1679235063
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_3
timestamp 1679235063
transform 1 0 1380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_9
timestamp 1679235063
transform 1 0 1932 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_13
timestamp 1679235063
transform 1 0 2300 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_23
timestamp 1679235063
transform 1 0 3220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1679235063
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1679235063
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_41
timestamp 1679235063
transform 1 0 4876 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1679235063
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1679235063
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1679235063
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_92
timestamp 1679235063
transform 1 0 9568 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_98
timestamp 1679235063
transform 1 0 10120 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1679235063
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_162
timestamp 1679235063
transform 1 0 16008 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_170
timestamp 1679235063
transform 1 0 16744 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1679235063
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_209
timestamp 1679235063
transform 1 0 20332 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_232
timestamp 1679235063
transform 1 0 22448 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1679235063
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_253
timestamp 1679235063
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_261
timestamp 1679235063
transform 1 0 25116 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_266
timestamp 1679235063
transform 1 0 25576 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_272
timestamp 1679235063
transform 1 0 26128 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_284
timestamp 1679235063
transform 1 0 27232 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1679235063
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1679235063
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_321
timestamp 1679235063
transform 1 0 30636 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_331
timestamp 1679235063
transform 1 0 31556 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_343
timestamp 1679235063
transform 1 0 32660 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_355
timestamp 1679235063
transform 1 0 33764 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1679235063
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1679235063
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_377
timestamp 1679235063
transform 1 0 35788 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_6
timestamp 1679235063
transform 1 0 1656 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_23
timestamp 1679235063
transform 1 0 3220 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_31
timestamp 1679235063
transform 1 0 3956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_43
timestamp 1679235063
transform 1 0 5060 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_51
timestamp 1679235063
transform 1 0 5796 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_57
timestamp 1679235063
transform 1 0 6348 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_74
timestamp 1679235063
transform 1 0 7912 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_86
timestamp 1679235063
transform 1 0 9016 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_98
timestamp 1679235063
transform 1 0 10120 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1679235063
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1679235063
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_121
timestamp 1679235063
transform 1 0 12236 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1679235063
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1679235063
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1679235063
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1679235063
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1679235063
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1679235063
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_181
timestamp 1679235063
transform 1 0 17756 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_225
timestamp 1679235063
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_233
timestamp 1679235063
transform 1 0 22540 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_250
timestamp 1679235063
transform 1 0 24104 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_258
timestamp 1679235063
transform 1 0 24840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_270
timestamp 1679235063
transform 1 0 25944 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1679235063
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_281
timestamp 1679235063
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_305
timestamp 1679235063
transform 1 0 29164 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_318
timestamp 1679235063
transform 1 0 30360 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1679235063
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1679235063
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1679235063
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1679235063
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1679235063
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_15
timestamp 1679235063
transform 1 0 2484 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_23
timestamp 1679235063
transform 1 0 3220 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_54
timestamp 1679235063
transform 1 0 6072 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_60
timestamp 1679235063
transform 1 0 6624 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_70
timestamp 1679235063
transform 1 0 7544 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1679235063
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_89
timestamp 1679235063
transform 1 0 9292 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_95
timestamp 1679235063
transform 1 0 9844 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_99
timestamp 1679235063
transform 1 0 10212 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_104
timestamp 1679235063
transform 1 0 10672 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_116
timestamp 1679235063
transform 1 0 11776 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_128
timestamp 1679235063
transform 1 0 12880 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_150
timestamp 1679235063
transform 1 0 14904 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_162
timestamp 1679235063
transform 1 0 16008 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_172
timestamp 1679235063
transform 1 0 16928 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_176
timestamp 1679235063
transform 1 0 17296 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_186
timestamp 1679235063
transform 1 0 18216 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1679235063
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1679235063
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1679235063
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1679235063
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1679235063
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1679235063
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1679235063
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_253
timestamp 1679235063
transform 1 0 24380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_275
timestamp 1679235063
transform 1 0 26404 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_279
timestamp 1679235063
transform 1 0 26772 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_296
timestamp 1679235063
transform 1 0 28336 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_304
timestamp 1679235063
transform 1 0 29072 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_328
timestamp 1679235063
transform 1 0 31280 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_340
timestamp 1679235063
transform 1 0 32384 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_352
timestamp 1679235063
transform 1 0 33488 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1679235063
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_377
timestamp 1679235063
transform 1 0 35788 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1679235063
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1679235063
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_27
timestamp 1679235063
transform 1 0 3588 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_35
timestamp 1679235063
transform 1 0 4324 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1679235063
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_57
timestamp 1679235063
transform 1 0 6348 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_76
timestamp 1679235063
transform 1 0 8096 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_116
timestamp 1679235063
transform 1 0 11776 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_134
timestamp 1679235063
transform 1 0 13432 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_195
timestamp 1679235063
transform 1 0 19044 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_199
timestamp 1679235063
transform 1 0 19412 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_213
timestamp 1679235063
transform 1 0 20700 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1679235063
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_234
timestamp 1679235063
transform 1 0 22632 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_244
timestamp 1679235063
transform 1 0 23552 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_255
timestamp 1679235063
transform 1 0 24564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_259
timestamp 1679235063
transform 1 0 24932 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_270
timestamp 1679235063
transform 1 0 25944 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1679235063
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1679235063
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_295
timestamp 1679235063
transform 1 0 28244 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_307
timestamp 1679235063
transform 1 0 29348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_319
timestamp 1679235063
transform 1 0 30452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_331
timestamp 1679235063
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1679235063
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1679235063
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1679235063
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1679235063
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_373
timestamp 1679235063
transform 1 0 35420 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_3
timestamp 1679235063
transform 1 0 1380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_12
timestamp 1679235063
transform 1 0 2208 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_22
timestamp 1679235063
transform 1 0 3128 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1679235063
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_41
timestamp 1679235063
transform 1 0 4876 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1679235063
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1679235063
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1679235063
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_109
timestamp 1679235063
transform 1 0 11132 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_117
timestamp 1679235063
transform 1 0 11868 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_134
timestamp 1679235063
transform 1 0 13432 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_144
timestamp 1679235063
transform 1 0 14352 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_156
timestamp 1679235063
transform 1 0 15456 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_168
timestamp 1679235063
transform 1 0 16560 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_174
timestamp 1679235063
transform 1 0 17112 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_179
timestamp 1679235063
transform 1 0 17572 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_191
timestamp 1679235063
transform 1 0 18676 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1679235063
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1679235063
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_215
timestamp 1679235063
transform 1 0 20884 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_235
timestamp 1679235063
transform 1 0 22724 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_256
timestamp 1679235063
transform 1 0 24656 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_260
timestamp 1679235063
transform 1 0 25024 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_282
timestamp 1679235063
transform 1 0 27048 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_294
timestamp 1679235063
transform 1 0 28152 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1679235063
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1679235063
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_320
timestamp 1679235063
transform 1 0 30544 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_338
timestamp 1679235063
transform 1 0 32200 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_350
timestamp 1679235063
transform 1 0 33304 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1679235063
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1679235063
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_377
timestamp 1679235063
transform 1 0 35788 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1679235063
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_21
timestamp 1679235063
transform 1 0 3036 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_42
timestamp 1679235063
transform 1 0 4968 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1679235063
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_57
timestamp 1679235063
transform 1 0 6348 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_63
timestamp 1679235063
transform 1 0 6900 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_73
timestamp 1679235063
transform 1 0 7820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_85
timestamp 1679235063
transform 1 0 8924 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1679235063
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1679235063
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1679235063
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1679235063
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1679235063
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1679235063
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1679235063
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1679235063
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1679235063
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1679235063
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_193
timestamp 1679235063
transform 1 0 18860 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_201
timestamp 1679235063
transform 1 0 19596 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1679235063
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1679235063
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1679235063
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1679235063
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_237
timestamp 1679235063
transform 1 0 22908 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_244
timestamp 1679235063
transform 1 0 23552 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_256
timestamp 1679235063
transform 1 0 24656 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_281
timestamp 1679235063
transform 1 0 26956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_296
timestamp 1679235063
transform 1 0 28336 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_304
timestamp 1679235063
transform 1 0 29072 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1679235063
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1679235063
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1679235063
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1679235063
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1679235063
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1679235063
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1679235063
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_29
timestamp 1679235063
transform 1 0 3772 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_39
timestamp 1679235063
transform 1 0 4692 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_68
timestamp 1679235063
transform 1 0 7360 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_76
timestamp 1679235063
transform 1 0 8096 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1679235063
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_88
timestamp 1679235063
transform 1 0 9200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_93
timestamp 1679235063
transform 1 0 9660 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_118
timestamp 1679235063
transform 1 0 11960 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_122
timestamp 1679235063
transform 1 0 12328 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_132
timestamp 1679235063
transform 1 0 13248 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_165
timestamp 1679235063
transform 1 0 16284 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1679235063
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1679235063
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1679235063
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1679235063
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1679235063
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1679235063
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1679235063
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1679235063
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1679235063
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_277
timestamp 1679235063
transform 1 0 26588 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_281
timestamp 1679235063
transform 1 0 26956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1679235063
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_309
timestamp 1679235063
transform 1 0 29532 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_313
timestamp 1679235063
transform 1 0 29900 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_321
timestamp 1679235063
transform 1 0 30636 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_331
timestamp 1679235063
transform 1 0 31556 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_343
timestamp 1679235063
transform 1 0 32660 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_355
timestamp 1679235063
transform 1 0 33764 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1679235063
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1679235063
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_377
timestamp 1679235063
transform 1 0 35788 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_7
timestamp 1679235063
transform 1 0 1748 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_12
timestamp 1679235063
transform 1 0 2208 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_22
timestamp 1679235063
transform 1 0 3128 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1679235063
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1679235063
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1679235063
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_57
timestamp 1679235063
transform 1 0 6348 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1679235063
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1679235063
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_113
timestamp 1679235063
transform 1 0 11500 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_133
timestamp 1679235063
transform 1 0 13340 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_158
timestamp 1679235063
transform 1 0 15640 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_169
timestamp 1679235063
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_194
timestamp 1679235063
transform 1 0 18952 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1679235063
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1679235063
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1679235063
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1679235063
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1679235063
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_281
timestamp 1679235063
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_308
timestamp 1679235063
transform 1 0 29440 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_320
timestamp 1679235063
transform 1 0 30544 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1679235063
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1679235063
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1679235063
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1679235063
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1679235063
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_3
timestamp 1679235063
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_22
timestamp 1679235063
transform 1 0 3128 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_45
timestamp 1679235063
transform 1 0 5244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_57
timestamp 1679235063
transform 1 0 6348 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_81
timestamp 1679235063
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1679235063
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_118
timestamp 1679235063
transform 1 0 11960 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_124
timestamp 1679235063
transform 1 0 12512 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1679235063
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1679235063
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_152
timestamp 1679235063
transform 1 0 15088 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_172
timestamp 1679235063
transform 1 0 16928 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_187
timestamp 1679235063
transform 1 0 18308 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_197
timestamp 1679235063
transform 1 0 19228 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_253
timestamp 1679235063
transform 1 0 24380 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_284
timestamp 1679235063
transform 1 0 27232 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_296
timestamp 1679235063
transform 1 0 28336 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1679235063
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1679235063
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1679235063
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1679235063
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1679235063
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1679235063
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1679235063
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_377
timestamp 1679235063
transform 1 0 35788 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1679235063
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1679235063
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1679235063
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_39
timestamp 1679235063
transform 1 0 4692 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_43
timestamp 1679235063
transform 1 0 5060 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_47
timestamp 1679235063
transform 1 0 5428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1679235063
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1679235063
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1679235063
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1679235063
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1679235063
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1679235063
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1679235063
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1679235063
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1679235063
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_137
timestamp 1679235063
transform 1 0 13708 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_146
timestamp 1679235063
transform 1 0 14536 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_158
timestamp 1679235063
transform 1 0 15640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1679235063
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1679235063
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_173
timestamp 1679235063
transform 1 0 17020 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_193
timestamp 1679235063
transform 1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_212
timestamp 1679235063
transform 1 0 20608 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_225
timestamp 1679235063
transform 1 0 21804 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_242
timestamp 1679235063
transform 1 0 23368 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_254
timestamp 1679235063
transform 1 0 24472 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_266
timestamp 1679235063
transform 1 0 25576 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_274
timestamp 1679235063
transform 1 0 26312 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1679235063
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_297
timestamp 1679235063
transform 1 0 28428 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_309
timestamp 1679235063
transform 1 0 29532 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_321
timestamp 1679235063
transform 1 0 30636 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1679235063
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1679235063
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1679235063
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1679235063
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_373
timestamp 1679235063
transform 1 0 35420 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1679235063
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1679235063
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1679235063
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_29
timestamp 1679235063
transform 1 0 3772 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_33
timestamp 1679235063
transform 1 0 4140 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_37
timestamp 1679235063
transform 1 0 4508 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_74
timestamp 1679235063
transform 1 0 7912 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1679235063
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_89
timestamp 1679235063
transform 1 0 9292 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_97
timestamp 1679235063
transform 1 0 10028 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_103
timestamp 1679235063
transform 1 0 10580 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_115
timestamp 1679235063
transform 1 0 11684 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_58_133
timestamp 1679235063
transform 1 0 13340 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1679235063
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_157
timestamp 1679235063
transform 1 0 15548 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_163
timestamp 1679235063
transform 1 0 16100 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_173
timestamp 1679235063
transform 1 0 17020 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_185
timestamp 1679235063
transform 1 0 18124 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 1679235063
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1679235063
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1679235063
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1679235063
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1679235063
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1679235063
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1679235063
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1679235063
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1679235063
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1679235063
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1679235063
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1679235063
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1679235063
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1679235063
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1679235063
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1679235063
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1679235063
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1679235063
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1679235063
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1679235063
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_377
timestamp 1679235063
transform 1 0 35788 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1679235063
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1679235063
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_27
timestamp 1679235063
transform 1 0 3588 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1679235063
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_57
timestamp 1679235063
transform 1 0 6348 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_79
timestamp 1679235063
transform 1 0 8372 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_116
timestamp 1679235063
transform 1 0 11776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_133
timestamp 1679235063
transform 1 0 13340 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_150
timestamp 1679235063
transform 1 0 14904 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_172
timestamp 1679235063
transform 1 0 16928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_199
timestamp 1679235063
transform 1 0 19412 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_207
timestamp 1679235063
transform 1 0 20148 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_219
timestamp 1679235063
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1679235063
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_234
timestamp 1679235063
transform 1 0 22632 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_246
timestamp 1679235063
transform 1 0 23736 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_256
timestamp 1679235063
transform 1 0 24656 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_260
timestamp 1679235063
transform 1 0 25024 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1679235063
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1679235063
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1679235063
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1679235063
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1679235063
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1679235063
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1679235063
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1679235063
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1679235063
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1679235063
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_7
timestamp 1679235063
transform 1 0 1748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 1679235063
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1679235063
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1679235063
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1679235063
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_53
timestamp 1679235063
transform 1 0 5980 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_64
timestamp 1679235063
transform 1 0 6992 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_76
timestamp 1679235063
transform 1 0 8096 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_89
timestamp 1679235063
transform 1 0 9292 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_95
timestamp 1679235063
transform 1 0 9844 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_107
timestamp 1679235063
transform 1 0 10948 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_119
timestamp 1679235063
transform 1 0 12052 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_131
timestamp 1679235063
transform 1 0 13156 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1679235063
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_150
timestamp 1679235063
transform 1 0 14904 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_162
timestamp 1679235063
transform 1 0 16008 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_174
timestamp 1679235063
transform 1 0 17112 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_191
timestamp 1679235063
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1679235063
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp 1679235063
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_201
timestamp 1679235063
transform 1 0 19596 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_214
timestamp 1679235063
transform 1 0 20792 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_234
timestamp 1679235063
transform 1 0 22632 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_256
timestamp 1679235063
transform 1 0 24656 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_276
timestamp 1679235063
transform 1 0 26496 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_288
timestamp 1679235063
transform 1 0 27600 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_300
timestamp 1679235063
transform 1 0 28704 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1679235063
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_320
timestamp 1679235063
transform 1 0 30544 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_332
timestamp 1679235063
transform 1 0 31648 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_344
timestamp 1679235063
transform 1 0 32752 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_356
timestamp 1679235063
transform 1 0 33856 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1679235063
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_377
timestamp 1679235063
transform 1 0 35788 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1679235063
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1679235063
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1679235063
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1679235063
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1679235063
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1679235063
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_60
timestamp 1679235063
transform 1 0 6624 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_72
timestamp 1679235063
transform 1 0 7728 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_84
timestamp 1679235063
transform 1 0 8832 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_96
timestamp 1679235063
transform 1 0 9936 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_108
timestamp 1679235063
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1679235063
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1679235063
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1679235063
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1679235063
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1679235063
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1679235063
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_178
timestamp 1679235063
transform 1 0 17480 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_190
timestamp 1679235063
transform 1 0 18584 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_198
timestamp 1679235063
transform 1 0 19320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_215
timestamp 1679235063
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1679235063
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1679235063
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1679235063
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1679235063
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1679235063
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1679235063
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1679235063
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1679235063
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_293
timestamp 1679235063
transform 1 0 28060 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_301
timestamp 1679235063
transform 1 0 28796 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_326
timestamp 1679235063
transform 1 0 31096 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1679235063
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1679235063
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1679235063
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1679235063
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1679235063
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1679235063
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1679235063
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1679235063
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1679235063
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_41
timestamp 1679235063
transform 1 0 4876 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_49
timestamp 1679235063
transform 1 0 5612 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_67
timestamp 1679235063
transform 1 0 7268 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_79
timestamp 1679235063
transform 1 0 8372 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1679235063
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1679235063
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1679235063
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1679235063
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1679235063
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1679235063
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1679235063
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1679235063
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_153
timestamp 1679235063
transform 1 0 15180 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_159
timestamp 1679235063
transform 1 0 15732 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_176
timestamp 1679235063
transform 1 0 17296 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_181
timestamp 1679235063
transform 1 0 17756 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1679235063
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_197
timestamp 1679235063
transform 1 0 19228 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_209
timestamp 1679235063
transform 1 0 20332 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_217
timestamp 1679235063
transform 1 0 21068 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_235
timestamp 1679235063
transform 1 0 22724 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1679235063
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1679235063
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1679235063
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1679235063
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1679235063
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1679235063
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1679235063
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1679235063
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_309
timestamp 1679235063
transform 1 0 29532 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1679235063
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1679235063
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1679235063
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1679235063
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1679235063
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_377
timestamp 1679235063
transform 1 0 35788 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1679235063
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1679235063
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1679235063
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1679235063
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1679235063
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1679235063
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_57
timestamp 1679235063
transform 1 0 6348 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_61
timestamp 1679235063
transform 1 0 6716 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_75
timestamp 1679235063
transform 1 0 8004 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_87
timestamp 1679235063
transform 1 0 9108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_99
timestamp 1679235063
transform 1 0 10212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1679235063
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1679235063
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1679235063
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1679235063
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1679235063
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_161
timestamp 1679235063
transform 1 0 15916 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_169
timestamp 1679235063
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_173
timestamp 1679235063
transform 1 0 17020 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_193
timestamp 1679235063
transform 1 0 18860 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_213
timestamp 1679235063
transform 1 0 20700 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_234
timestamp 1679235063
transform 1 0 22632 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_252
timestamp 1679235063
transform 1 0 24288 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_264
timestamp 1679235063
transform 1 0 25392 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1679235063
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1679235063
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1679235063
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_305
timestamp 1679235063
transform 1 0 29164 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_313
timestamp 1679235063
transform 1 0 29900 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_318
timestamp 1679235063
transform 1 0 30360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 1679235063
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1679235063
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1679235063
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1679235063
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1679235063
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1679235063
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1679235063
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1679235063
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_29
timestamp 1679235063
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_37
timestamp 1679235063
transform 1 0 4508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 1679235063
transform 1 0 5520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_57
timestamp 1679235063
transform 1 0 6348 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_65
timestamp 1679235063
transform 1 0 7084 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_70
timestamp 1679235063
transform 1 0 7544 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1679235063
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1679235063
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_97
timestamp 1679235063
transform 1 0 10028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_105
timestamp 1679235063
transform 1 0 10764 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1679235063
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_113
timestamp 1679235063
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_125
timestamp 1679235063
transform 1 0 12604 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_133
timestamp 1679235063
transform 1 0 13340 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1679235063
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_153
timestamp 1679235063
transform 1 0 15180 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_161
timestamp 1679235063
transform 1 0 15916 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_169
timestamp 1679235063
transform 1 0 16652 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_177
timestamp 1679235063
transform 1 0 17388 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_190
timestamp 1679235063
transform 1 0 18584 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1679235063
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1679235063
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_225
timestamp 1679235063
transform 1 0 21804 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_239
timestamp 1679235063
transform 1 0 23092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1679235063
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1679235063
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_265
timestamp 1679235063
transform 1 0 25484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_273
timestamp 1679235063
transform 1 0 26220 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1679235063
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_281
timestamp 1679235063
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 1679235063
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1679235063
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1679235063
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_321
timestamp 1679235063
transform 1 0 30636 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_329
timestamp 1679235063
transform 1 0 31372 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_337
timestamp 1679235063
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_349
timestamp 1679235063
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1679235063
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1679235063
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_370
timestamp 1679235063
transform 1 0 35144 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 36248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1679235063
transform 1 0 2116 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1679235063
transform 1 0 4600 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1679235063
transform 1 0 1380 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 21344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1679235063
transform 1 0 35604 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1679235063
transform 1 0 28428 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1679235063
transform 1 0 20148 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 36248 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1679235063
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 1380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1679235063
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1679235063
transform 1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1679235063
transform 1 0 36248 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1679235063
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1679235063
transform 1 0 35972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1679235063
transform 1 0 36156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1679235063
transform 1 0 36156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1679235063
transform 1 0 30452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1679235063
transform 1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1679235063
transform 1 0 10396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1679235063
transform 1 0 1564 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1679235063
transform 1 0 22724 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1679235063
transform 1 0 16192 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1679235063
transform 1 0 25852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1679235063
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1679235063
transform 1 0 36156 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1679235063
transform 1 0 36156 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1679235063
transform 1 0 35972 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1679235063
transform 1 0 31464 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1679235063
transform -1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1679235063
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1679235063
transform 1 0 36156 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1679235063
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1679235063
transform 1 0 36156 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1679235063
transform 1 0 7176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1679235063
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1679235063
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1679235063
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 36800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 36800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 36800 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 36800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 36800 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 36800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 36800 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 36800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 36800 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 36800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 36800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 36800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 36800 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 36800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 36800 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 36800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 36800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 36800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 36800 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 36800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 36800 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 36800 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 36800 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 36800 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 36800 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 36800 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 36800 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 36800 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 36800 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 36800 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 36800 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 36800 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 36800 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 36800 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 36800 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 36800 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 36800 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 36800 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 36800 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 36800 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 36800 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1679235063
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1679235063
transform -1 0 36800 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1679235063
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1679235063
transform -1 0 36800 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1679235063
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1679235063
transform -1 0 36800 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1679235063
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1679235063
transform -1 0 36800 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1679235063
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1679235063
transform -1 0 36800 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1679235063
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1679235063
transform -1 0 36800 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1679235063
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1679235063
transform -1 0 36800 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1679235063
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1679235063
transform -1 0 36800 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1679235063
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1679235063
transform -1 0 36800 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1679235063
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1679235063
transform -1 0 36800 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1679235063
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1679235063
transform -1 0 36800 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1679235063
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1679235063
transform -1 0 36800 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1679235063
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1679235063
transform -1 0 36800 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1679235063
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1679235063
transform -1 0 36800 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1679235063
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1679235063
transform -1 0 36800 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1679235063
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1679235063
transform -1 0 36800 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1679235063
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1679235063
transform -1 0 36800 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1679235063
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1679235063
transform -1 0 36800 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1679235063
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1679235063
transform -1 0 36800 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1679235063
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1679235063
transform -1 0 36800 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1679235063
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1679235063
transform -1 0 36800 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1679235063
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1679235063
transform -1 0 36800 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1679235063
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1679235063
transform -1 0 36800 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1679235063
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1679235063
transform -1 0 36800 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1679235063
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1679235063
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1679235063
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1679235063
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1679235063
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1679235063
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1679235063
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1679235063
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1679235063
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1679235063
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1679235063
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1679235063
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1679235063
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1679235063
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1679235063
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1679235063
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1679235063
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1679235063
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1679235063
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1679235063
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1679235063
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1679235063
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1679235063
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1679235063
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1679235063
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1679235063
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1679235063
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1679235063
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1679235063
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1679235063
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1679235063
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1679235063
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1679235063
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1679235063
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1679235063
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1679235063
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1679235063
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1679235063
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1679235063
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1679235063
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1679235063
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1679235063
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1679235063
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1679235063
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1679235063
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1679235063
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1679235063
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1679235063
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1679235063
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1679235063
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1679235063
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1679235063
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1679235063
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1679235063
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1679235063
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1679235063
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1679235063
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1679235063
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1679235063
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1679235063
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1679235063
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1679235063
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1679235063
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1679235063
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1679235063
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1679235063
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1679235063
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1679235063
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1679235063
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1679235063
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1679235063
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1679235063
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1679235063
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1679235063
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1679235063
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1679235063
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1679235063
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1679235063
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1679235063
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1679235063
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1679235063
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1679235063
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1679235063
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1679235063
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1679235063
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1679235063
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1679235063
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1679235063
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1679235063
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1679235063
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1679235063
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1679235063
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1679235063
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1679235063
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1679235063
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1679235063
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1679235063
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1679235063
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1679235063
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1679235063
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1679235063
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1679235063
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1679235063
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1679235063
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1679235063
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1679235063
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1679235063
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1679235063
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1679235063
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1679235063
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1679235063
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1679235063
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1679235063
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1679235063
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  vahid6i_110 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 35880 0 1 36992
box -38 -48 314 592
<< labels >>
flabel metal3 s 37136 7488 37936 7608 0 FreeSans 480 0 0 0 D_R_data[0]
port 0 nsew signal input
flabel metal2 s 1306 39280 1362 40080 0 FreeSans 224 90 0 0 D_R_data[1]
port 1 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 D_R_data[2]
port 2 nsew signal input
flabel metal2 s 4526 39280 4582 40080 0 FreeSans 224 90 0 0 D_R_data[3]
port 3 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 D_R_data[4]
port 4 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 D_R_data[5]
port 5 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 D_R_data[6]
port 6 nsew signal input
flabel metal2 s 28354 39280 28410 40080 0 FreeSans 224 90 0 0 D_R_data[7]
port 7 nsew signal input
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 D_W_data[0]
port 8 nsew signal tristate
flabel metal3 s 37136 1368 37936 1488 0 FreeSans 480 0 0 0 D_W_data[1]
port 9 nsew signal tristate
flabel metal3 s 37136 14288 37936 14408 0 FreeSans 480 0 0 0 D_W_data[2]
port 10 nsew signal tristate
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 D_W_data[3]
port 11 nsew signal tristate
flabel metal3 s 37136 4768 37936 4888 0 FreeSans 480 0 0 0 D_W_data[4]
port 12 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 D_W_data[5]
port 13 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 D_W_data[6]
port 14 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 D_W_data[7]
port 15 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 D_addr[0]
port 16 nsew signal tristate
flabel metal3 s 37136 36728 37936 36848 0 FreeSans 480 0 0 0 D_addr[1]
port 17 nsew signal tristate
flabel metal2 s 10322 39280 10378 40080 0 FreeSans 224 90 0 0 D_addr[2]
port 18 nsew signal tristate
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 D_addr[3]
port 19 nsew signal tristate
flabel metal2 s 22558 39280 22614 40080 0 FreeSans 224 90 0 0 D_addr[4]
port 20 nsew signal tristate
flabel metal2 s 16118 39280 16174 40080 0 FreeSans 224 90 0 0 D_addr[5]
port 21 nsew signal tristate
flabel metal2 s 25778 39280 25834 40080 0 FreeSans 224 90 0 0 D_addr[6]
port 22 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 D_addr[7]
port 23 nsew signal tristate
flabel metal3 s 37136 33328 37936 33448 0 FreeSans 480 0 0 0 D_rd
port 24 nsew signal tristate
flabel metal3 s 37136 27208 37936 27328 0 FreeSans 480 0 0 0 D_wr
port 25 nsew signal tristate
flabel metal3 s 37136 20408 37936 20528 0 FreeSans 480 0 0 0 I_addr[0]
port 26 nsew signal tristate
flabel metal2 s 31574 39280 31630 40080 0 FreeSans 224 90 0 0 I_addr[1]
port 27 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 I_addr[2]
port 28 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 I_addr[3]
port 29 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 I_addr[4]
port 30 nsew signal tristate
flabel metal3 s 37136 29928 37936 30048 0 FreeSans 480 0 0 0 I_addr[5]
port 31 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 I_addr[6]
port 32 nsew signal tristate
flabel metal3 s 37136 23808 37936 23928 0 FreeSans 480 0 0 0 I_addr[7]
port 33 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 I_data[0]
port 34 nsew signal input
flabel metal2 s 19338 39280 19394 40080 0 FreeSans 224 90 0 0 I_data[1]
port 35 nsew signal input
flabel metal3 s 37136 10888 37936 11008 0 FreeSans 480 0 0 0 I_data[2]
port 36 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 I_data[3]
port 37 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 I_data[4]
port 38 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 I_data[5]
port 39 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 I_data[6]
port 40 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 I_data[7]
port 41 nsew signal input
flabel metal2 s 37370 39280 37426 40080 0 FreeSans 224 90 0 0 I_rd
port 42 nsew signal tristate
flabel metal4 s 4868 2128 5188 37584 0 FreeSans 1920 90 0 0 VGND
port 43 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 37584 0 FreeSans 1920 90 0 0 VGND
port 43 nsew ground bidirectional
flabel metal5 s 1056 6006 36848 6326 0 FreeSans 2560 0 0 0 VGND
port 43 nsew ground bidirectional
flabel metal5 s 1056 36642 36848 36962 0 FreeSans 2560 0 0 0 VGND
port 43 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 VPWR
port 44 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 VPWR
port 44 nsew power bidirectional
flabel metal5 s 1056 5346 36848 5666 0 FreeSans 2560 0 0 0 VPWR
port 44 nsew power bidirectional
flabel metal5 s 1056 35982 36848 36302 0 FreeSans 2560 0 0 0 VPWR
port 44 nsew power bidirectional
flabel metal2 s 34794 39280 34850 40080 0 FreeSans 224 90 0 0 clock
port 45 nsew signal input
flabel metal2 s 7102 39280 7158 40080 0 FreeSans 224 90 0 0 led_clock
port 46 nsew signal tristate
flabel metal2 s 13542 39280 13598 40080 0 FreeSans 224 90 0 0 leds[0]
port 47 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 leds[1]
port 48 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 leds[2]
port 49 nsew signal tristate
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 leds[3]
port 50 nsew signal tristate
flabel metal3 s 37136 17008 37936 17128 0 FreeSans 480 0 0 0 reset
port 51 nsew signal input
rlabel metal1 18952 36992 18952 36992 0 VGND
rlabel metal1 18952 37536 18952 37536 0 VPWR
rlabel metal2 36478 7701 36478 7701 0 D_R_data[0]
rlabel metal1 1794 37162 1794 37162 0 D_R_data[1]
rlabel metal2 27094 1588 27094 1588 0 D_R_data[2]
rlabel metal2 4646 38335 4646 38335 0 D_R_data[3]
rlabel metal3 1050 25228 1050 25228 0 D_R_data[4]
rlabel metal2 21298 1588 21298 1588 0 D_R_data[5]
rlabel metal2 36110 1622 36110 1622 0 D_R_data[6]
rlabel metal2 28474 38335 28474 38335 0 D_R_data[7]
rlabel metal3 820 32028 820 32028 0 D_W_data[0]
rlabel metal3 36348 1428 36348 1428 0 D_W_data[1]
rlabel metal2 36386 14297 36386 14297 0 D_W_data[2]
rlabel metal3 820 22508 820 22508 0 D_W_data[3]
rlabel metal2 36386 4913 36386 4913 0 D_W_data[4]
rlabel metal1 1472 5882 1472 5882 0 D_W_data[5]
rlabel metal3 820 19108 820 19108 0 D_W_data[6]
rlabel metal3 1142 12308 1142 12308 0 D_W_data[7]
rlabel metal2 30314 1095 30314 1095 0 D_addr[0]
rlabel metal2 36386 36941 36386 36941 0 D_addr[1]
rlabel metal2 10626 38233 10626 38233 0 D_addr[2]
rlabel metal3 820 38148 820 38148 0 D_addr[3]
rlabel metal2 22954 38233 22954 38233 0 D_addr[4]
rlabel metal2 16422 38233 16422 38233 0 D_addr[5]
rlabel metal2 26082 38233 26082 38233 0 D_addr[6]
rlabel metal2 14858 1520 14858 1520 0 D_addr[7]
rlabel via2 36386 33371 36386 33371 0 D_rd
rlabel via2 36386 27285 36386 27285 0 D_wr
rlabel metal2 36386 20621 36386 20621 0 I_addr[0]
rlabel metal2 31786 37825 31786 37825 0 I_addr[1]
rlabel metal2 2622 1520 2622 1520 0 I_addr[2]
rlabel metal2 46 1554 46 1554 0 I_addr[3]
rlabel metal3 1142 9588 1142 9588 0 I_addr[4]
rlabel via2 36386 30005 36386 30005 0 I_addr[5]
rlabel metal2 11638 1520 11638 1520 0 I_addr[6]
rlabel metal2 36386 23953 36386 23953 0 I_addr[7]
rlabel metal2 32890 1588 32890 1588 0 I_data[0]
rlabel metal1 20010 37230 20010 37230 0 I_data[1]
rlabel metal2 36478 11033 36478 11033 0 I_data[2]
rlabel metal2 5842 1588 5842 1588 0 I_data[3]
rlabel metal2 9062 1588 9062 1588 0 I_data[4]
rlabel metal3 1142 28628 1142 28628 0 I_data[5]
rlabel metal3 820 2788 820 2788 0 I_data[6]
rlabel metal2 18078 1588 18078 1588 0 I_data[7]
rlabel metal1 32338 18088 32338 18088 0 _0000_
rlabel metal2 30406 18207 30406 18207 0 _0001_
rlabel metal1 29762 20434 29762 20434 0 _0002_
rlabel metal1 18032 20774 18032 20774 0 _0003_
rlabel metal2 23414 17510 23414 17510 0 _0004_
rlabel metal1 21712 18734 21712 18734 0 _0005_
rlabel metal1 22356 15674 22356 15674 0 _0006_
rlabel metal1 17802 13498 17802 13498 0 _0007_
rlabel metal1 33442 17850 33442 17850 0 _0008_
rlabel metal2 29486 17442 29486 17442 0 _0009_
rlabel metal2 32246 18530 32246 18530 0 _0010_
rlabel metal2 26358 16354 26358 16354 0 _0011_
rlabel metal2 22402 15096 22402 15096 0 _0012_
rlabel metal2 20102 15878 20102 15878 0 _0013_
rlabel metal1 20730 15402 20730 15402 0 _0014_
rlabel metal1 16744 12954 16744 12954 0 _0015_
rlabel metal1 14025 30294 14025 30294 0 _0016_
rlabel metal2 7866 30498 7866 30498 0 _0017_
rlabel metal1 17234 30294 17234 30294 0 _0018_
rlabel viali 4917 30226 4917 30226 0 _0019_
rlabel metal1 29516 29546 29516 29546 0 _0020_
rlabel metal1 24962 29546 24962 29546 0 _0021_
rlabel metal1 21282 30634 21282 30634 0 _0022_
rlabel via1 10253 30226 10253 30226 0 _0023_
rlabel metal2 12466 28764 12466 28764 0 _0024_
rlabel metal2 1794 27234 1794 27234 0 _0025_
rlabel via1 15497 27438 15497 27438 0 _0026_
rlabel metal2 2070 28934 2070 28934 0 _0027_
rlabel via1 27181 29614 27181 29614 0 _0028_
rlabel metal1 23000 28730 23000 28730 0 _0029_
rlabel metal1 19228 28730 19228 28730 0 _0030_
rlabel metal1 8827 28118 8827 28118 0 _0031_
rlabel metal2 12374 30498 12374 30498 0 _0032_
rlabel metal1 6378 29206 6378 29206 0 _0033_
rlabel metal1 16049 30226 16049 30226 0 _0034_
rlabel metal1 3756 29546 3756 29546 0 _0035_
rlabel metal1 30953 29206 30953 29206 0 _0036_
rlabel metal1 23777 30634 23777 30634 0 _0037_
rlabel via1 19729 30702 19729 30702 0 _0038_
rlabel metal2 9154 30022 9154 30022 0 _0039_
rlabel metal1 14520 22678 14520 22678 0 _0040_
rlabel metal1 1840 20026 1840 20026 0 _0041_
rlabel metal1 17234 21590 17234 21590 0 _0042_
rlabel metal2 1794 23970 1794 23970 0 _0043_
rlabel metal1 27722 23018 27722 23018 0 _0044_
rlabel metal1 25346 21896 25346 21896 0 _0045_
rlabel metal1 21114 21896 21114 21896 0 _0046_
rlabel metal2 9338 21658 9338 21658 0 _0047_
rlabel metal2 12374 24582 12374 24582 0 _0048_
rlabel metal2 1978 21794 1978 21794 0 _0049_
rlabel metal2 15686 23494 15686 23494 0 _0050_
rlabel via1 1789 25262 1789 25262 0 _0051_
rlabel via1 27917 25262 27917 25262 0 _0052_
rlabel via1 26261 25262 26261 25262 0 _0053_
rlabel metal1 19212 25194 19212 25194 0 _0054_
rlabel metal1 8697 23834 8697 23834 0 _0055_
rlabel metal2 11914 18530 11914 18530 0 _0056_
rlabel metal2 1886 17442 1886 17442 0 _0057_
rlabel metal2 15226 18530 15226 18530 0 _0058_
rlabel via1 2157 18734 2157 18734 0 _0059_
rlabel metal1 28929 20842 28929 20842 0 _0060_
rlabel metal2 23414 21318 23414 21318 0 _0061_
rlabel metal1 21650 19754 21650 19754 0 _0062_
rlabel via1 8321 19346 8321 19346 0 _0063_
rlabel metal1 12236 34170 12236 34170 0 _0064_
rlabel metal1 6251 36074 6251 36074 0 _0065_
rlabel metal1 16049 34646 16049 34646 0 _0066_
rlabel metal1 4462 34170 4462 34170 0 _0067_
rlabel metal2 29670 31518 29670 31518 0 _0068_
rlabel metal1 23777 34986 23777 34986 0 _0069_
rlabel metal2 19734 35462 19734 35462 0 _0070_
rlabel metal1 9011 34646 9011 34646 0 _0071_
rlabel metal1 12231 32470 12231 32470 0 _0072_
rlabel metal1 3756 32810 3756 32810 0 _0073_
rlabel metal2 16054 32300 16054 32300 0 _0074_
rlabel metal1 3526 31382 3526 31382 0 _0075_
rlabel metal1 27998 32470 27998 32470 0 _0076_
rlabel metal1 23731 32470 23731 32470 0 _0077_
rlabel metal2 18906 33286 18906 33286 0 _0078_
rlabel metal1 8592 32402 8592 32402 0 _0079_
rlabel metal1 13708 34170 13708 34170 0 _0080_
rlabel metal1 6785 34714 6785 34714 0 _0081_
rlabel metal2 17066 34850 17066 34850 0 _0082_
rlabel metal1 5244 33626 5244 33626 0 _0083_
rlabel metal2 31786 30906 31786 30906 0 _0084_
rlabel metal1 25054 34986 25054 34986 0 _0085_
rlabel metal1 21190 34986 21190 34986 0 _0086_
rlabel metal1 10350 34170 10350 34170 0 _0087_
rlabel metal1 14352 33626 14352 33626 0 _0088_
rlabel metal2 1978 32674 1978 32674 0 _0089_
rlabel metal1 17418 33558 17418 33558 0 _0090_
rlabel metal1 1932 30906 1932 30906 0 _0091_
rlabel metal1 27324 31450 27324 31450 0 _0092_
rlabel metal1 26894 33558 26894 33558 0 _0093_
rlabel metal1 22816 32538 22816 32538 0 _0094_
rlabel metal1 9460 31382 9460 31382 0 _0095_
rlabel metal1 34040 10234 34040 10234 0 _0096_
rlabel metal1 34904 7854 34904 7854 0 _0097_
rlabel metal1 32420 5678 32420 5678 0 _0098_
rlabel metal1 29752 5678 29752 5678 0 _0099_
rlabel metal1 27503 7446 27503 7446 0 _0100_
rlabel metal1 32972 5202 32972 5202 0 _0101_
rlabel metal1 29205 3094 29205 3094 0 _0102_
rlabel metal1 32972 3502 32972 3502 0 _0103_
rlabel metal1 14025 27030 14025 27030 0 _0104_
rlabel metal1 3066 27030 3066 27030 0 _0105_
rlabel metal2 17618 26962 17618 26962 0 _0106_
rlabel metal2 3910 27846 3910 27846 0 _0107_
rlabel metal1 27998 27370 27998 27370 0 _0108_
rlabel metal2 25990 27574 25990 27574 0 _0109_
rlabel via1 21758 28101 21758 28101 0 _0110_
rlabel via1 10253 26962 10253 26962 0 _0111_
rlabel metal1 25284 10710 25284 10710 0 _0112_
rlabel metal1 12611 16150 12611 16150 0 _0113_
rlabel via1 5377 14382 5377 14382 0 _0114_
rlabel metal1 16049 15062 16049 15062 0 _0115_
rlabel metal1 3629 13974 3629 13974 0 _0116_
rlabel metal1 27354 17238 27354 17238 0 _0117_
rlabel metal1 22938 16150 22938 16150 0 _0118_
rlabel metal2 18722 15878 18722 15878 0 _0119_
rlabel via1 9149 16082 9149 16082 0 _0120_
rlabel metal2 11822 21794 11822 21794 0 _0121_
rlabel metal1 3399 20502 3399 20502 0 _0122_
rlabel metal2 15318 20706 15318 20706 0 _0123_
rlabel metal2 3818 23494 3818 23494 0 _0124_
rlabel metal2 29210 23494 29210 23494 0 _0125_
rlabel metal1 23731 22678 23731 22678 0 _0126_
rlabel via1 18809 22678 18809 22678 0 _0127_
rlabel metal1 7912 22202 7912 22202 0 _0128_
rlabel metal2 11822 16966 11822 16966 0 _0129_
rlabel via1 4641 16150 4641 16150 0 _0130_
rlabel metal2 15318 16354 15318 16354 0 _0131_
rlabel metal2 2714 15878 2714 15878 0 _0132_
rlabel metal2 26266 17442 26266 17442 0 _0133_
rlabel via1 22765 17646 22765 17646 0 _0134_
rlabel metal1 19166 17578 19166 17578 0 _0135_
rlabel metal2 8050 16218 8050 16218 0 _0136_
rlabel metal1 13554 17238 13554 17238 0 _0137_
rlabel metal2 6394 16354 6394 16354 0 _0138_
rlabel metal2 17250 16966 17250 16966 0 _0139_
rlabel metal1 4048 17306 4048 17306 0 _0140_
rlabel via1 29757 19414 29757 19414 0 _0141_
rlabel metal1 25024 17850 25024 17850 0 _0142_
rlabel metal2 21022 17442 21022 17442 0 _0143_
rlabel via1 9977 17170 9977 17170 0 _0144_
rlabel metal1 24548 12138 24548 12138 0 _0145_
rlabel metal2 21850 12002 21850 12002 0 _0146_
rlabel metal1 26128 9690 26128 9690 0 _0147_
rlabel metal2 24150 7650 24150 7650 0 _0148_
rlabel via1 12185 26350 12185 26350 0 _0149_
rlabel metal2 4646 22406 4646 22406 0 _0150_
rlabel metal1 15962 25160 15962 25160 0 _0151_
rlabel metal1 3721 24854 3721 24854 0 _0152_
rlabel metal1 29516 25194 29516 25194 0 _0153_
rlabel via1 24421 25942 24421 25942 0 _0154_
rlabel via1 19637 26350 19637 26350 0 _0155_
rlabel metal1 9246 25466 9246 25466 0 _0156_
rlabel via1 29205 12818 29205 12818 0 _0157_
rlabel metal1 29654 35734 29654 35734 0 _0158_
rlabel metal1 17418 36822 17418 36822 0 _0159_
rlabel via1 16141 36142 16141 36142 0 _0160_
rlabel via1 21569 36142 21569 36142 0 _0161_
rlabel metal1 19258 36822 19258 36822 0 _0162_
rlabel metal1 24134 13974 24134 13974 0 _0163_
rlabel metal2 16238 3298 16238 3298 0 _0164_
rlabel metal1 34812 12818 34812 12818 0 _0165_
rlabel metal2 35374 18870 35374 18870 0 _0166_
rlabel metal2 15134 8262 15134 8262 0 _0167_
rlabel metal1 13795 6358 13795 6358 0 _0168_
rlabel metal1 20143 9962 20143 9962 0 _0169_
rlabel metal2 25162 15266 25162 15266 0 _0170_
rlabel metal1 31954 20502 31954 20502 0 _0171_
rlabel via1 22305 13974 22305 13974 0 _0172_
rlabel viali 18253 13905 18253 13905 0 _0173_
rlabel metal2 20286 13702 20286 13702 0 _0174_
rlabel metal1 16636 10710 16636 10710 0 _0175_
rlabel metal1 34081 16490 34081 16490 0 _0176_
rlabel metal1 29194 16150 29194 16150 0 _0177_
rlabel metal1 31832 16218 31832 16218 0 _0178_
rlabel metal2 27002 14178 27002 14178 0 _0179_
rlabel metal1 33340 20910 33340 20910 0 _0180_
rlabel metal2 31234 18530 31234 18530 0 _0181_
rlabel metal1 32522 24378 32522 24378 0 _0182_
rlabel metal2 33810 22882 33810 22882 0 _0183_
rlabel metal1 20286 24684 20286 24684 0 _0184_
rlabel metal2 16514 23902 16514 23902 0 _0185_
rlabel metal1 12604 24174 12604 24174 0 _0186_
rlabel metal1 2208 21522 2208 21522 0 _0187_
rlabel metal1 15916 23086 15916 23086 0 _0188_
rlabel metal1 2162 25874 2162 25874 0 _0189_
rlabel metal1 28014 24922 28014 24922 0 _0190_
rlabel metal1 26680 25874 26680 25874 0 _0191_
rlabel metal1 19504 24922 19504 24922 0 _0192_
rlabel via2 8418 23749 8418 23749 0 _0193_
rlabel metal2 31234 21012 31234 21012 0 _0194_
rlabel metal1 16790 19856 16790 19856 0 _0195_
rlabel metal1 16606 19924 16606 19924 0 _0196_
rlabel metal2 12098 18700 12098 18700 0 _0197_
rlabel metal2 2070 17612 2070 17612 0 _0198_
rlabel metal2 15410 18972 15410 18972 0 _0199_
rlabel metal1 2484 19346 2484 19346 0 _0200_
rlabel metal2 29762 21114 29762 21114 0 _0201_
rlabel metal1 24104 20910 24104 20910 0 _0202_
rlabel via1 21390 19820 21390 19820 0 _0203_
rlabel metal2 9062 18530 9062 18530 0 _0204_
rlabel metal1 32062 26350 32062 26350 0 _0205_
rlabel metal1 24518 34476 24518 34476 0 _0206_
rlabel metal2 6762 34816 6762 34816 0 _0207_
rlabel metal1 12512 33966 12512 33966 0 _0208_
rlabel metal2 6210 35462 6210 35462 0 _0209_
rlabel metal1 16560 34170 16560 34170 0 _0210_
rlabel metal1 4600 33966 4600 33966 0 _0211_
rlabel metal1 29808 30906 29808 30906 0 _0212_
rlabel metal1 23920 34714 23920 34714 0 _0213_
rlabel metal1 19964 35054 19964 35054 0 _0214_
rlabel metal1 9476 35122 9476 35122 0 _0215_
rlabel metal2 24334 32674 24334 32674 0 _0216_
rlabel metal1 4554 32266 4554 32266 0 _0217_
rlabel metal2 12466 32436 12466 32436 0 _0218_
rlabel metal1 3772 32538 3772 32538 0 _0219_
rlabel metal2 16238 31994 16238 31994 0 _0220_
rlabel metal1 3680 31654 3680 31654 0 _0221_
rlabel metal2 28566 32198 28566 32198 0 _0222_
rlabel metal2 24242 33082 24242 33082 0 _0223_
rlabel metal1 19228 32878 19228 32878 0 _0224_
rlabel metal1 8418 31824 8418 31824 0 _0225_
rlabel metal1 22494 34476 22494 34476 0 _0226_
rlabel metal2 11730 34850 11730 34850 0 _0227_
rlabel metal2 13846 34442 13846 34442 0 _0228_
rlabel metal1 7084 34170 7084 34170 0 _0229_
rlabel metal1 17756 34578 17756 34578 0 _0230_
rlabel metal1 5842 33490 5842 33490 0 _0231_
rlabel metal2 31970 31620 31970 31620 0 _0232_
rlabel metal1 25530 34714 25530 34714 0 _0233_
rlabel metal1 21482 34714 21482 34714 0 _0234_
rlabel metal1 11086 34034 11086 34034 0 _0235_
rlabel metal1 22724 32334 22724 32334 0 _0236_
rlabel metal1 2990 32368 2990 32368 0 _0237_
rlabel metal1 14398 33082 14398 33082 0 _0238_
rlabel metal1 2254 32402 2254 32402 0 _0239_
rlabel metal1 17434 33082 17434 33082 0 _0240_
rlabel metal1 2254 30702 2254 30702 0 _0241_
rlabel metal1 27508 31314 27508 31314 0 _0242_
rlabel metal1 26588 33082 26588 33082 0 _0243_
rlabel metal1 22816 32402 22816 32402 0 _0244_
rlabel metal1 9338 31824 9338 31824 0 _0245_
rlabel metal1 27784 10234 27784 10234 0 _0246_
rlabel metal1 28566 6324 28566 6324 0 _0247_
rlabel metal2 33810 7140 33810 7140 0 _0248_
rlabel metal1 33718 9554 33718 9554 0 _0249_
rlabel metal1 32338 8466 32338 8466 0 _0250_
rlabel metal1 33442 10132 33442 10132 0 _0251_
rlabel metal2 33994 6528 33994 6528 0 _0252_
rlabel metal2 34270 9316 34270 9316 0 _0253_
rlabel metal1 33764 9690 33764 9690 0 _0254_
rlabel metal1 34546 7344 34546 7344 0 _0255_
rlabel metal1 30682 8942 30682 8942 0 _0256_
rlabel metal1 31464 5882 31464 5882 0 _0257_
rlabel metal2 33626 11084 33626 11084 0 _0258_
rlabel metal1 33442 9622 33442 9622 0 _0259_
rlabel metal2 33902 8398 33902 8398 0 _0260_
rlabel metal2 33902 10081 33902 10081 0 _0261_
rlabel metal1 34592 7446 34592 7446 0 _0262_
rlabel metal1 34086 7344 34086 7344 0 _0263_
rlabel metal1 32154 3366 32154 3366 0 _0264_
rlabel metal1 33442 7514 33442 7514 0 _0265_
rlabel metal1 32208 8602 32208 8602 0 _0266_
rlabel metal1 28382 7344 28382 7344 0 _0267_
rlabel viali 31648 7306 31648 7306 0 _0268_
rlabel metal1 32154 7242 32154 7242 0 _0269_
rlabel metal1 32338 7412 32338 7412 0 _0270_
rlabel metal2 31786 11577 31786 11577 0 _0271_
rlabel metal2 32062 11594 32062 11594 0 _0272_
rlabel metal2 32246 10880 32246 10880 0 _0273_
rlabel metal1 32614 9588 32614 9588 0 _0274_
rlabel metal1 31602 11764 31602 11764 0 _0275_
rlabel metal1 31924 9894 31924 9894 0 _0276_
rlabel metal2 31786 9724 31786 9724 0 _0277_
rlabel metal2 32384 7378 32384 7378 0 _0278_
rlabel metal2 31970 5508 31970 5508 0 _0279_
rlabel metal2 30774 7684 30774 7684 0 _0280_
rlabel metal1 30820 7922 30820 7922 0 _0281_
rlabel metal1 32039 10506 32039 10506 0 _0282_
rlabel metal2 28566 10778 28566 10778 0 _0283_
rlabel metal1 28566 10642 28566 10642 0 _0284_
rlabel metal2 27646 8228 27646 8228 0 _0285_
rlabel metal1 29343 10438 29343 10438 0 _0286_
rlabel metal1 29394 9962 29394 9962 0 _0287_
rlabel metal1 30314 7922 30314 7922 0 _0288_
rlabel metal1 30544 7922 30544 7922 0 _0289_
rlabel via1 30487 7786 30487 7786 0 _0290_
rlabel metal2 29486 6732 29486 6732 0 _0291_
rlabel metal2 30958 3264 30958 3264 0 _0292_
rlabel metal1 30912 4046 30912 4046 0 _0293_
rlabel metal1 31234 7174 31234 7174 0 _0294_
rlabel metal1 31280 7922 31280 7922 0 _0295_
rlabel metal1 29946 7922 29946 7922 0 _0296_
rlabel metal1 28014 8058 28014 8058 0 _0297_
rlabel metal2 27554 8126 27554 8126 0 _0298_
rlabel metal1 28060 7718 28060 7718 0 _0299_
rlabel metal2 26818 8806 26818 8806 0 _0300_
rlabel metal2 30314 11900 30314 11900 0 _0301_
rlabel metal2 31050 11050 31050 11050 0 _0302_
rlabel metal2 31878 9656 31878 9656 0 _0303_
rlabel metal2 27830 9690 27830 9690 0 _0304_
rlabel metal2 27922 9860 27922 9860 0 _0305_
rlabel metal2 29210 8670 29210 8670 0 _0306_
rlabel via1 27738 7990 27738 7990 0 _0307_
rlabel metal1 28382 7718 28382 7718 0 _0308_
rlabel metal2 30038 8058 30038 8058 0 _0309_
rlabel metal1 31556 4726 31556 4726 0 _0310_
rlabel metal2 31418 6460 31418 6460 0 _0311_
rlabel metal2 31878 6018 31878 6018 0 _0312_
rlabel metal1 31326 5695 31326 5695 0 _0313_
rlabel metal2 25898 5882 25898 5882 0 _0314_
rlabel metal2 25990 5508 25990 5508 0 _0315_
rlabel metal1 27002 5576 27002 5576 0 _0316_
rlabel metal1 26818 5712 26818 5712 0 _0317_
rlabel metal1 28014 5712 28014 5712 0 _0318_
rlabel metal1 27968 5542 27968 5542 0 _0319_
rlabel metal2 27370 8772 27370 8772 0 _0320_
rlabel metal2 27462 6834 27462 6834 0 _0321_
rlabel metal1 27692 5678 27692 5678 0 _0322_
rlabel metal1 30498 5848 30498 5848 0 _0323_
rlabel metal2 26036 2516 26036 2516 0 _0324_
rlabel metal1 31188 3570 31188 3570 0 _0325_
rlabel metal1 30682 2992 30682 2992 0 _0326_
rlabel metal1 29806 3502 29806 3502 0 _0327_
rlabel metal1 28014 4794 28014 4794 0 _0328_
rlabel metal2 25070 3638 25070 3638 0 _0329_
rlabel metal2 26726 4386 26726 4386 0 _0330_
rlabel metal2 26542 4284 26542 4284 0 _0331_
rlabel metal1 28934 4590 28934 4590 0 _0332_
rlabel metal1 28520 4522 28520 4522 0 _0333_
rlabel metal2 29762 3910 29762 3910 0 _0334_
rlabel metal1 32384 3502 32384 3502 0 _0335_
rlabel metal1 27370 3026 27370 3026 0 _0336_
rlabel metal2 25714 3332 25714 3332 0 _0337_
rlabel metal1 25898 2618 25898 2618 0 _0338_
rlabel metal1 26450 4080 26450 4080 0 _0339_
rlabel metal2 26266 4556 26266 4556 0 _0340_
rlabel metal1 25438 3978 25438 3978 0 _0341_
rlabel metal2 26174 3740 26174 3740 0 _0342_
rlabel metal1 28382 3502 28382 3502 0 _0343_
rlabel metal1 27048 3162 27048 3162 0 _0344_
rlabel metal1 27278 3570 27278 3570 0 _0345_
rlabel metal1 28198 3570 28198 3570 0 _0346_
rlabel metal1 32292 3434 32292 3434 0 _0347_
rlabel metal1 32016 2958 32016 2958 0 _0348_
rlabel metal1 31050 3162 31050 3162 0 _0349_
rlabel metal2 31602 3298 31602 3298 0 _0350_
rlabel metal1 21850 27472 21850 27472 0 _0351_
rlabel metal1 14536 26418 14536 26418 0 _0352_
rlabel metal1 14214 26554 14214 26554 0 _0353_
rlabel metal1 3588 26554 3588 26554 0 _0354_
rlabel metal2 17802 26554 17802 26554 0 _0355_
rlabel metal1 4140 27438 4140 27438 0 _0356_
rlabel metal2 27922 27642 27922 27642 0 _0357_
rlabel metal1 26174 26996 26174 26996 0 _0358_
rlabel metal1 21390 27642 21390 27642 0 _0359_
rlabel viali 10166 26347 10166 26347 0 _0360_
rlabel via2 21574 9707 21574 9707 0 _0361_
rlabel metal1 34960 18190 34960 18190 0 _0362_
rlabel metal1 18722 15538 18722 15538 0 _0363_
rlabel metal2 16790 15708 16790 15708 0 _0364_
rlabel metal1 12696 15674 12696 15674 0 _0365_
rlabel metal1 5980 14994 5980 14994 0 _0366_
rlabel metal2 16882 15300 16882 15300 0 _0367_
rlabel metal2 4002 14586 4002 14586 0 _0368_
rlabel metal2 27738 17000 27738 17000 0 _0369_
rlabel metal2 22862 16252 22862 16252 0 _0370_
rlabel metal1 19090 15470 19090 15470 0 _0371_
rlabel metal1 9062 15504 9062 15504 0 _0372_
rlabel metal2 19642 23290 19642 23290 0 _0373_
rlabel metal1 16376 21454 16376 21454 0 _0374_
rlabel metal2 12926 21692 12926 21692 0 _0375_
rlabel metal1 3726 20910 3726 20910 0 _0376_
rlabel metal2 15502 20876 15502 20876 0 _0377_
rlabel metal1 3450 23086 3450 23086 0 _0378_
rlabel metal1 29486 23086 29486 23086 0 _0379_
rlabel metal1 24196 23086 24196 23086 0 _0380_
rlabel metal2 18998 23290 18998 23290 0 _0381_
rlabel metal1 8510 21930 8510 21930 0 _0382_
rlabel metal1 19458 17170 19458 17170 0 _0383_
rlabel metal2 16422 16796 16422 16796 0 _0384_
rlabel metal1 12052 16558 12052 16558 0 _0385_
rlabel metal2 4830 16116 4830 16116 0 _0386_
rlabel metal1 15962 16082 15962 16082 0 _0387_
rlabel metal2 3082 15946 3082 15946 0 _0388_
rlabel metal2 26450 17374 26450 17374 0 _0389_
rlabel metal1 22908 17306 22908 17306 0 _0390_
rlabel metal2 18906 17476 18906 17476 0 _0391_
rlabel metal1 8556 16150 8556 16150 0 _0392_
rlabel metal1 21022 18360 21022 18360 0 _0393_
rlabel metal1 14674 17680 14674 17680 0 _0394_
rlabel metal2 13478 17340 13478 17340 0 _0395_
rlabel metal2 6578 16524 6578 16524 0 _0396_
rlabel metal1 17250 16558 17250 16558 0 _0397_
rlabel metal1 4324 17170 4324 17170 0 _0398_
rlabel metal1 29900 18938 29900 18938 0 _0399_
rlabel metal1 25070 17646 25070 17646 0 _0400_
rlabel metal1 21528 17170 21528 17170 0 _0401_
rlabel metal1 10442 17714 10442 17714 0 _0402_
rlabel metal2 23782 11526 23782 11526 0 _0403_
rlabel metal1 24196 11594 24196 11594 0 _0404_
rlabel metal2 34914 12036 34914 12036 0 _0405_
rlabel metal1 22034 11696 22034 11696 0 _0406_
rlabel metal2 24058 9316 24058 9316 0 _0407_
rlabel metal1 32338 25772 32338 25772 0 _0408_
rlabel metal1 9154 25296 9154 25296 0 _0409_
rlabel metal2 12466 26486 12466 26486 0 _0410_
rlabel metal1 4600 22746 4600 22746 0 _0411_
rlabel metal1 16422 25262 16422 25262 0 _0412_
rlabel metal1 4048 25262 4048 25262 0 _0413_
rlabel metal1 29440 24922 29440 24922 0 _0414_
rlabel metal1 24564 25466 24564 25466 0 _0415_
rlabel metal2 19918 26486 19918 26486 0 _0416_
rlabel metal1 9936 25330 9936 25330 0 _0417_
rlabel metal1 22494 36652 22494 36652 0 _0418_
rlabel metal1 29486 12206 29486 12206 0 _0419_
rlabel metal2 29762 35462 29762 35462 0 _0420_
rlabel metal2 17986 36550 17986 36550 0 _0421_
rlabel metal2 16698 36278 16698 36278 0 _0422_
rlabel metal1 21758 36754 21758 36754 0 _0423_
rlabel metal1 19366 36346 19366 36346 0 _0424_
rlabel metal1 24242 13498 24242 13498 0 _0425_
rlabel metal1 16560 3026 16560 3026 0 _0426_
rlabel metal1 34638 18190 34638 18190 0 _0427_
rlabel metal2 15318 8330 15318 8330 0 _0428_
rlabel metal1 14444 6766 14444 6766 0 _0429_
rlabel metal1 32752 22134 32752 22134 0 _0430_
rlabel metal1 22080 13498 22080 13498 0 _0431_
rlabel metal1 18906 13498 18906 13498 0 _0432_
rlabel metal2 20470 13770 20470 13770 0 _0433_
rlabel metal2 16790 10438 16790 10438 0 _0434_
rlabel metal2 33810 16388 33810 16388 0 _0435_
rlabel metal2 29762 15878 29762 15878 0 _0436_
rlabel metal1 32062 16082 32062 16082 0 _0437_
rlabel metal2 27186 14348 27186 14348 0 _0438_
rlabel metal2 33166 16864 33166 16864 0 _0439_
rlabel metal1 33028 20026 33028 20026 0 _0440_
rlabel metal2 30590 17306 30590 17306 0 _0441_
rlabel metal2 31418 18190 31418 18190 0 _0442_
rlabel metal1 32798 16218 32798 16218 0 _0443_
rlabel metal1 32384 24174 32384 24174 0 _0444_
rlabel metal2 33442 18734 33442 18734 0 _0445_
rlabel metal1 33626 22610 33626 22610 0 _0446_
rlabel metal1 14214 7854 14214 7854 0 _0447_
rlabel metal2 11362 7616 11362 7616 0 _0448_
rlabel metal2 11822 5610 11822 5610 0 _0449_
rlabel metal2 14122 11934 14122 11934 0 _0450_
rlabel metal1 10856 7854 10856 7854 0 _0451_
rlabel metal1 15134 8942 15134 8942 0 _0452_
rlabel metal1 11408 6766 11408 6766 0 _0453_
rlabel metal1 10488 6426 10488 6426 0 _0454_
rlabel metal1 10258 5338 10258 5338 0 _0455_
rlabel metal1 12742 5168 12742 5168 0 _0456_
rlabel metal2 12558 5474 12558 5474 0 _0457_
rlabel metal1 10350 6970 10350 6970 0 _0458_
rlabel metal1 11730 6970 11730 6970 0 _0459_
rlabel metal1 13846 9146 13846 9146 0 _0460_
rlabel metal2 14858 9350 14858 9350 0 _0461_
rlabel metal1 17434 6256 17434 6256 0 _0462_
rlabel metal2 20194 5542 20194 5542 0 _0463_
rlabel metal1 20838 6256 20838 6256 0 _0464_
rlabel via1 20656 5678 20656 5678 0 _0465_
rlabel metal1 17296 6290 17296 6290 0 _0466_
rlabel metal2 20010 6052 20010 6052 0 _0467_
rlabel metal2 16790 4930 16790 4930 0 _0468_
rlabel metal2 16974 4896 16974 4896 0 _0469_
rlabel metal1 18308 5678 18308 5678 0 _0470_
rlabel metal1 20516 5202 20516 5202 0 _0471_
rlabel metal2 21114 3264 21114 3264 0 _0472_
rlabel metal2 19918 6358 19918 6358 0 _0473_
rlabel metal1 21666 7276 21666 7276 0 _0474_
rlabel metal1 21114 7990 21114 7990 0 _0475_
rlabel metal1 17572 8058 17572 8058 0 _0476_
rlabel metal1 16790 8534 16790 8534 0 _0477_
rlabel metal1 13202 11764 13202 11764 0 _0478_
rlabel metal2 12006 11050 12006 11050 0 _0479_
rlabel metal1 11730 11696 11730 11696 0 _0480_
rlabel metal2 15226 8636 15226 8636 0 _0481_
rlabel metal2 19090 8126 19090 8126 0 _0482_
rlabel metal2 18998 6256 18998 6256 0 _0483_
rlabel metal1 18906 6358 18906 6358 0 _0484_
rlabel metal2 20470 7140 20470 7140 0 _0485_
rlabel metal1 21068 8466 21068 8466 0 _0486_
rlabel metal1 24932 10574 24932 10574 0 _0487_
rlabel metal1 21482 5780 21482 5780 0 _0488_
rlabel metal2 20884 7854 20884 7854 0 _0489_
rlabel metal2 21206 5882 21206 5882 0 _0490_
rlabel metal1 21206 5882 21206 5882 0 _0491_
rlabel metal2 21942 8500 21942 8500 0 _0492_
rlabel metal1 24656 10438 24656 10438 0 _0493_
rlabel metal2 22126 7106 22126 7106 0 _0494_
rlabel metal2 22218 7548 22218 7548 0 _0495_
rlabel metal1 21988 7446 21988 7446 0 _0496_
rlabel metal2 14582 14076 14582 14076 0 _0497_
rlabel metal1 14030 13940 14030 13940 0 _0498_
rlabel metal1 15088 13838 15088 13838 0 _0499_
rlabel metal2 14858 24548 14858 24548 0 _0500_
rlabel metal1 21942 20298 21942 20298 0 _0501_
rlabel metal2 20470 23698 20470 23698 0 _0502_
rlabel metal2 11638 26146 11638 26146 0 _0503_
rlabel metal2 13846 23766 13846 23766 0 _0504_
rlabel metal2 14490 24242 14490 24242 0 _0505_
rlabel metal1 15042 24786 15042 24786 0 _0506_
rlabel metal1 17296 32266 17296 32266 0 _0507_
rlabel metal1 16445 31790 16445 31790 0 _0508_
rlabel metal1 15180 27302 15180 27302 0 _0509_
rlabel metal2 18998 25024 18998 25024 0 _0510_
rlabel metal2 21390 26146 21390 26146 0 _0511_
rlabel metal1 17848 25806 17848 25806 0 _0512_
rlabel metal2 14674 25194 14674 25194 0 _0513_
rlabel metal1 13156 24786 13156 24786 0 _0514_
rlabel metal2 20286 19006 20286 19006 0 _0515_
rlabel metal1 5888 21454 5888 21454 0 _0516_
rlabel metal1 14398 18394 14398 18394 0 _0517_
rlabel metal1 14398 24752 14398 24752 0 _0518_
rlabel metal1 15180 25194 15180 25194 0 _0519_
rlabel metal2 20194 25296 20194 25296 0 _0520_
rlabel metal2 14490 24956 14490 24956 0 _0521_
rlabel metal1 22724 32946 22724 32946 0 _0522_
rlabel metal2 6670 31892 6670 31892 0 _0523_
rlabel metal1 8556 32198 8556 32198 0 _0524_
rlabel metal2 20838 25568 20838 25568 0 _0525_
rlabel metal2 7406 24922 7406 24922 0 _0526_
rlabel metal1 6532 23562 6532 23562 0 _0527_
rlabel metal1 7176 23834 7176 23834 0 _0528_
rlabel via2 10166 18139 10166 18139 0 _0529_
rlabel metal1 21988 18938 21988 18938 0 _0530_
rlabel metal1 7820 17850 7820 17850 0 _0531_
rlabel metal2 7682 25772 7682 25772 0 _0532_
rlabel metal2 7130 24378 7130 24378 0 _0533_
rlabel metal1 18216 23834 18216 23834 0 _0534_
rlabel metal1 18032 24378 18032 24378 0 _0535_
rlabel metal1 18630 32742 18630 32742 0 _0536_
rlabel metal1 18216 24718 18216 24718 0 _0537_
rlabel metal2 18538 21352 18538 21352 0 _0538_
rlabel metal2 18630 24514 18630 24514 0 _0539_
rlabel metal1 18860 26010 18860 26010 0 _0540_
rlabel metal1 17802 24786 17802 24786 0 _0541_
rlabel metal1 7406 31790 7406 31790 0 _0542_
rlabel metal1 7084 24786 7084 24786 0 _0543_
rlabel metal1 7222 23562 7222 23562 0 _0544_
rlabel metal2 7590 24242 7590 24242 0 _0545_
rlabel metal1 6302 18394 6302 18394 0 _0546_
rlabel metal2 6854 26656 6854 26656 0 _0547_
rlabel metal2 6670 25228 6670 25228 0 _0548_
rlabel metal1 26220 24378 26220 24378 0 _0549_
rlabel metal2 23782 24412 23782 24412 0 _0550_
rlabel metal1 23690 25874 23690 25874 0 _0551_
rlabel metal1 23644 24378 23644 24378 0 _0552_
rlabel metal2 23414 23511 23414 23511 0 _0553_
rlabel metal1 23506 23834 23506 23834 0 _0554_
rlabel metal2 29118 27914 29118 27914 0 _0555_
rlabel metal2 23506 25466 23506 25466 0 _0556_
rlabel metal2 25714 32521 25714 32521 0 _0557_
rlabel metal2 22954 25534 22954 25534 0 _0558_
rlabel metal2 24058 23800 24058 23800 0 _0559_
rlabel metal1 24150 23664 24150 23664 0 _0560_
rlabel metal1 25024 18394 25024 18394 0 _0561_
rlabel metal1 24656 24922 24656 24922 0 _0562_
rlabel metal1 22678 24854 22678 24854 0 _0563_
rlabel metal2 21666 24072 21666 24072 0 _0564_
rlabel metal2 21850 24582 21850 24582 0 _0565_
rlabel metal2 22218 32963 22218 32963 0 _0566_
rlabel metal1 21482 24718 21482 24718 0 _0567_
rlabel metal2 21482 19635 21482 19635 0 _0568_
rlabel metal2 21298 24548 21298 24548 0 _0569_
rlabel metal2 21298 26384 21298 26384 0 _0570_
rlabel metal2 21206 25534 21206 25534 0 _0571_
rlabel metal1 11868 31994 11868 31994 0 _0572_
rlabel metal2 10718 25466 10718 25466 0 _0573_
rlabel metal2 11730 23800 11730 23800 0 _0574_
rlabel metal1 11408 24378 11408 24378 0 _0575_
rlabel metal1 11270 18394 11270 18394 0 _0576_
rlabel metal1 11684 25194 11684 25194 0 _0577_
rlabel metal1 10488 25262 10488 25262 0 _0578_
rlabel metal1 24840 19414 24840 19414 0 _0579_
rlabel metal2 25254 32079 25254 32079 0 _0580_
rlabel via2 25898 19363 25898 19363 0 _0581_
rlabel metal2 25806 32096 25806 32096 0 _0582_
rlabel metal1 15410 20910 15410 20910 0 _0583_
rlabel metal2 19642 20638 19642 20638 0 _0584_
rlabel metal1 14674 20876 14674 20876 0 _0585_
rlabel metal2 14214 21182 14214 21182 0 _0586_
rlabel metal1 14398 19822 14398 19822 0 _0587_
rlabel metal2 19458 20808 19458 20808 0 _0588_
rlabel via1 20102 19669 20102 19669 0 _0589_
rlabel metal2 20194 20604 20194 20604 0 _0590_
rlabel metal1 14076 21046 14076 21046 0 _0591_
rlabel metal1 13892 20026 13892 20026 0 _0592_
rlabel metal1 8234 19788 8234 19788 0 _0593_
rlabel via2 20309 19380 20309 19380 0 _0594_
rlabel metal1 14214 19278 14214 19278 0 _0595_
rlabel metal1 14582 19482 14582 19482 0 _0596_
rlabel via2 17066 18819 17066 18819 0 _0597_
rlabel metal2 17618 18938 17618 18938 0 _0598_
rlabel metal1 14858 20570 14858 20570 0 _0599_
rlabel via2 21022 21437 21022 21437 0 _0600_
rlabel metal1 13754 19822 13754 19822 0 _0601_
rlabel metal1 9062 32742 9062 32742 0 _0602_
rlabel metal1 9108 19822 9108 19822 0 _0603_
rlabel metal1 7084 21046 7084 21046 0 _0604_
rlabel metal2 8510 20400 8510 20400 0 _0605_
rlabel metal2 8234 19414 8234 19414 0 _0606_
rlabel metal2 8786 23936 8786 23936 0 _0607_
rlabel metal2 8326 20026 8326 20026 0 _0608_
rlabel metal1 18630 20978 18630 20978 0 _0609_
rlabel metal2 17894 20434 17894 20434 0 _0610_
rlabel metal2 17158 21454 17158 21454 0 _0611_
rlabel metal1 17664 20230 17664 20230 0 _0612_
rlabel metal2 18262 19686 18262 19686 0 _0613_
rlabel metal1 18630 20570 18630 20570 0 _0614_
rlabel metal1 17526 20366 17526 20366 0 _0615_
rlabel metal1 19918 29002 19918 29002 0 _0616_
rlabel metal1 11362 32946 11362 32946 0 _0617_
rlabel metal1 7636 21658 7636 21658 0 _0618_
rlabel metal1 7452 20910 7452 20910 0 _0619_
rlabel metal1 6440 18938 6440 18938 0 _0620_
rlabel metal1 7038 20026 7038 20026 0 _0621_
rlabel via3 7245 21828 7245 21828 0 _0622_
rlabel metal1 17158 21488 17158 21488 0 _0623_
rlabel metal2 6946 21114 6946 21114 0 _0624_
rlabel metal2 6946 23630 6946 23630 0 _0625_
rlabel metal2 7038 21386 7038 21386 0 _0626_
rlabel metal1 26542 20978 26542 20978 0 _0627_
rlabel metal1 27370 20944 27370 20944 0 _0628_
rlabel metal1 27876 21046 27876 21046 0 _0629_
rlabel metal1 27600 21114 27600 21114 0 _0630_
rlabel metal2 29210 19720 29210 19720 0 _0631_
rlabel metal1 28934 20570 28934 20570 0 _0632_
rlabel metal2 28106 20672 28106 20672 0 _0633_
rlabel metal1 26864 32198 26864 32198 0 _0634_
rlabel metal1 24794 20434 24794 20434 0 _0635_
rlabel metal1 25852 23494 25852 23494 0 _0636_
rlabel metal1 24932 20230 24932 20230 0 _0637_
rlabel metal2 26266 19720 26266 19720 0 _0638_
rlabel metal1 25576 20570 25576 20570 0 _0639_
rlabel metal1 24426 20400 24426 20400 0 _0640_
rlabel metal1 21528 21386 21528 21386 0 _0641_
rlabel metal1 20562 20910 20562 20910 0 _0642_
rlabel metal1 21344 21522 21344 21522 0 _0643_
rlabel metal2 20378 21216 20378 21216 0 _0644_
rlabel metal2 21206 19346 21206 19346 0 _0645_
rlabel metal1 20378 20570 20378 20570 0 _0646_
rlabel metal1 20884 20910 20884 20910 0 _0647_
rlabel metal1 20194 20944 20194 20944 0 _0648_
rlabel metal1 11132 23494 11132 23494 0 _0649_
rlabel metal2 11270 20706 11270 20706 0 _0650_
rlabel metal2 11500 32742 11500 32742 0 _0651_
rlabel metal1 11454 20366 11454 20366 0 _0652_
rlabel metal2 11270 19448 11270 19448 0 _0653_
rlabel metal1 10948 20026 10948 20026 0 _0654_
rlabel metal1 12144 20910 12144 20910 0 _0655_
rlabel metal1 10994 20468 10994 20468 0 _0656_
rlabel metal1 21574 10132 21574 10132 0 _0657_
rlabel metal1 33672 16014 33672 16014 0 _0658_
rlabel metal1 19826 13294 19826 13294 0 _0659_
rlabel metal1 19826 14382 19826 14382 0 _0660_
rlabel metal2 22310 14790 22310 14790 0 _0661_
rlabel metal1 19780 14586 19780 14586 0 _0662_
rlabel metal2 20746 14552 20746 14552 0 _0663_
rlabel metal1 16836 11322 16836 11322 0 _0664_
rlabel metal1 21804 8466 21804 8466 0 _0665_
rlabel metal1 18124 13226 18124 13226 0 _0666_
rlabel metal1 23828 9554 23828 9554 0 _0667_
rlabel metal2 23598 9350 23598 9350 0 _0668_
rlabel metal2 32706 15776 32706 15776 0 _0669_
rlabel metal1 34316 17102 34316 17102 0 _0670_
rlabel metal2 33626 17476 33626 17476 0 _0671_
rlabel metal1 29716 16762 29716 16762 0 _0672_
rlabel metal1 32292 17306 32292 17306 0 _0673_
rlabel metal2 27002 15878 27002 15878 0 _0674_
rlabel metal1 33580 14926 33580 14926 0 _0675_
rlabel metal1 32200 12410 32200 12410 0 _0676_
rlabel metal2 32982 12614 32982 12614 0 _0677_
rlabel metal2 29118 13362 29118 13362 0 _0678_
rlabel metal1 29440 10642 29440 10642 0 _0679_
rlabel metal1 30866 13498 30866 13498 0 _0680_
rlabel metal2 25622 12988 25622 12988 0 _0681_
rlabel metal1 22954 7514 22954 7514 0 _0682_
rlabel metal2 21390 4420 21390 4420 0 _0683_
rlabel metal2 19642 3468 19642 3468 0 _0684_
rlabel metal1 25714 2414 25714 2414 0 _0685_
rlabel metal2 22862 3468 22862 3468 0 _0686_
rlabel viali 17706 3502 17706 3502 0 _0687_
rlabel metal1 33810 14892 33810 14892 0 _0688_
rlabel metal2 33258 14586 33258 14586 0 _0689_
rlabel metal1 29486 14042 29486 14042 0 _0690_
rlabel metal2 30774 14756 30774 14756 0 _0691_
rlabel metal1 27140 12410 27140 12410 0 _0692_
rlabel metal1 23736 5338 23736 5338 0 _0693_
rlabel metal1 21942 5338 21942 5338 0 _0694_
rlabel metal2 21850 3638 21850 3638 0 _0695_
rlabel metal2 20102 3196 20102 3196 0 _0696_
rlabel metal1 15318 5202 15318 5202 0 _0697_
rlabel metal1 16054 5644 16054 5644 0 _0698_
rlabel metal1 15870 5712 15870 5712 0 _0699_
rlabel metal1 11776 13294 11776 13294 0 _0700_
rlabel metal1 10672 14042 10672 14042 0 _0701_
rlabel metal1 10534 14416 10534 14416 0 _0702_
rlabel metal1 11868 13838 11868 13838 0 _0703_
rlabel metal2 13938 14178 13938 14178 0 _0704_
rlabel metal1 10488 13158 10488 13158 0 _0705_
rlabel metal1 9108 12410 9108 12410 0 _0706_
rlabel metal1 9292 12886 9292 12886 0 _0707_
rlabel metal2 10350 11390 10350 11390 0 _0708_
rlabel metal1 8142 12954 8142 12954 0 _0709_
rlabel metal1 8280 12206 8280 12206 0 _0710_
rlabel metal2 8970 11084 8970 11084 0 _0711_
rlabel metal1 8648 9554 8648 9554 0 _0712_
rlabel metal2 9430 11322 9430 11322 0 _0713_
rlabel metal2 9062 10370 9062 10370 0 _0714_
rlabel metal1 7958 7412 7958 7412 0 _0715_
rlabel via1 7590 7378 7590 7378 0 _0716_
rlabel metal2 8602 9690 8602 9690 0 _0717_
rlabel metal1 8372 6290 8372 6290 0 _0718_
rlabel metal2 8694 5508 8694 5508 0 _0719_
rlabel metal1 9154 5712 9154 5712 0 _0720_
rlabel metal1 9798 5202 9798 5202 0 _0721_
rlabel metal1 7866 5542 7866 5542 0 _0722_
rlabel metal1 7222 7922 7222 7922 0 _0723_
rlabel metal1 7130 7412 7130 7412 0 _0724_
rlabel metal2 7682 8058 7682 8058 0 _0725_
rlabel metal1 6578 6358 6578 6358 0 _0726_
rlabel metal1 8142 5848 8142 5848 0 _0727_
rlabel metal1 8878 5202 8878 5202 0 _0728_
rlabel metal1 4876 10030 4876 10030 0 _0729_
rlabel metal1 4232 9962 4232 9962 0 _0730_
rlabel metal1 5014 9962 5014 9962 0 _0731_
rlabel metal1 5750 6256 5750 6256 0 _0732_
rlabel metal1 5566 6630 5566 6630 0 _0733_
rlabel metal1 6164 6222 6164 6222 0 _0734_
rlabel metal1 5474 7854 5474 7854 0 _0735_
rlabel metal1 5796 12750 5796 12750 0 _0736_
rlabel metal2 5290 8330 5290 8330 0 _0737_
rlabel metal1 4646 7820 4646 7820 0 _0738_
rlabel metal1 4462 7888 4462 7888 0 _0739_
rlabel metal1 16054 12818 16054 12818 0 _0740_
rlabel metal1 18586 12206 18586 12206 0 _0741_
rlabel metal1 18032 12614 18032 12614 0 _0742_
rlabel metal1 18768 11866 18768 11866 0 _0743_
rlabel metal1 12834 9486 12834 9486 0 _0744_
rlabel metal1 14398 8432 14398 8432 0 _0745_
rlabel metal1 14582 10778 14582 10778 0 _0746_
rlabel metal2 14122 10914 14122 10914 0 _0747_
rlabel via2 11638 8925 11638 8925 0 _0748_
rlabel metal1 16790 11254 16790 11254 0 _0749_
rlabel metal1 13340 21862 13340 21862 0 _0750_
rlabel metal1 14030 17578 14030 17578 0 _0751_
rlabel metal1 30452 21930 30452 21930 0 _0752_
rlabel metal2 31878 26622 31878 26622 0 _0753_
rlabel metal1 32246 25228 32246 25228 0 _0754_
rlabel metal2 31142 27234 31142 27234 0 _0755_
rlabel metal1 30728 22066 30728 22066 0 _0756_
rlabel metal1 18814 30158 18814 30158 0 _0757_
rlabel metal1 17986 29648 17986 29648 0 _0758_
rlabel metal1 14214 29818 14214 29818 0 _0759_
rlabel metal1 13846 13872 13846 13872 0 _0760_
rlabel metal1 14076 12818 14076 12818 0 _0761_
rlabel metal1 13938 8602 13938 8602 0 _0762_
rlabel metal2 14030 12682 14030 12682 0 _0763_
rlabel metal1 14352 11866 14352 11866 0 _0764_
rlabel metal1 13754 12954 13754 12954 0 _0765_
rlabel metal1 13478 12750 13478 12750 0 _0766_
rlabel metal1 6762 14926 6762 14926 0 _0767_
rlabel metal1 7406 33830 7406 33830 0 _0768_
rlabel metal2 8050 30668 8050 30668 0 _0769_
rlabel metal1 12696 11866 12696 11866 0 _0770_
rlabel metal2 12374 14076 12374 14076 0 _0771_
rlabel metal1 11914 13906 11914 13906 0 _0772_
rlabel metal1 11500 12138 11500 12138 0 _0773_
rlabel metal1 11868 12342 11868 12342 0 _0774_
rlabel metal1 17434 12206 17434 12206 0 _0775_
rlabel metal1 16790 15334 16790 15334 0 _0776_
rlabel metal1 17388 17646 17388 17646 0 _0777_
rlabel metal1 17296 29818 17296 29818 0 _0778_
rlabel metal2 9614 10948 9614 10948 0 _0779_
rlabel metal1 9752 9486 9752 9486 0 _0780_
rlabel metal1 11822 9588 11822 9588 0 _0781_
rlabel metal1 11224 9078 11224 9078 0 _0782_
rlabel metal1 12052 9690 12052 9690 0 _0783_
rlabel metal1 12190 9928 12190 9928 0 _0784_
rlabel metal1 15916 12614 15916 12614 0 _0785_
rlabel metal1 4692 14994 4692 14994 0 _0786_
rlabel metal1 4784 19142 4784 19142 0 _0787_
rlabel metal2 5290 30226 5290 30226 0 _0788_
rlabel metal2 8418 13498 8418 13498 0 _0789_
rlabel metal1 8510 13226 8510 13226 0 _0790_
rlabel metal1 7682 13430 7682 13430 0 _0791_
rlabel metal1 7820 11730 7820 11730 0 _0792_
rlabel metal1 7544 10574 7544 10574 0 _0793_
rlabel metal1 7268 11322 7268 11322 0 _0794_
rlabel metal1 7222 10676 7222 10676 0 _0795_
rlabel metal2 7498 10948 7498 10948 0 _0796_
rlabel metal1 14122 11560 14122 11560 0 _0797_
rlabel metal1 14260 9486 14260 9486 0 _0798_
rlabel metal2 16146 11900 16146 11900 0 _0799_
rlabel metal1 16974 11526 16974 11526 0 _0800_
rlabel metal1 29072 17510 29072 17510 0 _0801_
rlabel metal1 30038 18734 30038 18734 0 _0802_
rlabel metal1 29486 29274 29486 29274 0 _0803_
rlabel metal2 7866 7820 7866 7820 0 _0804_
rlabel metal1 8326 7820 8326 7820 0 _0805_
rlabel metal1 8142 7888 8142 7888 0 _0806_
rlabel metal1 12098 7888 12098 7888 0 _0807_
rlabel metal1 13294 7514 13294 7514 0 _0808_
rlabel metal2 11914 8058 11914 8058 0 _0809_
rlabel metal2 13570 8092 13570 8092 0 _0810_
rlabel metal1 20746 11152 20746 11152 0 _0811_
rlabel metal1 24012 17238 24012 17238 0 _0812_
rlabel metal1 24518 34578 24518 34578 0 _0813_
rlabel metal1 25024 29274 25024 29274 0 _0814_
rlabel metal1 7176 7514 7176 7514 0 _0815_
rlabel metal1 6900 9894 6900 9894 0 _0816_
rlabel metal2 6394 8806 6394 8806 0 _0817_
rlabel metal1 7084 9418 7084 9418 0 _0818_
rlabel metal1 6486 10098 6486 10098 0 _0819_
rlabel metal1 10304 9350 10304 9350 0 _0820_
rlabel metal1 13570 10132 13570 10132 0 _0821_
rlabel metal1 18906 11322 18906 11322 0 _0822_
rlabel metal1 19366 17068 19366 17068 0 _0823_
rlabel metal2 21620 20230 21620 20230 0 _0824_
rlabel metal1 21528 30362 21528 30362 0 _0825_
rlabel metal1 5198 10676 5198 10676 0 _0826_
rlabel metal1 5842 10608 5842 10608 0 _0827_
rlabel metal1 5428 9554 5428 9554 0 _0828_
rlabel metal1 5474 9622 5474 9622 0 _0829_
rlabel metal1 6992 10506 6992 10506 0 _0830_
rlabel metal1 11408 8058 11408 8058 0 _0831_
rlabel metal2 10994 9860 10994 9860 0 _0832_
rlabel via2 10350 10659 10350 10659 0 _0833_
rlabel metal1 8740 16218 8740 16218 0 _0834_
rlabel metal2 10350 34680 10350 34680 0 _0835_
rlabel metal1 10350 29648 10350 29648 0 _0836_
rlabel metal1 12834 19482 12834 19482 0 _0837_
rlabel metal1 31970 26384 31970 26384 0 _0838_
rlabel metal1 30682 21998 30682 21998 0 _0839_
rlabel metal1 20194 28628 20194 28628 0 _0840_
rlabel metal1 16560 27982 16560 27982 0 _0841_
rlabel metal2 12558 28662 12558 28662 0 _0842_
rlabel metal2 2714 19516 2714 19516 0 _0843_
rlabel metal2 2898 27132 2898 27132 0 _0844_
rlabel metal2 16238 32640 16238 32640 0 _0845_
rlabel metal1 15732 28050 15732 28050 0 _0846_
rlabel metal2 2990 19805 2990 19805 0 _0847_
rlabel metal1 2346 28526 2346 28526 0 _0848_
rlabel metal1 28566 31790 28566 31790 0 _0849_
rlabel metal1 27416 30226 27416 30226 0 _0850_
rlabel metal1 24150 33388 24150 33388 0 _0851_
rlabel metal1 23276 28526 23276 28526 0 _0852_
rlabel metal1 22287 32402 22287 32402 0 _0853_
rlabel metal1 19504 28526 19504 28526 0 _0854_
rlabel metal1 9338 21522 9338 21522 0 _0855_
rlabel metal1 9200 28458 9200 28458 0 _0856_
rlabel metal2 32338 24106 32338 24106 0 _0857_
rlabel metal2 32982 25568 32982 25568 0 _0858_
rlabel metal2 32062 26860 32062 26860 0 _0859_
rlabel metal1 16790 29716 16790 29716 0 _0860_
rlabel metal1 12604 30226 12604 30226 0 _0861_
rlabel metal2 6210 29308 6210 29308 0 _0862_
rlabel metal1 16514 29818 16514 29818 0 _0863_
rlabel metal1 3956 29274 3956 29274 0 _0864_
rlabel metal1 31004 28730 31004 28730 0 _0865_
rlabel metal1 24196 30362 24196 30362 0 _0866_
rlabel metal2 19918 30838 19918 30838 0 _0867_
rlabel metal1 9476 29682 9476 29682 0 _0868_
rlabel metal2 31786 24772 31786 24772 0 _0869_
rlabel metal1 32614 22950 32614 22950 0 _0870_
rlabel metal1 22678 21454 22678 21454 0 _0871_
rlabel metal2 2714 22372 2714 22372 0 _0872_
rlabel metal1 14352 22202 14352 22202 0 _0873_
rlabel metal2 2070 20298 2070 20298 0 _0874_
rlabel metal1 17158 21114 17158 21114 0 _0875_
rlabel metal1 2070 23698 2070 23698 0 _0876_
rlabel metal1 27830 22746 27830 22746 0 _0877_
rlabel metal1 25714 22950 25714 22950 0 _0878_
rlabel metal1 21574 21658 21574 21658 0 _0879_
rlabel metal1 10074 21590 10074 21590 0 _0880_
rlabel metal1 15042 9690 15042 9690 0 _0881_
rlabel metal1 14030 10234 14030 10234 0 _0882_
rlabel metal2 11822 9316 11822 9316 0 _0883_
rlabel metal1 10028 7514 10028 7514 0 _0884_
rlabel metal2 12466 5508 12466 5508 0 _0885_
rlabel metal1 12604 5338 12604 5338 0 _0886_
rlabel metal1 10258 5644 10258 5644 0 _0887_
rlabel metal2 10350 7684 10350 7684 0 _0888_
rlabel metal1 34960 37230 34960 37230 0 clock
rlabel metal2 7406 38233 7406 38233 0 led_clock
rlabel metal1 13708 37094 13708 37094 0 leds[0]
rlabel metal2 23874 1520 23874 1520 0 leds[1]
rlabel metal3 820 15708 820 15708 0 leds[2]
rlabel metal3 820 34748 820 34748 0 leds[3]
rlabel metal2 19826 9775 19826 9775 0 net1
rlabel metal2 20194 36958 20194 36958 0 net10
rlabel metal1 32384 24718 32384 24718 0 net100
rlabel metal1 32338 24786 32338 24786 0 net101
rlabel metal2 21298 36822 21298 36822 0 net102
rlabel metal1 22816 36754 22816 36754 0 net103
rlabel metal2 19458 29954 19458 29954 0 net104
rlabel metal1 27002 31790 27002 31790 0 net105
rlabel metal1 29670 35530 29670 35530 0 net106
rlabel metal1 23828 37162 23828 37162 0 net107
rlabel metal2 29946 36754 29946 36754 0 net108
rlabel via2 30866 36125 30866 36125 0 net109
rlabel metal2 36294 11526 36294 11526 0 net11
rlabel metal1 36662 37162 36662 37162 0 net110
rlabel metal1 6292 4114 6292 4114 0 net12
rlabel metal1 9374 4114 9374 4114 0 net13
rlabel via1 1697 6358 1697 6358 0 net14
rlabel metal1 1426 3128 1426 3128 0 net15
rlabel metal1 18027 3026 18027 3026 0 net16
rlabel metal2 30130 36958 30130 36958 0 net17
rlabel metal1 35236 14994 35236 14994 0 net18
rlabel metal2 1610 23055 1610 23055 0 net19
rlabel metal2 2346 25398 2346 25398 0 net2
rlabel metal1 34868 2958 34868 2958 0 net20
rlabel metal1 18170 14790 18170 14790 0 net21
rlabel metal1 1426 22644 1426 22644 0 net22
rlabel metal1 21298 9452 21298 9452 0 net23
rlabel metal2 5842 8126 5842 8126 0 net24
rlabel metal2 12466 19618 12466 19618 0 net25
rlabel metal1 11868 15334 11868 15334 0 net26
rlabel metal1 30130 2414 30130 2414 0 net27
rlabel metal2 36202 36516 36202 36516 0 net28
rlabel metal2 10442 36924 10442 36924 0 net29
rlabel metal1 22701 2346 22701 2346 0 net3
rlabel metal1 4278 37196 4278 37196 0 net30
rlabel metal2 22310 37060 22310 37060 0 net31
rlabel metal2 20654 37026 20654 37026 0 net32
rlabel metal3 25783 36516 25783 36516 0 net33
rlabel metal1 15502 2414 15502 2414 0 net34
rlabel metal1 36110 33490 36110 33490 0 net35
rlabel metal1 35834 27438 35834 27438 0 net36
rlabel metal1 36202 20842 36202 20842 0 net37
rlabel metal1 31556 37162 31556 37162 0 net38
rlabel metal1 31096 10030 31096 10030 0 net39
rlabel metal1 5198 37230 5198 37230 0 net4
rlabel metal2 2254 2142 2254 2142 0 net40
rlabel metal2 1518 9112 1518 9112 0 net41
rlabel metal1 36386 30226 36386 30226 0 net42
rlabel metal1 11730 2448 11730 2448 0 net43
rlabel metal1 36156 24174 36156 24174 0 net44
rlabel metal2 6854 37060 6854 37060 0 net45
rlabel metal1 13248 37230 13248 37230 0 net46
rlabel metal1 23920 2414 23920 2414 0 net47
rlabel metal1 1656 16082 1656 16082 0 net48
rlabel metal2 2024 21556 2024 21556 0 net49
rlabel metal2 1840 19924 1840 19924 0 net5
rlabel metal2 12650 9078 12650 9078 0 net50
rlabel metal1 8004 12750 8004 12750 0 net51
rlabel metal2 15502 14212 15502 14212 0 net52
rlabel metal2 17342 14722 17342 14722 0 net53
rlabel metal1 4554 13294 4554 13294 0 net54
rlabel metal1 15364 13362 15364 13362 0 net55
rlabel metal1 31280 4590 31280 4590 0 net56
rlabel metal1 3128 2414 3128 2414 0 net57
rlabel metal2 21298 8704 21298 8704 0 net58
rlabel metal1 21942 5644 21942 5644 0 net59
rlabel metal1 20470 2618 20470 2618 0 net6
rlabel metal1 21758 8976 21758 8976 0 net60
rlabel metal1 33166 13362 33166 13362 0 net61
rlabel metal2 33350 14620 33350 14620 0 net62
rlabel metal1 18124 9894 18124 9894 0 net63
rlabel metal2 9338 4828 9338 4828 0 net64
rlabel metal1 1702 18734 1702 18734 0 net65
rlabel metal1 7406 16694 7406 16694 0 net66
rlabel metal1 4922 14382 4922 14382 0 net67
rlabel metal2 14858 19108 14858 19108 0 net68
rlabel metal1 16698 19312 16698 19312 0 net69
rlabel metal2 35926 2465 35926 2465 0 net7
rlabel metal1 14858 19278 14858 19278 0 net70
rlabel metal2 28566 4352 28566 4352 0 net71
rlabel metal2 19274 10302 19274 10302 0 net72
rlabel metal2 34730 6800 34730 6800 0 net73
rlabel metal2 22034 14501 22034 14501 0 net74
rlabel metal1 20104 16014 20104 16014 0 net75
rlabel metal1 22494 17612 22494 17612 0 net76
rlabel metal2 25898 17697 25898 17697 0 net77
rlabel metal2 32430 19040 32430 19040 0 net78
rlabel metal1 32890 16626 32890 16626 0 net79
rlabel metal1 28704 37230 28704 37230 0 net8
rlabel metal1 34638 12682 34638 12682 0 net80
rlabel metal1 34776 19754 34776 19754 0 net81
rlabel metal1 2162 21998 2162 21998 0 net82
rlabel metal1 1518 25228 1518 25228 0 net83
rlabel metal1 8924 22066 8924 22066 0 net84
rlabel metal1 15226 27404 15226 27404 0 net85
rlabel metal2 14996 20910 14996 20910 0 net86
rlabel metal2 15134 26316 15134 26316 0 net87
rlabel metal1 1610 31348 1610 31348 0 net88
rlabel metal1 9844 32334 9844 32334 0 net89
rlabel metal1 33028 2618 33028 2618 0 net9
rlabel metal1 4830 36142 4830 36142 0 net90
rlabel metal1 6992 36754 6992 36754 0 net91
rlabel metal1 11960 32402 11960 32402 0 net92
rlabel metal1 11914 34544 11914 34544 0 net93
rlabel metal1 17480 36006 17480 36006 0 net94
rlabel via1 15502 32861 15502 32861 0 net95
rlabel metal1 7130 36788 7130 36788 0 net96
rlabel metal1 18538 22474 18538 22474 0 net97
rlabel metal2 19366 25857 19366 25857 0 net98
rlabel metal1 33212 23086 33212 23086 0 net99
rlabel metal1 14490 14382 14490 14382 0 po_0._1_\[0\]
rlabel metal2 12558 14144 12558 14144 0 po_0._1_\[1\]
rlabel metal2 9430 13158 9430 13158 0 po_0._1_\[2\]
rlabel metal2 7406 12988 7406 12988 0 po_0._1_\[3\]
rlabel metal1 8188 14246 8188 14246 0 po_0._1_\[4\]
rlabel metal1 5934 7956 5934 7956 0 po_0._1_\[5\]
rlabel metal1 4278 10064 4278 10064 0 po_0._1_\[6\]
rlabel metal2 5474 12988 5474 12988 0 po_0._1_\[7\]
rlabel metal1 14950 10778 14950 10778 0 po_0.alu_0._10_\[0\]
rlabel metal2 13110 12546 13110 12546 0 po_0.alu_0._10_\[1\]
rlabel metal2 11638 11356 11638 11356 0 po_0.alu_0._10_\[2\]
rlabel metal1 9568 8466 9568 8466 0 po_0.alu_0._10_\[3\]
rlabel metal1 10994 5066 10994 5066 0 po_0.alu_0._10_\[4\]
rlabel metal1 9568 5338 9568 5338 0 po_0.alu_0._10_\[5\]
rlabel via2 9246 5763 9246 5763 0 po_0.alu_0._10_\[6\]
rlabel metal2 9890 7548 9890 7548 0 po_0.alu_0._10_\[7\]
rlabel metal1 15042 10234 15042 10234 0 po_0.alu_0._11_\[0\]
rlabel metal1 14214 11696 14214 11696 0 po_0.alu_0._11_\[1\]
rlabel metal2 12558 11526 12558 11526 0 po_0.alu_0._11_\[2\]
rlabel metal2 10442 8772 10442 8772 0 po_0.alu_0._11_\[3\]
rlabel metal1 12972 5882 12972 5882 0 po_0.alu_0._11_\[4\]
rlabel metal2 12834 6528 12834 6528 0 po_0.alu_0._11_\[5\]
rlabel metal1 10810 5882 10810 5882 0 po_0.alu_0._11_\[6\]
rlabel metal1 10764 8058 10764 8058 0 po_0.alu_0._11_\[7\]
rlabel metal1 14168 7310 14168 7310 0 po_0.alu_0.s0
rlabel metal1 14030 8500 14030 8500 0 po_0.alu_0.s1
rlabel metal1 33856 12954 33856 12954 0 po_0.muxf_0.rf_w_data\[0\]
rlabel metal2 14950 13022 14950 13022 0 po_0.muxf_0.rf_w_data\[1\]
rlabel metal2 18400 13804 18400 13804 0 po_0.muxf_0.rf_w_data\[2\]
rlabel metal1 15594 12784 15594 12784 0 po_0.muxf_0.rf_w_data\[3\]
rlabel metal1 22402 36754 22402 36754 0 po_0.muxf_0.rf_w_data\[4\]
rlabel metal1 19642 14450 19642 14450 0 po_0.muxf_0.rf_w_data\[5\]
rlabel metal2 21206 13804 21206 13804 0 po_0.muxf_0.rf_w_data\[6\]
rlabel metal1 18722 3366 18722 3366 0 po_0.muxf_0.rf_w_data\[7\]
rlabel metal1 18354 12750 18354 12750 0 po_0.muxf_0.s0
rlabel metal1 18860 12274 18860 12274 0 po_0.muxf_0.s1
rlabel metal2 13386 20230 13386 20230 0 po_0.regf_0._3_\[0\]
rlabel metal2 8142 17340 8142 17340 0 po_0.regf_0._3_\[1\]
rlabel metal1 17572 14994 17572 14994 0 po_0.regf_0._3_\[2\]
rlabel metal1 7360 20434 7360 20434 0 po_0.regf_0._3_\[3\]
rlabel metal1 26082 14382 26082 14382 0 po_0.regf_0._3_\[4\]
rlabel metal2 18446 14756 18446 14756 0 po_0.regf_0._3_\[5\]
rlabel metal1 19228 19346 19228 19346 0 po_0.regf_0._3_\[6\]
rlabel metal2 10810 17850 10810 17850 0 po_0.regf_0._3_\[7\]
rlabel metal1 14168 24582 14168 24582 0 po_0.regf_0._5_\[0\]
rlabel metal1 6992 13974 6992 13974 0 po_0.regf_0._5_\[1\]
rlabel metal1 16606 13498 16606 13498 0 po_0.regf_0._5_\[2\]
rlabel metal1 6348 24582 6348 24582 0 po_0.regf_0._5_\[3\]
rlabel metal2 17250 14824 17250 14824 0 po_0.regf_0._5_\[4\]
rlabel metal2 21114 12359 21114 12359 0 po_0.regf_0._5_\[5\]
rlabel metal2 20930 18173 20930 18173 0 po_0.regf_0._5_\[6\]
rlabel metal2 10028 17748 10028 17748 0 po_0.regf_0._5_\[7\]
rlabel metal2 13110 18768 13110 18768 0 po_0.regf_0.rf\[0\]\[0\]
rlabel metal1 6900 17102 6900 17102 0 po_0.regf_0.rf\[0\]\[1\]
rlabel metal1 17572 17510 17572 17510 0 po_0.regf_0.rf\[0\]\[2\]
rlabel metal2 4554 18496 4554 18496 0 po_0.regf_0.rf\[0\]\[3\]
rlabel metal1 30590 18734 30590 18734 0 po_0.regf_0.rf\[0\]\[4\]
rlabel metal1 24610 18700 24610 18700 0 po_0.regf_0.rf\[0\]\[5\]
rlabel metal1 19826 18190 19826 18190 0 po_0.regf_0.rf\[0\]\[6\]
rlabel metal2 10902 17476 10902 17476 0 po_0.regf_0.rf\[0\]\[7\]
rlabel metal1 13478 21998 13478 21998 0 po_0.regf_0.rf\[10\]\[0\]
rlabel via1 5670 20978 5670 20978 0 po_0.regf_0.rf\[10\]\[1\]
rlabel via1 17262 22066 17262 22066 0 po_0.regf_0.rf\[10\]\[2\]
rlabel metal1 4554 23494 4554 23494 0 po_0.regf_0.rf\[10\]\[3\]
rlabel via1 28026 23698 28026 23698 0 po_0.regf_0.rf\[10\]\[4\]
rlabel via1 25726 23698 25726 23698 0 po_0.regf_0.rf\[10\]\[5\]
rlabel metal1 20574 23630 20574 23630 0 po_0.regf_0.rf\[10\]\[6\]
rlabel metal1 9246 22576 9246 22576 0 po_0.regf_0.rf\[10\]\[7\]
rlabel metal1 13386 23630 13386 23630 0 po_0.regf_0.rf\[11\]\[0\]
rlabel via1 5290 21539 5290 21539 0 po_0.regf_0.rf\[11\]\[1\]
rlabel metal2 17618 23902 17618 23902 0 po_0.regf_0.rf\[11\]\[2\]
rlabel metal1 4646 24922 4646 24922 0 po_0.regf_0.rf\[11\]\[3\]
rlabel metal1 30452 24786 30452 24786 0 po_0.regf_0.rf\[11\]\[4\]
rlabel metal1 25254 25262 25254 25262 0 po_0.regf_0.rf\[11\]\[5\]
rlabel metal1 20562 26010 20562 26010 0 po_0.regf_0.rf\[11\]\[6\]
rlabel metal2 10442 23562 10442 23562 0 po_0.regf_0.rf\[11\]\[7\]
rlabel metal1 14950 32878 14950 32878 0 po_0.regf_0.rf\[12\]\[0\]
rlabel metal1 6762 32402 6762 32402 0 po_0.regf_0.rf\[12\]\[1\]
rlabel metal1 18354 32878 18354 32878 0 po_0.regf_0.rf\[12\]\[2\]
rlabel metal1 5566 30770 5566 30770 0 po_0.regf_0.rf\[12\]\[3\]
rlabel metal2 27922 31552 27922 31552 0 po_0.regf_0.rf\[12\]\[4\]
rlabel metal1 24702 32980 24702 32980 0 po_0.regf_0.rf\[12\]\[5\]
rlabel metal2 22310 33116 22310 33116 0 po_0.regf_0.rf\[12\]\[6\]
rlabel metal2 10258 32334 10258 32334 0 po_0.regf_0.rf\[12\]\[7\]
rlabel metal1 14720 34714 14720 34714 0 po_0.regf_0.rf\[13\]\[0\]
rlabel metal1 6670 32980 6670 32980 0 po_0.regf_0.rf\[13\]\[1\]
rlabel metal2 18722 34782 18722 34782 0 po_0.regf_0.rf\[13\]\[2\]
rlabel metal1 5428 31790 5428 31790 0 po_0.regf_0.rf\[13\]\[3\]
rlabel metal2 25162 30532 25162 30532 0 po_0.regf_0.rf\[13\]\[4\]
rlabel metal1 24610 32470 24610 32470 0 po_0.regf_0.rf\[13\]\[5\]
rlabel metal2 22126 33014 22126 33014 0 po_0.regf_0.rf\[13\]\[6\]
rlabel metal2 10074 32368 10074 32368 0 po_0.regf_0.rf\[13\]\[7\]
rlabel via1 14778 32402 14778 32402 0 po_0.regf_0.rf\[14\]\[0\]
rlabel metal2 4278 32640 4278 32640 0 po_0.regf_0.rf\[14\]\[1\]
rlabel metal2 16882 32640 16882 32640 0 po_0.regf_0.rf\[14\]\[2\]
rlabel via1 6498 31790 6498 31790 0 po_0.regf_0.rf\[14\]\[3\]
rlabel metal1 29164 31722 29164 31722 0 po_0.regf_0.rf\[14\]\[4\]
rlabel metal1 24472 32266 24472 32266 0 po_0.regf_0.rf\[14\]\[5\]
rlabel metal1 22862 32980 22862 32980 0 po_0.regf_0.rf\[14\]\[6\]
rlabel via1 11098 31858 11098 31858 0 po_0.regf_0.rf\[14\]\[7\]
rlabel metal2 13018 34204 13018 34204 0 po_0.regf_0.rf\[15\]\[0\]
rlabel metal1 7498 32946 7498 32946 0 po_0.regf_0.rf\[15\]\[1\]
rlabel metal2 16698 34204 16698 34204 0 po_0.regf_0.rf\[15\]\[2\]
rlabel metal1 5474 34714 5474 34714 0 po_0.regf_0.rf\[15\]\[3\]
rlabel metal1 30222 30804 30222 30804 0 po_0.regf_0.rf\[15\]\[4\]
rlabel metal2 24334 34816 24334 34816 0 po_0.regf_0.rf\[15\]\[5\]
rlabel metal2 22126 32640 22126 32640 0 po_0.regf_0.rf\[15\]\[6\]
rlabel metal2 10994 32368 10994 32368 0 po_0.regf_0.rf\[15\]\[7\]
rlabel metal1 12696 19346 12696 19346 0 po_0.regf_0.rf\[1\]\[0\]
rlabel metal1 6210 17714 6210 17714 0 po_0.regf_0.rf\[1\]\[1\]
rlabel metal1 16284 18938 16284 18938 0 po_0.regf_0.rf\[1\]\[2\]
rlabel metal1 3082 18938 3082 18938 0 po_0.regf_0.rf\[1\]\[3\]
rlabel metal2 28658 21318 28658 21318 0 po_0.regf_0.rf\[1\]\[4\]
rlabel metal1 24012 18734 24012 18734 0 po_0.regf_0.rf\[1\]\[5\]
rlabel metal1 19504 18734 19504 18734 0 po_0.regf_0.rf\[1\]\[6\]
rlabel metal2 9430 18972 9430 18972 0 po_0.regf_0.rf\[1\]\[7\]
rlabel via1 13950 18258 13950 18258 0 po_0.regf_0.rf\[2\]\[0\]
rlabel metal2 5750 15674 5750 15674 0 po_0.regf_0.rf\[2\]\[1\]
rlabel metal1 16560 16490 16560 16490 0 po_0.regf_0.rf\[2\]\[2\]
rlabel metal2 4186 16320 4186 16320 0 po_0.regf_0.rf\[2\]\[3\]
rlabel metal1 27600 17646 27600 17646 0 po_0.regf_0.rf\[2\]\[4\]
rlabel metal2 23874 18360 23874 18360 0 po_0.regf_0.rf\[2\]\[5\]
rlabel metal2 20654 17408 20654 17408 0 po_0.regf_0.rf\[2\]\[6\]
rlabel via1 10546 18258 10546 18258 0 po_0.regf_0.rf\[2\]\[7\]
rlabel metal2 13846 18768 13846 18768 0 po_0.regf_0.rf\[3\]\[0\]
rlabel metal2 6946 17952 6946 17952 0 po_0.regf_0.rf\[3\]\[1\]
rlabel metal2 16514 15232 16514 15232 0 po_0.regf_0.rf\[3\]\[2\]
rlabel metal1 4554 15062 4554 15062 0 po_0.regf_0.rf\[3\]\[3\]
rlabel metal2 28290 18938 28290 18938 0 po_0.regf_0.rf\[3\]\[4\]
rlabel metal2 23966 18428 23966 18428 0 po_0.regf_0.rf\[3\]\[5\]
rlabel metal2 20286 18428 20286 18428 0 po_0.regf_0.rf\[3\]\[6\]
rlabel via1 10442 18275 10442 18275 0 po_0.regf_0.rf\[3\]\[7\]
rlabel metal1 14122 28526 14122 28526 0 po_0.regf_0.rf\[4\]\[0\]
rlabel metal1 6946 26962 6946 26962 0 po_0.regf_0.rf\[4\]\[1\]
rlabel metal1 17112 27982 17112 27982 0 po_0.regf_0.rf\[4\]\[2\]
rlabel metal1 5198 28186 5198 28186 0 po_0.regf_0.rf\[4\]\[3\]
rlabel metal1 28842 28118 28842 28118 0 po_0.regf_0.rf\[4\]\[4\]
rlabel metal1 24150 27506 24150 27506 0 po_0.regf_0.rf\[4\]\[5\]
rlabel metal2 20746 28458 20746 28458 0 po_0.regf_0.rf\[4\]\[6\]
rlabel metal1 10350 27506 10350 27506 0 po_0.regf_0.rf\[4\]\[7\]
rlabel metal1 14536 29614 14536 29614 0 po_0.regf_0.rf\[5\]\[0\]
rlabel metal2 7406 31110 7406 31110 0 po_0.regf_0.rf\[5\]\[1\]
rlabel via1 17802 29563 17802 29563 0 po_0.regf_0.rf\[5\]\[2\]
rlabel metal1 5520 29614 5520 29614 0 po_0.regf_0.rf\[5\]\[3\]
rlabel metal2 29946 29376 29946 29376 0 po_0.regf_0.rf\[5\]\[4\]
rlabel metal2 25530 29376 25530 29376 0 po_0.regf_0.rf\[5\]\[5\]
rlabel metal1 20608 28526 20608 28526 0 po_0.regf_0.rf\[5\]\[6\]
rlabel metal1 10166 28526 10166 28526 0 po_0.regf_0.rf\[5\]\[7\]
rlabel metal1 14076 28662 14076 28662 0 po_0.regf_0.rf\[6\]\[0\]
rlabel metal1 3266 27336 3266 27336 0 po_0.regf_0.rf\[6\]\[1\]
rlabel via1 17906 28050 17906 28050 0 po_0.regf_0.rf\[6\]\[2\]
rlabel via1 6222 28526 6222 28526 0 po_0.regf_0.rf\[6\]\[3\]
rlabel metal1 28060 29818 28060 29818 0 po_0.regf_0.rf\[6\]\[4\]
rlabel metal1 24794 28934 24794 28934 0 po_0.regf_0.rf\[6\]\[5\]
rlabel metal2 19918 28730 19918 28730 0 po_0.regf_0.rf\[6\]\[6\]
rlabel metal2 9798 28356 9798 28356 0 po_0.regf_0.rf\[6\]\[7\]
rlabel metal1 13248 30362 13248 30362 0 po_0.regf_0.rf\[7\]\[0\]
rlabel metal2 7866 29376 7866 29376 0 po_0.regf_0.rf\[7\]\[1\]
rlabel metal2 16606 29852 16606 29852 0 po_0.regf_0.rf\[7\]\[2\]
rlabel metal1 6026 28594 6026 28594 0 po_0.regf_0.rf\[7\]\[3\]
rlabel metal2 31970 28730 31970 28730 0 po_0.regf_0.rf\[7\]\[4\]
rlabel metal1 24334 30226 24334 30226 0 po_0.regf_0.rf\[7\]\[5\]
rlabel metal2 20746 28866 20746 28866 0 po_0.regf_0.rf\[7\]\[6\]
rlabel metal2 11086 28526 11086 28526 0 po_0.regf_0.rf\[7\]\[7\]
rlabel metal1 14444 21998 14444 21998 0 po_0.regf_0.rf\[8\]\[0\]
rlabel metal2 2990 20740 2990 20740 0 po_0.regf_0.rf\[8\]\[1\]
rlabel metal1 17572 20910 17572 20910 0 po_0.regf_0.rf\[8\]\[2\]
rlabel metal2 2530 24072 2530 24072 0 po_0.regf_0.rf\[8\]\[3\]
rlabel metal1 27186 23732 27186 23732 0 po_0.regf_0.rf\[8\]\[4\]
rlabel metal2 26266 22576 26266 22576 0 po_0.regf_0.rf\[8\]\[5\]
rlabel metal1 20056 23154 20056 23154 0 po_0.regf_0.rf\[8\]\[6\]
rlabel metal1 10764 22066 10764 22066 0 po_0.regf_0.rf\[8\]\[7\]
rlabel metal2 13018 24378 13018 24378 0 po_0.regf_0.rf\[9\]\[0\]
rlabel metal1 4370 21420 4370 21420 0 po_0.regf_0.rf\[9\]\[1\]
rlabel metal1 16284 22950 16284 22950 0 po_0.regf_0.rf\[9\]\[2\]
rlabel metal2 2898 25670 2898 25670 0 po_0.regf_0.rf\[9\]\[3\]
rlabel metal2 28290 25024 28290 25024 0 po_0.regf_0.rf\[9\]\[4\]
rlabel metal2 27370 25670 27370 25670 0 po_0.regf_0.rf\[9\]\[5\]
rlabel metal2 20010 25024 20010 25024 0 po_0.regf_0.rf\[9\]\[6\]
rlabel metal1 9706 23698 9706 23698 0 po_0.regf_0.rf\[9\]\[7\]
rlabel metal1 34500 16762 34500 16762 0 po_0.regf_0.rp_addr\[0\]
rlabel metal1 30360 16218 30360 16218 0 po_0.regf_0.rp_addr\[1\]
rlabel metal1 32752 16762 32752 16762 0 po_0.regf_0.rp_addr\[2\]
rlabel metal2 27462 14790 27462 14790 0 po_0.regf_0.rp_addr\[3\]
rlabel metal1 25944 15334 25944 15334 0 po_0.regf_0.rp_rd
rlabel metal1 23046 14042 23046 14042 0 po_0.regf_0.rq_addr\[0\]
rlabel metal1 19504 14042 19504 14042 0 po_0.regf_0.rq_addr\[1\]
rlabel metal1 21114 14042 21114 14042 0 po_0.regf_0.rq_addr\[2\]
rlabel metal2 17158 10506 17158 10506 0 po_0.regf_0.rq_addr\[3\]
rlabel metal1 19504 9894 19504 9894 0 po_0.regf_0.rq_rd
rlabel metal1 32476 22610 32476 22610 0 po_0.regf_0.w_addr\[0\]
rlabel metal2 32338 22406 32338 22406 0 po_0.regf_0.w_addr\[1\]
rlabel metal1 33810 25262 33810 25262 0 po_0.regf_0.w_addr\[2\]
rlabel metal1 32798 23256 32798 23256 0 po_0.regf_0.w_addr\[3\]
rlabel metal1 32200 22610 32200 22610 0 po_0.regf_0.w_wr
rlabel metal2 36478 17119 36478 17119 0 reset
rlabel metal2 27186 10234 27186 10234 0 uc_0._00_
rlabel metal1 33626 9996 33626 9996 0 uc_0._01_
rlabel metal2 29210 8024 29210 8024 0 uc_0._02_
rlabel metal1 34132 10642 34132 10642 0 uc_0._21_\[0\]
rlabel metal1 33258 11764 33258 11764 0 uc_0._21_\[1\]
rlabel metal1 32246 11696 32246 11696 0 uc_0._21_\[2\]
rlabel metal1 12420 3944 12420 3944 0 uc_0._21_\[3\]
rlabel metal1 18538 4114 18538 4114 0 uc_0._21_\[4\]
rlabel metal1 24794 5678 24794 5678 0 uc_0._21_\[5\]
rlabel via2 4278 2907 4278 2907 0 uc_0._21_\[6\]
rlabel metal1 18860 3162 18860 3162 0 uc_0._21_\[7\]
rlabel metal1 33626 14348 33626 14348 0 uc_0.bc_0.358$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:960$35.$result\[0\]
rlabel metal1 29854 14348 29854 14348 0 uc_0.bc_0.358$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:960$35.$result\[1\]
rlabel metal2 31878 14586 31878 14586 0 uc_0.bc_0.358$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:960$35.$result\[2\]
rlabel metal2 27278 12988 27278 12988 0 uc_0.bc_0.358$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:960$35.$result\[3\]
rlabel metal1 23598 5678 23598 5678 0 uc_0.bc_0.358$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:960$35.$result\[4\]
rlabel via1 22217 5678 22217 5678 0 uc_0.bc_0.358$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:960$35.$result\[5\]
rlabel metal2 21574 3706 21574 3706 0 uc_0.bc_0.358$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:960$35.$result\[6\]
rlabel metal1 20470 3060 20470 3060 0 uc_0.bc_0.358$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:960$35.$result\[7\]
rlabel metal1 33350 12852 33350 12852 0 uc_0.bc_0.359$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:987$36.$result\[0\]
rlabel metal1 28704 13498 28704 13498 0 uc_0.bc_0.359$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:987$36.$result\[1\]
rlabel metal1 31142 13940 31142 13940 0 uc_0.bc_0.359$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:987$36.$result\[2\]
rlabel metal1 25990 12852 25990 12852 0 uc_0.bc_0.359$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:987$36.$result\[3\]
rlabel metal1 23138 7820 23138 7820 0 uc_0.bc_0.359$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:987$36.$result\[4\]
rlabel metal2 19458 3332 19458 3332 0 uc_0.bc_0.359$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:987$36.$result\[5\]
rlabel metal2 22678 3332 22678 3332 0 uc_0.bc_0.359$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:987$36.$result\[6\]
rlabel via2 18078 3485 18078 3485 0 uc_0.bc_0.359$func$\/openlane\/designs\/vahid6i\/src\/vahid6i.v:987$36.$result\[7\]
rlabel metal1 18538 7820 18538 7820 0 uc_0.bc_0._12_\[0\]
rlabel metal1 16974 5814 16974 5814 0 uc_0.bc_0._12_\[1\]
rlabel metal2 18446 7786 18446 7786 0 uc_0.bc_0._12_\[2\]
rlabel metal2 18906 8840 18906 8840 0 uc_0.bc_0._12_\[3\]
rlabel metal1 34178 16150 34178 16150 0 uc_0.bc_0._14_\[0\]
rlabel metal1 30590 16490 30590 16490 0 uc_0.bc_0._14_\[1\]
rlabel metal2 32614 15130 32614 15130 0 uc_0.bc_0._14_\[2\]
rlabel metal2 27554 14858 27554 14858 0 uc_0.bc_0._14_\[3\]
rlabel metal2 24242 6052 24242 6052 0 uc_0.bc_0._14_\[4\]
rlabel metal2 22586 6086 22586 6086 0 uc_0.bc_0._14_\[5\]
rlabel metal2 22034 3434 22034 3434 0 uc_0.bc_0._14_\[6\]
rlabel metal2 20838 3264 20838 3264 0 uc_0.bc_0._14_\[7\]
rlabel metal2 20930 9248 20930 9248 0 uc_0.bc_0._85_\[0\]
rlabel metal1 18487 7446 18487 7446 0 uc_0.bc_0._85_\[1\]
rlabel metal2 21114 8058 21114 8058 0 uc_0.bc_0._85_\[2\]
rlabel metal1 20930 9486 20930 9486 0 uc_0.bc_0._85_\[3\]
<< properties >>
string FIXED_BBOX 0 0 37936 40080
<< end >>
