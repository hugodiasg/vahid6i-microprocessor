* NGSPICE file created from vahid6i.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_2 abstract view
.subckt sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt vahid6i D_R_data[0] D_R_data[1] D_R_data[2] D_R_data[3] D_R_data[4] D_R_data[5]
+ D_R_data[6] D_R_data[7] D_W_data[0] D_W_data[1] D_W_data[2] D_W_data[3] D_W_data[4]
+ D_W_data[5] D_W_data[6] D_W_data[7] D_addr[0] D_addr[1] D_addr[2] D_addr[3] D_addr[4]
+ D_addr[5] D_addr[6] D_addr[7] D_rd D_wr I_addr[0] I_addr[1] I_addr[2] I_addr[3]
+ I_addr[4] I_addr[5] I_addr[6] I_addr[7] I_data[0] I_data[1] I_data[2] I_data[3]
+ I_data[4] I_data[5] I_data[6] I_data[7] I_rd VGND VPWR clock led_clock leds[0] leds[1]
+ leds[2] leds[3] reset
XFILLER_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2037_ net99 _0183_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1270_ _0760_ _0704_ _0498_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__o21bai_1
XFILLER_44_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0985_ _0004_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__clkbuf_4
X_1606_ _0316_ _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__or2_1
XFILLER_59_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1468_ _0212_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
Xfanout105 net106 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlymetal6s2s_1
X_1399_ po_0.regf_0.w_addr\[0\] VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__buf_2
X_1537_ _0252_ _0253_ _0250_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
XFILLER_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1253_ _0479_ _0450_ _0447_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__or3_1
X_1322_ net6 _0741_ _0743_ po_0.muxf_0.rf_w_data\[5\] VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__a22oi_1
XFILLER_49_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1184_ uc_0.bc_0._14_\[4\] uc_0._21_\[4\] _0688_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__mux2_1
X_0968_ _0509_ _0511_ _0512_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__a21bo_1
X_0899_ _0455_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1871_ net82 _0049_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1940_ net64 net15 VGND VGND VPWR VPWR uc_0._21_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1236_ _0731_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__clkbuf_2
X_1305_ _0710_ po_0._1_\[2\] _0480_ _0792_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a31o_1
XFILLER_64_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1098_ po_0.regf_0.rf\[0\]\[4\] po_0.regf_0.rf\[1\]\[4\] po_0.regf_0.rf\[2\]\[4\]
+ po_0.regf_0.rf\[3\]\[4\] _0597_ _0598_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__mux4_1
X_1167_ uc_0._21_\[5\] VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__clkbuf_2
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1021_ po_0.regf_0.rf\[0\]\[5\] po_0.regf_0.rf\[1\]\[5\] po_0.regf_0.rf\[2\]\[5\]
+ po_0.regf_0.rf\[3\]\[5\] _0529_ _0530_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__mux4_1
X_1854_ net106 _0036_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1923_ net71 _0101_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dfxtp_1
X_1785_ _0429_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1219_ po_0._1_\[3\] net51 VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__or2b_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_5 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1570_ uc_0._21_\[3\] net40 _0271_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__o21ai_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1004_ po_0.regf_0.rf\[0\]\[3\] po_0.regf_0.rf\[1\]\[3\] po_0.regf_0.rf\[2\]\[3\]
+ po_0.regf_0.rf\[3\]\[3\] _0529_ _0530_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__mux4_1
XFILLER_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1768_ _0421_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
X_1906_ net105 _0084_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1837_ po_0.regf_0._3_\[3\] net52 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlxtp_1
XFILLER_57_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1699_ po_0.regf_0.w_addr\[0\] _0752_ po_0.regf_0.w_wr _0194_ VGND VGND VPWR VPWR
+ _0383_ sky130_fd_sc_hd__and4b_2
XFILLER_1_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput31 net31 VGND VGND VPWR VPWR D_addr[4] sky130_fd_sc_hd__buf_2
Xoutput42 net42 VGND VGND VPWR VPWR I_addr[5] sky130_fd_sc_hd__buf_2
Xoutput20 net20 VGND VGND VPWR VPWR D_W_data[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1622_ _0330_ _0331_ _0321_ _0319_ _0317_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__a221o_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1484_ _0221_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1553_ _0250_ _0255_ _0266_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a21oi_1
X_2036_ net100 _0182_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0984_ _0514_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__and2b_1
X_1605_ _0292_ uc_0._21_\[4\] _0314_ _0315_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__o22a_1
X_1536_ uc_0._01_ uc_0._00_ uc_0._02_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__nor3_2
Xfanout106 net107 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1467_ _0802_ po_0.regf_0.rf\[15\]\[4\] _0206_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__mux2_1
X_1398_ _0860_ _0835_ _0868_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2019_ _2019_/D net58 VGND VGND VPWR VPWR uc_0.bc_0._14_\[6\] sky130_fd_sc_hd__dlxtn_1
XFILLER_12_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1321_ _0807_ _0809_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__nand2_1
X_1252_ po_0.alu_0._10_\[0\] po_0.alu_0._11_\[0\] _0745_ VGND VGND VPWR VPWR _0746_
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1183_ _0692_ VGND VGND VPWR VPWR _2016_/D sky130_fd_sc_hd__clkbuf_1
X_0967_ _0007_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__clkbuf_2
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1519_ po_0.regf_0.rf\[12\]\[3\] _0847_ _0237_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__mux2_1
X_0898_ _0449_ _0453_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__or2b_1
XFILLER_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1870_ net85 _0048_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1166_ _0682_ VGND VGND VPWR VPWR _1999_/D sky130_fd_sc_hd__clkbuf_1
X_1235_ _0729_ _0730_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__or2_1
X_1304_ _0480_ _0710_ po_0._1_\[2\] _0792_ _0793_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__a311o_1
XFILLER_60_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1097_ _0600_ _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__and2b_1
X_1999_ _1999_/D net59 VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[4\] sky130_fd_sc_hd__dlxtn_2
XFILLER_47_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1020_ _0500_ _0559_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__and2b_1
XFILLER_19_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1922_ net72 _0100_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_1
X_1853_ net88 _0035_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1784_ _0448_ _0464_ _0659_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__mux2_1
X_1149_ _0672_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__clkbuf_1
X_1218_ net50 po_0._1_\[4\] VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__nor2_1
XFILLER_43_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1003_ _0514_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__and2b_1
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1905_ net90 _0083_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1767_ po_0.muxf_0.rf_w_data\[2\] net29 _0418_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux2_1
X_1698_ _0834_ _0374_ _0382_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__a21oi_1
X_1836_ po_0.regf_0._3_\[2\] net53 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlxtp_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput32 net32 VGND VGND VPWR VPWR D_addr[5] sky130_fd_sc_hd__buf_2
Xoutput43 net43 VGND VGND VPWR VPWR I_addr[6] sky130_fd_sc_hd__buf_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput21 net21 VGND VGND VPWR VPWR D_W_data[2] sky130_fd_sc_hd__buf_2
XFILLER_0_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1621_ _0317_ _0328_ _0330_ _0331_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__o211ai_1
XFILLER_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1552_ _0247_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__inv_2
X_1483_ po_0.regf_0.rf\[14\]\[3\] _0847_ _0217_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__mux2_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2035_ net79 _0181_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1819_ net88 _0017_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0983_ po_0.regf_0.rf\[8\]\[1\] po_0.regf_0.rf\[9\]\[1\] po_0.regf_0.rf\[10\]\[1\]
+ po_0.regf_0.rf\[11\]\[1\] _0515_ _0516_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__mux4_1
Xfanout107 net108 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlymetal6s2s_1
X_1604_ _0292_ uc_0._21_\[4\] _0314_ _0315_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__nor4_1
X_1535_ _0247_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__clkbuf_2
X_1466_ _0211_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
X_1397_ _0860_ po_0.regf_0.rf\[7\]\[7\] VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__nand2_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2018_ _2018_/D net59 VGND VGND VPWR VPWR uc_0.bc_0._14_\[5\] sky130_fd_sc_hd__dlxtn_1
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1320_ net24 _0451_ _0447_ _0808_ _0748_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__o311a_1
X_1251_ po_0.alu_0.s1 po_0.alu_0.s0 VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__nand2b_2
X_1182_ uc_0.bc_0._14_\[3\] uc_0._21_\[3\] _0688_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__mux2_1
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0966_ _0510_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__clkbuf_2
XFILLER_32_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0897_ _0454_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1518_ _0240_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
X_1449_ _0201_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1303_ _0715_ _0716_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__nor2_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1096_ po_0.regf_0.rf\[8\]\[4\] po_0.regf_0.rf\[9\]\[4\] po_0.regf_0.rf\[10\]\[4\]
+ po_0.regf_0.rf\[11\]\[4\] _0594_ _0595_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__mux4_1
X_1165_ po_0.muxf_0.rf_w_data\[4\] uc_0._21_\[4\] _0676_ VGND VGND VPWR VPWR _0682_
+ sky130_fd_sc_hd__mux2_1
X_1234_ net25 po_0._1_\[6\] VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__nor2_1
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0949_ _0494_ _0495_ _0475_ _0482_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__o31a_2
X_1998_ _1998_/D net61 VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[3\] sky130_fd_sc_hd__dlxtn_2
XFILLER_20_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1852_ net95 _0034_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1921_ net71 _0099_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_2
X_1783_ _0428_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1079_ po_0.regf_0.rf\[4\]\[2\] po_0.regf_0.rf\[5\]\[2\] po_0.regf_0.rf\[6\]\[2\]
+ po_0.regf_0.rf\[7\]\[2\] _0597_ _0598_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__mux4_1
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1148_ po_0.regf_0.rp_addr\[1\] uc_0.bc_0._14_\[1\] _0670_ VGND VGND VPWR VPWR _0672_
+ sky130_fd_sc_hd__mux2_1
X_1217_ net50 po_0._1_\[4\] VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__and2_1
XFILLER_40_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1002_ po_0.regf_0.rf\[8\]\[3\] po_0.regf_0.rf\[9\]\[3\] po_0.regf_0.rf\[10\]\[3\]
+ po_0.regf_0.rf\[11\]\[3\] _0515_ _0516_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__mux4_1
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1904_ net93 _0082_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1835_ po_0.regf_0._3_\[1\] net52 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlxtp_1
X_1766_ _0420_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
X_1697_ po_0.regf_0.rf\[10\]\[7\] _0374_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__nor2_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput33 net33 VGND VGND VPWR VPWR D_addr[6] sky130_fd_sc_hd__buf_2
Xoutput44 net44 VGND VGND VPWR VPWR I_addr[7] sky130_fd_sc_hd__buf_2
Xoutput22 net22 VGND VGND VPWR VPWR D_W_data[3] sky130_fd_sc_hd__buf_2
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1482_ _0220_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
X_1620_ net56 _0683_ _0329_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__or3_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1551_ net57 VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ net99 _0180_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[0\] sky130_fd_sc_hd__dfxtp_1
X_1818_ net92 _0016_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1749_ _0411_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0982_ _0524_ _0525_ _0007_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout108 net109 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlymetal6s2s_1
X_1465_ _0787_ po_0.regf_0.rf\[15\]\[3\] _0207_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__mux2_1
X_1603_ net56 uc_0._21_\[5\] VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__and2_1
X_1534_ _0250_ _0675_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__xnor2_1
X_1396_ _0867_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
X_2017_ _2017_/D net59 VGND VGND VPWR VPWR uc_0.bc_0._14_\[4\] sky130_fd_sc_hd__dlxtn_1
XFILLER_50_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1181_ _0691_ VGND VGND VPWR VPWR _2015_/D sky130_fd_sc_hd__clkbuf_1
X_1250_ _0450_ _0447_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__nor2_2
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0965_ _0006_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__buf_2
X_0896_ _0449_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__or2b_1
X_1517_ po_0.regf_0.rf\[12\]\[2\] _0845_ _0237_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_1
X_1448_ po_0.regf_0.rf\[1\]\[4\] _0849_ _0195_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_1
X_1379_ po_0.regf_0.w_addr\[0\] po_0.regf_0.w_addr\[1\] po_0.regf_0.w_wr VGND VGND
+ VPWR VPWR _0857_ sky130_fd_sc_hd__nand3_1
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout90 net91 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1233_ net25 po_0._1_\[6\] VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__and2_1
X_1302_ net51 po_0._1_\[3\] VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__and2_1
XFILLER_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1095_ _0627_ _0585_ _0003_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__a21bo_1
X_1164_ _0681_ VGND VGND VPWR VPWR _1998_/D sky130_fd_sc_hd__clkbuf_1
X_0948_ _0464_ uc_0.bc_0._14_\[6\] VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__nor2_1
X_1997_ _1997_/D net61 VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[2\] sky130_fd_sc_hd__dlxtn_2
XFILLER_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1851_ net89 _0033_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1920_ net71 _0098_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_1
X_1782_ _0452_ uc_0.bc_0._85_\[1\] _0660_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__mux2_1
X_1216_ _0712_ _0714_ VGND VGND VPWR VPWR po_0.alu_0._10_\[3\] sky130_fd_sc_hd__xor2_1
XFILLER_52_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1078_ po_0.regf_0.rf\[0\]\[2\] po_0.regf_0.rf\[1\]\[2\] po_0.regf_0.rf\[2\]\[2\]
+ po_0.regf_0.rf\[3\]\[2\] _0597_ _0598_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__mux4_1
X_1147_ _0671_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _0542_ _0525_ _0007_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__a21bo_1
XFILLER_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1765_ po_0.muxf_0.rf_w_data\[1\] net28 _0418_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__mux2_1
X_1903_ net91 _0081_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1834_ po_0.regf_0._3_\[0\] net52 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlxtp_1
X_1696_ _0381_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput34 net34 VGND VGND VPWR VPWR D_addr[7] sky130_fd_sc_hd__buf_2
Xoutput23 net23 VGND VGND VPWR VPWR D_W_data[4] sky130_fd_sc_hd__buf_2
Xoutput45 net45 VGND VGND VPWR VPWR led_clock sky130_fd_sc_hd__buf_2
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1481_ po_0.regf_0.rf\[14\]\[2\] _0845_ _0217_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__mux2_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1550_ _0255_ _0257_ _0265_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__o21a_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2033_ net77 _0179_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1748_ _0768_ po_0.regf_0.rf\[11\]\[1\] _0409_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux2_1
X_1817_ _0446_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
X_1679_ po_0.regf_0.rf\[3\]\[7\] _0364_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__nor2_1
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0981_ _0510_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__clkbuf_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1602_ net56 _0683_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__nor2_1
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout109 net17 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
X_1464_ _0210_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
X_1395_ _0824_ po_0.regf_0.rf\[7\]\[6\] _0859_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__mux2_1
X_1533_ _0249_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__clkbuf_2
X_2016_ _2016_/D net61 VGND VGND VPWR VPWR uc_0.bc_0._14_\[3\] sky130_fd_sc_hd__dlxtn_1
XFILLER_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1180_ uc_0.bc_0._14_\[2\] _0679_ _0688_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__mux2_1
X_0964_ po_0.regf_0.rf\[12\]\[0\] po_0.regf_0.rf\[13\]\[0\] po_0.regf_0.rf\[14\]\[0\]
+ po_0.regf_0.rf\[15\]\[0\] _0507_ _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__mux4_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1516_ _0239_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
X_0895_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1378_ _0855_ _0841_ _0856_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__a21oi_1
X_1447_ _0200_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout91 net96 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout80 net81 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1232_ _0728_ VGND VGND VPWR VPWR po_0.alu_0._10_\[5\] sky130_fd_sc_hd__clkbuf_1
X_1301_ _0763_ _0789_ _0790_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1094_ po_0.regf_0.rf\[12\]\[4\] po_0.regf_0.rf\[13\]\[4\] po_0.regf_0.rf\[14\]\[4\]
+ po_0.regf_0.rf\[15\]\[4\] _0580_ _0582_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__mux4_1
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1163_ po_0.muxf_0.rf_w_data\[3\] uc_0._21_\[3\] _0676_ VGND VGND VPWR VPWR _0681_
+ sky130_fd_sc_hd__mux2_1
X_0947_ _0464_ uc_0.bc_0._14_\[6\] uc_0.bc_0._14_\[7\] VGND VGND VPWR VPWR _0494_
+ sky130_fd_sc_hd__a21o_1
X_1996_ _1996_/D net61 VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[1\] sky130_fd_sc_hd__dlxtn_2
XFILLER_50_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1850_ net92 _0032_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1781_ _0362_ net36 _0427_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__a21bo_1
XFILLER_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1146_ po_0.regf_0.rp_addr\[0\] uc_0.bc_0._14_\[0\] _0670_ VGND VGND VPWR VPWR _0671_
+ sky130_fd_sc_hd__mux2_1
X_1215_ _0705_ _0708_ _0713_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1077_ _0588_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__and2b_1
XFILLER_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1979_ net74 _0145_ VGND VGND VPWR VPWR po_0.muxf_0.s1 sky130_fd_sc_hd__dfxtp_1
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1000_ po_0.regf_0.rf\[12\]\[3\] po_0.regf_0.rf\[13\]\[3\] po_0.regf_0.rf\[14\]\[3\]
+ po_0.regf_0.rf\[15\]\[3\] _0522_ _0523_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__mux4_1
X_1902_ net93 _0080_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1764_ _0419_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
X_1833_ po_0.regf_0._5_\[7\] net54 VGND VGND VPWR VPWR po_0._1_\[7\] sky130_fd_sc_hd__dlxtp_1
X_1695_ po_0.regf_0.rf\[10\]\[6\] _0823_ _0373_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__mux2_1
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1129_ _0657_ _0492_ uc_0.bc_0._85_\[3\] VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__and3_2
XFILLER_31_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput46 net46 VGND VGND VPWR VPWR leds[0] sky130_fd_sc_hd__buf_2
Xoutput35 net35 VGND VGND VPWR VPWR D_rd sky130_fd_sc_hd__buf_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput24 net24 VGND VGND VPWR VPWR D_W_data[5] sky130_fd_sc_hd__buf_2
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1480_ _0219_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2032_ net79 _0178_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1747_ _0410_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
X_1816_ _0754_ _0445_ _0430_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__mux2_1
X_1678_ _0371_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0980_ po_0.regf_0.rf\[12\]\[1\] po_0.regf_0.rf\[13\]\[1\] po_0.regf_0.rf\[14\]\[1\]
+ po_0.regf_0.rf\[15\]\[1\] _0522_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__mux4_1
X_1601_ _0311_ _0252_ _0312_ _0264_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__a31o_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1532_ net37 VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__clkbuf_2
X_1463_ _0777_ po_0.regf_0.rf\[15\]\[2\] _0207_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__mux2_1
X_1394_ _0866_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2015_ _2015_/D net62 VGND VGND VPWR VPWR uc_0.bc_0._14_\[2\] sky130_fd_sc_hd__dlxtn_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0963_ _0503_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__buf_2
XFILLER_32_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0894_ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1515_ po_0.regf_0.rf\[12\]\[1\] _0843_ _0237_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__mux2_1
X_1377_ po_0.regf_0.rf\[6\]\[7\] _0841_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__nor2_1
X_1446_ po_0.regf_0.rf\[1\]\[3\] _0847_ _0196_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux2_1
XFILLER_23_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout92 net95 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
Xfanout81 net109 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
Xfanout70 net109 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1231_ _0726_ _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__and2b_1
X_1300_ _0706_ _0707_ _0709_ _0710_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__nand4_1
X_1162_ _0680_ VGND VGND VPWR VPWR _1997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1093_ _0619_ _0621_ _0624_ _0626_ VGND VGND VPWR VPWR po_0.regf_0._3_\[3\] sky130_fd_sc_hd__o22a_1
X_0946_ _0487_ _0493_ VGND VGND VPWR VPWR uc_0.bc_0._85_\[0\] sky130_fd_sc_hd__nor2_1
X_1995_ _1995_/D net61 VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[0\] sky130_fd_sc_hd__dlxtn_1
X_1429_ po_0.regf_0.rf\[9\]\[4\] _0849_ _0184_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__mux2_1
XFILLER_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1780_ _0487_ _0493_ _0666_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__or3_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1145_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__buf_2
X_1214_ po_0._1_\[2\] _0480_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__and2b_1
XFILLER_60_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1076_ po_0.regf_0.rf\[8\]\[2\] po_0.regf_0.rf\[9\]\[2\] po_0.regf_0.rf\[10\]\[2\]
+ po_0.regf_0.rf\[11\]\[2\] _0589_ _0590_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__mux4_1
X_1978_ net66 _0144_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0929_ net20 VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__clkbuf_2
XFILLER_43_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1901_ net89 _0079_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1832_ po_0.regf_0._5_\[6\] net54 VGND VGND VPWR VPWR po_0._1_\[6\] sky130_fd_sc_hd__dlxtp_1
X_1694_ _0380_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1763_ po_0.muxf_0.rf_w_data\[0\] net27 _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
X_1059_ po_0.regf_0.rf\[0\]\[0\] po_0.regf_0.rf\[1\]\[0\] po_0.regf_0.rf\[2\]\[0\]
+ po_0.regf_0.rf\[3\]\[0\] _0594_ _0595_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__mux4_1
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1128_ _0486_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput36 net36 VGND VGND VPWR VPWR D_wr sky130_fd_sc_hd__buf_2
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput25 net25 VGND VGND VPWR VPWR D_W_data[6] sky130_fd_sc_hd__clkbuf_4
Xoutput47 net47 VGND VGND VPWR VPWR leds[1] sky130_fd_sc_hd__buf_2
XFILLER_56_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2031_ net78 _0177_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1815_ uc_0.bc_0._14_\[3\] po_0.muxf_0.rf_w_data\[3\] _0658_ VGND VGND VPWR VPWR
+ _0445_ sky130_fd_sc_hd__mux2_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1746_ _0751_ po_0.regf_0.rf\[11\]\[0\] _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__mux2_1
X_1677_ po_0.regf_0.rf\[3\]\[6\] _0823_ _0363_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__mux2_1
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1462_ _0209_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
X_1600_ _0279_ _0293_ _0310_ _0269_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__nand4_1
X_1531_ _0246_ _0247_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__nor2_2
X_1393_ _0813_ po_0.regf_0.rf\[7\]\[5\] _0859_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__mux2_1
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2014_ _2014_/D net61 VGND VGND VPWR VPWR uc_0.bc_0._14_\[1\] sky130_fd_sc_hd__dlxtn_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1729_ _0813_ po_0.regf_0.rf\[0\]\[5\] _0393_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux2_1
XFILLER_58_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0962_ _0501_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0893_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1514_ _0238_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
X_1445_ _0199_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1376_ _0834_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__clkbuf_2
XFILLER_23_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout93 net95 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout82 net84 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
Xfanout71 net73 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout60 net18 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlymetal6s2s_1
X_1092_ _0623_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__and2b_1
X_1230_ _0719_ _0725_ _0722_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__nand3_1
X_1161_ po_0.muxf_0.rf_w_data\[2\] _0679_ _0676_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__mux2_1
X_1994_ net84 _0156_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_0945_ _0492_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__clkbuf_2
X_1428_ _0189_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1359_ po_0.regf_0.rf\[6\]\[1\] _0843_ _0841_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__mux2_1
XFILLER_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1213_ _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1075_ _0609_ _0585_ _0003_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__a21bo_1
X_1144_ _0487_ _0493_ _0666_ _0667_ _0668_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__o32ai_4
X_1977_ net75 _0143_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_0928_ net24 net50 net26 net25 VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__nor4_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1900_ net102 _0078_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1831_ po_0.regf_0._5_\[5\] net54 VGND VGND VPWR VPWR po_0._1_\[5\] sky130_fd_sc_hd__dlxtp_1
X_1693_ po_0.regf_0.rf\[10\]\[5\] _0812_ _0373_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__mux2_1
X_1762_ _0666_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__clkbuf_4
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1127_ _0650_ _0652_ _0654_ _0656_ VGND VGND VPWR VPWR po_0.regf_0._3_\[7\] sky130_fd_sc_hd__o22a_1
X_1058_ _0581_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__buf_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput37 net37 VGND VGND VPWR VPWR I_addr[0] sky130_fd_sc_hd__clkbuf_4
Xoutput48 net48 VGND VGND VPWR VPWR leds[2] sky130_fd_sc_hd__buf_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput26 net26 VGND VGND VPWR VPWR D_W_data[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_56_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ net79 _0176_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1745_ _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__buf_2
X_1814_ _0444_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1676_ _0370_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1461_ _0768_ po_0.regf_0.rf\[15\]\[1\] _0207_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__mux2_1
X_1392_ _0865_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
X_1530_ uc_0._02_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__clkbuf_2
X_2013_ _2013_/D net62 VGND VGND VPWR VPWR uc_0.bc_0._14_\[0\] sky130_fd_sc_hd__dlxtn_1
XFILLER_50_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1728_ _0399_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1659_ _0834_ _0352_ _0360_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0961_ _0500_ _0505_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__and2b_1
XFILLER_32_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0892_ po_0.alu_0.s1 VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__clkbuf_2
X_1513_ po_0.regf_0.rf\[12\]\[0\] _0837_ _0237_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux2_1
X_1375_ _0854_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
X_1444_ po_0.regf_0.rf\[1\]\[2\] _0845_ _0196_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__mux2_1
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout94 net95 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
Xfanout83 net84 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
Xfanout50 net23 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout72 net81 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
Xfanout61 net62 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1091_ po_0.regf_0.rf\[8\]\[3\] po_0.regf_0.rf\[9\]\[3\] po_0.regf_0.rf\[10\]\[3\]
+ po_0.regf_0.rf\[11\]\[3\] _0580_ _0582_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__mux4_1
X_1160_ uc_0._21_\[2\] VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__clkbuf_2
X_1993_ net98 _0155_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_0944_ _0475_ _0482_ _0489_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__a31oi_2
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1427_ po_0.regf_0.rf\[9\]\[3\] _0847_ _0185_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux2_1
X_1358_ _0767_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__clkbuf_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1289_ _0779_ _0712_ _0745_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1212_ _0709_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__and2_1
X_1074_ po_0.regf_0.rf\[12\]\[2\] po_0.regf_0.rf\[13\]\[2\] po_0.regf_0.rf\[14\]\[2\]
+ po_0.regf_0.rf\[15\]\[2\] _0580_ _0582_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__mux4_1
X_1143_ net60 _0496_ _0486_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__or3b_1
XFILLER_18_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1976_ net76 _0142_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_0927_ uc_0.bc_0._12_\[2\] uc_0.bc_0._12_\[3\] uc_0.bc_0._12_\[1\] uc_0.bc_0._12_\[0\]
+ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__and4b_1
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1761_ _0409_ _0835_ _0417_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__o21ai_1
X_1830_ po_0.regf_0._5_\[4\] net54 VGND VGND VPWR VPWR po_0._1_\[4\] sky130_fd_sc_hd__dlxtp_1
X_1692_ _0379_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
X_1126_ _0655_ _0623_ _0586_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__a21o_1
X_1057_ _0579_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__clkbuf_4
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1959_ net99 _0125_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xoutput38 net38 VGND VGND VPWR VPWR I_addr[1] sky130_fd_sc_hd__clkbuf_4
Xoutput49 net49 VGND VGND VPWR VPWR leds[3] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR D_addr[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1744_ _0857_ _0858_ _0754_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__or3b_4
X_1813_ _0858_ _0443_ _0430_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__mux2_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1675_ po_0.regf_0.rf\[3\]\[5\] _0812_ _0363_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__mux2_1
XFILLER_53_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1109_ _0635_ _0637_ _0593_ _0640_ VGND VGND VPWR VPWR po_0.regf_0._3_\[5\] sky130_fd_sc_hd__o22a_1
XFILLER_26_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1460_ _0208_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
X_1391_ _0802_ po_0.regf_0.rf\[7\]\[4\] _0859_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__mux2_1
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2012_ net79 _0166_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_1
X_1658_ po_0.regf_0.rf\[4\]\[7\] _0352_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__nor2_1
X_1727_ _0802_ po_0.regf_0.rf\[0\]\[4\] _0393_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__mux2_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1589_ _0275_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__nor2_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0960_ po_0.regf_0.rf\[8\]\[0\] po_0.regf_0.rf\[9\]\[0\] po_0.regf_0.rf\[10\]\[0\]
+ po_0.regf_0.rf\[11\]\[0\] _0502_ _0504_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__mux4_1
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1512_ _0236_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__buf_2
X_0891_ _0448_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1374_ po_0.regf_0.rf\[6\]\[6\] _0853_ _0840_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__mux2_1
X_1443_ _0198_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout62 net18 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
Xfanout73 net81 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
Xfanout51 net22 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout95 net96 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout84 net87 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1090_ _0622_ _0623_ _0586_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__a21bo_1
X_1992_ net98 _0154_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_0943_ _0463_ _0490_ _0488_ _0471_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__a211o_1
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1357_ _0842_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
X_1426_ _0188_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
X_1288_ _0708_ _0772_ _0706_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__o21ai_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1142_ net60 _0665_ _0492_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__nor3_2
X_1211_ net51 po_0._1_\[3\] VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__or2_1
XFILLER_60_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1073_ _0603_ _0605_ _0593_ _0608_ VGND VGND VPWR VPWR po_0.regf_0._3_\[1\] sky130_fd_sc_hd__o22a_1
XFILLER_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1975_ net78 _0141_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_0926_ uc_0.bc_0._12_\[1\] uc_0.bc_0._12_\[3\] uc_0.bc_0._12_\[2\] uc_0.bc_0._12_\[0\]
+ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__or4bb_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1409_ po_0.regf_0.rf\[8\]\[3\] _0847_ _0872_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__mux2_1
XFILLER_45_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1760_ _0409_ po_0.regf_0.rf\[11\]\[7\] VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__nand2_1
X_1691_ po_0.regf_0.rf\[10\]\[4\] _0801_ _0373_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__mux2_1
XFILLER_30_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1125_ po_0.regf_0.rf\[4\]\[7\] po_0.regf_0.rf\[5\]\[7\] po_0.regf_0.rf\[6\]\[7\]
+ po_0.regf_0.rf\[7\]\[7\] _0616_ _0617_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux4_1
X_1056_ _0003_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__buf_2
XFILLER_21_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput28 net28 VGND VGND VPWR VPWR D_addr[1] sky130_fd_sc_hd__buf_2
X_1889_ net90 _0067_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1958_ net82 _0124_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xoutput39 net57 VGND VGND VPWR VPWR I_addr[2] sky130_fd_sc_hd__clkbuf_4
X_0909_ _0460_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1674_ _0369_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
X_1812_ uc_0.bc_0._14_\[2\] po_0.muxf_0.rf_w_data\[2\] _0658_ VGND VGND VPWR VPWR
+ _0443_ sky130_fd_sc_hd__mux2_1
X_1743_ _0489_ _0267_ _0487_ _0688_ _0676_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__a2111oi_1
XFILLER_53_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1039_ po_0.regf_0.rf\[4\]\[7\] po_0.regf_0.rf\[5\]\[7\] po_0.regf_0.rf\[6\]\[7\]
+ po_0.regf_0.rf\[7\]\[7\] _0501_ _0503_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__mux4_1
X_1108_ _0638_ _0639_ _0584_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__mux2_1
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1390_ _0864_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2011_ net80 _0165_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfxtp_1
X_1657_ _0359_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
X_1726_ _0398_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
X_1588_ _0679_ net39 _0259_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__o21ai_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0890_ _0447_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1511_ _0869_ po_0.regf_0.w_addr\[1\] _0839_ _0205_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__and4bb_2
X_1442_ po_0.regf_0.rf\[1\]\[1\] _0843_ _0196_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__mux2_1
X_1373_ _0823_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__clkbuf_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1709_ po_0.regf_0.rf\[2\]\[4\] _0801_ _0383_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__mux2_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout96 net108 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout85 net86 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout52 po_0.regf_0.rp_rd VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
Xfanout63 net64 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xfanout74 net77 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1991_ net100 _0153_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_0942_ _0464_ uc_0.bc_0._14_\[6\] uc_0.bc_0._14_\[7\] uc_0.bc_0._14_\[4\] VGND VGND
+ VPWR VPWR _0490_ sky130_fd_sc_hd__a211o_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1425_ po_0.regf_0.rf\[9\]\[2\] _0845_ _0185_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux2_1
X_1287_ _0778_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
X_1356_ po_0.regf_0.rf\[6\]\[0\] _0837_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__mux2_1
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1072_ _0606_ _0607_ _0600_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__mux2_1
X_1141_ uc_0.bc_0._85_\[2\] _0496_ _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__nand3_4
X_1210_ net51 po_0._1_\[3\] VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__nand2_1
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1974_ net65 _0140_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_0925_ uc_0.bc_0._14_\[5\] uc_0.bc_0._14_\[7\] VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__or2_1
X_1408_ _0875_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1339_ _0736_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__inv_2
XFILLER_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1690_ _0378_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1055_ _0588_ _0591_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__and2b_1
X_1124_ _0588_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__and2b_1
X_1957_ net86 _0123_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput29 net29 VGND VGND VPWR VPWR D_addr[2] sky130_fd_sc_hd__buf_2
X_1888_ net93 _0066_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0908_ _0448_ _0452_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__or2b_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1811_ _0442_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1673_ po_0.regf_0.rf\[3\]\[4\] _0801_ _0363_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux2_1
XFILLER_7_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1742_ _0362_ uc_0._01_ _0407_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__a21bo_1
X_1107_ po_0.regf_0.rf\[4\]\[5\] po_0.regf_0.rf\[5\]\[5\] po_0.regf_0.rf\[6\]\[5\]
+ po_0.regf_0.rf\[7\]\[5\] _0579_ _0581_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__mux4_1
X_1038_ po_0.regf_0.rf\[0\]\[7\] po_0.regf_0.rf\[1\]\[7\] po_0.regf_0.rf\[2\]\[7\]
+ po_0.regf_0.rf\[3\]\[7\] _0529_ _0530_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__mux4_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2010_ net63 _0164_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfxtp_1
XFILLER_43_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1725_ _0787_ po_0.regf_0.rf\[0\]\[3\] _0394_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__mux2_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1656_ po_0.regf_0.rf\[4\]\[6\] _0823_ _0351_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux2_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1587_ _0297_ _0298_ _0285_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__o21ai_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1510_ _0227_ _0835_ _0235_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__o21ai_1
X_1441_ _0197_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1372_ _0852_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
X_1708_ _0388_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1639_ _0292_ _0310_ _0324_ _0281_ net44 VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__a41o_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout86 net87 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
Xfanout97 net101 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
Xfanout75 net77 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout64 net70 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
Xfanout53 po_0.regf_0.rp_rd VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1990_ net83 _0152_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_0941_ _0469_ _0467_ _0483_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__a211oi_2
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1355_ _0840_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__buf_2
X_1424_ _0187_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1286_ po_0.regf_0.rf\[5\]\[2\] _0777_ _0758_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__mux2_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1071_ po_0.regf_0.rf\[4\]\[1\] po_0.regf_0.rf\[5\]\[1\] po_0.regf_0.rf\[6\]\[1\]
+ po_0.regf_0.rf\[7\]\[1\] _0597_ _0598_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__mux4_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1140_ _0463_ _0465_ _0467_ _0469_ _0472_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__a221o_2
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1973_ net69 _0139_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_0924_ net58 _0473_ VGND VGND VPWR VPWR uc_0.bc_0._85_\[1\] sky130_fd_sc_hd__nor2_1
X_1338_ _0825_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
X_1407_ po_0.regf_0.rf\[8\]\[2\] _0845_ _0872_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__mux2_1
XFILLER_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1269_ po_0.alu_0.s1 _0447_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__and2b_1
XFILLER_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1054_ po_0.regf_0.rf\[8\]\[0\] po_0.regf_0.rf\[9\]\[0\] po_0.regf_0.rf\[10\]\[0\]
+ po_0.regf_0.rf\[11\]\[0\] _0589_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__mux4_1
X_1123_ po_0.regf_0.rf\[0\]\[7\] po_0.regf_0.rf\[1\]\[7\] po_0.regf_0.rf\[2\]\[7\]
+ po_0.regf_0.rf\[3\]\[7\] _0589_ _0590_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__mux4_1
X_1887_ net90 _0065_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1956_ net82 _0122_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_0907_ _0459_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput19 net19 VGND VGND VPWR VPWR D_W_data[0] sky130_fd_sc_hd__buf_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1810_ _0838_ _0441_ _0430_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__mux2_1
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1741_ _0487_ _0657_ _0496_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__or3_1
XFILLER_15_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1672_ _0368_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1106_ po_0.regf_0.rf\[0\]\[5\] po_0.regf_0.rf\[1\]\[5\] po_0.regf_0.rf\[2\]\[5\]
+ po_0.regf_0.rf\[3\]\[5\] _0597_ _0598_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__mux4_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1037_ _0500_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__and2b_1
X_1939_ net64 net14 VGND VGND VPWR VPWR uc_0._21_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1724_ _0397_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1655_ _0358_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1586_ _0285_ _0297_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__or3_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1371_ po_0.regf_0.rf\[6\]\[5\] _0851_ _0840_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__mux2_1
X_1440_ po_0.regf_0.rf\[1\]\[0\] _0837_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1707_ po_0.regf_0.rf\[2\]\[3\] _0786_ _0384_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__mux2_1
X_1638_ _0335_ _0326_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__or2_1
XFILLER_58_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ uc_0._21_\[3\] net40 VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__and2_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout98 net101 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
Xfanout87 net96 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
Xfanout65 net67 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_2
Xfanout76 net77 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
Xfanout54 po_0.regf_0.rq_rd VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0940_ _0484_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__clkbuf_2
XFILLER_9_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1354_ _0756_ _0838_ _0839_ _0755_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__and4b_2
X_1285_ _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__clkbuf_2
X_1423_ po_0.regf_0.rf\[9\]\[1\] _0843_ _0185_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux2_1
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1070_ po_0.regf_0.rf\[0\]\[1\] po_0.regf_0.rf\[1\]\[1\] po_0.regf_0.rf\[2\]\[1\]
+ po_0.regf_0.rf\[3\]\[1\] _0594_ _0595_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__mux4_1
XFILLER_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1972_ net66 _0138_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_0923_ _0463_ _0465_ _0467_ _0469_ _0472_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__a221oi_1
X_1337_ po_0.regf_0.rf\[5\]\[6\] _0824_ _0757_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__mux2_1
X_1406_ _0874_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1268_ _0479_ po_0._1_\[0\] _0760_ _0704_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__a211o_1
XFILLER_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1199_ _0479_ po_0._1_\[0\] VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__and2b_1
XFILLER_15_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1122_ _0651_ _0623_ _0586_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__a21bo_1
XFILLER_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1053_ _0581_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__buf_2
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1886_ net93 _0064_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1955_ net86 _0121_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_0906_ _0449_ _0453_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__or2b_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1671_ po_0.regf_0.rf\[3\]\[3\] _0786_ _0364_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__mux2_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1740_ po_0.muxf_0.s0 _0405_ _0406_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__o21ba_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1105_ _0600_ _0636_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__and2b_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1036_ po_0.regf_0.rf\[8\]\[7\] po_0.regf_0.rf\[9\]\[7\] po_0.regf_0.rf\[10\]\[7\]
+ po_0.regf_0.rf\[11\]\[7\] _0502_ _0504_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__mux4_1
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1869_ net75 _0011_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__dfxtp_2
X_1938_ net64 net13 VGND VGND VPWR VPWR uc_0._21_\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1654_ po_0.regf_0.rf\[4\]\[5\] _0812_ _0351_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__mux2_1
X_1723_ _0777_ po_0.regf_0.rf\[0\]\[2\] _0394_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__mux2_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1585_ uc_0._21_\[4\] _0292_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__and2b_1
X_1019_ po_0.regf_0.rf\[8\]\[5\] po_0.regf_0.rf\[9\]\[5\] po_0.regf_0.rf\[10\]\[5\]
+ po_0.regf_0.rf\[11\]\[5\] _0502_ _0504_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__mux4_1
XFILLER_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1370_ _0812_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__clkbuf_2
X_1706_ _0387_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
X_1637_ _0343_ _0248_ _0346_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__nand3_1
X_1499_ _0777_ po_0.regf_0.rf\[13\]\[2\] _0227_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__mux2_1
XFILLER_58_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ _0249_ _0675_ _0258_ _0259_ _0273_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__o221ai_2
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout55 po_0.regf_0.rq_rd VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout88 net91 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout99 net101 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
Xfanout77 net81 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout66 net67 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1422_ _0186_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1353_ po_0.regf_0.w_wr VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1284_ net3 _0741_ _0743_ po_0.muxf_0.rf_w_data\[2\] _0775_ VGND VGND VPWR VPWR _0776_
+ sky130_fd_sc_hd__a221o_2
XFILLER_63_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0999_ _0535_ _0537_ _0539_ _0541_ VGND VGND VPWR VPWR po_0.regf_0._5_\[2\] sky130_fd_sc_hd__o22a_1
XFILLER_46_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1971_ net68 _0137_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_0922_ _0471_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__clkbuf_2
X_1405_ po_0.regf_0.rf\[8\]\[1\] _0843_ _0872_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__mux2_1
X_1336_ _0823_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__clkbuf_2
XFILLER_36_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1198_ _0470_ _0468_ _0466_ _0462_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__a31o_2
Xinput1 D_R_data[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_1267_ po_0._1_\[1\] _0478_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__and2b_1
XFILLER_3_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1121_ po_0.regf_0.rf\[12\]\[7\] po_0.regf_0.rf\[13\]\[7\] po_0.regf_0.rf\[14\]\[7\]
+ po_0.regf_0.rf\[15\]\[7\] _0616_ _0617_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__mux4_1
X_1052_ _0579_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__clkbuf_4
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1954_ net66 _0120_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1885_ net65 _0063_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_0905_ _0458_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1319_ po_0.alu_0._11_\[5\] _0450_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__or2b_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1670_ _0367_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1035_ _0572_ _0525_ _0007_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__a21bo_1
X_1104_ po_0.regf_0.rf\[8\]\[5\] po_0.regf_0.rf\[9\]\[5\] po_0.regf_0.rf\[10\]\[5\]
+ po_0.regf_0.rf\[11\]\[5\] _0594_ _0595_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__mux4_1
XFILLER_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1937_ net64 net12 VGND VGND VPWR VPWR uc_0._21_\[3\] sky130_fd_sc_hd__dfxtp_2
X_1868_ net78 _0010_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__dfxtp_1
X_1799_ _0435_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1653_ _0357_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _0396_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
X_1584_ net41 uc_0._21_\[4\] VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__and2b_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1018_ _0557_ _0525_ _0007_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__a21bo_1
XFILLER_1_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1705_ po_0.regf_0.rf\[2\]\[2\] _0776_ _0384_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__mux2_1
X_1636_ _0344_ _0345_ _0339_ _0340_ _0330_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__o221ai_1
X_1567_ _0249_ net38 _0266_ _0279_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__and4_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1498_ _0229_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout89 net91 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout78 net80 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
Xfanout67 net70 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout56 net42 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1421_ po_0.regf_0.rf\[9\]\[0\] _0837_ _0185_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux2_1
XFILLER_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1352_ po_0.regf_0.w_addr\[1\] VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__clkbuf_2
X_1283_ _0770_ _0774_ _0748_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__o21a_1
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0998_ _0540_ _0511_ _0520_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__a21o_1
X_1619_ net56 _0683_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__o21ai_2
XFILLER_27_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1970_ net66 _0136_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_0921_ _0470_ _0462_ _0466_ _0468_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__nor4b_1
XFILLER_18_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1404_ _0873_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1335_ _0799_ _0821_ _0822_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__o21ai_4
Xinput2 D_R_data[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
X_1266_ _0759_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1197_ _0698_ _0699_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__nor2_1
XFILLER_51_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1051_ _0584_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__clkbuf_2
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1120_ _0600_ _0649_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__and2b_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1884_ net97 _0062_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1953_ net75 _0119_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_0904_ _0449_ _0453_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__or2b_1
X_1318_ _0805_ _0806_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__nand2_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1249_ _0742_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__clkbuf_2
XFILLER_62_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1034_ po_0.regf_0.rf\[12\]\[7\] po_0.regf_0.rf\[13\]\[7\] po_0.regf_0.rf\[14\]\[7\]
+ po_0.regf_0.rf\[15\]\[7\] _0522_ _0523_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__mux4_1
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1103_ _0634_ _0585_ _0003_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__a21bo_1
X_1867_ net78 _0009_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__dfxtp_1
X_1936_ net80 net11 VGND VGND VPWR VPWR uc_0._21_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1798_ po_0.regf_0.rp_addr\[0\] uc_0.bc_0._14_\[0\] _0670_ VGND VGND VPWR VPWR _0435_
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1721_ _0768_ po_0.regf_0.rf\[0\]\[1\] _0394_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux2_1
X_1652_ po_0.regf_0.rf\[4\]\[4\] _0801_ _0351_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__mux2_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1583_ _0294_ _0252_ _0295_ _0264_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__a31o_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ po_0.regf_0.rf\[12\]\[5\] po_0.regf_0.rf\[13\]\[5\] po_0.regf_0.rf\[14\]\[5\]
+ po_0.regf_0.rf\[15\]\[5\] _0522_ _0523_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__mux4_1
X_1919_ net73 _0097_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_2
XFILLER_1_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1704_ _0386_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1497_ _0768_ po_0.regf_0.rf\[13\]\[1\] _0227_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__mux2_1
X_1635_ _0685_ _0324_ _0336_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__nor3_1
X_1566_ _0279_ _0269_ _0247_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__o21ai_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout68 net69 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout79 net80 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout57 net39 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_2
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1351_ _0750_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__clkbuf_2
X_1420_ _0184_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__buf_2
X_1282_ _0708_ _0772_ _0773_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0997_ po_0.regf_0.rf\[4\]\[2\] po_0.regf_0.rf\[5\]\[2\] po_0.regf_0.rf\[6\]\[2\]
+ po_0.regf_0.rf\[7\]\[2\] _0507_ _0508_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__mux4_1
X_1618_ uc_0._21_\[6\] net43 VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1549_ _0260_ _0248_ _0261_ _0263_ _0264_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__a311o_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0920_ uc_0.bc_0._12_\[0\] VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__clkbuf_2
X_1265_ po_0.regf_0.rf\[5\]\[0\] _0751_ _0758_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__mux2_1
X_1403_ po_0.regf_0.rf\[8\]\[0\] _0837_ _0872_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__mux2_1
XFILLER_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1334_ net7 _0741_ _0743_ po_0.muxf_0.rf_w_data\[6\] VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__a22oi_2
XFILLER_51_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput3 D_R_data[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_1196_ _0470_ _0468_ _0466_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1050_ _0583_ _0585_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__a21bo_1
XFILLER_33_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1883_ net97 _0061_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1952_ net76 _0118_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_0903_ _0457_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1317_ _0804_ _0796_ _0725_ _0745_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__a31oi_1
X_1248_ po_0.muxf_0.s0 po_0.muxf_0.s1 VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__and2b_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1179_ _0690_ VGND VGND VPWR VPWR _2014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1102_ po_0.regf_0.rf\[12\]\[5\] po_0.regf_0.rf\[13\]\[5\] po_0.regf_0.rf\[14\]\[5\]
+ po_0.regf_0.rf\[15\]\[5\] _0580_ _0582_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__mux4_1
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1033_ _0565_ _0567_ _0569_ _0571_ VGND VGND VPWR VPWR po_0.regf_0._5_\[6\] sky130_fd_sc_hd__o22a_1
X_1935_ net103 net10 VGND VGND VPWR VPWR uc_0._21_\[1\] sky130_fd_sc_hd__dfxtp_2
X_1866_ net78 _0008_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__dfxtp_1
X_1797_ _0434_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1651_ _0356_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
X_1720_ _0395_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ _0250_ _0255_ _0266_ _0279_ _0293_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a41o_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1016_ _0550_ _0552_ _0554_ _0556_ VGND VGND VPWR VPWR po_0.regf_0._5_\[4\] sky130_fd_sc_hd__o22a_1
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1849_ net89 _0031_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1918_ net73 _0096_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfxtp_1
XFILLER_57_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1703_ po_0.regf_0.rf\[2\]\[1\] _0767_ _0384_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__mux2_1
X_1634_ _0685_ net43 _0336_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__o21a_1
X_1496_ _0228_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ net40 VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_2
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout69 net70 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout58 net60 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1350_ _0758_ _0835_ _0836_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__a21oi_1
X_1281_ _0708_ _0772_ _0762_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__o21ai_1
XFILLER_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0996_ _0514_ _0538_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__and2b_1
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1617_ _0299_ _0308_ _0318_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__a21oi_1
X_1479_ po_0.regf_0.rf\[14\]\[1\] _0843_ _0217_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__mux2_1
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1548_ _0253_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__clkbuf_2
XFILLER_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1402_ _0871_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__buf_2
Xinput4 D_R_data[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dlymetal6s2s_1
X_1264_ _0757_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__clkbuf_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1333_ _0818_ _0819_ _0820_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__a21oi_2
X_1195_ _0462_ _0466_ _0470_ _0468_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__and4b_1
X_0979_ _0503_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__buf_2
XFILLER_59_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1882_ net99 _0060_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1951_ net78 _0117_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_0902_ _0449_ _0453_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__or2b_1
X_1316_ _0723_ _0724_ _0796_ _0804_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__a2bb2o_1
X_1247_ _0740_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__clkbuf_2
X_1178_ uc_0.bc_0._14_\[1\] uc_0._21_\[1\] _0688_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__mux2_1
XFILLER_64_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1032_ _0570_ _0511_ _0512_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__a21o_1
XFILLER_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1101_ _0628_ _0630_ _0593_ _0633_ VGND VGND VPWR VPWR po_0.regf_0._3_\[4\] sky130_fd_sc_hd__o22a_1
X_1934_ net71 net9 VGND VGND VPWR VPWR uc_0._21_\[0\] sky130_fd_sc_hd__dfxtp_1
X_1865_ net84 _0047_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1796_ po_0.regf_0.rq_addr\[3\] po_0.muxf_0.rf_w_data\[7\] _0659_ VGND VGND VPWR
+ VPWR _0434_ sky130_fd_sc_hd__mux2_1
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1650_ po_0.regf_0.rf\[4\]\[3\] _0786_ _0352_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux2_1
X_1581_ _0293_ _0281_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__nand2_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1015_ _0555_ _0511_ _0512_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__a21o_1
XFILLER_34_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1917_ net89 _0095_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1848_ net104 _0030_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1779_ _0362_ net35 _0405_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__a21o_1
XFILLER_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1702_ _0385_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
X_1633_ _0337_ _0338_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o21ai_1
X_1564_ _0266_ _0257_ _0270_ _0278_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__o22a_1
X_1495_ _0751_ po_0.regf_0.rf\[13\]\[0\] _0227_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__mux2_1
XFILLER_39_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2047_ po_0.alu_0._10_\[7\] _0888_ VGND VGND VPWR VPWR po_0.alu_0._11_\[7\] sky130_fd_sc_hd__ebufn_1
Xfanout59 net60 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1280_ _0703_ po_0._1_\[0\] _0479_ _0771_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__a31oi_2
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0995_ po_0.regf_0.rf\[0\]\[2\] po_0.regf_0.rf\[1\]\[2\] po_0.regf_0.rf\[2\]\[2\]
+ po_0.regf_0.rf\[3\]\[2\] _0515_ _0516_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__mux4_1
X_1616_ _0325_ _0326_ _0252_ _0264_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__a31oi_1
X_1547_ _0250_ _0255_ _0262_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a21oi_1
X_1478_ _0218_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1401_ _0869_ _0752_ _0839_ _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__and4bb_2
X_1263_ _0752_ _0753_ _0755_ _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__and4b_2
Xinput5 D_R_data[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1194_ net46 _0468_ _0469_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__a21o_1
X_1332_ _0451_ po_0.alu_0._11_\[6\] _0744_ net25 VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__a22o_1
X_0978_ _0501_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1950_ net67 _0116_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1881_ net65 _0059_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_0901_ _0456_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1315_ net50 po_0._1_\[4\] VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__nand2_1
XFILLER_24_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1246_ po_0.muxf_0.s1 po_0.muxf_0.s0 VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__and2b_1
X_1177_ _0689_ VGND VGND VPWR VPWR _2013_/D sky130_fd_sc_hd__clkbuf_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1031_ po_0.regf_0.rf\[4\]\[6\] po_0.regf_0.rf\[5\]\[6\] po_0.regf_0.rf\[6\]\[6\]
+ po_0.regf_0.rf\[7\]\[6\] _0507_ _0508_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__mux4_1
XFILLER_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1100_ _0631_ _0632_ _0584_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__mux2_1
X_1933_ net85 _0111_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1864_ net97 _0046_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1795_ _0433_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__clkbuf_1
X_1229_ _0719_ _0722_ _0725_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1580_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_2
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1014_ po_0.regf_0.rf\[4\]\[4\] po_0.regf_0.rf\[5\]\[4\] po_0.regf_0.rf\[6\]\[4\]
+ po_0.regf_0.rf\[7\]\[4\] _0507_ _0508_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__mux4_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1916_ net102 _0094_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1847_ net104 _0029_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1778_ _0426_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1701_ po_0.regf_0.rf\[2\]\[0\] _0750_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__mux2_1
X_1494_ _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__buf_2
X_1632_ _0339_ _0340_ _0341_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o21bai_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1563_ _0274_ _0276_ _0252_ _0246_ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__a2111oi_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2046_ po_0.alu_0._10_\[6\] _0887_ VGND VGND VPWR VPWR po_0.alu_0._11_\[6\] sky130_fd_sc_hd__ebufn_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0994_ _0536_ _0511_ _0512_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__a21bo_1
X_1477_ po_0.regf_0.rf\[14\]\[0\] _0837_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__mux2_1
X_1615_ _0292_ _0310_ net43 _0281_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__nand4_1
X_1546_ _0249_ _0255_ _0247_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2029_ net64 _0175_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1400_ _0858_ po_0.regf_0.w_addr\[3\] VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__and2b_1
XFILLER_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1331_ _0816_ _0817_ _0732_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__a21o_1
X_1262_ po_0.regf_0.w_addr\[0\] VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1193_ _0697_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xinput6 D_R_data[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_0977_ _0506_ _0513_ _0518_ _0521_ VGND VGND VPWR VPWR po_0.regf_0._5_\[0\] sky130_fd_sc_hd__o22a_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1529_ uc_0._00_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__clkbuf_2
XFILLER_42_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ net68 _0058_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_0900_ _0449_ _0453_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__or2b_1
X_1314_ _0803_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1176_ uc_0.bc_0._14_\[0\] _0675_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__mux2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1245_ _0738_ _0739_ VGND VGND VPWR VPWR po_0.alu_0._10_\[7\] sky130_fd_sc_hd__nand2_1
XFILLER_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1030_ _0514_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__and2b_1
X_1932_ net98 _0110_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1863_ net97 _0045_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1794_ po_0.regf_0.rq_addr\[2\] po_0.muxf_0.rf_w_data\[6\] _0659_ VGND VGND VPWR
+ VPWR _0433_ sky130_fd_sc_hd__mux2_1
X_1228_ _0723_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__nor2_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1159_ _0678_ VGND VGND VPWR VPWR _1996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1013_ _0514_ _0553_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__and2b_1
X_1915_ net103 _0093_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1846_ net105 _0028_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1777_ po_0.muxf_0.rf_w_data\[7\] net34 _0666_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1700_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__buf_2
X_1631_ net56 _0683_ _0329_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__o21a_1
X_1493_ _0838_ _0753_ _0205_ _0869_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__nand4b_4
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1562_ _0276_ _0273_ _0261_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__a21boi_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2045_ po_0.alu_0._10_\[5\] _0886_ VGND VGND VPWR VPWR po_0.alu_0._11_\[5\] sky130_fd_sc_hd__ebufn_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1829_ po_0.regf_0._5_\[3\] net54 VGND VGND VPWR VPWR po_0._1_\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0993_ po_0.regf_0.rf\[12\]\[2\] po_0.regf_0.rf\[13\]\[2\] po_0.regf_0.rf\[14\]\[2\]
+ po_0.regf_0.rf\[15\]\[2\] _0507_ _0508_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__mux4_1
XFILLER_51_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1614_ _0293_ _0310_ _0281_ _0324_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a31o_1
X_1476_ _0216_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__buf_2
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1545_ net37 uc_0._21_\[0\] _0258_ _0259_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__o22ai_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2028_ net74 _0174_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1261_ _0754_ po_0.regf_0.w_addr\[2\] VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__and2b_1
X_1330_ _0732_ _0816_ _0817_ _0745_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__a31oi_1
XFILLER_51_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1192_ _0462_ _0466_ _0470_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__a21bo_1
Xinput7 D_R_data[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
X_0976_ _0519_ _0511_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__a21o_1
XFILLER_32_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1459_ _0751_ po_0.regf_0.rf\[15\]\[0\] _0207_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__mux2_1
X_1528_ _0855_ _0237_ _0245_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__a21oi_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1313_ po_0.regf_0.rf\[5\]\[4\] _0802_ _0757_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__mux2_1
X_1244_ _0735_ _0737_ _0736_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__a21o_1
X_1175_ _0472_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__buf_2
X_0959_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__clkbuf_2
XFILLER_20_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput10 I_data[1] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
X_1931_ net98 _0109_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1862_ net99 _0044_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1793_ _0432_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1227_ net24 po_0._1_\[5\] VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__nor2_1
X_1158_ po_0.muxf_0.rf_w_data\[1\] uc_0._21_\[1\] _0676_ VGND VGND VPWR VPWR _0678_
+ sky130_fd_sc_hd__mux2_1
X_1089_ _0584_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__clkbuf_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1012_ po_0.regf_0.rf\[0\]\[4\] po_0.regf_0.rf\[1\]\[4\] po_0.regf_0.rf\[2\]\[4\]
+ po_0.regf_0.rf\[3\]\[4\] _0515_ _0516_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__mux4_1
X_1914_ net105 _0092_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1845_ net88 _0027_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1776_ _0425_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1630_ _0321_ _0319_ _0317_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__a21oi_1
X_1492_ _0855_ _0217_ _0225_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1561_ net38 uc_0._21_\[1\] _0271_ _0275_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__o22ai_4
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2044_ po_0.alu_0._10_\[4\] _0885_ VGND VGND VPWR VPWR po_0.alu_0._11_\[4\] sky130_fd_sc_hd__ebufn_1
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1759_ _0416_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
X_1828_ po_0.regf_0._5_\[2\] net55 VGND VGND VPWR VPWR po_0._1_\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0992_ _0500_ _0534_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__and2b_1
XFILLER_5_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1613_ net43 VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__clkbuf_2
XFILLER_8_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1544_ _0249_ _0675_ _0258_ _0259_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__or4_1
X_1475_ _0756_ _0838_ _0839_ _0205_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__and4b_2
XFILLER_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2027_ net69 _0173_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput8 D_R_data[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
X_1260_ po_0.regf_0.w_addr\[3\] VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1191_ _0696_ VGND VGND VPWR VPWR _2020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0975_ _0007_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__clkbuf_2
XFILLER_32_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1527_ po_0.regf_0.rf\[12\]\[7\] _0237_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__nor2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1458_ _0206_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__buf_2
X_1389_ _0787_ po_0.regf_0.rf\[7\]\[3\] _0860_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__mux2_1
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1312_ _0801_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__clkbuf_2
X_1174_ _0687_ VGND VGND VPWR VPWR _2002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1243_ _0735_ _0736_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__nand3_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xvahid6i_110 VGND VGND VPWR VPWR I_rd vahid6i_110/LO sky130_fd_sc_hd__conb_1
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0958_ _0005_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__buf_2
X_0889_ po_0.alu_0.s0 VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1930_ net100 _0108_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1861_ net82 _0043_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xinput11 I_data[2] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_1792_ po_0.regf_0.rq_addr\[1\] po_0.muxf_0.rf_w_data\[5\] _0659_ VGND VGND VPWR
+ VPWR _0432_ sky130_fd_sc_hd__mux2_1
X_1226_ net24 po_0._1_\[5\] VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__and2_1
X_1157_ _0677_ VGND VGND VPWR VPWR _1995_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1088_ po_0.regf_0.rf\[12\]\[3\] po_0.regf_0.rf\[13\]\[3\] po_0.regf_0.rf\[14\]\[3\]
+ po_0.regf_0.rf\[15\]\[3\] _0616_ _0617_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__mux4_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1011_ _0551_ _0525_ _0512_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__a21bo_1
X_1913_ net88 _0091_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1844_ net85 _0026_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_1775_ po_0.muxf_0.rf_w_data\[6\] net33 _0666_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__mux2_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1209_ _0705_ _0708_ VGND VGND VPWR VPWR po_0.alu_0._10_\[2\] sky130_fd_sc_hd__xor2_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1560_ uc_0._21_\[2\] net57 VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__and2_1
X_1491_ po_0.regf_0.rf\[14\]\[7\] _0217_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__nor2_1
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2043_ po_0.alu_0._10_\[3\] _0884_ VGND VGND VPWR VPWR po_0.alu_0._11_\[3\] sky130_fd_sc_hd__ebufn_1
X_1827_ po_0.regf_0._5_\[1\] net54 VGND VGND VPWR VPWR po_0._1_\[1\] sky130_fd_sc_hd__dlxtp_1
X_1758_ _0824_ po_0.regf_0.rf\[11\]\[6\] _0408_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux2_1
X_1689_ po_0.regf_0.rf\[10\]\[3\] _0786_ _0374_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__mux2_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0991_ po_0.regf_0.rf\[8\]\[2\] po_0.regf_0.rf\[9\]\[2\] po_0.regf_0.rf\[10\]\[2\]
+ po_0.regf_0.rf\[11\]\[2\] _0502_ _0504_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__mux4_1
X_1474_ _0207_ _0835_ _0215_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__o21ai_1
XFILLER_5_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1612_ _0310_ _0257_ _0313_ _0323_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__o22a_1
XFILLER_8_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1543_ net38 uc_0._21_\[1\] VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__nor2_2
XFILLER_27_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2026_ net74 _0172_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1190_ uc_0.bc_0._14_\[7\] uc_0._21_\[7\] _0472_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__mux2_1
Xinput9 I_data[0] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_44_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0974_ po_0.regf_0.rf\[4\]\[0\] po_0.regf_0.rf\[5\]\[0\] po_0.regf_0.rf\[6\]\[0\]
+ po_0.regf_0.rf\[7\]\[0\] _0507_ _0508_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__mux4_1
XFILLER_59_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1526_ _0244_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
X_1457_ _0869_ _0838_ _0753_ _0205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__nand4_4
X_1388_ _0863_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2009_ net74 _0163_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dfxtp_1
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1311_ net5 _0741_ _0743_ po_0.muxf_0.rf_w_data\[4\] _0800_ VGND VGND VPWR VPWR _0801_
+ sky130_fd_sc_hd__a221o_2
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1173_ po_0.muxf_0.rf_w_data\[7\] uc_0._21_\[7\] _0488_ VGND VGND VPWR VPWR _0687_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1242_ po_0._1_\[6\] net25 VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__or2b_1
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0957_ _0501_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__buf_2
XFILLER_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1509_ _0227_ po_0.regf_0.rf\[13\]\[7\] VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__nand2_1
XFILLER_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1860_ net86 _0042_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xinput12 I_data[3] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
X_1791_ _0431_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1087_ _0588_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__and2b_1
X_1225_ po_0._1_\[4\] net50 VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__or2b_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1156_ po_0.muxf_0.rf_w_data\[0\] _0675_ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__mux2_1
X_1989_ net87 _0151_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ po_0.regf_0.rf\[12\]\[4\] po_0.regf_0.rf\[13\]\[4\] po_0.regf_0.rf\[14\]\[4\]
+ po_0.regf_0.rf\[15\]\[4\] _0522_ _0523_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__mux4_1
X_1912_ net94 _0090_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_1843_ net83 _0025_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1774_ _0424_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1208_ _0706_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__nand2_2
X_1139_ _0664_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1490_ _0224_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2042_ po_0.alu_0._10_\[2\] _0883_ VGND VGND VPWR VPWR po_0.alu_0._11_\[2\] sky130_fd_sc_hd__ebufn_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1826_ po_0.regf_0._5_\[0\] net55 VGND VGND VPWR VPWR po_0._1_\[0\] sky130_fd_sc_hd__dlxtp_1
X_1757_ _0415_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
X_1688_ _0377_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0990_ _0526_ _0528_ _0520_ _0533_ VGND VGND VPWR VPWR po_0.regf_0._5_\[1\] sky130_fd_sc_hd__o22a_1
X_1611_ _0319_ _0321_ _0322_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1473_ _0207_ po_0.regf_0.rf\[15\]\[7\] VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__nand2_1
X_1542_ net38 uc_0._21_\[1\] VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__and2_1
XFILLER_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2025_ net99 _0171_ VGND VGND VPWR VPWR po_0.regf_0.w_wr sky130_fd_sc_hd__dfxtp_1
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1809_ uc_0.bc_0._14_\[1\] po_0.muxf_0.rf_w_data\[1\] _0658_ VGND VGND VPWR VPWR
+ _0441_ sky130_fd_sc_hd__mux2_1
XFILLER_60_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0973_ _0514_ _0517_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__and2b_1
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1525_ po_0.regf_0.rf\[12\]\[6\] _0853_ _0236_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__mux2_1
X_1387_ _0777_ po_0.regf_0.rf\[7\]\[2\] _0860_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__mux2_1
X_1456_ _0858_ _0754_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__and2_2
X_2008_ net102 _0162_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfxtp_1
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1310_ _0797_ _0798_ _0799_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__a21oi_1
X_1241_ net26 po_0._1_\[7\] VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__xnor2_2
XFILLER_64_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1172_ _0686_ VGND VGND VPWR VPWR _2001_/D sky130_fd_sc_hd__clkbuf_1
X_0956_ _0004_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__buf_2
XFILLER_32_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1508_ _0234_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
X_1439_ _0195_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__buf_2
XFILLER_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput13 I_data[4] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
X_1790_ po_0.regf_0.rq_addr\[0\] po_0.muxf_0.rf_w_data\[4\] _0659_ VGND VGND VPWR
+ VPWR _0431_ sky130_fd_sc_hd__mux2_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1224_ _0721_ VGND VGND VPWR VPWR po_0.alu_0._10_\[4\] sky130_fd_sc_hd__clkbuf_1
X_1086_ po_0.regf_0.rf\[0\]\[3\] po_0.regf_0.rf\[1\]\[3\] po_0.regf_0.rf\[2\]\[3\]
+ po_0.regf_0.rf\[3\]\[3\] _0589_ _0590_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__mux4_1
X_1155_ _0488_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__buf_2
X_1988_ net82 _0150_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0939_ net59 VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__clkbuf_2
XFILLER_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1773_ po_0.muxf_0.rf_w_data\[5\] net32 _0418_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux2_1
X_1911_ net90 _0089_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1842_ net92 _0024_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1207_ net21 po_0._1_\[2\] VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__or2_1
XFILLER_33_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1069_ _0588_ _0604_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__and2b_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1138_ po_0.regf_0.rq_addr\[3\] po_0.muxf_0.rf_w_data\[7\] _0660_ VGND VGND VPWR
+ VPWR _0664_ sky130_fd_sc_hd__mux2_1
XFILLER_17_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2041_ po_0.alu_0._10_\[1\] _0882_ VGND VGND VPWR VPWR po_0.alu_0._11_\[1\] sky130_fd_sc_hd__ebufn_1
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1825_ net92 _0023_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1756_ _0813_ po_0.regf_0.rf\[11\]\[5\] _0408_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__mux2_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1687_ po_0.regf_0.rf\[10\]\[2\] _0776_ _0374_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__mux2_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1610_ _0299_ _0308_ _0318_ _0247_ _0246_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__a311o_1
XFILLER_8_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1472_ _0214_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
X_1541_ _0256_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__clkbuf_2
X_2024_ net77 _0170_ VGND VGND VPWR VPWR po_0.regf_0.rp_rd sky130_fd_sc_hd__dfxtp_1
XFILLER_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1808_ _0440_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
X_1739_ _0657_ uc_0.bc_0._85_\[3\] _0667_ _0660_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__a31o_1
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0972_ po_0.regf_0.rf\[0\]\[0\] po_0.regf_0.rf\[1\]\[0\] po_0.regf_0.rf\[2\]\[0\]
+ po_0.regf_0.rf\[3\]\[0\] _0515_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__mux4_1
X_1524_ _0243_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
X_1386_ _0862_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
X_1455_ _0855_ _0196_ _0204_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__a21oi_1
X_2007_ net102 _0161_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfxtp_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1171_ po_0.muxf_0.rf_w_data\[6\] _0685_ _0488_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__mux2_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1240_ _0726_ _0733_ _0732_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0955_ _0006_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1507_ _0824_ po_0.regf_0.rf\[13\]\[6\] _0226_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__mux2_1
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1369_ _0850_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
X_1438_ _0752_ _0839_ _0194_ _0756_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__and4b_2
XFILLER_62_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 I_data[5] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1223_ _0719_ _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__and2_1
X_1154_ uc_0._21_\[0\] VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__clkbuf_2
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1085_ _0618_ _0585_ _0586_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__a21o_1
X_1987_ net85 _0149_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_0938_ net58 _0486_ VGND VGND VPWR VPWR uc_0.bc_0._85_\[2\] sky130_fd_sc_hd__nor2_1
XFILLER_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1910_ net93 _0088_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1772_ _0423_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
X_1841_ po_0.regf_0._3_\[7\] net52 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlxtp_1
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1137_ _0663_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
X_1206_ _0480_ po_0._1_\[2\] VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__nand2_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1068_ po_0.regf_0.rf\[8\]\[1\] po_0.regf_0.rf\[9\]\[1\] po_0.regf_0.rf\[10\]\[1\]
+ po_0.regf_0.rf\[11\]\[1\] _0589_ _0590_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__mux4_1
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2040_ po_0.alu_0._10_\[0\] _0881_ VGND VGND VPWR VPWR po_0.alu_0._11_\[0\] sky130_fd_sc_hd__ebufn_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1824_ net104 _0022_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1755_ _0414_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
X_1686_ _0376_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1540_ uc_0._01_ _0246_ uc_0._02_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__or3_1
X_1471_ _0824_ po_0.regf_0.rf\[15\]\[6\] _0206_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__mux2_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2023_ net72 _0169_ VGND VGND VPWR VPWR po_0.regf_0.rq_rd sky130_fd_sc_hd__dfxtp_1
XFILLER_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1807_ _0869_ _0439_ _0430_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__mux2_1
X_1669_ po_0.regf_0.rf\[3\]\[2\] _0776_ _0364_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__mux2_1
X_1738_ _0493_ _0403_ _0404_ _0405_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__a211oi_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0971_ _0503_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__buf_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1523_ po_0.regf_0.rf\[12\]\[5\] _0851_ _0236_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__mux2_1
X_1454_ po_0.regf_0.rf\[1\]\[7\] _0196_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__nor2_1
X_1385_ _0768_ po_0.regf_0.rf\[7\]\[1\] _0860_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__mux2_1
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2006_ net94 _0160_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1170_ uc_0._21_\[6\] VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__clkbuf_2
XFILLER_64_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0954_ _0499_ VGND VGND VPWR VPWR po_0.alu_0._10_\[0\] sky130_fd_sc_hd__clkbuf_1
X_1506_ _0233_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
X_1437_ _0858_ _0754_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__nor2_1
X_1368_ po_0.regf_0.rf\[6\]\[4\] _0849_ _0840_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__mux2_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1299_ _0478_ po_0._1_\[1\] VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__nand2_1
XFILLER_7_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput15 I_data[6] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
X_1084_ po_0.regf_0.rf\[4\]\[3\] po_0.regf_0.rf\[5\]\[3\] po_0.regf_0.rf\[6\]\[3\]
+ po_0.regf_0.rf\[7\]\[3\] _0616_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__mux4_1
X_1153_ _0674_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
X_1222_ _0715_ _0716_ _0718_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__or3_1
X_1986_ net72 _0148_ VGND VGND VPWR VPWR uc_0._02_ sky130_fd_sc_hd__dfxtp_1
X_0937_ _0474_ uc_0.bc_0._14_\[6\] _0475_ _0482_ _0485_ VGND VGND VPWR VPWR _0486_
+ sky130_fd_sc_hd__o311a_1
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1840_ po_0.regf_0._3_\[6\] net53 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlxtp_1
X_1771_ po_0.muxf_0.rf_w_data\[4\] net31 _0418_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux2_1
X_1067_ _0602_ _0585_ _0003_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__a21bo_1
X_1205_ _0700_ _0704_ _0701_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__o21ai_1
X_1136_ po_0.regf_0.rq_addr\[2\] po_0.muxf_0.rf_w_data\[6\] _0660_ VGND VGND VPWR
+ VPWR _0663_ sky130_fd_sc_hd__mux2_1
X_1969_ net75 _0135_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1823_ net104 _0021_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1754_ _0802_ po_0.regf_0.rf\[11\]\[4\] _0408_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux2_1
X_1685_ po_0.regf_0.rf\[10\]\[1\] _0767_ _0374_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__mux2_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1119_ po_0.regf_0.rf\[8\]\[7\] po_0.regf_0.rf\[9\]\[7\] po_0.regf_0.rf\[10\]\[7\]
+ po_0.regf_0.rf\[11\]\[7\] _0594_ _0595_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__mux4_1
XFILLER_44_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1470_ _0213_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2022_ net63 _0168_ VGND VGND VPWR VPWR po_0.alu_0.s0 sky130_fd_sc_hd__dfxtp_1
X_1806_ uc_0.bc_0._14_\[0\] po_0.muxf_0.rf_w_data\[0\] _0658_ VGND VGND VPWR VPWR
+ _0439_ sky130_fd_sc_hd__mux2_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1668_ _0366_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
X_1599_ _0279_ _0293_ _0269_ _0310_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__a31o_1
X_1737_ _0657_ _0493_ _0496_ uc_0.bc_0._85_\[1\] VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__and4b_1
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0970_ _0501_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1522_ _0242_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_1453_ _0203_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2005_ net94 _0159_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfxtp_1
X_1384_ _0861_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0953_ _0497_ _0498_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__and2_1
X_1505_ _0813_ po_0.regf_0.rf\[13\]\[5\] _0226_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__mux2_1
X_1367_ _0801_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__clkbuf_2
X_1436_ _0855_ _0185_ _0193_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__a21oi_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1298_ _0788_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput16 I_data[7] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1221_ _0715_ _0716_ _0718_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__o21ai_1
X_1083_ _0581_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__buf_2
XFILLER_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1152_ po_0.regf_0.rp_addr\[3\] uc_0.bc_0._14_\[3\] _0670_ VGND VGND VPWR VPWR _0674_
+ sky130_fd_sc_hd__mux2_1
X_0936_ _0470_ _0483_ _0484_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a21oi_1
X_1985_ net72 _0147_ VGND VGND VPWR VPWR uc_0._01_ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1419_ _0752_ _0753_ _0870_ _0756_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__and4b_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1770_ _0422_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1204_ _0478_ po_0._1_\[1\] VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__and2b_1
X_1066_ po_0.regf_0.rf\[12\]\[1\] po_0.regf_0.rf\[13\]\[1\] po_0.regf_0.rf\[14\]\[1\]
+ po_0.regf_0.rf\[15\]\[1\] _0580_ _0582_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__mux4_1
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1135_ _0662_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1899_ net103 _0077_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1968_ net76 _0134_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_0919_ _0468_ uc_0.bc_0._12_\[0\] VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1822_ net105 _0020_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1753_ _0413_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
X_1684_ _0375_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
X_1118_ _0642_ _0644_ _0646_ _0648_ VGND VGND VPWR VPWR po_0.regf_0._3_\[6\] sky130_fd_sc_hd__o22a_1
X_1049_ _0003_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2021_ net70 _0167_ VGND VGND VPWR VPWR po_0.alu_0.s1 sky130_fd_sc_hd__dfxtp_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1736_ _0403_ _0667_ po_0.muxf_0.s1 VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__a21oi_1
X_1805_ _0438_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1667_ po_0.regf_0.rf\[3\]\[1\] _0767_ _0364_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__mux2_1
X_1598_ net56 VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__clkbuf_2
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1521_ po_0.regf_0.rf\[12\]\[4\] _0849_ _0236_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__mux2_1
X_1383_ _0751_ po_0.regf_0.rf\[7\]\[0\] _0860_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__mux2_1
X_1452_ po_0.regf_0.rf\[1\]\[6\] _0853_ _0195_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__mux2_1
XFILLER_4_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2004_ net106 _0158_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfxtp_1
XFILLER_35_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1719_ _0751_ po_0.regf_0.rf\[0\]\[0\] _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__mux2_1
XFILLER_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0952_ _0479_ po_0._1_\[0\] VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__nand2_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1504_ _0232_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
X_1366_ _0848_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
X_1435_ po_0.regf_0.rf\[9\]\[7\] _0185_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__nor2_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1297_ po_0.regf_0.rf\[5\]\[3\] _0787_ _0758_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__mux2_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput17 clock VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1151_ _0673_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
X_1220_ _0712_ _0714_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__o21ai_1
X_1082_ _0579_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__clkbuf_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0935_ uc_0.bc_0._12_\[0\] uc_0.bc_0._12_\[1\] uc_0.bc_0._12_\[3\] uc_0.bc_0._12_\[2\]
+ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nor4b_1
X_1984_ net63 uc_0.bc_0._85_\[3\] VGND VGND VPWR VPWR uc_0.bc_0._12_\[3\] sky130_fd_sc_hd__dfxtp_1
X_1349_ po_0.regf_0.rf\[5\]\[7\] _0758_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__nor2_1
X_1418_ _0855_ _0872_ _0880_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__a21oi_1
XFILLER_28_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1203_ _0700_ _0703_ VGND VGND VPWR VPWR po_0.alu_0._10_\[1\] sky130_fd_sc_hd__xor2_1
X_1134_ po_0.regf_0.rq_addr\[1\] po_0.muxf_0.rf_w_data\[5\] _0660_ VGND VGND VPWR
+ VPWR _0662_ sky130_fd_sc_hd__mux2_1
X_1065_ _0587_ _0592_ _0593_ _0601_ VGND VGND VPWR VPWR po_0.regf_0._3_\[0\] sky130_fd_sc_hd__o22a_1
XFILLER_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1898_ net105 _0076_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1967_ net76 _0133_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_0918_ uc_0.bc_0._12_\[1\] VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1821_ net88 _0019_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1752_ _0787_ po_0.regf_0.rf\[11\]\[3\] _0409_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux2_1
X_1683_ po_0.regf_0.rf\[10\]\[0\] _0750_ _0374_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__mux2_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1117_ _0647_ _0623_ _0593_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__a21o_1
X_1048_ _0584_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__clkbuf_2
XFILLER_21_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2020_ _2020_/D net58 VGND VGND VPWR VPWR uc_0.bc_0._14_\[7\] sky130_fd_sc_hd__dlxtn_1
XFILLER_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1666_ _0365_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
X_1804_ po_0.regf_0.rp_addr\[3\] uc_0.bc_0._14_\[3\] _0669_ VGND VGND VPWR VPWR _0438_
+ sky130_fd_sc_hd__mux2_1
X_1735_ _0657_ uc_0.bc_0._85_\[3\] VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__and2_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ _0293_ _0257_ _0296_ _0309_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__o22a_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1520_ _0241_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
X_1382_ _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__buf_2
X_1451_ _0202_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2003_ net80 _0157_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfxtp_1
X_1649_ _0355_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
X_1718_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__buf_2
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0951_ net19 po_0._1_\[0\] VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__or2_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1503_ _0802_ po_0.regf_0.rf\[13\]\[4\] _0226_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__mux2_1
XFILLER_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1365_ po_0.regf_0.rf\[6\]\[3\] _0847_ _0841_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__mux2_1
X_1434_ _0192_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
X_1296_ _0786_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__clkbuf_2
XFILLER_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 reset VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1150_ po_0.regf_0.rp_addr\[2\] uc_0.bc_0._14_\[2\] _0670_ VGND VGND VPWR VPWR _0673_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1081_ _0610_ _0612_ _0593_ _0615_ VGND VGND VPWR VPWR po_0.regf_0._3_\[2\] sky130_fd_sc_hd__o22a_1
X_0934_ uc_0.bc_0._12_\[3\] uc_0.bc_0._12_\[2\] uc_0.bc_0._12_\[1\] VGND VGND VPWR
+ VPWR _0483_ sky130_fd_sc_hd__nor3b_1
X_1983_ net72 uc_0.bc_0._85_\[2\] VGND VGND VPWR VPWR uc_0.bc_0._12_\[2\] sky130_fd_sc_hd__dfxtp_1
X_1417_ po_0.regf_0.rf\[8\]\[7\] _0872_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__nor2_1
X_1348_ _0834_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__clkbuf_2
X_1279_ _0478_ po_0._1_\[1\] VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__and2_1
XFILLER_36_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1064_ _0596_ _0599_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__mux2_1
X_1133_ _0661_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
X_1202_ _0701_ _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__nand2_1
X_1966_ net65 _0132_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1897_ net88 _0075_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_0917_ _0462_ _0466_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__nor2_1
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1820_ net92 _0018_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1751_ _0412_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
X_1682_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__buf_2
X_1116_ po_0.regf_0.rf\[4\]\[6\] po_0.regf_0.rf\[5\]\[6\] po_0.regf_0.rf\[6\]\[6\]
+ po_0.regf_0.rf\[7\]\[6\] _0616_ _0617_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__mux4_1
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1047_ _0002_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1949_ net69 _0115_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1803_ _0437_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
X_1734_ _0394_ _0835_ _0402_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__o21ai_1
X_1665_ po_0.regf_0.rf\[3\]\[0\] _0750_ _0364_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux2_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1596_ _0306_ _0248_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__and3_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ po_0.regf_0.rf\[1\]\[5\] _0851_ _0195_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1381_ _0754_ _0857_ _0858_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__or3b_2
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2002_ _2002_/D net58 VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[7\] sky130_fd_sc_hd__dlxtn_1
XFILLER_16_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1648_ po_0.regf_0.rf\[4\]\[2\] _0776_ _0352_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux2_1
X_1717_ po_0.regf_0.w_addr\[0\] po_0.regf_0.w_addr\[1\] po_0.regf_0.w_wr _0194_ VGND
+ VGND VPWR VPWR _0393_ sky130_fd_sc_hd__or4bb_4
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ net41 VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_2
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0950_ net60 _0496_ VGND VGND VPWR VPWR uc_0.bc_0._85_\[3\] sky130_fd_sc_hd__nor2_2
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1502_ _0231_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
X_1433_ po_0.regf_0.rf\[9\]\[6\] _0853_ _0184_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1364_ _0786_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__clkbuf_2
X_1295_ _0783_ _0784_ _0748_ _0785_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__a31o_2
XFILLER_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1080_ _0613_ _0614_ _0584_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__mux2_1
X_1982_ net63 uc_0.bc_0._85_\[1\] VGND VGND VPWR VPWR uc_0.bc_0._12_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0933_ _0476_ _0477_ _0481_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__nand3_1
X_1416_ _0879_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
X_1347_ _0830_ _0832_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__a21oi_4
XFILLER_36_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1278_ _0450_ po_0.alu_0._11_\[2\] _0744_ _0480_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__a22o_1
XFILLER_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1201_ net20 po_0._1_\[1\] VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__or2b_1
X_1063_ _0002_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__clkbuf_2
X_1132_ po_0.regf_0.rq_addr\[0\] po_0.muxf_0.rf_w_data\[4\] _0660_ VGND VGND VPWR
+ VPWR _0661_ sky130_fd_sc_hd__mux2_1
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1965_ net68 _0131_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_0916_ uc_0.bc_0._12_\[2\] VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__clkbuf_2
X_1896_ net95 _0074_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1750_ _0777_ po_0.regf_0.rf\[11\]\[2\] _0409_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__mux2_1
X_1681_ po_0.regf_0.w_addr\[0\] _0752_ po_0.regf_0.w_wr _0870_ VGND VGND VPWR VPWR
+ _0373_ sky130_fd_sc_hd__and4b_2
X_1046_ po_0.regf_0.rf\[12\]\[0\] po_0.regf_0.rf\[13\]\[0\] po_0.regf_0.rf\[14\]\[0\]
+ po_0.regf_0.rf\[15\]\[0\] _0580_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__mux4_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1115_ _0588_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__and2b_1
X_1879_ net65 _0057_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1948_ net67 _0114_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1733_ _0394_ po_0.regf_0.rf\[0\]\[7\] VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__nand2_1
X_1802_ po_0.regf_0.rp_addr\[2\] uc_0.bc_0._14_\[2\] _0669_ VGND VGND VPWR VPWR _0437_
+ sky130_fd_sc_hd__mux2_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1664_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__buf_2
X_1595_ _0305_ _0288_ _0307_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__o21bai_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1029_ po_0.regf_0.rf\[0\]\[6\] po_0.regf_0.rf\[1\]\[6\] po_0.regf_0.rf\[2\]\[6\]
+ po_0.regf_0.rf\[3\]\[6\] _0515_ _0516_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__mux4_1
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1380_ po_0.regf_0.w_addr\[2\] VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2001_ _2001_/D net59 VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[6\] sky130_fd_sc_hd__dlxtn_1
XFILLER_50_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1716_ _0834_ _0384_ _0392_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__a21oi_1
X_1647_ _0354_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _0291_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1501_ _0787_ po_0.regf_0.rf\[13\]\[3\] _0227_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__mux2_1
X_1363_ _0846_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
X_1432_ _0191_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
X_1294_ net4 _0740_ _0742_ po_0.muxf_0.rf_w_data\[3\] VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__a22o_1
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1981_ net63 uc_0.bc_0._85_\[0\] VGND VGND VPWR VPWR uc_0.bc_0._12_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0932_ _0478_ _0479_ net51 _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__nor4_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1415_ po_0.regf_0.rf\[8\]\[6\] _0853_ _0871_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__mux2_1
XFILLER_28_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1346_ net8 _0741_ _0743_ po_0.muxf_0.rf_w_data\[7\] VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__a22o_1
XFILLER_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1277_ _0769_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1200_ po_0._1_\[1\] net20 VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__or2b_1
X_1062_ po_0.regf_0.rf\[4\]\[0\] po_0.regf_0.rf\[5\]\[0\] po_0.regf_0.rf\[6\]\[0\]
+ po_0.regf_0.rf\[7\]\[0\] _0597_ _0598_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__mux4_1
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1131_ _0659_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__buf_2
X_1895_ net90 _0073_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1964_ net65 _0130_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_0915_ _0464_ uc_0.bc_0._14_\[7\] VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__nor2_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1329_ _0804_ _0724_ _0723_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__o21ba_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1680_ _0834_ _0364_ _0372_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1114_ po_0.regf_0.rf\[0\]\[6\] po_0.regf_0.rf\[1\]\[6\] po_0.regf_0.rf\[2\]\[6\]
+ po_0.regf_0.rf\[3\]\[6\] _0589_ _0590_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__mux4_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1045_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__buf_2
X_1878_ net68 _0056_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1947_ net68 _0113_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1663_ _0869_ _0838_ _0753_ _0194_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__and4_2
X_1732_ _0401_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
X_1801_ _0436_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _0299_ _0300_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__nand2_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1028_ _0566_ _0525_ _0512_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__a21bo_1
XFILLER_39_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2000_ _2000_/D net58 VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[5\] sky130_fd_sc_hd__dlxtn_2
XFILLER_50_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1646_ po_0.regf_0.rf\[4\]\[1\] _0767_ _0352_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux2_1
X_1715_ po_0.regf_0.rf\[2\]\[7\] _0384_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__nor2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1577_ _0290_ _0279_ _0253_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__mux2_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1500_ _0230_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
X_1362_ po_0.regf_0.rf\[6\]\[2\] _0845_ _0841_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__mux2_1
X_1431_ po_0.regf_0.rf\[9\]\[5\] _0851_ _0184_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux2_1
X_1293_ net51 _0451_ _0447_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__or3_1
XFILLER_63_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1629_ _0330_ _0331_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__nand2_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0931_ net21 VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1980_ net74 _0146_ VGND VGND VPWR VPWR po_0.muxf_0.s0 sky130_fd_sc_hd__dfxtp_1
XFILLER_20_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1276_ po_0.regf_0.rf\[5\]\[1\] _0768_ _0758_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__mux2_1
X_1414_ _0878_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
X_1345_ net26 _0452_ _0448_ _0831_ _0748_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__o311a_1
XFILLER_51_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1130_ _0658_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__buf_2
XFILLER_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1061_ _0001_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__buf_2
X_1894_ net92 _0072_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1963_ net68 _0129_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_0914_ uc_0.bc_0._14_\[5\] VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__clkbuf_2
X_1259_ po_0.regf_0.w_wr VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__buf_2
X_1328_ _0795_ _0791_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__o21ai_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1113_ _0643_ _0623_ _0586_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__a21bo_1
X_1044_ _0001_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__clkbuf_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1877_ net83 _0055_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1946_ net69 _0015_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__dfxtp_2
XFILLER_52_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1800_ po_0.regf_0.rp_addr\[1\] uc_0.bc_0._14_\[1\] _0669_ VGND VGND VPWR VPWR _0436_
+ sky130_fd_sc_hd__mux2_1
X_1731_ _0824_ po_0.regf_0.rf\[0\]\[6\] _0393_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__mux2_1
X_1662_ _0487_ _0246_ _0362_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__o21a_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ _0299_ _0300_ _0303_ _0304_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a221o_1
X_1027_ po_0.regf_0.rf\[12\]\[6\] po_0.regf_0.rf\[13\]\[6\] po_0.regf_0.rf\[14\]\[6\]
+ po_0.regf_0.rf\[15\]\[6\] _0522_ _0523_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__mux4_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1929_ net83 _0107_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1645_ _0353_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_1714_ _0391_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1576_ _0280_ _0281_ _0288_ _0289_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__o22ai_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1430_ _0190_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1361_ _0776_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__clkbuf_2
X_1292_ _0452_ _0448_ _0781_ _0782_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__o211ai_1
XFILLER_63_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1628_ _0685_ _0324_ _0336_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__nor3b_1
X_1559_ _0250_ _0675_ _0258_ _0259_ _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__o221a_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0930_ net19 VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__clkbuf_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1413_ po_0.regf_0.rf\[8\]\[5\] _0851_ _0871_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__mux2_1
XFILLER_5_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1275_ _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__clkbuf_2
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1344_ po_0.alu_0._11_\[7\] _0451_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__or2b_1
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout100 net101 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1060_ _0000_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__clkbuf_4
X_1962_ net84 _0128_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1893_ net90 _0071_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_0913_ uc_0.bc_0._12_\[1\] _0462_ uc_0.bc_0._12_\[2\] uc_0.bc_0._12_\[0\] VGND VGND
+ VPWR VPWR _0463_ sky130_fd_sc_hd__and4bb_1
XFILLER_64_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1258_ po_0.regf_0.w_addr\[1\] VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1189_ _0695_ VGND VGND VPWR VPWR _2019_/D sky130_fd_sc_hd__clkbuf_1
X_1327_ _0715_ _0716_ _0723_ _0724_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__nor4_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1112_ po_0.regf_0.rf\[12\]\[6\] po_0.regf_0.rf\[13\]\[6\] po_0.regf_0.rf\[14\]\[6\]
+ po_0.regf_0.rf\[15\]\[6\] _0616_ _0617_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__mux4_1
X_1043_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1945_ net75 _0014_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__dfxtp_1
X_1876_ net98 _0054_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1730_ _0400_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1661_ _0361_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__buf_2
X_1592_ _0679_ _0266_ _0285_ _0283_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__o22a_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1026_ _0500_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__and2b_1
XFILLER_26_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1928_ net85 _0106_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_1859_ net82 _0041_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1713_ po_0.regf_0.rf\[2\]\[6\] _0823_ _0383_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__mux2_1
X_1644_ po_0.regf_0.rf\[4\]\[0\] _0750_ _0352_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__mux2_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1575_ _0276_ _0282_ _0287_ uc_0._02_ _0246_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__a311o_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1009_ _0500_ _0549_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__and2b_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1360_ _0844_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1291_ _0745_ po_0.alu_0._11_\[3\] VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__nand2_1
XFILLER_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1489_ po_0.regf_0.rf\[14\]\[6\] _0853_ _0216_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__mux2_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1627_ _0685_ _0324_ _0336_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__o21ba_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1558_ _0271_ _0272_ _0259_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__nand3b_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1412_ _0877_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1343_ _0827_ _0762_ _0829_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__nand3_1
XFILLER_51_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1274_ _0765_ _0748_ _0766_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__a21o_2
X_0989_ _0531_ _0532_ _0510_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__mux2_1
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout101 net108 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1892_ net102 _0070_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1961_ net97 _0127_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0912_ uc_0.bc_0._12_\[3\] VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1326_ _0814_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
X_1257_ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__clkbuf_2
XFILLER_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1188_ uc_0.bc_0._14_\[6\] _0685_ _0472_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__mux2_1
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1111_ _0600_ _0641_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__and2b_1
X_1042_ _0000_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__buf_2
X_1875_ net98 _0053_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1944_ net75 _0013_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1309_ _0740_ _0742_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__or2_1
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ _0665_ uc_0.bc_0._85_\[2\] uc_0.bc_0._85_\[3\] uc_0.bc_0._85_\[0\] VGND VGND
+ VPWR VPWR _0361_ sky130_fd_sc_hd__or4b_1
X_1591_ _0283_ _0284_ _0286_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__o21a_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1025_ po_0.regf_0.rf\[8\]\[6\] po_0.regf_0.rf\[9\]\[6\] po_0.regf_0.rf\[10\]\[6\]
+ po_0.regf_0.rf\[11\]\[6\] _0502_ _0504_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__mux4_1
XFILLER_34_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1927_ net83 _0105_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1858_ net86 _0040_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1789_ _0362_ _0753_ _0430_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__a21o_1
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1643_ _0351_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__buf_2
X_1712_ _0390_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 po_0.muxf_0.rf_w_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1574_ _0276_ _0282_ _0287_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__a21oi_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1008_ po_0.regf_0.rf\[8\]\[4\] po_0.regf_0.rf\[9\]\[4\] po_0.regf_0.rf\[10\]\[4\]
+ po_0.regf_0.rf\[11\]\[4\] _0502_ _0504_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__mux4_1
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1290_ _0712_ _0779_ _0780_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__o21ai_1
XFILLER_31_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1626_ uc_0._21_\[7\] net44 VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__xnor2_1
X_1488_ _0223_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1557_ _0679_ net57 VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__nand2_1
XFILLER_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1411_ po_0.regf_0.rf\[8\]\[4\] _0849_ _0871_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__mux2_1
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1342_ _0729_ _0828_ _0736_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__o21ai_1
X_1273_ net2 _0740_ _0742_ po_0.muxf_0.rf_w_data\[1\] VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__a22o_1
X_0988_ po_0.regf_0.rf\[4\]\[1\] po_0.regf_0.rf\[5\]\[1\] po_0.regf_0.rf\[6\]\[1\]
+ po_0.regf_0.rf\[7\]\[1\] _0529_ _0530_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__mux4_1
Xfanout102 net107 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
X_1609_ _0285_ _0297_ _0298_ _0307_ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__o32ai_4
XFILLER_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1891_ net103 _0069_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1960_ net97 _0126_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_0911_ _0461_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1325_ po_0.regf_0.rf\[5\]\[5\] _0813_ _0757_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__mux2_1
X_1256_ net1 _0741_ _0743_ po_0.muxf_0.rf_w_data\[0\] _0749_ VGND VGND VPWR VPWR _0750_
+ sky130_fd_sc_hd__a221o_2
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1187_ _0694_ VGND VGND VPWR VPWR _2018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ po_0.regf_0.rf\[8\]\[6\] po_0.regf_0.rf\[9\]\[6\] po_0.regf_0.rf\[10\]\[6\]
+ po_0.regf_0.rf\[11\]\[6\] _0594_ _0595_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__mux4_1
X_1041_ _0573_ _0575_ _0520_ _0578_ VGND VGND VPWR VPWR po_0.regf_0._5_\[7\] sky130_fd_sc_hd__o22a_1
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1874_ net100 _0052_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1943_ net74 _0012_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1239_ _0732_ _0734_ VGND VGND VPWR VPWR po_0.alu_0._10_\[6\] sky130_fd_sc_hd__xnor2_1
X_1308_ _0451_ po_0.alu_0._11_\[4\] _0744_ net50 VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__a22oi_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1590_ _0261_ _0302_ _0276_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__o21ai_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1024_ _0558_ _0560_ _0520_ _0563_ VGND VGND VPWR VPWR po_0.regf_0._5_\[5\] sky130_fd_sc_hd__o22a_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1857_ net89 _0039_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1926_ net85 _0104_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1788_ _0403_ _0667_ _0405_ _0658_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__a211o_2
XFILLER_25_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1642_ _0756_ po_0.regf_0.w_addr\[1\] _0839_ _0755_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__and4bb_2
X_1711_ po_0.regf_0.rf\[2\]\[5\] _0812_ _0383_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux2_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_2 po_0.regf_0._5_\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ _0283_ _0284_ _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__o21ai_1
X_1007_ _0543_ _0545_ _0520_ _0548_ VGND VGND VPWR VPWR po_0.regf_0._5_\[3\] sky130_fd_sc_hd__o22a_1
XFILLER_26_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1909_ net93 _0087_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1625_ net44 VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__inv_2
X_1556_ uc_0._21_\[2\] net57 VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__nor2_2
X_1487_ po_0.regf_0.rf\[14\]\[5\] _0851_ _0216_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__mux2_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2039_ net91 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1410_ _0876_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
X_1341_ _0816_ _0817_ _0732_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__a21oi_1
X_1272_ _0761_ _0762_ _0763_ _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__a31o_1
XFILLER_51_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0987_ po_0.regf_0.rf\[0\]\[1\] po_0.regf_0.rf\[1\]\[1\] po_0.regf_0.rf\[2\]\[1\]
+ po_0.regf_0.rf\[3\]\[1\] _0529_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__mux4_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout103 net107 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlymetal6s2s_1
X_1539_ net38 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__clkbuf_2
X_1608_ _0303_ _0304_ _0305_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1890_ net105 _0068_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0910_ _0448_ _0452_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__or2b_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1324_ _0812_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__clkbuf_2
X_1186_ _0464_ _0683_ _0472_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__mux2_1
X_1255_ _0744_ _0746_ _0747_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__o211a_1
XFILLER_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1040_ _0576_ _0577_ _0510_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1942_ net72 _0112_ VGND VGND VPWR VPWR uc_0._00_ sky130_fd_sc_hd__dfxtp_1
X_1873_ net83 _0051_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1169_ _0684_ VGND VGND VPWR VPWR _2000_/D sky130_fd_sc_hd__clkbuf_1
X_1238_ _0726_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__nor2_1
X_1307_ _0791_ _0794_ _0762_ _0796_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__o211ai_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1023_ _0561_ _0562_ _0510_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__mux2_1
XFILLER_19_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1925_ net71 _0103_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dfxtp_2
X_1856_ net104 _0038_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1787_ _0362_ net52 _0670_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__a21o_1
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1710_ _0389_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
X_1641_ _0335_ _0264_ _0347_ _0350_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__a22oi_1
XANTENNA_3 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1572_ _0679_ net57 _0285_ _0283_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__o22ai_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1006_ _0546_ _0547_ _0510_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1908_ net102 _0086_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1839_ po_0.regf_0._3_\[5\] net52 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlxtp_1
XFILLER_57_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput40 net40 VGND VGND VPWR VPWR I_addr[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_63_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1624_ _0327_ _0334_ _0257_ _0324_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__o2bb2a_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1555_ _0267_ _0268_ _0269_ _0257_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__o31ai_1
X_1486_ _0222_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1340_ _0729_ _0826_ _0819_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__nand3b_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1271_ _0450_ po_0.alu_0._11_\[1\] _0744_ _0478_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__a22o_1
X_0986_ _0005_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__buf_2
XFILLER_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1469_ _0813_ po_0.regf_0.rf\[15\]\[5\] _0206_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__mux2_1
Xfanout104 net107 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlymetal6s2s_1
X_1607_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__inv_2
X_1538_ uc_0._01_ _0248_ _0251_ _0254_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__a31o_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1323_ _0810_ _0811_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__nand2_2
X_1185_ _0693_ VGND VGND VPWR VPWR _2017_/D sky130_fd_sc_hd__clkbuf_1
X_1254_ _0740_ _0742_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__nor2_2
X_0969_ _0006_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__clkbuf_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1872_ net86 _0050_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_1941_ net63 net16 VGND VGND VPWR VPWR uc_0._21_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1306_ _0795_ _0791_ _0793_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__o21ai_1
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1099_ po_0.regf_0.rf\[4\]\[4\] po_0.regf_0.rf\[5\]\[4\] po_0.regf_0.rf\[6\]\[4\]
+ po_0.regf_0.rf\[7\]\[4\] _0579_ _0581_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__mux4_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1168_ po_0.muxf_0.rf_w_data\[5\] _0683_ _0488_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__mux2_1
X_1237_ po_0._1_\[5\] net24 VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__and2b_1
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1022_ po_0.regf_0.rf\[4\]\[5\] po_0.regf_0.rf\[5\]\[5\] po_0.regf_0.rf\[6\]\[5\]
+ po_0.regf_0.rf\[7\]\[5\] _0501_ _0503_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__mux4_1
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1855_ net104 _0037_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1924_ net71 _0102_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dfxtp_2
X_1786_ _0657_ _0493_ uc_0.bc_0._85_\[3\] _0361_ net55 VGND VGND VPWR VPWR _0169_
+ sky130_fd_sc_hd__a32o_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1640_ _0348_ _0349_ _0252_ _0264_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__a31oi_1
XANTENNA_4 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1571_ uc_0._21_\[3\] net40 VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__nor2_2
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1005_ po_0.regf_0.rf\[4\]\[3\] po_0.regf_0.rf\[5\]\[3\] po_0.regf_0.rf\[6\]\[3\]
+ po_0.regf_0.rf\[7\]\[3\] _0529_ _0530_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__mux4_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1907_ net103 _0085_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1838_ po_0.regf_0._3_\[4\] net53 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlxtp_1
X_1769_ po_0.muxf_0.rf_w_data\[3\] net30 _0418_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__mux2_1
XFILLER_57_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput30 net30 VGND VGND VPWR VPWR D_addr[3] sky130_fd_sc_hd__clkbuf_4
Xoutput41 net41 VGND VGND VPWR VPWR I_addr[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_48_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1485_ po_0.regf_0.rf\[14\]\[4\] _0849_ _0216_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__mux2_1
X_1623_ _0332_ _0248_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__nand3_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1554_ _0249_ _0255_ _0266_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__and3_1
.ends

