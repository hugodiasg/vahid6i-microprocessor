* NGSPICE file created from vahid6i.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

.subckt vahid6i D_R_data[0] D_R_data[10] D_R_data[11] D_R_data[12] D_R_data[13] D_R_data[14]
+ D_R_data[15] D_R_data[1] D_R_data[2] D_R_data[3] D_R_data[4] D_R_data[5] D_R_data[6]
+ D_R_data[7] D_R_data[8] D_R_data[9] D_W_data[0] D_W_data[10] D_W_data[11] D_W_data[12]
+ D_W_data[13] D_W_data[14] D_W_data[15] D_W_data[1] D_W_data[2] D_W_data[3] D_W_data[4]
+ D_W_data[5] D_W_data[6] D_W_data[7] D_W_data[8] D_W_data[9] D_addr[0] D_addr[1]
+ D_addr[2] D_addr[3] D_addr[4] D_addr[5] D_addr[6] D_addr[7] D_rd D_wr I_addr[0]
+ I_addr[10] I_addr[11] I_addr[12] I_addr[13] I_addr[14] I_addr[15] I_addr[1] I_addr[2]
+ I_addr[3] I_addr[4] I_addr[5] I_addr[6] I_addr[7] I_addr[8] I_addr[9] I_data[0]
+ I_data[10] I_data[11] I_data[12] I_data[13] I_data[14] I_data[15] I_data[1] I_data[2]
+ I_data[3] I_data[4] I_data[5] I_data[6] I_data[7] I_data[8] I_data[9] I_rd VGND
+ VPWR clock led_clock leds[0] leds[1] leds[2] leds[3] reset
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3155_ _0862_ po_0.regf_0.rf\[0\]\[11\] _1386_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__mux2_1
X_3086_ _1353_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__clkbuf_1
X_2106_ _1524_ po_0._1_\[2\] VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__nor2_1
X_2037_ _0511_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__and2b_1
XFILLER_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2939_ _1242_ _1241_ _1120_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__o21a_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2724_ po_0.regf_0.rf\[12\]\[10\] _0972_ _1070_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__mux2_1
X_2655_ _0862_ po_0.regf_0.rf\[14\]\[11\] _1031_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__mux2_1
X_2586_ po_0.regf_0.rf\[1\]\[12\] _0976_ _0984_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__mux2_1
Xfanout127 net130 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout138 net141 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
Xfanout105 net106 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
Xfanout116 net117 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout149 net152 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3207_ _1420_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3138_ _0778_ po_0.regf_0.rf\[0\]\[3\] _1379_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__mux2_1
XFILLER_67_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3069_ _1555_ net28 _1344_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__mux2_1
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2440_ _0911_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
X_2371_ _0773_ po_0.alu_0._11_\[10\] _0746_ _1522_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__a22o_1
XFILLER_68_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2707_ po_0.regf_0.rf\[12\]\[2\] _0955_ _1063_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__mux2_1
X_3687_ net182 _0335_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dfxtp_1
X_2638_ _0778_ po_0.regf_0.rf\[14\]\[3\] _1024_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__mux2_1
X_2569_ po_0.regf_0.rf\[1\]\[4\] _0959_ _0985_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__mux2_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1940_ _0459_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__clkbuf_4
XFILLER_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1871_ po_0.regf_0.rf\[8\]\[11\] po_0.regf_0.rf\[9\]\[11\] po_0.regf_0.rf\[10\]\[11\]
+ po_0.regf_0.rf\[11\]\[11\] _1597_ _1598_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux4_1
X_3610_ net137 _0258_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3541_ net183 _0193_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfxtp_1
X_3472_ net100 _0124_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2423_ _0897_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
X_2354_ net15 _0823_ _0834_ _0753_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__a22o_2
XFILLER_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2285_ _0770_ _0761_ _0621_ _0619_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__a211oi_1
XFILLER_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2070_ po_0.regf_0.rf\[4\]\[14\] po_0.regf_0.rf\[5\]\[14\] po_0.regf_0.rf\[6\]\[14\]
+ po_0.regf_0.rf\[7\]\[14\] _0444_ _0445_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__mux4_1
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2972_ _1247_ _1263_ _1269_ _1237_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__and4_1
X_1923_ _0000_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__buf_4
X_1854_ _1603_ _0388_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__and2b_1
X_1785_ po_0.regf_0.rf\[12\]\[2\] po_0.regf_0.rf\[13\]\[2\] po_0.regf_0.rf\[14\]\[2\]
+ po_0.regf_0.rf\[15\]\[2\] _1562_ _1564_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__mux4_1
X_3524_ net145 _0176_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3455_ net122 _0107_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_2406_ _0880_ _0752_ _0881_ _0823_ net5 VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__a32o_2
X_3386_ net158 _0042_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_2337_ _0658_ _0763_ _1488_ _0732_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__o311a_1
X_2268_ _0755_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2199_ _0691_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__clkbuf_2
XFILLER_65_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_5 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _1437_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__buf_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ po_0.regf_0.rf\[2\]\[2\] _0767_ _1398_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__mux2_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2122_ _0611_ _0612_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__nand2_1
XFILLER_66_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2053_ _0450_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__and2b_1
XFILLER_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2955_ _1249_ _1253_ _1242_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__o21a_1
X_1906_ po_0.regf_0.rf\[0\]\[15\] po_0.regf_0.rf\[1\]\[15\] po_0.regf_0.rf\[2\]\[15\]
+ po_0.regf_0.rf\[3\]\[15\] _1600_ _1601_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__mux4_1
X_2886_ uc_0._21_\[5\] _1193_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__nand2_1
X_1837_ po_0.regf_0.rf\[0\]\[7\] po_0.regf_0.rf\[1\]\[7\] po_0.regf_0.rf\[2\]\[7\]
+ po_0.regf_0.rf\[3\]\[7\] _1592_ _1593_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__mux4_1
X_3507_ net107 _0159_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_1768_ _1582_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__buf_2
X_1699_ net83 net84 net41 net40 VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__nor4_1
X_3438_ net159 _0090_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ po_0.regf_0._3_\[9\] net89 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlxtp_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput42 net42 VGND VGND VPWR VPWR D_W_data[1] sky130_fd_sc_hd__buf_2
Xoutput75 net75 VGND VGND VPWR VPWR I_addr[8] sky130_fd_sc_hd__clkbuf_4
Xoutput53 net53 VGND VGND VPWR VPWR D_addr[2] sky130_fd_sc_hd__buf_2
Xoutput64 net96 VGND VGND VPWR VPWR I_addr[12] sky130_fd_sc_hd__buf_2
XFILLER_0_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2740_ po_0.regf_0.rf\[11\]\[1\] _0953_ _1082_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__mux2_1
X_2671_ _0768_ po_0.regf_0.rf\[13\]\[2\] _1043_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__mux2_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3223_ po_0.regf_0.rf\[8\]\[10\] _0852_ _1424_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__mux2_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3154_ _1391_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__clkbuf_1
X_3085_ uc_0._21_\[13\] net21 _1343_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__mux2_1
X_2105_ _1524_ po_0._1_\[2\] VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__and2_1
X_2036_ po_0.regf_0.rf\[8\]\[10\] po_0.regf_0.rf\[9\]\[10\] po_0.regf_0.rf\[10\]\[10\]
+ po_0.regf_0.rf\[11\]\[10\] _0512_ _0513_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__mux4_1
XFILLER_35_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2938_ _1241_ _1242_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__nand2_1
X_2869_ _1161_ _1135_ _1178_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__o21ba_1
XFILLER_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2723_ _1074_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2654_ _1036_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
X_2585_ _0998_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
Xfanout128 net130 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
Xfanout106 net126 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout117 net125 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout139 net141 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlymetal6s2s_1
X_3206_ po_0.regf_0.rf\[8\]\[2\] _0767_ _1417_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__mux2_1
X_3137_ _1382_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3068_ _1343_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__buf_2
XFILLER_23_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2019_ po_0.regf_0.rf\[8\]\[8\] po_0.regf_0.rf\[9\]\[8\] po_0.regf_0.rf\[10\]\[8\]
+ po_0.regf_0.rf\[11\]\[8\] _0512_ _0513_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__mux4_1
XFILLER_23_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2370_ _0847_ _0678_ _0677_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__nand3_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2706_ _1065_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
X_3686_ net175 _0334_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfxtp_2
X_2637_ _1027_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
X_2568_ _0989_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2499_ _0944_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1870_ _0402_ _1571_ _1589_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__a21o_1
X_3540_ net181 _0192_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfxtp_1
X_3471_ net120 _0123_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_2422_ po_0.regf_0.rf\[5\]\[14\] _0896_ _0743_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__mux2_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2353_ net86 _0747_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__a21o_1
X_2284_ _1524_ po_0._1_\[2\] VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__nand2_1
X_1999_ _0520_ _0462_ _0493_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__a21bo_1
X_3669_ net175 _0317_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2971_ _1271_ _1270_ _1262_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__nand3b_1
X_1922_ _0449_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__buf_2
X_1853_ po_0.regf_0.rf\[0\]\[9\] po_0.regf_0.rf\[1\]\[9\] po_0.regf_0.rf\[2\]\[9\]
+ po_0.regf_0.rf\[3\]\[9\] _1597_ _1598_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__mux4_1
X_1784_ _1590_ _1595_ _1596_ _1604_ VGND VGND VPWR VPWR po_0.regf_0._5_\[1\] sky130_fd_sc_hd__o22a_1
X_3523_ net108 _0175_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_3454_ net164 _0106_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_2405_ net83 _0763_ _1487_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__or3_1
XFILLER_69_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3385_ net115 _0041_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2336_ _0813_ _0816_ _0817_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__o21ai_1
X_2267_ _0751_ _0753_ _0754_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__a21o_2
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2198_ _0689_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__nor2_1
XFILLER_52_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_6 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _1400_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2121_ _0614_ _0615_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__nand2_1
X_2052_ po_0.regf_0.rf\[8\]\[12\] po_0.regf_0.rf\[9\]\[12\] po_0.regf_0.rf\[10\]\[12\]
+ po_0.regf_0.rf\[11\]\[12\] _0472_ _0473_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__mux4_1
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2954_ net98 net62 VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__xnor2_1
X_1905_ _1603_ _0433_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__and2b_1
X_2885_ net72 VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__clkbuf_2
X_1836_ _0372_ _1567_ _0007_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__a21o_1
X_1767_ po_0.regf_0.rf\[12\]\[1\] po_0.regf_0.rf\[13\]\[1\] po_0.regf_0.rf\[14\]\[1\]
+ po_0.regf_0.rf\[15\]\[1\] _1562_ _1564_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__mux4_1
X_3506_ net112 _0158_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_1698_ net46 net45 net48 _1526_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__nor4_1
X_3437_ net116 _0089_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ po_0.regf_0._3_\[8\] net88 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlxtp_1
XFILLER_66_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _0784_ _0800_ _0801_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__a21oi_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3299_ _1472_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__buf_2
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput43 net43 VGND VGND VPWR VPWR D_W_data[2] sky130_fd_sc_hd__buf_2
Xoutput76 net76 VGND VGND VPWR VPWR I_addr[9] sky130_fd_sc_hd__clkbuf_4
Xoutput65 net95 VGND VGND VPWR VPWR I_addr[13] sky130_fd_sc_hd__buf_2
Xoutput54 net54 VGND VGND VPWR VPWR D_addr[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2670_ _1045_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
X_3222_ _1428_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3153_ _0853_ po_0.regf_0.rf\[0\]\[10\] _1386_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__mux2_1
X_2104_ _0604_ _0607_ VGND VGND VPWR VPWR po_0.alu_0._10_\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3084_ _1352_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2035_ _0552_ _0530_ _0493_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__a21bo_1
XFILLER_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2937_ net75 _1221_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__xor2_1
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2868_ _1173_ _1174_ _1177_ _1134_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__o211a_1
X_2799_ _1115_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__clkbuf_1
X_1819_ po_0.regf_0.rf\[0\]\[5\] po_0.regf_0.rf\[1\]\[5\] po_0.regf_0.rf\[2\]\[5\]
+ po_0.regf_0.rf\[3\]\[5\] _1609_ _1610_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__mux4_1
XFILLER_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2722_ po_0.regf_0.rf\[12\]\[9\] _0970_ _1070_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__mux2_1
XFILLER_8_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2653_ _0853_ po_0.regf_0.rf\[14\]\[10\] _1031_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__mux2_1
X_2584_ po_0.regf_0.rf\[1\]\[11\] _0974_ _0992_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__mux2_1
XFILLER_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout107 net111 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout129 net130 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout118 net121 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlymetal6s2s_1
X_3205_ _1419_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__clkbuf_1
X_3136_ _0768_ po_0.regf_0.rf\[0\]\[2\] _1379_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__mux2_1
XFILLER_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3067_ uc_0._03_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_82_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2018_ _0537_ _0530_ _0493_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__a21bo_1
XFILLER_42_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3685_ net184 _0333_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfxtp_2
X_2705_ po_0.regf_0.rf\[12\]\[1\] _0953_ _1063_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__mux2_1
X_2636_ _0768_ po_0.regf_0.rf\[14\]\[2\] _1024_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__mux2_1
X_2567_ po_0.regf_0.rf\[1\]\[3\] _0957_ _0985_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__mux2_1
X_2498_ _0862_ po_0.regf_0.rf\[7\]\[11\] _0938_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__mux2_1
XFILLER_59_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3119_ _1372_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3470_ net159 _0122_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_2421_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2352_ _0831_ _0832_ _0763_ po_0.alu_0._11_\[8\] VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__a2bb2o_1
X_2283_ _0769_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1998_ po_0.regf_0.rf\[12\]\[6\] po_0.regf_0.rf\[13\]\[6\] po_0.regf_0.rf\[14\]\[6\]
+ po_0.regf_0.rf\[15\]\[6\] _0458_ _0460_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__mux4_1
X_3668_ net174 _0316_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[2\] sky130_fd_sc_hd__dfxtp_1
X_2619_ po_0.regf_0.rf\[15\]\[11\] _0974_ _1011_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__mux2_1
X_3599_ net159 _0247_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2970_ _1262_ _1270_ _1271_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__a21bo_1
X_1921_ _0002_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1852_ _0381_ _0383_ _0385_ _0387_ VGND VGND VPWR VPWR po_0.regf_0._5_\[8\] sky130_fd_sc_hd__o22a_1
X_1783_ _1599_ _1602_ _1603_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__mux2_1
X_3522_ net112 _0174_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_3453_ net124 _0105_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_2404_ _0877_ _0878_ _0762_ _0879_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__a31o_1
X_3384_ net118 _0040_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_2335_ _1491_ po_0.alu_0._11_\[7\] _0731_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__o21ai_1
X_2266_ po_0.muxf_0.rf_w_data\[1\] _0725_ _0727_ net8 VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__a22o_1
XFILLER_37_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2197_ net84 po_0._1_\[12\] VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__nor2_1
XFILLER_25_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_7 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2120_ _0615_ _0613_ _0619_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__o2bb2ai_1
X_2051_ _0566_ _0530_ _0003_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__a21bo_1
XFILLER_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2953_ _1247_ _1134_ _1251_ _1256_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__o22a_1
X_1904_ po_0.regf_0.rf\[8\]\[15\] po_0.regf_0.rf\[9\]\[15\] po_0.regf_0.rf\[10\]\[15\]
+ po_0.regf_0.rf\[11\]\[15\] _1597_ _1598_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux4_1
X_2884_ uc_0._21_\[5\] net72 VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__or2_1
X_1835_ po_0.regf_0.rf\[4\]\[7\] po_0.regf_0.rf\[5\]\[7\] po_0.regf_0.rf\[6\]\[7\]
+ po_0.regf_0.rf\[7\]\[7\] _0352_ _0353_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__mux4_1
X_1766_ _1569_ _1577_ _1584_ _1587_ VGND VGND VPWR VPWR po_0.regf_0._5_\[0\] sky130_fd_sc_hd__o22a_1
X_3505_ net127 _0157_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_1697_ net47 VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__clkbuf_2
X_3436_ net120 _0088_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ po_0.regf_0._3_\[7\] net88 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlxtp_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _0650_ _0647_ _0648_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__or3_1
X_3298_ _1439_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__clkbuf_4
X_2249_ po_0.regf_0.w_wr VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__clkbuf_2
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput66 net94 VGND VGND VPWR VPWR I_addr[14] sky130_fd_sc_hd__clkbuf_4
Xoutput44 net44 VGND VGND VPWR VPWR D_W_data[3] sky130_fd_sc_hd__clkbuf_4
Xoutput55 net55 VGND VGND VPWR VPWR D_addr[4] sky130_fd_sc_hd__buf_2
Xoutput77 net77 VGND VGND VPWR VPWR I_rd sky130_fd_sc_hd__clkbuf_4
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3221_ po_0.regf_0.rf\[8\]\[9\] _0843_ _1424_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__mux2_1
X_3152_ _1390_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2103_ _0605_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__nor2_1
X_3083_ uc_0._21_\[12\] net20 _1343_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__mux2_1
X_2034_ po_0.regf_0.rf\[12\]\[10\] po_0.regf_0.rf\[13\]\[10\] po_0.regf_0.rf\[14\]\[10\]
+ po_0.regf_0.rf\[15\]\[10\] _0458_ _0460_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__mux4_1
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2936_ _1238_ _1217_ _1240_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__o21ai_4
X_2867_ _1123_ _1133_ _1144_ _1161_ _1176_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__a41o_1
X_1818_ _1591_ _0356_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__and2b_1
X_2798_ po_0.regf_0.rf\[10\]\[12\] _0976_ _1100_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__mux2_1
X_1749_ _1570_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__clkbuf_2
XFILLER_77_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3419_ net162 _0071_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2721_ _1073_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2652_ _1035_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
X_2583_ _0997_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
Xfanout108 net111 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
Xfanout119 net121 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_1
X_3204_ po_0.regf_0.rf\[8\]\[1\] _0755_ _1417_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__mux2_1
X_3135_ _1381_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3066_ _1342_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__clkbuf_1
X_2017_ po_0.regf_0.rf\[12\]\[8\] po_0.regf_0.rf\[13\]\[8\] po_0.regf_0.rf\[14\]\[8\]
+ po_0.regf_0.rf\[15\]\[8\] _0458_ _0460_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__mux4_1
XFILLER_35_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2919_ uc_0._21_\[7\] _1222_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__or2_1
XFILLER_5_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3684_ net184 _0332_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfxtp_1
X_2704_ _1064_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__clkbuf_1
X_2635_ _1026_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
X_2566_ _0988_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
X_2497_ _0943_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3118_ po_0.regf_0.rf\[3\]\[10\] _0852_ _1367_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__mux2_1
XFILLER_55_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3049_ _1333_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout90 po_0.regf_0.rp_rd VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_2
X_2420_ net6 _0728_ _0894_ _0752_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__a22o_2
X_2351_ _0668_ _0827_ _0830_ _0730_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__a31o_1
X_2282_ po_0.regf_0.rf\[5\]\[2\] _0768_ _0744_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__mux2_1
XFILLER_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1997_ _0510_ _0515_ _0517_ _0519_ VGND VGND VPWR VPWR po_0.regf_0._3_\[5\] sky130_fd_sc_hd__o22a_1
X_3667_ net167 _0315_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[1\] sky130_fd_sc_hd__dfxtp_1
X_3598_ net144 _0246_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2618_ _1016_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
X_2549_ _0977_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1920_ _0446_ _0447_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__nand2_1
X_1851_ _1585_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__and2b_1
X_3521_ net128 _0173_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_1782_ _0006_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__buf_2
X_3452_ net122 _0104_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_3383_ net154 _0039_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2403_ _0773_ po_0.alu_0._11_\[13\] _0746_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__a21o_1
X_2334_ _0647_ _0802_ _0814_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__o211a_1
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2265_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__clkbuf_2
X_2196_ net84 po_0._1_\[12\] VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__and2_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_8 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2050_ po_0.regf_0.rf\[12\]\[12\] po_0.regf_0.rf\[13\]\[12\] po_0.regf_0.rf\[14\]\[12\]
+ po_0.regf_0.rf\[15\]\[12\] _0488_ _0489_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__mux4_1
XFILLER_81_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2952_ _1252_ _1254_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__a21boi_1
X_1903_ _0431_ _1571_ _1582_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__a21o_1
X_2883_ _1179_ _1135_ _1182_ _1191_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__o22a_1
X_1834_ _0371_ VGND VGND VPWR VPWR po_0.regf_0._5_\[6\] sky130_fd_sc_hd__clkbuf_1
X_1765_ _1585_ _1586_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__and2b_1
X_3504_ net107 _0156_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3435_ net156 _0087_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1696_ _1513_ net87 net44 _1524_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__nor4_1
X_3366_ po_0.regf_0._3_\[6\] net89 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlxtp_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _0629_ _0630_ _0651_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__a21oi_1
X_3297_ _1435_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__inv_2
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ po_0.regf_0.w_addr\[3\] VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2179_ po_0._1_\[8\] net86 VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__or2b_1
XFILLER_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput56 net56 VGND VGND VPWR VPWR D_addr[5] sky130_fd_sc_hd__buf_2
Xoutput45 net45 VGND VGND VPWR VPWR D_W_data[4] sky130_fd_sc_hd__clkbuf_4
Xoutput67 net67 VGND VGND VPWR VPWR I_addr[15] sky130_fd_sc_hd__buf_2
Xoutput78 net78 VGND VGND VPWR VPWR led_clock sky130_fd_sc_hd__clkbuf_4
XFILLER_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3220_ _1427_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__clkbuf_1
X_3151_ _0844_ po_0.regf_0.rf\[0\]\[9\] _1386_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__mux2_1
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2102_ net87 po_0._1_\[1\] VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__nor2_1
X_3082_ _1351_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__clkbuf_1
X_2033_ _0545_ _0547_ _0549_ _0551_ VGND VGND VPWR VPWR po_0.regf_0._3_\[9\] sky130_fd_sc_hd__o22a_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2935_ _1239_ _1226_ _1224_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__a21bo_1
X_2866_ _1161_ _1175_ _1126_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__o21ai_1
X_1817_ po_0.regf_0.rf\[8\]\[5\] po_0.regf_0.rf\[9\]\[5\] po_0.regf_0.rf\[10\]\[5\]
+ po_0.regf_0.rf\[11\]\[5\] _1592_ _1593_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux4_1
X_2797_ _1114_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1748_ _0006_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__buf_2
X_1679_ _1511_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__clkbuf_1
X_3418_ net166 _0070_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3349_ po_0.regf_0._5_\[5\] po_0.regf_0.rq_rd VGND VGND VPWR VPWR po_0._1_\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2720_ po_0.regf_0.rf\[12\]\[8\] _0968_ _1070_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__mux2_1
X_2651_ _0844_ po_0.regf_0.rf\[14\]\[9\] _1031_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__mux2_1
X_2582_ po_0.regf_0.rf\[1\]\[10\] _0972_ _0992_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__mux2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout109 net110 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlymetal6s2s_1
X_3203_ _1418_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__clkbuf_1
X_3134_ _0756_ po_0.regf_0.rf\[0\]\[1\] _1379_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__mux2_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3065_ _1549_ net27 _1337_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__mux2_1
X_2016_ _0531_ _0533_ _0471_ _0536_ VGND VGND VPWR VPWR po_0.regf_0._3_\[7\] sky130_fd_sc_hd__o22a_1
XFILLER_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2918_ uc_0._21_\[6\] net73 _1221_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__or4b_2
XFILLER_31_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2849_ _1144_ _1135_ _1148_ _1159_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__o22a_1
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2703_ po_0.regf_0.rf\[12\]\[0\] _0949_ _1063_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__mux2_1
X_3683_ net188 _0331_ VGND VGND VPWR VPWR po_0.muxf_0.s1 sky130_fd_sc_hd__dfxtp_1
X_2634_ _0756_ po_0.regf_0.rf\[14\]\[1\] _1024_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__mux2_1
X_2565_ po_0.regf_0.rf\[1\]\[2\] _0955_ _0985_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__mux2_1
X_2496_ _0853_ po_0.regf_0.rf\[7\]\[10\] _0938_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__mux2_1
XFILLER_59_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3117_ _1371_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3048_ po_0.regf_0.rf\[4\]\[12\] _0873_ _1318_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__mux2_1
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout91 net93 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2350_ _0827_ _0830_ _0668_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__a21oi_2
X_2281_ _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__clkbuf_2
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1996_ _0487_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__and2b_1
X_3666_ net179 _0314_ VGND VGND VPWR VPWR po_0.regf_0.rp_addr\[0\] sky130_fd_sc_hd__dfxtp_1
X_3597_ net138 _0245_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2617_ po_0.regf_0.rf\[15\]\[10\] _0972_ _1011_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__mux2_1
X_2548_ po_0.regf_0.rf\[9\]\[12\] _0976_ _0950_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__mux2_1
X_2479_ _0768_ po_0.regf_0.rf\[7\]\[2\] _0931_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__mux2_1
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1850_ po_0.regf_0.rf\[8\]\[8\] po_0.regf_0.rf\[9\]\[8\] po_0.regf_0.rf\[10\]\[8\]
+ po_0.regf_0.rf\[11\]\[8\] _1573_ _1575_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__mux4_1
X_1781_ po_0.regf_0.rf\[4\]\[1\] po_0.regf_0.rf\[5\]\[1\] po_0.regf_0.rf\[6\]\[1\]
+ po_0.regf_0.rf\[7\]\[1\] _1600_ _1601_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__mux4_1
X_3520_ net110 _0172_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3451_ net162 _0103_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2402_ _0869_ _0692_ _0689_ _0701_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__a211o_1
X_3382_ net155 _0038_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2333_ net48 po_0._1_\[7\] VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__or2_1
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2264_ _0732_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__clkbuf_2
XFILLER_57_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2195_ _0685_ _0688_ VGND VGND VPWR VPWR po_0.alu_0._10_\[11\] sky130_fd_sc_hd__xnor2_1
XFILLER_25_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1979_ po_0.regf_0.rf\[0\]\[4\] po_0.regf_0.rf\[1\]\[4\] po_0.regf_0.rf\[2\]\[4\]
+ po_0.regf_0.rf\[3\]\[4\] _0466_ _0467_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__mux4_1
X_3718_ po_0.alu_0._10_\[15\] _1639_ VGND VGND VPWR VPWR po_0.alu_0._11_\[15\] sky130_fd_sc_hd__ebufn_1
XFILLER_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3649_ net178 _0297_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2951_ _1252_ _1254_ _1120_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__o21a_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1902_ po_0.regf_0.rf\[12\]\[15\] po_0.regf_0.rf\[13\]\[15\] po_0.regf_0.rf\[14\]\[15\]
+ po_0.regf_0.rf\[15\]\[15\] _0352_ _0353_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__mux4_1
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2882_ _1183_ _1188_ _1190_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__o21ba_1
X_1833_ _0365_ _0370_ _1582_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__mux2_1
X_1764_ po_0.regf_0.rf\[8\]\[0\] po_0.regf_0.rf\[9\]\[0\] po_0.regf_0.rf\[10\]\[0\]
+ po_0.regf_0.rf\[11\]\[0\] _1573_ _1575_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__mux4_1
X_3503_ net122 _0155_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_1695_ net43 VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__clkbuf_2
X_3434_ net159 _0086_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3365_ po_0.regf_0._3_\[5\] net90 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlxtp_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _1470_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__clkbuf_1
X_2316_ _0773_ po_0.alu_0._11_\[6\] _0746_ _1526_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__a22o_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2178_ _0673_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__inv_2
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput35 net35 VGND VGND VPWR VPWR D_W_data[0] sky130_fd_sc_hd__buf_2
Xoutput46 net46 VGND VGND VPWR VPWR D_W_data[5] sky130_fd_sc_hd__buf_2
Xoutput57 net57 VGND VGND VPWR VPWR D_addr[6] sky130_fd_sc_hd__clkbuf_4
Xoutput79 net79 VGND VGND VPWR VPWR leds[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput68 net99 VGND VGND VPWR VPWR I_addr[1] sky130_fd_sc_hd__buf_2
XFILLER_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3150_ _1389_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2101_ net87 po_0._1_\[1\] VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__and2_1
X_3081_ uc_0._21_\[11\] net19 _1343_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__mux2_1
X_2032_ _0550_ _0447_ _0443_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__a21o_1
X_2934_ _1555_ _1193_ _1210_ _1211_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__a2bb2o_1
X_2865_ _1122_ net68 _1144_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__and3_1
X_1816_ _0354_ _1567_ _1589_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__a21o_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2796_ po_0.regf_0.rf\[10\]\[11\] _0974_ _1108_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__mux2_1
X_1747_ _1565_ _1567_ _1568_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__a21o_1
X_1678_ _1499_ _1492_ VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__or2_1
X_3417_ net150 _0069_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3348_ po_0.regf_0._5_\[4\] po_0.regf_0.rq_rd VGND VGND VPWR VPWR po_0._1_\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _1461_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2650_ _1034_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
X_2581_ _0996_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3202_ po_0.regf_0.rf\[8\]\[0\] _0735_ _1417_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__mux2_1
X_3133_ _1380_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3064_ _1341_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__clkbuf_1
X_2015_ _0534_ _0535_ _0499_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__mux2_1
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2917_ _1559_ _1222_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__nand2_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2848_ _1149_ _1153_ _1154_ _1158_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__a31oi_1
X_2779_ po_0.regf_0.rf\[10\]\[3\] _0957_ _1101_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__mux2_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2702_ _1062_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__buf_2
X_3682_ net187 _0330_ VGND VGND VPWR VPWR po_0.muxf_0.s0 sky130_fd_sc_hd__dfxtp_1
X_2633_ _1025_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
X_2564_ _0987_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
X_2495_ _0942_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
X_3116_ po_0.regf_0.rf\[3\]\[9\] _0843_ _1367_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__mux2_1
XFILLER_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3047_ _1332_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout92 net93 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2280_ _0765_ _0753_ _0766_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__a21o_2
XFILLER_69_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1995_ po_0.regf_0.rf\[8\]\[5\] po_0.regf_0.rf\[9\]\[5\] po_0.regf_0.rf\[10\]\[5\]
+ po_0.regf_0.rf\[11\]\[5\] _0488_ _0489_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__mux4_1
X_3665_ net165 _0313_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[3\] sky130_fd_sc_hd__dfxtp_1
X_2616_ _1015_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
X_3596_ net144 _0244_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2547_ _0873_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__clkbuf_2
X_2478_ _0933_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1780_ _1574_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__buf_2
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3450_ net164 _0102_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3381_ net135 _0037_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2401_ _0876_ _0701_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__nand2_1
X_2332_ net48 _0659_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__nand2_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2263_ _0729_ po_0.alu_0._11_\[1\] _0747_ net87 _0750_ VGND VGND VPWR VPWR _0751_
+ sky130_fd_sc_hd__a221o_1
X_2194_ _0681_ _0686_ _0687_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1978_ _0501_ _0462_ _0470_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__a21o_1
X_3717_ po_0.alu_0._10_\[14\] _1638_ VGND VGND VPWR VPWR po_0.alu_0._11_\[14\] sky130_fd_sc_hd__ebufn_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3648_ net163 _0296_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3579_ net172 _0231_ VGND VGND VPWR VPWR uc_0._21_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2950_ _1249_ _1253_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__nor2_1
XFILLER_15_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1901_ _0430_ VGND VGND VPWR VPWR po_0.regf_0._5_\[14\] sky130_fd_sc_hd__clkbuf_1
X_2881_ _1128_ _1126_ _1189_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__or3_1
X_1832_ _0368_ _0369_ _1570_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__mux2_1
X_1763_ _1566_ VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__clkbuf_2
X_3502_ net164 _0154_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_1694_ net50 net86 net85 _1522_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__or4_1
X_3433_ net148 _0085_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ po_0.regf_0._3_\[4\] net90 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlxtp_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _0798_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
X_3295_ _1460_ _1469_ _1436_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__and3b_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ po_0.muxf_0.rf_w_data\[0\] _0725_ _0728_ net1 _0734_ VGND VGND VPWR VPWR _0735_
+ sky130_fd_sc_hd__a221o_2
X_2177_ _0672_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__clkbuf_2
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput36 net36 VGND VGND VPWR VPWR D_W_data[10] sky130_fd_sc_hd__clkbuf_4
Xoutput58 net58 VGND VGND VPWR VPWR D_addr[7] sky130_fd_sc_hd__buf_2
Xoutput47 net47 VGND VGND VPWR VPWR D_W_data[6] sky130_fd_sc_hd__buf_2
Xoutput69 net69 VGND VGND VPWR VPWR I_addr[2] sky130_fd_sc_hd__buf_2
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2100_ _1513_ po_0._1_\[0\] VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__and2b_1
X_3080_ _1350_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__clkbuf_1
X_2031_ po_0.regf_0.rf\[4\]\[9\] po_0.regf_0.rf\[5\]\[9\] po_0.regf_0.rf\[6\]\[9\]
+ po_0.regf_0.rf\[7\]\[9\] _0444_ _0445_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__mux4_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2933_ _1212_ _1213_ _1224_ _1226_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__o211ai_2
X_2864_ _1172_ _1170_ _1128_ _1126_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__a211o_1
X_1815_ po_0.regf_0.rf\[12\]\[5\] po_0.regf_0.rf\[13\]\[5\] po_0.regf_0.rf\[14\]\[5\]
+ po_0.regf_0.rf\[15\]\[5\] _0352_ _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux4_1
X_2795_ _1113_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__clkbuf_1
X_1746_ _0007_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__buf_2
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1677_ _1510_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__clkbuf_1
X_3416_ net149 _0068_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3347_ po_0.regf_0._5_\[3\] net93 VGND VGND VPWR VPWR po_0._1_\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ po_0.muxf_0.rf_w_data\[0\] _1124_ _1460_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__mux2_1
X_2229_ _0707_ po_0._1_\[14\] VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__nor2_1
XFILLER_53_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2580_ po_0.regf_0.rf\[1\]\[9\] _0970_ _0992_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__mux2_1
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3201_ _1416_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__buf_2
X_3132_ _0736_ po_0.regf_0.rf\[0\]\[0\] _1379_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__mux2_1
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3063_ _1163_ net26 _1337_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__mux2_1
XFILLER_35_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2014_ po_0.regf_0.rf\[4\]\[7\] po_0.regf_0.rf\[5\]\[7\] po_0.regf_0.rf\[6\]\[7\]
+ po_0.regf_0.rf\[7\]\[7\] _0475_ _0476_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__mux4_1
X_2916_ net74 VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2847_ _1140_ _1155_ _1156_ _1157_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__a211o_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2778_ _1104_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
X_1729_ _1554_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2701_ _0929_ _0927_ _0738_ _1061_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__and4_4
X_3681_ net187 _0329_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[7\] sky130_fd_sc_hd__dfxtp_1
X_2632_ _0736_ po_0.regf_0.rf\[14\]\[0\] _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2563_ po_0.regf_0.rf\[1\]\[1\] _0953_ _0985_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__mux2_1
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2494_ _0844_ po_0.regf_0.rf\[7\]\[9\] _0938_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__mux2_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3115_ _1370_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3046_ po_0.regf_0.rf\[4\]\[11\] _0861_ _1326_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__mux2_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout93 po_0.regf_0.rq_rd VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1994_ _0516_ _0487_ _0463_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__a21bo_1
XFILLER_9_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3664_ net160 _0312_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[2\] sky130_fd_sc_hd__dfxtp_1
X_2615_ po_0.regf_0.rf\[15\]\[9\] _0970_ _1011_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__mux2_1
X_3595_ net148 _0243_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2546_ _0975_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
X_2477_ _0756_ po_0.regf_0.rf\[7\]\[1\] _0931_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__mux2_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3029_ po_0.regf_0.rf\[4\]\[3\] _0777_ _1319_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__mux2_1
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2400_ _0869_ _0692_ _0689_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__a21o_1
X_3380_ net134 _0036_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2331_ _0647_ _0812_ _0802_ _0748_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__o31ai_1
X_2262_ _1515_ _0605_ _0606_ _0748_ _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__o311a_1
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2193_ _1522_ po_0._1_\[10\] VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__and2b_1
XFILLER_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1977_ po_0.regf_0.rf\[4\]\[4\] po_0.regf_0.rf\[5\]\[4\] po_0.regf_0.rf\[6\]\[4\]
+ po_0.regf_0.rf\[7\]\[4\] _0479_ _0480_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__mux4_1
X_3716_ po_0.alu_0._10_\[13\] _1637_ VGND VGND VPWR VPWR po_0.alu_0._11_\[13\] sky130_fd_sc_hd__ebufn_1
X_3647_ net163 _0295_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3578_ net174 _0230_ VGND VGND VPWR VPWR uc_0._21_\[6\] sky130_fd_sc_hd__dfxtp_1
X_2529_ _0950_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__buf_2
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1900_ _0426_ _0429_ _1582_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux2_1
X_2880_ _1183_ _1188_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__and2_1
X_1831_ po_0.regf_0.rf\[4\]\[6\] po_0.regf_0.rf\[5\]\[6\] po_0.regf_0.rf\[6\]\[6\]
+ po_0.regf_0.rf\[7\]\[6\] _0366_ _0367_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux4_1
X_1762_ _1580_ _1581_ _1583_ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__a21o_1
X_3501_ net124 _0153_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_1693_ net36 VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__clkbuf_2
X_3432_ net140 _0084_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3363_ po_0.regf_0._3_\[3\] net89 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlxtp_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ po_0.regf_0.rf\[5\]\[5\] _0797_ _0744_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__mux2_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ uc_0.bc_0._70_\[2\] _0593_ _1435_ po_0.muxf_0.s0 VGND VGND VPWR VPWR _1469_
+ sky130_fd_sc_hd__a31o_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _1513_ _0729_ _1488_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__o31a_1
X_2176_ _0671_ po_0._1_\[9\] VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__xor2_1
XFILLER_80_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput48 net48 VGND VGND VPWR VPWR D_W_data[7] sky130_fd_sc_hd__buf_2
XFILLER_0_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput37 net37 VGND VGND VPWR VPWR D_W_data[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput59 net59 VGND VGND VPWR VPWR D_rd sky130_fd_sc_hd__buf_2
XFILLER_16_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2030_ _0465_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__and2b_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2932_ _1206_ _1222_ net75 _1201_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__and4_1
XFILLER_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2863_ _1170_ _1172_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__nor2_1
X_1814_ _1563_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__buf_4
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2794_ po_0.regf_0.rf\[10\]\[10\] _0972_ _1108_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__mux2_1
X_1745_ _1566_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__buf_2
X_1676_ _1499_ _1492_ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__or2_1
X_3415_ net145 _0067_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3346_ po_0.regf_0._5_\[2\] net93 VGND VGND VPWR VPWR po_0._1_\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _1441_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__clkbuf_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2228_ _0707_ po_0._1_\[14\] VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__and2_1
X_2159_ _0657_ VGND VGND VPWR VPWR po_0.alu_0._10_\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_26_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3200_ po_0.regf_0.w_addr\[2\] _0737_ po_0.regf_0.w_wr _1061_ VGND VGND VPWR VPWR
+ _1416_ sky130_fd_sc_hd__and4b_4
X_3131_ _1378_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__buf_2
XFILLER_67_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3062_ _1340_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2013_ po_0.regf_0.rf\[0\]\[7\] po_0.regf_0.rf\[1\]\[7\] po_0.regf_0.rf\[2\]\[7\]
+ po_0.regf_0.rf\[3\]\[7\] _0524_ _0525_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__mux4_1
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2915_ uc_0._21_\[7\] net74 VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__nor2_1
X_2846_ _1129_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__clkbuf_2
X_2777_ po_0.regf_0.rf\[10\]\[2\] _0955_ _1101_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__mux2_1
X_1728_ po_0.regf_0.rq_addr\[0\] _1549_ _1553_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__mux2_1
X_1659_ _1500_ _1493_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__or2_1
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ net129 _0017_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2700_ _0740_ _0739_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__nor2_1
X_3680_ net179 _0328_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[6\] sky130_fd_sc_hd__dfxtp_1
X_2631_ _1023_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__buf_2
X_2562_ _0986_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
X_2493_ _0941_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3114_ po_0.regf_0.rf\[3\]\[8\] _0835_ _1367_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__mux2_1
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3045_ _1331_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2829_ _1122_ net99 _1129_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__a21boi_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout83 net39 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
Xfanout94 net66 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_4
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1993_ po_0.regf_0.rf\[12\]\[5\] po_0.regf_0.rf\[13\]\[5\] po_0.regf_0.rf\[14\]\[5\]
+ po_0.regf_0.rf\[15\]\[5\] _0479_ _0480_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__mux4_1
XFILLER_9_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3663_ net172 _0311_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[1\] sky130_fd_sc_hd__dfxtp_1
X_2614_ _1014_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_3594_ net131 _0242_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2545_ po_0.regf_0.rf\[9\]\[11\] _0974_ _0964_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__mux2_1
X_2476_ _0932_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3028_ _1322_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2330_ _0660_ _0661_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__nor2_1
X_2261_ _0605_ _0606_ po_0._1_\[0\] _1513_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_84_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2192_ _0675_ _0673_ _0680_ _0677_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__o211a_1
XFILLER_65_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1976_ _0494_ _0496_ _0471_ _0500_ VGND VGND VPWR VPWR po_0.regf_0._3_\[3\] sky130_fd_sc_hd__o22a_1
XFILLER_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3715_ po_0.alu_0._10_\[12\] _1636_ VGND VGND VPWR VPWR po_0.alu_0._11_\[12\] sky130_fd_sc_hd__ebufn_1
X_3646_ net151 _0294_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3577_ net172 _0229_ VGND VGND VPWR VPWR uc_0._21_\[5\] sky130_fd_sc_hd__dfxtp_1
X_2528_ _0808_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__clkbuf_2
X_2459_ _0921_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1830_ po_0.regf_0.rf\[0\]\[6\] po_0.regf_0.rf\[1\]\[6\] po_0.regf_0.rf\[2\]\[6\]
+ po_0.regf_0.rf\[3\]\[6\] _0366_ _0367_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__mux4_1
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1761_ _1582_ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__clkbuf_2
X_3500_ net123 _0152_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_1692_ _1521_ VGND VGND VPWR VPWR uc_0.bc_0._70_\[2\] sky130_fd_sc_hd__clkbuf_2
X_3431_ net143 _0083_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3362_ po_0.regf_0._3_\[2\] net90 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlxtp_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _0796_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _1468_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__clkbuf_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _1491_ po_0.alu_0._11_\[0\] _0731_ po_0.alu_0._10_\[0\] _0732_ VGND VGND VPWR
+ VPWR _0733_ sky130_fd_sc_hd__o221a_1
X_2175_ net50 VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__clkbuf_2
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1959_ po_0.regf_0.rf\[12\]\[2\] po_0.regf_0.rf\[13\]\[2\] po_0.regf_0.rf\[14\]\[2\]
+ po_0.regf_0.rf\[15\]\[2\] _0444_ _0445_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__mux4_1
X_3629_ net137 _0277_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xoutput49 net86 VGND VGND VPWR VPWR D_W_data[8] sky130_fd_sc_hd__buf_2
Xoutput38 net84 VGND VGND VPWR VPWR D_W_data[12] sky130_fd_sc_hd__buf_2
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2931_ _1235_ _1230_ _1126_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__o21ai_1
XFILLER_43_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2862_ _1149_ _1154_ _1171_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__a21oi_2
X_1813_ _1561_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__buf_4
X_2793_ _1112_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1744_ _0006_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__clkbuf_2
X_3414_ net150 _0066_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_1675_ _1509_ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__clkbuf_1
X_3345_ po_0.regf_0._5_\[1\] net93 VGND VGND VPWR VPWR po_0._1_\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3276_ _1459_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__clkbuf_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ po_0._1_\[14\] _0707_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__or2b_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2158_ _0653_ _0656_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__and2b_1
X_2089_ po_0.regf_0.rp_addr\[2\] uc_0._21_\[10\] _0596_ VGND VGND VPWR VPWR _0599_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3130_ _0929_ _0737_ _0738_ _1061_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__or4bb_4
XFILLER_79_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3061_ _1151_ net25 _1337_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__mux2_1
X_2012_ _0511_ _0532_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__and2b_1
XFILLER_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2914_ _1206_ _1134_ _1209_ _1220_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__o22a_1
X_2845_ _1128_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__buf_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2776_ _1103_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__clkbuf_1
X_1727_ _1552_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__buf_2
X_1658_ _1499_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__dlymetal6s2s_1
X_3328_ net127 _0016_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3259_ po_0.regf_0.rp_addr\[1\] uc_0._21_\[9\] _0595_ VGND VGND VPWR VPWR _1449_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2630_ _1022_ _0740_ _0739_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__or3b_4
X_2561_ po_0.regf_0.rf\[1\]\[0\] _0949_ _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__mux2_1
X_2492_ _0836_ po_0.regf_0.rf\[7\]\[8\] _0938_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__mux2_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3113_ _1369_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__clkbuf_1
X_3044_ po_0.regf_0.rf\[4\]\[10\] _0852_ _1326_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__mux2_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2828_ _1122_ uc_0._21_\[0\] _1137_ _1138_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__o22ai_1
X_2759_ po_0.regf_0.rf\[11\]\[10\] _0972_ _1089_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__mux2_1
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout95 net65 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
Xfanout84 net38 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_4
XFILLER_69_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1992_ _0511_ _0514_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__and2b_1
X_3662_ net174 _0310_ VGND VGND VPWR VPWR po_0.regf_0.rq_addr\[0\] sky130_fd_sc_hd__dfxtp_1
X_3593_ net143 _0241_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2613_ po_0.regf_0.rf\[15\]\[8\] _0968_ _1011_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__mux2_1
X_2544_ _0861_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__clkbuf_2
XFILLER_5_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2475_ _0736_ po_0.regf_0.rf\[7\]\[0\] _0931_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__mux2_1
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3027_ po_0.regf_0.rf\[4\]\[2\] _0767_ _1319_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__mux2_1
XFILLER_24_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2260_ _1490_ _1487_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__and2_2
XFILLER_77_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2191_ _0683_ _0684_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__nor2_2
XFILLER_65_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1975_ _0497_ _0498_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__mux2_1
X_3714_ po_0.alu_0._10_\[11\] _1635_ VGND VGND VPWR VPWR po_0.alu_0._11_\[11\] sky130_fd_sc_hd__ebufn_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3645_ net152 _0293_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3576_ net179 _0228_ VGND VGND VPWR VPWR uc_0._21_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2527_ _0962_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
X_2458_ po_0.regf_0.rf\[6\]\[10\] _0853_ _0916_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__mux2_1
XFILLER_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2389_ _0695_ _0672_ _0679_ _0685_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__nand4_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1760_ _0007_ VGND VGND VPWR VPWR _1582_ sky130_fd_sc_hd__clkinv_2
X_1691_ _1517_ _1520_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__and2b_1
X_3430_ net149 _0082_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3361_ po_0.regf_0._3_\[1\] net89 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlxtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2312_ po_0.muxf_0.rf_w_data\[5\] _0725_ _0728_ net12 _0795_ VGND VGND VPWR VPWR
+ _0796_ sky130_fd_sc_hd__a221o_4
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ po_0.muxf_0.rf_w_data\[7\] _1559_ _1441_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__mux2_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _0724_ _0726_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__nor2_2
X_2174_ _0668_ _0670_ VGND VGND VPWR VPWR po_0.alu_0._10_\[8\] sky130_fd_sc_hd__xor2_1
XFILLER_80_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1958_ _0465_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__and2b_1
X_1889_ _1603_ _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__and2b_1
X_3628_ net144 _0276_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xoutput39 net39 VGND VGND VPWR VPWR D_W_data[13] sky130_fd_sc_hd__clkbuf_4
X_3559_ net130 _0211_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2930_ net75 VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__clkbuf_2
X_2861_ _1150_ _1152_ _1137_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2792_ po_0.regf_0.rf\[10\]\[9\] _0970_ _1108_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__mux2_1
X_1812_ _0346_ _0348_ _1596_ _0351_ VGND VGND VPWR VPWR po_0.regf_0._5_\[4\] sky130_fd_sc_hd__o22a_1
X_1743_ po_0.regf_0.rf\[4\]\[0\] po_0.regf_0.rf\[5\]\[0\] po_0.regf_0.rf\[6\]\[0\]
+ po_0.regf_0.rf\[7\]\[0\] _1562_ _1564_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__mux4_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1674_ _1499_ _1492_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__or2_1
X_3413_ net151 _0065_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3344_ po_0.regf_0._5_\[0\] net93 VGND VGND VPWR VPWR po_0._1_\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _1458_ _0927_ _1443_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__mux2_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2226_ _0714_ _0715_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__or2_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2157_ _0652_ _0654_ _0655_ _0649_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__nand4_1
X_2088_ _0598_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3060_ _1339_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2011_ po_0.regf_0.rf\[8\]\[7\] po_0.regf_0.rf\[9\]\[7\] po_0.regf_0.rf\[10\]\[7\]
+ po_0.regf_0.rf\[11\]\[7\] _0512_ _0513_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__mux4_1
XFILLER_75_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2913_ _1218_ _1219_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__nor2_1
X_2844_ _1153_ _1154_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__nand2_1
X_2775_ po_0.regf_0.rf\[10\]\[1\] _0953_ _1101_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__mux2_1
X_1726_ _1550_ _1551_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__nand2_2
X_1657_ _1488_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3327_ _1548_ _1486_ _1119_ _1438_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__a2bb2o_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3258_ _1448_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2209_ _0700_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__clkbuf_2
X_3189_ _1410_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2560_ _0984_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__clkbuf_4
X_2491_ _0940_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3112_ po_0.regf_0.rf\[3\]\[7\] _0820_ _1367_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__mux2_1
X_3043_ _1330_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2827_ _1122_ _1124_ _1137_ _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__or4_1
X_2758_ _1093_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_1
X_1709_ _1533_ _1534_ _1537_ net34 VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__a31o_1
X_2689_ _1055_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout96 net64 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout85 net37 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
XFILLER_45_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1991_ po_0.regf_0.rf\[0\]\[5\] po_0.regf_0.rf\[1\]\[5\] po_0.regf_0.rf\[2\]\[5\]
+ po_0.regf_0.rf\[3\]\[5\] _0512_ _0513_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__mux4_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3661_ net145 _0309_ VGND VGND VPWR VPWR po_0.regf_0.w_wr sky130_fd_sc_hd__dfxtp_1
X_2612_ _1013_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3592_ net167 _0015_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__dfxtp_1
X_2543_ _0973_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
X_2474_ _0930_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__buf_2
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3026_ _1321_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2190_ net85 po_0._1_\[11\] VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__and2_1
XFILLER_77_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1974_ _0449_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__clkbuf_4
X_3713_ po_0.alu_0._10_\[10\] _1634_ VGND VGND VPWR VPWR po_0.alu_0._11_\[10\] sky130_fd_sc_hd__ebufn_1
X_3644_ net146 _0292_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3575_ net174 _0227_ VGND VGND VPWR VPWR uc_0._21_\[3\] sky130_fd_sc_hd__dfxtp_1
X_2526_ po_0.regf_0.rf\[9\]\[5\] _0961_ _0951_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__mux2_1
X_2457_ _0920_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
X_2388_ _1522_ po_0._1_\[10\] po_0._1_\[11\] net85 _0864_ VGND VGND VPWR VPWR _0865_
+ sky130_fd_sc_hd__a221oi_4
XFILLER_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3009_ _1306_ _1303_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__nand2_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1690_ uc_0._21_\[15\] uc_0._21_\[14\] _1518_ _1519_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__nor4b_2
X_3360_ po_0.regf_0._3_\[0\] net89 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlxtp_1
X_2311_ _0640_ _0763_ _1488_ _0732_ _0794_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__o311a_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _1467_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__clkbuf_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2242_ _0730_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__buf_2
X_2173_ _0663_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__nand2_1
XFILLER_65_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1957_ po_0.regf_0.rf\[0\]\[2\] po_0.regf_0.rf\[1\]\[2\] po_0.regf_0.rf\[2\]\[2\]
+ po_0.regf_0.rf\[3\]\[2\] _0466_ _0467_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__mux4_1
X_1888_ po_0.regf_0.rf\[8\]\[13\] po_0.regf_0.rf\[9\]\[13\] po_0.regf_0.rf\[10\]\[13\]
+ po_0.regf_0.rf\[11\]\[13\] _1597_ _1598_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux4_1
X_3627_ net148 _0275_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3558_ net136 _0210_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2509_ _0742_ _0927_ _0906_ _0741_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__and4b_4
X_3489_ net110 _0141_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2860_ _1166_ _1169_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__nand2_1
X_1811_ _0349_ _0350_ _1613_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__mux2_1
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2791_ _1111_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1742_ _1563_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__clkbuf_4
X_1673_ _1508_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__clkbuf_1
X_3412_ net145 _0064_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ net100 _0031_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ uc_0._21_\[11\] _1163_ _1552_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__mux2_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2225_ net41 po_0._1_\[15\] VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__and2b_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2156_ net47 po_0._1_\[6\] VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__or2_1
XFILLER_53_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2087_ po_0.regf_0.rp_addr\[1\] uc_0._21_\[9\] _0596_ VGND VGND VPWR VPWR _0598_
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2989_ _1119_ _1156_ _1248_ _1278_ _1289_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__o41a_1
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2010_ _0529_ _0530_ _0493_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__a21bo_1
XFILLER_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2912_ _1217_ _1214_ _1156_ _1127_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__a211o_1
X_2843_ _1150_ _1152_ _1137_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__nand3_1
X_2774_ _1102_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__clkbuf_1
X_1725_ _1521_ uc_0.bc_0._70_\[1\] _1546_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__nand3_1
X_1656_ _1498_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__clkbuf_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _1533_ _1534_ _1537_ _1356_ _1471_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__a311o_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ po_0.regf_0.rp_addr\[0\] uc_0._21_\[8\] _0596_ VGND VGND VPWR VPWR _1448_
+ sky130_fd_sc_hd__mux2_1
X_2208_ net83 po_0._1_\[13\] VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__xor2_1
X_3188_ po_0.regf_0.rf\[2\]\[10\] _0852_ _1405_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__mux2_1
X_2139_ _0630_ _0629_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__and2b_1
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2490_ _0821_ po_0.regf_0.rf\[7\]\[7\] _0938_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__mux2_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3111_ _1368_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3042_ po_0.regf_0.rf\[4\]\[9\] _0843_ _1326_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__mux2_1
XFILLER_36_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2826_ net99 uc_0._21_\[1\] VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__and2_1
X_2757_ po_0.regf_0.rf\[11\]\[9\] _0970_ _1089_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__mux2_1
X_1708_ _1536_ _1519_ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__nand2_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2688_ _0853_ po_0.regf_0.rf\[13\]\[10\] _1050_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__mux2_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _1163_ net54 _1472_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__mux2_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout97 net63 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout86 net49 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_2
XFILLER_10_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1990_ _0459_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__buf_2
XFILLER_60_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3660_ net189 _0308_ VGND VGND VPWR VPWR po_0.regf_0.rp_rd sky130_fd_sc_hd__dfxtp_1
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2611_ po_0.regf_0.rf\[15\]\[7\] _0966_ _1011_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__mux2_1
X_3591_ net165 _0014_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__dfxtp_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2542_ po_0.regf_0.rf\[9\]\[10\] _0972_ _0964_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__mux2_1
X_2473_ _0927_ _0738_ _0928_ _0929_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__nand4b_4
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3025_ po_0.regf_0.rf\[4\]\[1\] _0755_ _1319_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__mux2_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2809_ net61 VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__clkbuf_2
XFILLER_3_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1973_ po_0.regf_0.rf\[4\]\[3\] po_0.regf_0.rf\[5\]\[3\] po_0.regf_0.rf\[6\]\[3\]
+ po_0.regf_0.rf\[7\]\[3\] _0475_ _0476_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__mux4_1
XFILLER_60_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3712_ po_0.alu_0._10_\[9\] _1633_ VGND VGND VPWR VPWR po_0.alu_0._11_\[9\] sky130_fd_sc_hd__ebufn_1
X_3643_ net152 _0291_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3574_ net179 _0226_ VGND VGND VPWR VPWR uc_0._21_\[2\] sky130_fd_sc_hd__dfxtp_1
X_2525_ _0796_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__clkbuf_2
X_2456_ po_0.regf_0.rf\[6\]\[9\] _0844_ _0916_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__mux2_1
X_2387_ _0671_ po_0._1_\[9\] _0846_ _0679_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__o211a_1
XFILLER_83_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3008_ _1303_ _1306_ _1120_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__o21a_1
XFILLER_43_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2310_ _0791_ _0748_ _0792_ _0793_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__a31o_1
X_3290_ po_0.muxf_0.rf_w_data\[6\] _1557_ _1441_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__mux2_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _1490_ po_0.alu_0.s0 VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__nand2_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2172_ _0659_ _0658_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__or2b_1
XFILLER_18_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1956_ _0481_ _0462_ _0470_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__a21o_1
X_1887_ _0417_ _1571_ _1589_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__a21o_1
X_3626_ net131 _0274_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3557_ net135 _0209_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2508_ _0735_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__clkbuf_2
X_3488_ net100 _0140_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_2439_ po_0.regf_0.rf\[6\]\[1\] _0756_ _0909_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__mux2_1
XFILLER_29_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1810_ po_0.regf_0.rf\[4\]\[4\] po_0.regf_0.rf\[5\]\[4\] po_0.regf_0.rf\[6\]\[4\]
+ po_0.regf_0.rf\[7\]\[4\] _1600_ _1601_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__mux4_1
XFILLER_30_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2790_ po_0.regf_0.rf\[10\]\[8\] _0968_ _1108_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__mux2_1
X_1741_ _0005_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__buf_2
X_1672_ _1499_ _1502_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__or2_1
X_3411_ net164 _0011_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__dfxtp_2
X_3342_ net105 _0030_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _1457_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkbuf_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2224_ po_0._1_\[15\] net41 VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__and2b_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _1526_ po_0._1_\[6\] VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__nand2_1
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2086_ _0597_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2988_ _1284_ _1286_ _1121_ _1288_ _1131_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__a311o_1
X_1939_ _0457_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__clkbuf_4
X_3609_ net132 _0257_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2911_ _1214_ _1217_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__nor2_1
X_2842_ net99 _1136_ _1150_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__a2bb2o_1
X_2773_ po_0.regf_0.rf\[10\]\[0\] _0949_ _1101_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__mux2_1
X_1724_ _1517_ _1545_ _1538_ uc_0.bc_0._70_\[3\] VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__o211ai_2
XFILLER_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1655_ _1489_ _1493_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__or2_1
X_3325_ _1538_ _1435_ _0594_ _1473_ _1485_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__o311a_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _1447_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__clkbuf_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _0689_ _0690_ _0698_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__o21ai_1
X_3187_ _1409_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2138_ _0638_ VGND VGND VPWR VPWR po_0.alu_0._10_\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_66_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2069_ _0465_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__and2b_1
XFILLER_22_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3110_ po_0.regf_0.rf\[3\]\[6\] _0808_ _1367_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__mux2_1
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3041_ _1329_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2825_ net99 _1136_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__nor2_1
X_2756_ _1092_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
X_1707_ uc_0.bc_0._05_\[0\] _1535_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__xor2_1
X_2687_ _1054_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _1476_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3239_ _1356_ _1357_ _1546_ _0594_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__or4_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout98 net76 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
Xfanout87 net42 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2610_ _1012_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
X_3590_ net159 _0013_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__dfxtp_1
X_2541_ _0852_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2472_ po_0.regf_0.w_addr\[2\] VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__clkbuf_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3024_ _1320_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2808_ _1120_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__clkbuf_2
X_2739_ _1083_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1972_ po_0.regf_0.rf\[0\]\[3\] po_0.regf_0.rf\[1\]\[3\] po_0.regf_0.rf\[2\]\[3\]
+ po_0.regf_0.rf\[3\]\[3\] _0472_ _0473_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__mux4_1
X_3711_ po_0.alu_0._10_\[8\] _1632_ VGND VGND VPWR VPWR po_0.alu_0._11_\[8\] sky130_fd_sc_hd__ebufn_1
X_3642_ net151 _0290_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3573_ net181 _0225_ VGND VGND VPWR VPWR uc_0._21_\[1\] sky130_fd_sc_hd__dfxtp_1
X_2524_ _0960_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_2455_ _0919_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
X_2386_ _0863_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3007_ net95 _1282_ _1304_ _1305_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__o22ai_2
XFILLER_71_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ po_0.alu_0.s1 VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__buf_2
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2171_ _0666_ _0667_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__or2_2
XFILLER_65_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1955_ po_0.regf_0.rf\[4\]\[2\] po_0.regf_0.rf\[5\]\[2\] po_0.regf_0.rf\[6\]\[2\]
+ po_0.regf_0.rf\[7\]\[2\] _0479_ _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__mux4_1
X_1886_ po_0.regf_0.rf\[12\]\[13\] po_0.regf_0.rf\[13\]\[13\] po_0.regf_0.rf\[14\]\[13\]
+ po_0.regf_0.rf\[15\]\[13\] _0352_ _0353_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__mux4_1
X_3625_ net143 _0273_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3556_ net131 _0208_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2507_ _0948_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
X_3487_ net120 _0139_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_2438_ _0910_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_1
X_2369_ _0677_ _0678_ _0847_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__a21o_1
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1740_ _1561_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__clkbuf_4
X_1671_ _1507_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__clkbuf_1
X_3410_ net166 _0010_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__dfxtp_1
X_3341_ net109 _0029_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3272_ _1456_ _0929_ _1443_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__mux2_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _0712_ _0713_ VGND VGND VPWR VPWR po_0.alu_0._10_\[14\] sky130_fd_sc_hd__nor2_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _0647_ _0648_ _0649_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2085_ po_0.regf_0.rp_addr\[0\] uc_0._21_\[8\] _0596_ VGND VGND VPWR VPWR _0597_
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2987_ _1278_ _1274_ _1157_ _1287_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__o211a_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1938_ _0449_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__clkbuf_2
X_1869_ po_0.regf_0.rf\[12\]\[11\] po_0.regf_0.rf\[13\]\[11\] po_0.regf_0.rf\[14\]\[11\]
+ po_0.regf_0.rf\[15\]\[11\] _0352_ _0353_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux4_1
X_3608_ net108 _0256_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_3539_ net107 _0191_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2910_ _1183_ _1188_ _1198_ _1216_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__a31oi_4
XFILLER_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2841_ net69 _1151_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__nand2_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2772_ _1100_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__buf_2
X_1723_ uc_0._21_\[4\] VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__clkbuf_2
XFILLER_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1654_ _1497_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__clkbuf_1
X_3324_ _1248_ _1484_ _1356_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__o21ba_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ po_0.regf_0.rq_addr\[3\] _1559_ _1442_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__mux2_1
XFILLER_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2206_ _0692_ _0698_ VGND VGND VPWR VPWR po_0.alu_0._10_\[12\] sky130_fd_sc_hd__xnor2_1
X_3186_ po_0.regf_0.rf\[2\]\[9\] _0843_ _1405_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__mux2_1
X_2137_ _0634_ _0637_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__and2b_1
XFILLER_66_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2068_ po_0.regf_0.rf\[0\]\[14\] po_0.regf_0.rf\[1\]\[14\] po_0.regf_0.rf\[2\]\[14\]
+ po_0.regf_0.rf\[3\]\[14\] _0466_ _0467_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__mux4_1
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3040_ po_0.regf_0.rf\[4\]\[8\] _0835_ _1326_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__mux2_1
XFILLER_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2824_ uc_0._21_\[1\] VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__clkbuf_2
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2755_ po_0.regf_0.rf\[11\]\[8\] _0968_ _1089_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__mux2_1
X_1706_ uc_0.bc_0._05_\[1\] VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2686_ _0844_ po_0.regf_0.rf\[13\]\[9\] _1050_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__mux2_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ _1151_ net53 _1473_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__mux2_1
XFILLER_86_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _1520_ uc_0.bc_0._70_\[1\] _1435_ _1436_ _1489_ VGND VGND VPWR VPWR _0306_
+ sky130_fd_sc_hd__a32o_1
X_3169_ po_0.regf_0.rf\[2\]\[1\] _0755_ _1398_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__mux2_1
XFILLER_54_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout99 net68 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_4
Xfanout88 net89 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2540_ _0971_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2471_ po_0.regf_0.w_addr\[0\] po_0.regf_0.w_addr\[1\] VGND VGND VPWR VPWR _0928_
+ sky130_fd_sc_hd__and2_2
XFILLER_83_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3023_ po_0.regf_0.rf\[4\]\[0\] _0735_ _1319_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__mux2_1
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2807_ uc_0._00_ uc_0._02_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__nor2_2
X_2738_ po_0.regf_0.rf\[11\]\[0\] _0949_ _1082_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__mux2_1
X_2669_ _0756_ po_0.regf_0.rf\[13\]\[1\] _1043_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__mux2_1
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1971_ _0465_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__and2b_1
X_3710_ po_0.alu_0._10_\[7\] _1631_ VGND VGND VPWR VPWR po_0.alu_0._11_\[7\] sky130_fd_sc_hd__ebufn_1
X_3641_ net145 _0289_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3572_ net181 _0224_ VGND VGND VPWR VPWR uc_0._21_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2523_ po_0.regf_0.rf\[9\]\[4\] _0959_ _0951_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__mux2_1
X_2454_ po_0.regf_0.rf\[6\]\[8\] _0836_ _0916_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__mux2_1
X_2385_ po_0.regf_0.rf\[5\]\[11\] _0862_ _0810_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__mux2_1
XFILLER_68_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput1 D_R_data[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3006_ net63 _1280_ _1279_ _1241_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2170_ net86 po_0._1_\[8\] VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__nor2_1
XFILLER_65_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1954_ _0440_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__clkbuf_4
XFILLER_21_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3624_ net108 _0272_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_1885_ _0410_ _0412_ _0416_ VGND VGND VPWR VPWR po_0.regf_0._5_\[12\] sky130_fd_sc_hd__o21a_1
X_3555_ net181 _0207_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfxtp_2
X_2506_ _0904_ po_0.regf_0.rf\[7\]\[15\] _0930_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__mux2_1
X_3486_ net159 _0138_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_2437_ po_0.regf_0.rf\[6\]\[0\] _0736_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__mux2_1
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2368_ _0671_ po_0._1_\[9\] _0846_ _0831_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__o22ai_1
X_2299_ _0620_ _0618_ _0635_ _0636_ _0782_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__o2111ai_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1670_ _1500_ _1502_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__or2_1
X_3340_ net102 _0028_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ uc_0._21_\[10\] _1151_ _1552_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__mux2_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2222_ _0705_ _0708_ _0709_ _0711_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__and4_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ _0650_ _0651_ _0639_ _0634_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__o22ai_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2084_ _0595_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__buf_2
XFILLER_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2986_ _1264_ _1283_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__nand2_1
X_1937_ _0461_ _0462_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__a21bo_1
X_1868_ _0401_ VGND VGND VPWR VPWR po_0.regf_0._5_\[10\] sky130_fd_sc_hd__clkbuf_1
X_3607_ net116 _0255_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_3538_ net112 _0190_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_1799_ _1617_ _1585_ _1583_ VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__a21o_1
X_3469_ net116 _0121_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2840_ uc_0._21_\[2\] VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__clkbuf_2
XFILLER_31_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2771_ po_0.regf_0.w_addr\[2\] _0737_ po_0.regf_0.w_wr _0907_ VGND VGND VPWR VPWR
+ _1100_ sky130_fd_sc_hd__and4b_4
X_1722_ _1517_ _1548_ VGND VGND VPWR VPWR uc_0.bc_0._70_\[3\] sky130_fd_sc_hd__nor2_1
X_1653_ _1489_ _1493_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__or2_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _1535_ _1519_ _1539_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__and3b_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3254_ _1446_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__clkbuf_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _0694_ _0697_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__or2_1
X_3185_ _1408_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2136_ _0622_ _0635_ _0636_ _0633_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__nand4_1
XFILLER_66_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2067_ _0580_ _0487_ _0463_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__a21bo_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2969_ net62 net97 VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2823_ _1134_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__clkbuf_2
X_2754_ _1091_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
X_1705_ uc_0._21_\[13\] _1520_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__nand2_1
X_2685_ _1053_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
X_3306_ _1475_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__clkbuf_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _1550_ _1551_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__and2_1
X_3168_ _1399_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2119_ _0620_ _0618_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__nor2_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3099_ po_0.regf_0.rf\[3\]\[1\] _0755_ _1360_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__mux2_1
XFILLER_54_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout89 po_0.regf_0.rp_rd VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2470_ po_0.regf_0.w_addr\[3\] VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3022_ _1318_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__buf_2
XFILLER_51_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2806_ uc_0._01_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__clkbuf_2
X_2737_ _1081_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__clkbuf_4
X_2668_ _1044_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
X_2599_ _1006_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1970_ po_0.regf_0.rf\[8\]\[3\] po_0.regf_0.rf\[9\]\[3\] po_0.regf_0.rf\[10\]\[3\]
+ po_0.regf_0.rf\[11\]\[3\] _0466_ _0467_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__mux4_1
XFILLER_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ net101 _0288_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_3571_ net101 _0223_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_2522_ _0788_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__clkbuf_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2453_ _0918_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
X_2384_ _0861_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__clkbuf_2
XFILLER_68_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput2 D_R_data[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
X_3005_ _1283_ _1282_ _1292_ _1293_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1953_ _0439_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__clkbuf_4
X_1884_ _0413_ _1581_ _1568_ _0415_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a211o_1
X_3623_ net104 _0271_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_3554_ net181 _0206_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfxtp_1
X_2505_ _0947_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
X_3485_ net116 _0137_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_2436_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__buf_2
XFILLER_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2367_ net49 po_0._1_\[8\] po_0._1_\[9\] net50 VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__a22o_1
X_2298_ _0620_ _0618_ _0782_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__o21a_1
XFILLER_56_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _1455_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__clkbuf_1
X_2221_ _0708_ _0709_ _0705_ _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__a22oi_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2152_ _0640_ _0641_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__and2_1
XFILLER_26_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2083_ _0593_ uc_0.bc_0._70_\[0\] _0594_ _1552_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__a31o_2
XFILLER_19_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2985_ _1283_ _1282_ _1285_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__o21ai_1
X_1936_ _0003_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__clkbuf_2
X_1867_ _0397_ _0400_ _1582_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__mux2_1
X_3606_ net113 _0254_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_1798_ po_0.regf_0.rf\[12\]\[3\] po_0.regf_0.rf\[13\]\[3\] po_0.regf_0.rf\[14\]\[3\]
+ po_0.regf_0.rf\[15\]\[3\] _1562_ _1564_ VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__mux4_1
X_3537_ net128 _0189_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3468_ net120 _0120_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3399_ net154 _0055_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2419_ _0889_ _0892_ _0762_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__a31o_1
XFILLER_69_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2770_ _1099_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_1
X_1721_ _1541_ _1542_ _1518_ _1547_ _1533_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__o41a_1
X_1652_ _1496_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__clkbuf_1
X_3322_ _0594_ _1483_ _1482_ _1337_ _1473_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o221a_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ po_0.regf_0.rq_addr\[2\] _1557_ _1442_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__mux2_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ po_0.regf_0.rf\[2\]\[8\] _0835_ _1405_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__mux2_1
X_2204_ _0663_ _0669_ _0696_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__a21oi_1
X_2135_ net45 po_0._1_\[4\] VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__or2_1
XFILLER_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2066_ po_0.regf_0.rf\[12\]\[14\] po_0.regf_0.rf\[13\]\[14\] po_0.regf_0.rf\[14\]\[14\]
+ po_0.regf_0.rf\[15\]\[14\] _0479_ _0480_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__mux4_1
XFILLER_81_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2968_ _1263_ _1247_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__or2b_1
X_1919_ _0438_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__buf_2
X_2899_ net73 VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2822_ _1119_ _1128_ _1126_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__or3_2
X_2753_ po_0.regf_0.rf\[11\]\[7\] _0966_ _1089_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__mux2_1
X_1704_ _1530_ _1532_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__nand2_1
X_2684_ _0836_ po_0.regf_0.rf\[13\]\[8\] _1050_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__mux2_1
X_3305_ _1136_ net52 _1473_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__mux2_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3236_ _1546_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__clkbuf_2
X_3167_ po_0.regf_0.rf\[2\]\[0\] _0735_ _1398_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__mux2_1
X_3098_ _1361_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__clkbuf_1
X_2118_ net44 VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__clkbuf_2
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2049_ _0560_ _0562_ _0443_ _0565_ VGND VGND VPWR VPWR po_0.regf_0._3_\[11\] sky130_fd_sc_hd__o22a_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3021_ _0737_ _0906_ _1061_ _0742_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__and4b_4
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2805_ _1118_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__clkbuf_1
X_2736_ po_0.regf_0.w_addr\[2\] _0927_ po_0.regf_0.w_wr _0928_ VGND VGND VPWR VPWR
+ _1081_ sky130_fd_sc_hd__and4b_4
X_2667_ _0736_ po_0.regf_0.rf\[13\]\[0\] _1043_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__mux2_1
X_2598_ po_0.regf_0.rf\[15\]\[1\] _0953_ _1004_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__mux2_1
XFILLER_86_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3219_ po_0.regf_0.rf\[8\]\[8\] _0835_ _1424_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__mux2_1
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3570_ net105 _0222_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_2521_ _0958_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
X_2452_ po_0.regf_0.rf\[6\]\[7\] _0821_ _0916_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__mux2_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2383_ net3 _0823_ _0858_ _0860_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__a22o_2
X_3004_ net65 net94 VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__xnor2_1
Xinput3 D_R_data[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2719_ _1072_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
X_3699_ net184 uc_0.bc_0._70_\[1\] VGND VGND VPWR VPWR uc_0.bc_0._05_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1952_ _0464_ _0469_ _0471_ _0478_ VGND VGND VPWR VPWR po_0.regf_0._3_\[1\] sky130_fd_sc_hd__o22a_1
X_1883_ _1566_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__and2b_1
X_3622_ net128 _0270_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3553_ net177 _0205_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfxtp_1
X_2504_ _0896_ po_0.regf_0.rf\[7\]\[14\] _0930_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__mux2_1
X_3484_ net120 _0136_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_2435_ _0737_ _0906_ _0907_ _0742_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__and4b_4
XFILLER_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2366_ _0845_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
X_2297_ _0623_ _0760_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__a21o_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _0702_ _0701_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__o21a_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2151_ _0640_ _0641_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__nor2_1
XFILLER_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2082_ uc_0.bc_0._70_\[2\] uc_0.bc_0._70_\[3\] VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__or2_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2984_ _1241_ _1279_ _1281_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__a21o_1
X_1935_ _0449_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__buf_2
X_1866_ _0398_ _0399_ _1570_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux2_1
X_3605_ net103 _0253_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_1797_ _1603_ _1615_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__and2b_1
X_3536_ net109 _0188_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3467_ net156 _0119_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2418_ _0773_ po_0.alu_0._11_\[14\] _0746_ _0707_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__a22o_1
X_3398_ net155 _0054_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2349_ _0658_ _0659_ _0828_ _0829_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1720_ uc_0._21_\[13\] uc_0._21_\[15\] uc_0._21_\[14\] VGND VGND VPWR VPWR _1547_
+ sky130_fd_sc_hd__or3b_1
X_1651_ _1489_ _1493_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__or2_1
X_3321_ _1356_ _0593_ _1435_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__or3_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _1445_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__clkbuf_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _1407_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__clkbuf_1
X_2203_ _0695_ _0673_ _0679_ _0685_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__or4_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2134_ _0629_ _0630_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__nand2_2
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2065_ _0450_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__and2b_1
XFILLER_81_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2967_ net97 VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__clkbuf_2
X_1918_ po_0.regf_0.rf\[12\]\[0\] po_0.regf_0.rf\[13\]\[0\] po_0.regf_0.rf\[14\]\[0\]
+ po_0.regf_0.rf\[15\]\[0\] _0444_ _0445_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__mux4_1
X_2898_ _1205_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__clkbuf_1
X_1849_ _0384_ _1581_ _1583_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__a21o_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3519_ net122 _0171_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2821_ net99 VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__clkbuf_2
X_2752_ _1090_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
X_1703_ uc_0.bc_0._05_\[0\] uc_0.bc_0._05_\[3\] _1531_ VGND VGND VPWR VPWR _1532_
+ sky130_fd_sc_hd__and3_1
X_2683_ _1052_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ _1474_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _1551_ _0729_ _1550_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__a21bo_1
XFILLER_86_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _1397_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3097_ po_0.regf_0.rf\[3\]\[0\] _0735_ _1360_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__mux2_1
X_2117_ net44 _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__and2_1
XFILLER_54_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2048_ _0563_ _0564_ _0499_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__mux2_1
XFILLER_42_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3020_ net67 _1135_ _1313_ _1317_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2804_ po_0.regf_0.rf\[10\]\[15\] _0982_ _1100_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__mux2_1
X_2735_ _1080_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
X_2666_ _1042_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__buf_2
X_2597_ _1005_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3218_ _1426_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3149_ _0836_ po_0.regf_0.rf\[0\]\[8\] _1386_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__mux2_1
XFILLER_42_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2520_ po_0.regf_0.rf\[9\]\[3\] _0957_ _0951_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__mux2_1
X_2451_ _0917_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2382_ _1491_ po_0.alu_0._11_\[11\] _0859_ net85 _0752_ VGND VGND VPWR VPWR _0860_
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3003_ _1300_ _1301_ _1248_ _1147_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__a31oi_1
Xinput4 D_R_data[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2718_ po_0.regf_0.rf\[12\]\[7\] _0966_ _1070_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__mux2_1
X_3698_ net184 uc_0.bc_0._70_\[0\] VGND VGND VPWR VPWR uc_0.bc_0._05_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2649_ _0836_ po_0.regf_0.rf\[14\]\[8\] _1031_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__mux2_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1951_ _0474_ _0477_ _0450_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__mux2_1
X_1882_ po_0.regf_0.rf\[0\]\[12\] po_0.regf_0.rf\[1\]\[12\] po_0.regf_0.rf\[2\]\[12\]
+ po_0.regf_0.rf\[3\]\[12\] _1572_ _1574_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux4_1
X_3621_ net103 _0269_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3552_ net176 _0204_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfxtp_1
X_2503_ _0946_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
X_3483_ net156 _0135_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_2434_ _0740_ _0739_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__and2b_1
X_2365_ po_0.regf_0.rf\[5\]\[9\] _0844_ _0810_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__mux2_1
X_2296_ _1524_ po_0._1_\[2\] po_0._1_\[3\] net44 VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__a22o_1
XFILLER_24_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2150_ _0641_ _0640_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__or2b_1
X_2081_ _1533_ _1534_ _1537_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__and3_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2983_ _1241_ _1279_ _1281_ _1282_ _1283_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__a2111o_1
XFILLER_61_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1934_ po_0.regf_0.rf\[12\]\[1\] po_0.regf_0.rf\[13\]\[1\] po_0.regf_0.rf\[14\]\[1\]
+ po_0.regf_0.rf\[15\]\[1\] _0458_ _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__mux4_1
X_1865_ po_0.regf_0.rf\[4\]\[10\] po_0.regf_0.rf\[5\]\[10\] po_0.regf_0.rf\[6\]\[10\]
+ po_0.regf_0.rf\[7\]\[10\] _0366_ _0367_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__mux4_1
X_3604_ net118 _0252_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_1796_ po_0.regf_0.rf\[8\]\[3\] po_0.regf_0.rf\[9\]\[3\] po_0.regf_0.rf\[10\]\[3\]
+ po_0.regf_0.rf\[11\]\[3\] _1597_ _1598_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__mux4_1
X_3535_ net122 _0187_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_3466_ net162 _0118_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2417_ _0890_ _0891_ _0888_ _0887_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__o211ai_1
X_3397_ net134 _0053_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2348_ _0640_ _0641_ _0654_ _0655_ _0803_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__o2111ai_2
X_2279_ po_0.muxf_0.rf_w_data\[2\] _0724_ _0727_ net9 VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__a22o_1
XFILLER_25_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1650_ _1495_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__clkbuf_1
X_3320_ uc_0.bc_0._70_\[2\] _0593_ _1482_ net77 VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o2bb2a_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ po_0.regf_0.rq_addr\[1\] _1555_ _1442_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__mux2_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3182_ po_0.regf_0.rf\[2\]\[7\] _0820_ _1405_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__mux2_1
X_2202_ _0666_ _0667_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__nor2_1
XFILLER_78_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2133_ _0631_ _0632_ _0633_ _0622_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__a2bb2oi_2
X_2064_ po_0.regf_0.rf\[8\]\[14\] po_0.regf_0.rf\[9\]\[14\] po_0.regf_0.rf\[10\]\[14\]
+ po_0.regf_0.rf\[11\]\[14\] _0472_ _0473_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__mux4_1
XFILLER_19_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2966_ _1268_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__clkbuf_1
X_1917_ _0440_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__clkbuf_4
X_2897_ _1204_ _1193_ _1131_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__mux2_1
X_1848_ po_0.regf_0.rf\[12\]\[8\] po_0.regf_0.rf\[13\]\[8\] po_0.regf_0.rf\[14\]\[8\]
+ po_0.regf_0.rf\[15\]\[8\] _1578_ _1579_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__mux4_1
X_1779_ _1572_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__clkbuf_4
X_3518_ net164 _0170_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_3449_ net137 _0101_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2820_ _1119_ _1121_ _1125_ _1132_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__a31o_1
X_2751_ po_0.regf_0.rf\[11\]\[6\] _0963_ _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__mux2_1
X_1702_ uc_0.bc_0._05_\[1\] uc_0.bc_0._05_\[2\] VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__nor2_1
X_2682_ _0821_ po_0.regf_0.rf\[13\]\[7\] _1050_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__mux2_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3303_ _1124_ net51 _1473_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__mux2_1
X_3234_ _1434_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__clkbuf_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _0742_ po_0.regf_0.w_addr\[3\] _0906_ _0907_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__and4bb_4
XFILLER_39_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3096_ _1359_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2116_ po_0._1_\[3\] VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__clkbuf_2
XFILLER_54_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2047_ po_0.regf_0.rf\[4\]\[11\] po_0.regf_0.rf\[5\]\[11\] po_0.regf_0.rf\[6\]\[11\]
+ po_0.regf_0.rf\[7\]\[11\] _0451_ _0452_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__mux4_1
XFILLER_54_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2949_ net75 net98 VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__nor2_1
XFILLER_77_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2803_ _1117_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_1
X_2734_ po_0.regf_0.rf\[12\]\[15\] _0982_ _1062_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__mux2_1
X_2665_ _0739_ _1022_ _0740_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__or3b_4
X_2596_ po_0.regf_0.rf\[15\]\[0\] _0949_ _1004_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__mux2_1
XFILLER_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3217_ po_0.regf_0.rf\[8\]\[7\] _0820_ _1424_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__mux2_1
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3148_ _1388_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3079_ uc_0._21_\[10\] net18 _1344_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__mux2_1
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2450_ po_0.regf_0.rf\[6\]\[6\] _0809_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__mux2_1
X_2381_ po_0.alu_0.s1 _1487_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__or2_1
X_3002_ _1278_ _1290_ net94 _1274_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__nand4_1
Xinput5 D_R_data[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2717_ _1071_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
X_3697_ net183 _0345_ VGND VGND VPWR VPWR uc_0._01_ sky130_fd_sc_hd__dfxtp_1
X_2648_ _1033_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
X_2579_ _0995_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1950_ po_0.regf_0.rf\[4\]\[1\] po_0.regf_0.rf\[5\]\[1\] po_0.regf_0.rf\[6\]\[1\]
+ po_0.regf_0.rf\[7\]\[1\] _0475_ _0476_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__mux4_1
X_1881_ po_0.regf_0.rf\[4\]\[12\] po_0.regf_0.rf\[5\]\[12\] po_0.regf_0.rf\[6\]\[12\]
+ po_0.regf_0.rf\[7\]\[12\] _1578_ _1579_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux4_1
X_3620_ net116 _0268_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_3551_ net176 _0203_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfxtp_1
X_2502_ _0883_ po_0.regf_0.rf\[7\]\[13\] _0930_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__mux2_1
X_3482_ net156 _0134_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2433_ po_0.regf_0.w_wr VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__clkbuf_2
X_2364_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2295_ _0631_ _0632_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__nor2_1
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_10 net191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2080_ _0587_ _0589_ _0443_ _0592_ VGND VGND VPWR VPWR po_0.regf_0._3_\[15\] sky130_fd_sc_hd__o22a_1
XFILLER_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2982_ net97 net96 VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__and2_1
XFILLER_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1933_ _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__buf_2
XFILLER_61_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput30 I_data[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
X_1864_ po_0.regf_0.rf\[0\]\[10\] po_0.regf_0.rf\[1\]\[10\] po_0.regf_0.rf\[2\]\[10\]
+ po_0.regf_0.rf\[3\]\[10\] _0366_ _0367_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__mux4_1
X_3603_ net158 _0251_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_1795_ _1606_ _1608_ _1596_ _1614_ VGND VGND VPWR VPWR po_0.regf_0._5_\[2\] sky130_fd_sc_hd__o22a_1
X_3534_ net165 _0186_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_3465_ net137 _0117_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2416_ _0683_ _0865_ _0866_ _0868_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__o22a_1
X_3396_ net134 _0052_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2347_ _0658_ _0659_ _0647_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2278_ _0758_ _0761_ _0762_ _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__a31o_1
XFILLER_25_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _1444_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__clkbuf_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _0687_ _0685_ _0686_ po_0._1_\[11\] _0693_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__o32ai_2
X_3181_ _1406_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2132_ _0618_ _0620_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__or2b_1
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2063_ _0577_ VGND VGND VPWR VPWR po_0.regf_0._3_\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2965_ _1267_ _1263_ _1131_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__mux2_1
X_1916_ _0439_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__clkbuf_4
X_2896_ _1199_ _1120_ _1200_ _1203_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__a31o_1
X_1847_ _1591_ _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__and2b_1
X_1778_ po_0.regf_0.rf\[0\]\[1\] po_0.regf_0.rf\[1\]\[1\] po_0.regf_0.rf\[2\]\[1\]
+ po_0.regf_0.rf\[3\]\[1\] _1597_ _1598_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__mux4_1
X_3517_ net124 _0169_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_3448_ net140 _0100_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ net129 _0035_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2750_ _1081_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__buf_2
X_2681_ _1051_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
X_1701_ _1523_ _1529_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__nor2_1
X_3302_ uc_0.bc_0._70_\[2\] _0593_ _1435_ _1438_ net59 VGND VGND VPWR VPWR _0333_
+ sky130_fd_sc_hd__a32o_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3233_ po_0.regf_0.rf\[8\]\[15\] _0903_ _1416_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__mux2_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3164_ _1396_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__clkbuf_1
X_3095_ _0742_ po_0.regf_0.w_addr\[3\] _0906_ _0928_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__and4bb_4
X_2115_ _0617_ VGND VGND VPWR VPWR po_0.alu_0._10_\[2\] sky130_fd_sc_hd__clkbuf_1
X_2046_ po_0.regf_0.rf\[0\]\[11\] po_0.regf_0.rf\[1\]\[11\] po_0.regf_0.rf\[2\]\[11\]
+ po_0.regf_0.rf\[3\]\[11\] _0524_ _0525_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__mux4_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2948_ _1235_ _1221_ _1243_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__o21a_1
X_2879_ _1186_ _1187_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__nor2_2
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2802_ po_0.regf_0.rf\[10\]\[14\] _0980_ _1100_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__mux2_1
X_2733_ _1079_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
X_2664_ _1041_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
X_2595_ _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__buf_2
XFILLER_86_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3216_ _1425_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__clkbuf_1
X_3147_ _0821_ po_0.regf_0.rf\[0\]\[7\] _1386_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__mux2_1
XFILLER_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3078_ _1349_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__clkbuf_1
X_2029_ po_0.regf_0.rf\[0\]\[9\] po_0.regf_0.rf\[1\]\[9\] po_0.regf_0.rf\[2\]\[9\]
+ po_0.regf_0.rf\[3\]\[9\] _0466_ _0467_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__mux4_1
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2380_ _0685_ _0856_ _0857_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3001_ _1278_ _1290_ _1274_ net94 VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__a31o_1
Xinput6 D_R_data[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3696_ net183 _0344_ VGND VGND VPWR VPWR uc_0._02_ sky130_fd_sc_hd__dfxtp_1
X_2716_ po_0.regf_0.rf\[12\]\[6\] _0963_ _1070_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__mux2_1
X_2647_ _0821_ po_0.regf_0.rf\[14\]\[7\] _1031_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__mux2_1
X_2578_ po_0.regf_0.rf\[1\]\[8\] _0968_ _0992_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__mux2_1
XFILLER_55_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _0411_ _1581_ _1583_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__a21o_1
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3550_ net173 _0202_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfxtp_4
X_2501_ _0945_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
X_3481_ net138 _0133_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2432_ _0905_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2363_ _0841_ _0842_ _0752_ _0823_ net16 VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__a32o_2
X_2294_ _0779_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_11 net191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3679_ net180 _0327_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2981_ net97 net96 VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__nor2_1
X_1932_ _0001_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__clkbuf_2
X_1863_ _0395_ _0396_ _1570_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__mux2_1
Xinput20 I_data[12] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
X_3602_ net117 _0250_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xinput31 I_data[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
X_1794_ _1611_ _1612_ _1613_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__mux2_1
X_3533_ net124 _0185_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_3464_ net139 _0116_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2415_ _0689_ _0690_ _0700_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__or3b_1
X_3395_ net129 _0051_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2346_ _0826_ _0782_ _0626_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__nand3_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2277_ _0763_ po_0.alu_0._11_\[2\] _0747_ _1524_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__a22o_1
XFILLER_84_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ net85 VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__inv_2
X_3180_ po_0.regf_0.rf\[2\]\[6\] _0808_ _1405_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__mux2_1
X_2131_ _0629_ _0630_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__nor2_1
XFILLER_81_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2062_ _0573_ _0574_ _0575_ _0576_ _0438_ _0470_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__mux4_1
X_2964_ _1261_ _1120_ _1262_ _1266_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__a31o_1
X_1915_ _0003_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__buf_2
X_2895_ _1201_ _1202_ _1129_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__and3b_1
X_1846_ po_0.regf_0.rf\[0\]\[8\] po_0.regf_0.rf\[1\]\[8\] po_0.regf_0.rf\[2\]\[8\]
+ po_0.regf_0.rf\[3\]\[8\] _1592_ _1593_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux4_1
X_1777_ _1574_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__clkbuf_4
X_3516_ net162 _0168_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3447_ net143 _0099_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ net134 _0034_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2329_ _0811_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2680_ _0809_ po_0.regf_0.rf\[13\]\[6\] _1050_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__mux2_1
X_1700_ _1525_ _1527_ _1528_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__nand3_2
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3301_ uc_0.bc_0._70_\[0\] _1440_ _1438_ net60 VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__a22o_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _1433_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__clkbuf_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _0904_ po_0.regf_0.rf\[0\]\[15\] _1378_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__mux2_1
XFILLER_66_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2114_ _0613_ _0616_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__and2_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3094_ uc_0.bc_0._70_\[2\] uc_0.bc_0._70_\[3\] _1358_ _1156_ _1356_ VGND VGND VPWR
+ VPWR _0240_ sky130_fd_sc_hd__o32a_1
X_2045_ _0511_ _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__and2b_1
XFILLER_22_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2947_ _1248_ _1250_ _1147_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__a21o_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2878_ _1185_ _1167_ _1184_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__and3_1
X_1829_ _0005_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__buf_2
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2801_ _1116_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__clkbuf_1
X_2732_ po_0.regf_0.rf\[12\]\[14\] _0980_ _1062_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__mux2_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2663_ _0904_ po_0.regf_0.rf\[14\]\[15\] _1023_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__mux2_1
X_2594_ _0929_ _0927_ _0738_ _0928_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__and4_4
X_3215_ po_0.regf_0.rf\[8\]\[6\] _0808_ _1424_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__mux2_1
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3146_ _1387_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3077_ uc_0._21_\[9\] net32 _1344_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__mux2_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2028_ _0546_ _0487_ _0463_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__a21bo_1
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3000_ _1119_ _1156_ _1248_ _1290_ _1299_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__o41a_1
Xinput7 D_R_data[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3695_ net185 _0343_ VGND VGND VPWR VPWR uc_0._03_ sky130_fd_sc_hd__dfxtp_1
X_2715_ _1062_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__buf_2
X_2646_ _1032_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
X_2577_ _0994_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3129_ _1377_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3480_ net139 _0132_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2500_ _0874_ po_0.regf_0.rf\[7\]\[12\] _0930_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__mux2_1
X_2431_ po_0.regf_0.rf\[5\]\[15\] _0904_ _0743_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__mux2_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2362_ _0671_ _0763_ _1487_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__or3_1
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2293_ po_0.regf_0.rf\[5\]\[3\] _0778_ _0744_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__mux2_1
XFILLER_64_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 _0930_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3678_ net187 _0326_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[4\] sky130_fd_sc_hd__dfxtp_1
X_2629_ po_0.regf_0.w_addr\[2\] po_0.regf_0.w_addr\[3\] po_0.regf_0.w_wr VGND VGND
+ VPWR VPWR _1022_ sky130_fd_sc_hd__nand3_1
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2980_ net97 _1280_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__nor2_1
X_1931_ _0457_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__clkbuf_4
X_1862_ po_0.regf_0.rf\[12\]\[10\] po_0.regf_0.rf\[13\]\[10\] po_0.regf_0.rf\[14\]\[10\]
+ po_0.regf_0.rf\[15\]\[10\] _0361_ _0362_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux4_1
Xinput21 I_data[13] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput10 D_R_data[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
X_3601_ net119 _0249_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xinput32 I_data[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
X_1793_ _0006_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__clkbuf_4
X_3532_ net162 _0184_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_3463_ net133 _0115_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2414_ _0885_ _0887_ _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__a21o_1
XFILLER_69_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3394_ net134 _0050_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2345_ _0824_ _0825_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__nor2_1
XFILLER_69_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2276_ po_0.alu_0.s1 VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__clkbuf_2
XFILLER_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2130_ _0629_ _0630_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__and2_1
X_2061_ po_0.regf_0.rf\[12\]\[13\] po_0.regf_0.rf\[13\]\[13\] po_0.regf_0.rf\[14\]\[13\]
+ po_0.regf_0.rf\[15\]\[13\] _0439_ _0440_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__mux4_1
XFILLER_66_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2963_ _1264_ _1129_ _1265_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__and3b_1
X_1914_ _0438_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__or2b_1
X_2894_ _1160_ _1179_ _1175_ _1193_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__a31o_1
XFILLER_8_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1845_ _0380_ _1571_ _0007_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__a21o_1
X_1776_ _1572_ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__buf_4
X_3515_ net163 _0167_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3446_ net149 _0098_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ net129 _0033_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ po_0.regf_0.rf\[5\]\[6\] _0809_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__mux2_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2259_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__clkbuf_2
XFILLER_80_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3300_ _1471_ _1473_ _1460_ po_0.muxf_0.s1 _1436_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__o221a_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ po_0.regf_0.rf\[8\]\[14\] _0895_ _1416_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__mux2_1
X_3162_ _1395_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__clkbuf_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2113_ _0614_ _0615_ _0611_ _0612_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__a22o_1
XFILLER_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3093_ _1356_ _1357_ _1546_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__or3_2
X_2044_ po_0.regf_0.rf\[8\]\[11\] po_0.regf_0.rf\[9\]\[11\] po_0.regf_0.rf\[10\]\[11\]
+ po_0.regf_0.rf\[11\]\[11\] _0512_ _0513_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__mux4_1
XFILLER_62_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2946_ _1230_ _1249_ _1237_ _1247_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2877_ _1184_ _1185_ _1167_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__a21oi_2
X_1828_ _0004_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__clkbuf_4
X_1759_ _1566_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__buf_2
X_3429_ net131 _0081_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2800_ po_0.regf_0.rf\[10\]\[13\] _0978_ _1100_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__mux2_1
X_2731_ _1078_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2662_ _1040_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2593_ _1002_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
X_3214_ _1416_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__buf_2
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3145_ _0809_ po_0.regf_0.rf\[0\]\[6\] _1386_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__mux2_1
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3076_ _1348_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2027_ po_0.regf_0.rf\[12\]\[9\] po_0.regf_0.rf\[13\]\[9\] po_0.regf_0.rf\[14\]\[9\]
+ po_0.regf_0.rf\[15\]\[9\] _0479_ _0480_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__mux4_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2929_ _1234_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput8 D_R_data[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3694_ net184 _0342_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfxtp_1
X_2714_ _1069_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
X_2645_ _0809_ po_0.regf_0.rf\[14\]\[6\] _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__mux2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2576_ po_0.regf_0.rf\[1\]\[7\] _0966_ _0992_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__mux2_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3128_ po_0.regf_0.rf\[3\]\[15\] _0903_ _1359_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__mux2_1
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3059_ _1136_ net24 _1337_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__mux2_1
XFILLER_82_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2430_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2361_ _0838_ _0839_ _0762_ _0840_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__a31o_1
X_2292_ _0777_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_13 _1559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3677_ net180 _0325_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[3\] sky130_fd_sc_hd__dfxtp_1
X_2628_ _1021_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
X_2559_ _0929_ po_0.regf_0.w_addr\[3\] _0906_ _0741_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__and4bb_4
XFILLER_28_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1930_ _0000_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__clkbuf_2
X_1861_ po_0.regf_0.rf\[8\]\[10\] po_0.regf_0.rf\[9\]\[10\] po_0.regf_0.rf\[10\]\[10\]
+ po_0.regf_0.rf\[11\]\[10\] _0361_ _0362_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__mux4_1
Xinput22 I_data[14] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlymetal6s2s_1
X_3600_ net156 _0248_ VGND VGND VPWR VPWR po_0.regf_0.rf\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xinput11 D_R_data[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
Xinput33 clock VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
X_1792_ po_0.regf_0.rf\[4\]\[2\] po_0.regf_0.rf\[5\]\[2\] po_0.regf_0.rf\[6\]\[2\]
+ po_0.regf_0.rf\[7\]\[2\] _1600_ _1601_ VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__mux4_1
X_3531_ net163 _0183_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3462_ net139 _0114_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3393_ net129 _0049_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2413_ _0708_ _0709_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__nand2_1
X_2344_ _0635_ _0636_ _0643_ _0642_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__nand4_1
XFILLER_69_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2275_ _0748_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__buf_2
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2060_ po_0.regf_0.rf\[8\]\[13\] po_0.regf_0.rf\[9\]\[13\] po_0.regf_0.rf\[10\]\[13\]
+ po_0.regf_0.rf\[11\]\[13\] _0439_ _0440_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__mux4_1
XFILLER_66_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2962_ _1235_ _1247_ _1230_ _1263_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__a31o_1
X_1913_ po_0.regf_0.rf\[8\]\[0\] po_0.regf_0.rf\[9\]\[0\] po_0.regf_0.rf\[10\]\[0\]
+ po_0.regf_0.rf\[11\]\[0\] _0439_ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__mux4_1
X_2893_ _1160_ _1179_ _1193_ _1175_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__and4_1
X_1844_ po_0.regf_0.rf\[4\]\[8\] po_0.regf_0.rf\[5\]\[8\] po_0.regf_0.rf\[6\]\[8\]
+ po_0.regf_0.rf\[7\]\[8\] _0352_ _0353_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__mux4_1
X_1775_ _1568_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__buf_2
X_3514_ net166 _0166_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3445_ net148 _0097_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ net127 _0032_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _0743_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__buf_2
XFILLER_57_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2258_ po_0.alu_0.s1 _1487_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__nor2_2
XFILLER_72_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2189_ net85 po_0._1_\[11\] VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__nor2_2
XFILLER_65_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _1432_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__clkbuf_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3161_ _0896_ po_0.regf_0.rf\[0\]\[14\] _1378_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__mux2_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2112_ po_0._1_\[2\] net43 VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__or2b_1
X_3092_ _1533_ _1534_ _1537_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__nand3_1
X_2043_ _0559_ _0530_ _0493_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__a21bo_1
XFILLER_54_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2945_ net75 net98 VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__and2_1
X_2876_ uc_0._21_\[4\] net71 VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__or2_1
X_1827_ _0363_ _0364_ _1570_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux2_1
X_1758_ po_0.regf_0.rf\[12\]\[0\] po_0.regf_0.rf\[13\]\[0\] po_0.regf_0.rf\[14\]\[0\]
+ po_0.regf_0.rf\[15\]\[0\] _1578_ _1579_ VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__mux4_1
X_1689_ uc_0.bc_0._05_\[2\] uc_0.bc_0._05_\[3\] VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__nor2_1
X_3428_ net143 _0080_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3359_ po_0.regf_0._5_\[15\] net91 VGND VGND VPWR VPWR po_0._1_\[15\] sky130_fd_sc_hd__dlxtp_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2730_ po_0.regf_0.rf\[12\]\[13\] _0978_ _1062_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__mux2_1
X_2661_ _0896_ po_0.regf_0.rf\[14\]\[14\] _1023_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__mux2_1
X_2592_ po_0.regf_0.rf\[1\]\[15\] _0982_ _0984_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__mux2_1
X_3213_ _1423_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3144_ _1378_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__buf_2
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3075_ uc_0._21_\[8\] net31 _1344_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__mux2_1
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2026_ _0450_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__and2b_1
XFILLER_24_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2928_ _1233_ _1222_ _1131_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__mux2_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2859_ _1167_ _1168_ _1150_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__o21ai_1
XFILLER_49_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 D_R_data[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2713_ po_0.regf_0.rf\[12\]\[5\] _0961_ _1063_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__mux2_1
X_3693_ net160 _0341_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfxtp_1
X_2644_ _1023_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__buf_2
X_2575_ _0993_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
X_3127_ _1376_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3058_ _1338_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2009_ _0449_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__buf_2
XFILLER_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2360_ _0773_ po_0.alu_0._11_\[9\] _0747_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__a21o_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2291_ po_0.muxf_0.rf_w_data\[3\] _0725_ _0728_ net10 _0776_ VGND VGND VPWR VPWR
+ _0777_ sky130_fd_sc_hd__a221o_2
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3676_ net187 _0324_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[2\] sky130_fd_sc_hd__dfxtp_1
X_2627_ po_0.regf_0.rf\[15\]\[15\] _0982_ _1003_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__mux2_1
X_2558_ _0983_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
X_2489_ _0939_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1860_ _0389_ _0391_ _1583_ _0394_ VGND VGND VPWR VPWR po_0.regf_0._5_\[9\] sky130_fd_sc_hd__o22a_1
Xinput12 D_R_data[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
X_1791_ po_0.regf_0.rf\[0\]\[2\] po_0.regf_0.rf\[1\]\[2\] po_0.regf_0.rf\[2\]\[2\]
+ po_0.regf_0.rf\[3\]\[2\] _1609_ _1610_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__mux4_1
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput23 I_data[15] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xinput34 reset VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
X_3530_ net166 _0182_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3461_ net131 _0113_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3392_ net127 _0048_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2412_ net83 po_0._1_\[13\] _0886_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2343_ _0654_ _0655_ _0815_ _0814_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__nand4_1
X_2274_ _0608_ _0609_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__or3b_1
XFILLER_84_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1989_ _0457_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__clkbuf_4
X_3659_ net178 _0307_ VGND VGND VPWR VPWR po_0.regf_0.rq_rd sky130_fd_sc_hd__dfxtp_1
XFILLER_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2961_ net98 _1263_ _1237_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__and3_2
X_1912_ _0001_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__buf_2
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2892_ _1196_ _1197_ _1183_ _1188_ _1186_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__a221o_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1843_ _0373_ _0375_ _0377_ _0379_ VGND VGND VPWR VPWR po_0.regf_0._5_\[7\] sky130_fd_sc_hd__o22a_1
X_1774_ _1591_ _1594_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__and2b_1
X_3513_ net151 _0165_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3444_ net132 _0096_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ po_0.regf_0._3_\[15\] net90 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlxtp_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _0808_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2257_ _0745_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2188_ _0679_ _0682_ VGND VGND VPWR VPWR po_0.alu_0._10_\[10\] sky130_fd_sc_hd__xor2_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3160_ _1394_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__clkbuf_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2111_ net43 po_0._1_\[2\] VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__or2b_1
X_3091_ _1517_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2042_ po_0.regf_0.rf\[12\]\[11\] po_0.regf_0.rf\[13\]\[11\] po_0.regf_0.rf\[14\]\[11\]
+ po_0.regf_0.rf\[15\]\[11\] _0488_ _0489_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__mux4_1
XFILLER_66_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2944_ _1157_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__buf_2
X_2875_ uc_0._21_\[4\] net71 VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__nand2_1
X_1826_ po_0.regf_0.rf\[12\]\[6\] po_0.regf_0.rf\[13\]\[6\] po_0.regf_0.rf\[14\]\[6\]
+ po_0.regf_0.rf\[15\]\[6\] _0361_ _0362_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__mux4_1
X_1757_ _1563_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__clkbuf_4
X_1688_ uc_0.bc_0._05_\[0\] uc_0.bc_0._05_\[1\] VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__nand2_1
X_3427_ net109 _0079_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3358_ po_0.regf_0._5_\[14\] net91 VGND VGND VPWR VPWR po_0._1_\[14\] sky130_fd_sc_hd__dlxtp_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2309_ _1491_ po_0.alu_0._11_\[5\] _0731_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__o21a_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ _1466_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2660_ _1039_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2591_ _1001_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3212_ po_0.regf_0.rf\[8\]\[5\] _0796_ _1417_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3143_ _1385_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3074_ _1347_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2025_ po_0.regf_0.rf\[8\]\[9\] po_0.regf_0.rf\[9\]\[9\] po_0.regf_0.rf\[10\]\[9\]
+ po_0.regf_0.rf\[11\]\[9\] _0472_ _0473_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__mux4_1
XFILLER_35_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2927_ _1128_ _1157_ _1228_ _1229_ _1232_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__o41ai_1
X_2858_ _1160_ uc_0._21_\[3\] VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__and2_1
X_1809_ po_0.regf_0.rf\[0\]\[4\] po_0.regf_0.rf\[1\]\[4\] po_0.regf_0.rf\[2\]\[4\]
+ po_0.regf_0.rf\[3\]\[4\] _1609_ _1610_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__mux4_1
X_2789_ _1110_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2712_ _1068_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
X_3692_ net160 _0340_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfxtp_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2643_ _1030_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
X_2574_ po_0.regf_0.rf\[1\]\[6\] _0963_ _0992_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__mux2_1
X_3126_ po_0.regf_0.rf\[3\]\[14\] _0895_ _1359_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__mux2_1
XFILLER_67_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3057_ _1124_ net17 _1337_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__mux2_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2008_ po_0.regf_0.rf\[12\]\[7\] po_0.regf_0.rf\[13\]\[7\] po_0.regf_0.rf\[14\]\[7\]
+ po_0.regf_0.rf\[15\]\[7\] _0458_ _0460_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__mux4_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2290_ _0620_ _0729_ _1488_ _0732_ _0775_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__o311a_1
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3675_ net187 _0323_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[1\] sky130_fd_sc_hd__dfxtp_1
X_2626_ _1020_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
X_2557_ po_0.regf_0.rf\[9\]\[15\] _0982_ _0950_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__mux2_1
X_2488_ _0809_ po_0.regf_0.rf\[7\]\[6\] _0938_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__mux2_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3109_ _1359_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__buf_2
XFILLER_43_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1790_ _1574_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__clkbuf_4
Xinput13 D_R_data[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput24 I_data[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3460_ net132 _0112_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3391_ net101 _0047_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_2411_ net83 po_0._1_\[13\] po_0._1_\[12\] net38 VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__o211a_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2342_ _0727_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__clkbuf_2
X_2273_ _1515_ _0606_ _0759_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1988_ _0449_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__buf_2
X_3658_ net180 _0306_ VGND VGND VPWR VPWR po_0.alu_0.s0 sky130_fd_sc_hd__dfxtp_1
X_2609_ po_0.regf_0.rf\[15\]\[6\] _0963_ _1011_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__mux2_1
X_3589_ net165 _0012_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout190 net191 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2960_ net62 VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1911_ _0000_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__buf_2
X_2891_ _1186_ _1189_ _1198_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__o21ai_1
X_1842_ _1585_ _0378_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__and2b_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1773_ po_0.regf_0.rf\[8\]\[1\] po_0.regf_0.rf\[9\]\[1\] po_0.regf_0.rf\[10\]\[1\]
+ po_0.regf_0.rf\[11\]\[1\] _1592_ _1593_ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__mux4_1
X_3512_ net150 _0164_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3443_ net107 _0095_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ po_0.regf_0._3_\[14\] net88 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlxtp_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ po_0.muxf_0.rf_w_data\[6\] _0725_ _0728_ net13 _0807_ VGND VGND VPWR VPWR
+ _0808_ sky130_fd_sc_hd__a221o_2
XFILLER_84_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2256_ po_0.regf_0.rf\[5\]\[0\] _0736_ _0744_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__mux2_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2187_ _0673_ _0675_ _0680_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__o211a_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2110_ _0608_ _0609_ _0611_ _0612_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__o211ai_1
X_3090_ _1355_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__clkbuf_1
X_2041_ _0553_ _0555_ _0471_ _0558_ VGND VGND VPWR VPWR po_0.regf_0._3_\[10\] sky130_fd_sc_hd__o22a_1
XFILLER_66_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2943_ net98 VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2874_ _1165_ _1162_ _1164_ _1170_ _1172_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__o32ai_4
X_1825_ po_0.regf_0.rf\[8\]\[6\] po_0.regf_0.rf\[9\]\[6\] po_0.regf_0.rf\[10\]\[6\]
+ po_0.regf_0.rf\[11\]\[6\] _0361_ _0362_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__mux4_1
X_1756_ _1561_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__buf_4
X_1687_ net34 VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__clkbuf_2
X_3426_ net112 _0078_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_3357_ po_0.regf_0._5_\[13\] net91 VGND VGND VPWR VPWR po_0._1_\[13\] sky130_fd_sc_hd__dlxtp_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _0643_ _0642_ _0783_ _0780_ _0631_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__a221o_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3288_ po_0.muxf_0.rf_w_data\[5\] _1555_ _1441_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__mux2_1
X_2239_ _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__buf_2
XFILLER_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2590_ po_0.regf_0.rf\[1\]\[14\] _0980_ _0984_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__mux2_1
XFILLER_5_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3211_ _1422_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_1
X_3142_ _0797_ po_0.regf_0.rf\[0\]\[5\] _1379_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__mux2_1
XFILLER_39_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3073_ _1559_ net30 _1344_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__mux2_1
X_2024_ _0538_ _0540_ _0471_ _0543_ VGND VGND VPWR VPWR po_0.regf_0._3_\[8\] sky130_fd_sc_hd__o22a_1
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2926_ _1230_ _1231_ _1129_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__or3b_1
X_2857_ _1160_ _1163_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__nor2_1
X_1808_ _1591_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__and2b_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2788_ po_0.regf_0.rf\[10\]\[7\] _0966_ _1108_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__mux2_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1739_ _0004_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__clkbuf_4
X_3409_ net166 _0009_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__dfxtp_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2711_ po_0.regf_0.rf\[12\]\[4\] _0959_ _1063_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__mux2_1
XFILLER_71_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3691_ net174 _0339_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfxtp_1
X_2642_ _0797_ po_0.regf_0.rf\[14\]\[5\] _1024_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__mux2_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2573_ _0984_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__buf_2
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3125_ _1375_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3056_ uc_0._03_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__buf_2
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2007_ _0521_ _0523_ _0471_ _0528_ VGND VGND VPWR VPWR po_0.regf_0._3_\[6\] sky130_fd_sc_hd__o22a_1
XFILLER_23_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2909_ _1186_ _1215_ _1197_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__o21a_1
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3674_ net180 _0322_ VGND VGND VPWR VPWR po_0.muxf_0.rf_w_data\[0\] sky130_fd_sc_hd__dfxtp_1
X_2625_ po_0.regf_0.rf\[15\]\[14\] _0980_ _1003_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__mux2_1
X_2556_ _0903_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__clkbuf_2
X_2487_ _0930_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__buf_2
X_3108_ _1366_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3039_ _1328_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput14 D_R_data[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
Xinput25 I_data[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
X_2410_ _0869_ _0700_ _0691_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__nand3_1
X_3390_ net105 _0046_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_2341_ _0822_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
X_2272_ net87 po_0._1_\[1\] VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__nand2_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1987_ _0509_ _0462_ _0470_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__a21o_1
X_3657_ net179 _0305_ VGND VGND VPWR VPWR po_0.alu_0.s1 sky130_fd_sc_hd__dfxtp_2
X_3588_ net181 _0240_ VGND VGND VPWR VPWR uc_0._00_ sky130_fd_sc_hd__dfxtp_1
X_2608_ _1003_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__buf_2
X_2539_ po_0.regf_0.rf\[9\]\[9\] _0970_ _0964_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__mux2_1
XFILLER_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout191 net33 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout180 net186 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1910_ _0002_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__buf_2
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2890_ _1196_ _1197_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__and2_1
X_1841_ po_0.regf_0.rf\[8\]\[7\] po_0.regf_0.rf\[9\]\[7\] po_0.regf_0.rf\[10\]\[7\]
+ po_0.regf_0.rf\[11\]\[7\] _1573_ _1575_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__mux4_1
XFILLER_30_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1772_ _1574_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__clkbuf_4
X_3511_ net146 _0163_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3442_ net103 _0094_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ po_0.regf_0._3_\[13\] net90 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlxtp_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _0799_ _0806_ _0752_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__o21a_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__buf_2
X_2186_ _0666_ _0667_ _0670_ _0674_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__o211ai_1
XFILLER_53_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3709_ po_0.alu_0._10_\[6\] _1630_ VGND VGND VPWR VPWR po_0.alu_0._11_\[6\] sky130_fd_sc_hd__ebufn_1
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2040_ _0556_ _0557_ _0499_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__mux2_1
XFILLER_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2942_ _1246_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2873_ _1180_ _1127_ _1181_ _1147_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__a31o_1
X_1824_ _0005_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__buf_2
X_1755_ _1571_ _1576_ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__and2b_1
X_1686_ _1516_ VGND VGND VPWR VPWR po_0.alu_0._10_\[0\] sky130_fd_sc_hd__clkbuf_1
X_3425_ net127 _0077_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3356_ po_0.regf_0._5_\[12\] net91 VGND VGND VPWR VPWR po_0._1_\[12\] sky130_fd_sc_hd__dlxtp_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2307_ _0635_ _0784_ _0651_ _0650_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__a211o_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _1465_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__clkbuf_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2238_ _0726_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__clkbuf_2
X_2169_ net86 po_0._1_\[8\] VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__and2_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3210_ po_0.regf_0.rf\[8\]\[4\] _0788_ _1417_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__mux2_1
X_3141_ _1384_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3072_ _1346_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__clkbuf_1
X_2023_ _0541_ _0542_ _0499_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__mux2_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2925_ _1206_ _1201_ _1222_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__a21oi_1
X_2856_ _1162_ _1164_ _1165_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__o21ai_1
X_1807_ po_0.regf_0.rf\[8\]\[4\] po_0.regf_0.rf\[9\]\[4\] po_0.regf_0.rf\[10\]\[4\]
+ po_0.regf_0.rf\[11\]\[4\] _1592_ _1593_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__mux4_1
X_2787_ _1109_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
X_1738_ _1560_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
X_1669_ _1506_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__clkbuf_1
X_3408_ net178 _0008_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__dfxtp_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ net118 _0027_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2710_ _1067_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3690_ net187 _0338_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dfxtp_1
X_2641_ _1029_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
X_2572_ _0991_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3124_ po_0.regf_0.rf\[3\]\[13\] _0882_ _1359_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__mux2_1
XFILLER_82_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3055_ _1336_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2006_ _0526_ _0527_ _0499_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__mux2_1
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2908_ _1549_ net71 _1195_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__o21a_1
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2839_ net69 uc_0._21_\[2\] VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__or2_1
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3673_ net125 _0321_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[3\] sky130_fd_sc_hd__dfxtp_1
X_2624_ _1019_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
X_2555_ _0981_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
X_2486_ _0937_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3107_ po_0.regf_0.rf\[3\]\[5\] _0796_ _1360_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__mux2_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3038_ po_0.regf_0.rf\[4\]\[7\] _0820_ _1326_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__mux2_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput26 I_data[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput15 D_R_data[8] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2340_ po_0.regf_0.rf\[5\]\[7\] _0821_ _0810_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__mux2_1
X_2271_ po_0._1_\[0\] _1513_ _0607_ _0623_ _0605_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__a311o_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1986_ po_0.regf_0.rf\[4\]\[5\] po_0.regf_0.rf\[5\]\[5\] po_0.regf_0.rf\[6\]\[5\]
+ po_0.regf_0.rf\[7\]\[5\] _0479_ _0480_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__mux4_1
X_3656_ net110 _0304_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_2607_ _1010_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
X_3587_ net179 _0239_ VGND VGND VPWR VPWR uc_0._21_\[15\] sky130_fd_sc_hd__dfxtp_1
X_2538_ _0843_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__clkbuf_2
X_2469_ _0926_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout181 net183 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout170 net190 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1840_ _0376_ _1581_ _1583_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__a21o_1
XFILLER_42_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1771_ _1572_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__clkbuf_4
X_3510_ net150 _0162_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3441_ net113 _0093_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ po_0.regf_0._3_\[12\] net90 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlxtp_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _0802_ _0748_ _0805_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__and3b_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _0737_ _0738_ _0741_ _0742_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__and4b_4
X_2185_ po_0._1_\[9\] _0671_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__or2b_1
XFILLER_18_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1969_ _0492_ _0462_ _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__a21bo_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3708_ po_0.alu_0._10_\[5\] _1629_ VGND VGND VPWR VPWR po_0.alu_0._11_\[5\] sky130_fd_sc_hd__ebufn_1
X_3639_ net104 _0287_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2941_ _1245_ _1235_ _1131_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__mux2_1
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2872_ _1122_ _1133_ _1144_ _1161_ _1179_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__a41o_1
XFILLER_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1823_ _0004_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__clkbuf_4
X_1754_ po_0.regf_0.rf\[0\]\[0\] po_0.regf_0.rf\[1\]\[0\] po_0.regf_0.rf\[2\]\[0\]
+ po_0.regf_0.rf\[3\]\[0\] _1573_ _1575_ VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__mux4_1
X_3424_ net109 _0076_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_1685_ _1514_ _1515_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__and2_1
X_3355_ po_0.regf_0._5_\[11\] net91 VGND VGND VPWR VPWR po_0._1_\[11\] sky130_fd_sc_hd__dlxtp_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _0790_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ po_0.muxf_0.rf_w_data\[4\] _1549_ _1441_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__mux2_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ po_0.muxf_0.s1 po_0.muxf_0.s0 VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__and2b_1
XFILLER_26_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2168_ _0665_ VGND VGND VPWR VPWR po_0.alu_0._10_\[7\] sky130_fd_sc_hd__clkbuf_1
X_2099_ _1539_ _1535_ _1541_ _1542_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__a31o_1
XFILLER_53_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3140_ _0789_ po_0.regf_0.rf\[0\]\[4\] _1379_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__mux2_1
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3071_ _1557_ net29 _1344_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__mux2_1
X_2022_ po_0.regf_0.rf\[4\]\[8\] po_0.regf_0.rf\[5\]\[8\] po_0.regf_0.rf\[6\]\[8\]
+ po_0.regf_0.rf\[7\]\[8\] _0475_ _0476_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__mux4_1
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2924_ _1206_ _1222_ _1201_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__and3_1
X_2855_ net69 _1151_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__nor2_1
X_1806_ _1623_ _1567_ _1589_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__a21o_1
X_2786_ po_0.regf_0.rf\[10\]\[6\] _0963_ _1108_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__mux2_1
X_1737_ po_0.regf_0.rq_addr\[3\] _1559_ _1553_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__mux2_1
X_1668_ _1500_ _1502_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__or2_1
X_3407_ net100 _0063_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ net158 _0026_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3269_ _1454_ _0739_ _1443_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__mux2_1
XFILLER_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2640_ _0789_ po_0.regf_0.rf\[14\]\[4\] _1024_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__mux2_1
X_2571_ po_0.regf_0.rf\[1\]\[5\] _0961_ _0985_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__mux2_1
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3123_ _1374_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3054_ po_0.regf_0.rf\[4\]\[15\] _0903_ _1318_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__mux2_1
XFILLER_82_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2005_ po_0.regf_0.rf\[4\]\[6\] po_0.regf_0.rf\[5\]\[6\] po_0.regf_0.rf\[6\]\[6\]
+ po_0.regf_0.rf\[7\]\[6\] _0475_ _0476_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__mux4_1
XFILLER_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2907_ _1212_ _1213_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__nor2_1
X_2838_ net61 uc_0._21_\[0\] _1137_ _1138_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__o22a_1
X_2769_ po_0.regf_0.rf\[11\]\[15\] _0982_ _1081_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__mux2_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ net123 _0320_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2623_ po_0.regf_0.rf\[15\]\[13\] _0978_ _1003_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__mux2_1
X_2554_ po_0.regf_0.rf\[9\]\[14\] _0980_ _0950_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__mux2_1
X_2485_ _0797_ po_0.regf_0.rf\[7\]\[5\] _0931_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__mux2_1
X_3106_ _1365_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3037_ _1327_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput16 D_R_data[9] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 I_data[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2270_ _0757_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1985_ _0502_ _0504_ _0506_ _0508_ VGND VGND VPWR VPWR po_0.regf_0._3_\[4\] sky130_fd_sc_hd__o22a_1
X_3655_ net113 _0303_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_2606_ po_0.regf_0.rf\[15\]\[5\] _0961_ _1004_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__mux2_1
X_3586_ net171 _0238_ VGND VGND VPWR VPWR uc_0._21_\[14\] sky130_fd_sc_hd__dfxtp_1
X_2537_ _0969_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
X_2468_ po_0.regf_0.rf\[6\]\[15\] _0904_ _0908_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__mux2_1
X_2399_ _0875_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout182 net183 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout160 net161 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
Xfanout171 net173 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1770_ _1566_ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__clkbuf_2
X_3440_ net112 _0092_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3371_ po_0.regf_0._3_\[11\] net88 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlxtp_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2322_ _0654_ _0655_ _0804_ _0643_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__a22o_1
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2253_ po_0.regf_0.w_addr\[2\] VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2184_ _0677_ _0678_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__nand2_2
XFILLER_21_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1968_ _0003_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__buf_2
X_1899_ _0427_ _0428_ _0006_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__mux2_1
X_3707_ po_0.alu_0._10_\[4\] _1628_ VGND VGND VPWR VPWR po_0.alu_0._11_\[4\] sky130_fd_sc_hd__ebufn_1
X_3638_ net113 _0286_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3569_ net110 _0221_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2940_ _1236_ _1237_ _1243_ _1244_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2871_ _1161_ _1179_ _1175_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__nand3_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1822_ _0355_ _0357_ _1596_ _0360_ VGND VGND VPWR VPWR po_0.regf_0._5_\[5\] sky130_fd_sc_hd__o22a_1
X_1753_ _1574_ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__buf_2
X_1684_ po_0._1_\[0\] net35 VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__nand2_1
X_3423_ net123 _0075_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ po_0.regf_0._5_\[10\] net92 VGND VGND VPWR VPWR po_0._1_\[10\] sky130_fd_sc_hd__dlxtp_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ po_0.regf_0.rf\[5\]\[4\] _0789_ _0744_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__mux2_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _1464_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__clkbuf_1
X_2236_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__buf_2
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2167_ _0663_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__and2_1
X_2098_ _0602_ _0603_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__nor2_2
XFILLER_13_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3070_ _1345_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2021_ po_0.regf_0.rf\[0\]\[8\] po_0.regf_0.rf\[1\]\[8\] po_0.regf_0.rf\[2\]\[8\]
+ po_0.regf_0.rf\[3\]\[8\] _0524_ _0525_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__mux4_1
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2923_ _1227_ _1218_ _1224_ _1226_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__o211a_1
X_2854_ _1163_ _1160_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__and2b_1
X_1805_ po_0.regf_0.rf\[12\]\[4\] po_0.regf_0.rf\[13\]\[4\] po_0.regf_0.rf\[14\]\[4\]
+ po_0.regf_0.rf\[15\]\[4\] _1562_ _1564_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__mux4_1
X_2785_ _1100_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__buf_2
X_1736_ uc_0._21_\[7\] VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__buf_2
X_1667_ _1505_ VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__clkbuf_1
X_3406_ net105 _0062_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_3337_ net115 _0025_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ uc_0._21_\[9\] _1136_ _1442_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__mux2_1
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3199_ _1415_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2219_ po_0._1_\[13\] net83 VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__or2b_1
XFILLER_38_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2570_ _0990_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
X_3122_ po_0.regf_0.rf\[3\]\[12\] _0873_ _1359_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__mux2_1
XFILLER_82_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3053_ _1335_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2004_ po_0.regf_0.rf\[0\]\[6\] po_0.regf_0.rf\[1\]\[6\] po_0.regf_0.rf\[2\]\[6\]
+ po_0.regf_0.rf\[3\]\[6\] _0524_ _0525_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__mux4_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2906_ _1192_ _1210_ _1211_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__and3_1
X_2837_ _1145_ _1146_ _1127_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__a31o_1
X_2768_ _1098_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2699_ _1060_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
X_1719_ _1517_ _1546_ VGND VGND VPWR VPWR uc_0.bc_0._70_\[0\] sky130_fd_sc_hd__nor2_1
XFILLER_86_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3671_ net178 _0319_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[1\] sky130_fd_sc_hd__dfxtp_1
X_2622_ _1018_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2553_ _0895_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2484_ _0936_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3105_ po_0.regf_0.rf\[3\]\[4\] _0788_ _1360_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__mux2_1
XFILLER_28_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3036_ po_0.regf_0.rf\[4\]\[6\] _0808_ _1326_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__mux2_1
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput17 I_data[0] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 I_data[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1984_ _0487_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__and2b_1
X_3654_ net128 _0302_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_2605_ _1009_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
X_3585_ net184 _0237_ VGND VGND VPWR VPWR uc_0._21_\[13\] sky130_fd_sc_hd__dfxtp_1
X_2536_ po_0.regf_0.rf\[9\]\[8\] _0968_ _0964_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__mux2_1
X_2467_ _0925_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2398_ po_0.regf_0.rf\[5\]\[12\] _0874_ _0743_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__mux2_1
XFILLER_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3019_ _1315_ _1121_ _1316_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__nand3_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout183 net185 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout150 net151 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout161 net170 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout172 net173 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3370_ po_0.regf_0._3_\[10\] net88 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlxtp_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _0626_ _0782_ _0780_ _0803_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__a31o_1
XFILLER_69_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ _0739_ _0740_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__and2b_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2183_ net36 po_0._1_\[10\] VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__or2b_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1967_ po_0.regf_0.rf\[12\]\[3\] po_0.regf_0.rf\[13\]\[3\] po_0.regf_0.rf\[14\]\[3\]
+ po_0.regf_0.rf\[15\]\[3\] _0458_ _0460_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__mux4_1
X_3706_ po_0.alu_0._10_\[3\] _1627_ VGND VGND VPWR VPWR po_0.alu_0._11_\[3\] sky130_fd_sc_hd__ebufn_1
X_1898_ po_0.regf_0.rf\[4\]\[14\] po_0.regf_0.rf\[5\]\[14\] po_0.regf_0.rf\[6\]\[14\]
+ po_0.regf_0.rf\[7\]\[14\] _0366_ _0367_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__mux4_1
X_3637_ net103 _0285_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_3568_ net103 _0220_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_2519_ _0777_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__clkbuf_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3499_ net162 _0151_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2870_ net71 VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1821_ _0358_ _0359_ _1613_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__mux2_1
X_1752_ _0005_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__clkbuf_2
XFILLER_7_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1683_ po_0._1_\[0\] _1513_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__or2_1
X_3422_ net164 _0074_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ po_0.regf_0._5_\[9\] net92 VGND VGND VPWR VPWR po_0._1_\[9\] sky130_fd_sc_hd__dlxtp_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2304_ _0788_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__clkbuf_2
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ po_0.muxf_0.rf_w_data\[3\] _1163_ _1460_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__mux2_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ po_0.muxf_0.s0 po_0.muxf_0.s1 VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__and2b_1
X_2166_ _0653_ _0660_ _0661_ _0662_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__or4_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2097_ _1539_ _1535_ _1541_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2999_ _1294_ _1121_ _1295_ _1298_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__a31o_1
XFILLER_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2020_ _0511_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__and2b_1
XFILLER_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2922_ _1224_ _1226_ _1227_ _1218_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__a211oi_1
X_2853_ uc_0._21_\[3\] VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__clkbuf_2
X_1804_ _1616_ _1618_ _1620_ _1622_ VGND VGND VPWR VPWR po_0.regf_0._5_\[3\] sky130_fd_sc_hd__o22a_1
X_2784_ _1107_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
X_1735_ _1558_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
X_1666_ _1500_ _1502_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__or2_1
X_3405_ net109 _0061_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3336_ net118 _0024_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _1453_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3198_ po_0.regf_0.rf\[2\]\[15\] _0903_ _1397_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__mux2_1
X_2218_ net40 po_0._1_\[14\] VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__or2_1
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2149_ _1526_ po_0._1_\[6\] VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__nor2_1
XFILLER_14_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3121_ _1373_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__clkbuf_1
X_3052_ po_0.regf_0.rf\[4\]\[14\] _0895_ _1318_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__mux2_1
XFILLER_75_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2003_ _0459_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__buf_2
XFILLER_63_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2905_ _1210_ _1211_ _1192_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__a21oi_1
X_2836_ _1130_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__clkbuf_2
X_2767_ po_0.regf_0.rf\[11\]\[14\] _0980_ _1081_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__mux2_1
X_2698_ _0904_ po_0.regf_0.rf\[13\]\[15\] _1042_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__mux2_1
X_1718_ _1545_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__clkbuf_2
X_1649_ _1489_ _1493_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__or2_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _0594_ _1358_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__nor2_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3670_ net178 _0318_ VGND VGND VPWR VPWR po_0.regf_0.w_addr\[0\] sky130_fd_sc_hd__dfxtp_1
X_2621_ po_0.regf_0.rf\[15\]\[12\] _0976_ _1003_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__mux2_1
X_2552_ _0979_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2483_ _0789_ po_0.regf_0.rf\[7\]\[4\] _0931_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__mux2_1
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3104_ _1364_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3035_ _1318_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__buf_2
X_2819_ _1127_ _1131_ _1123_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__mux2_1
XFILLER_86_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput18 I_data[10] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 I_data[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1983_ po_0.regf_0.rf\[8\]\[4\] po_0.regf_0.rf\[9\]\[4\] po_0.regf_0.rf\[10\]\[4\]
+ po_0.regf_0.rf\[11\]\[4\] _0488_ _0489_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__mux4_1
X_3653_ net113 _0301_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_2604_ po_0.regf_0.rf\[15\]\[4\] _0959_ _1004_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__mux2_1
X_3584_ net171 _0236_ VGND VGND VPWR VPWR uc_0._21_\[12\] sky130_fd_sc_hd__dfxtp_1
X_2535_ _0835_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__clkbuf_2
X_2466_ po_0.regf_0.rf\[6\]\[14\] _0896_ _0908_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__mux2_1
X_2397_ _0873_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__clkbuf_2
XFILLER_56_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3018_ _1314_ _1308_ _1310_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__nand3_1
XFILLER_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout140 net141 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
Xfanout173 net177 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xfanout151 net152 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout162 net169 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
Xfanout184 net185 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ net45 _0630_ _0641_ net46 VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__a22o_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ po_0.regf_0.w_addr\[0\] VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__clkbuf_2
XFILLER_38_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2182_ po_0._1_\[10\] _1522_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__or2b_1
XFILLER_65_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1966_ _0482_ _0484_ _0486_ _0491_ VGND VGND VPWR VPWR po_0.regf_0._3_\[2\] sky130_fd_sc_hd__o22a_1
X_3705_ po_0.alu_0._10_\[2\] _1626_ VGND VGND VPWR VPWR po_0.alu_0._11_\[2\] sky130_fd_sc_hd__ebufn_1
X_1897_ po_0.regf_0.rf\[0\]\[14\] po_0.regf_0.rf\[1\]\[14\] po_0.regf_0.rf\[2\]\[14\]
+ po_0.regf_0.rf\[3\]\[14\] _0366_ _0367_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__mux4_1
X_3636_ net118 _0284_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_3567_ net118 _0219_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_2518_ _0956_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3498_ net165 _0150_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2449_ _0908_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__buf_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1820_ po_0.regf_0.rf\[4\]\[5\] po_0.regf_0.rf\[5\]\[5\] po_0.regf_0.rf\[6\]\[5\]
+ po_0.regf_0.rf\[7\]\[5\] _1600_ _1601_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux4_1
XFILLER_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1751_ _1572_ VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1682_ net35 VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__clkbuf_2
X_3421_ net124 _0073_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ po_0.regf_0._5_\[8\] net92 VGND VGND VPWR VPWR po_0._1_\[8\] sky130_fd_sc_hd__dlxtp_1
X_2303_ _0786_ _0753_ _0787_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__a21o_2
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _1463_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__clkbuf_1
X_2234_ _0721_ _0723_ VGND VGND VPWR VPWR po_0.alu_0._10_\[15\] sky130_fd_sc_hd__nand2_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2165_ _0660_ _0661_ _0662_ _0653_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__o22ai_2
XFILLER_80_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2096_ _1542_ _1541_ _1535_ _1539_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__and4b_1
XFILLER_65_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2998_ _1296_ _1297_ _1157_ _1130_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__a31o_1
XFILLER_21_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1949_ _0001_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__clkbuf_4
X_3619_ net158 _0267_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2921_ _1210_ _1211_ _1192_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__a21boi_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2852_ net70 uc_0._21_\[3\] VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__and2b_1
X_1803_ _1621_ _1581_ _1568_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__a21o_1
X_2783_ po_0.regf_0.rf\[10\]\[5\] _0961_ _1101_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__mux2_1
X_1734_ po_0.regf_0.rq_addr\[2\] _1557_ _1553_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__mux2_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3404_ net105 _0060_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_1665_ _1504_ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__clkbuf_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ net154 _0023_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _1452_ _0740_ _1443_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__mux2_1
X_2217_ _0707_ po_0._1_\[14\] VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__nand2_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ _1414_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2148_ _1526_ po_0._1_\[6\] VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__and2_1
X_2079_ _0590_ _0591_ _0438_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__mux2_1
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3120_ po_0.regf_0.rf\[3\]\[11\] _0861_ _1367_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__mux2_1
XFILLER_67_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3051_ _1334_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__clkbuf_1
X_2002_ _0457_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2904_ uc_0._21_\[6\] net73 VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__or2_1
X_2835_ _1123_ _1133_ _1144_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__nand3_1
XFILLER_31_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2766_ _1097_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
X_2697_ _1059_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
X_1717_ _1519_ _1531_ _1539_ _1540_ _1544_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__o2111a_1
X_1648_ _1494_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ _1481_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__clkbuf_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3249_ po_0.regf_0.rq_addr\[0\] _1549_ _1553_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__mux2_1
XFILLER_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2620_ _1017_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
X_2551_ po_0.regf_0.rf\[9\]\[13\] _0978_ _0950_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__mux2_1
X_2482_ _0935_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3103_ po_0.regf_0.rf\[3\]\[3\] _0777_ _1360_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__mux2_1
X_3034_ _1325_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2818_ _1130_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__buf_2
X_2749_ _1088_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 I_data[11] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1982_ _0505_ _0447_ _0463_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__a21bo_1
X_3652_ net123 _0300_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_2603_ _1008_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
X_3583_ net171 _0235_ VGND VGND VPWR VPWR uc_0._21_\[11\] sky130_fd_sc_hd__dfxtp_1
X_2534_ _0967_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
X_2465_ _0924_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
X_2396_ net4 _0823_ _0872_ _0753_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__a22o_2
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3017_ _1314_ _1308_ _1310_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__a21o_1
XFILLER_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout130 net133 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
Xfanout141 net142 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout152 net153 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
Xfanout163 net169 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
Xfanout174 net176 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout185 net186 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ po_0.regf_0.w_addr\[1\] VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__clkbuf_2
X_2181_ _0674_ _0676_ VGND VGND VPWR VPWR po_0.alu_0._10_\[9\] sky130_fd_sc_hd__xor2_1
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1965_ _0487_ _0490_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__and2b_1
X_3704_ po_0.alu_0._10_\[1\] _1625_ VGND VGND VPWR VPWR po_0.alu_0._11_\[1\] sky130_fd_sc_hd__ebufn_1
X_1896_ _0424_ _0425_ _1570_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
X_3635_ net161 _0283_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_3566_ net158 _0218_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_3497_ net148 _0149_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2517_ po_0.regf_0.rf\[9\]\[2\] _0955_ _0951_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__mux2_1
X_2448_ _0915_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
X_2379_ _0685_ _0856_ _0731_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1750_ _0004_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__clkbuf_2
XFILLER_11_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1681_ _1512_ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__clkbuf_1
X_3420_ net122 _0072_ VGND VGND VPWR VPWR po_0.regf_0.rf\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_3351_ po_0.regf_0._5_\[7\] net92 VGND VGND VPWR VPWR po_0._1_\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2302_ po_0.muxf_0.rf_w_data\[4\] _0724_ _0727_ net11 VGND VGND VPWR VPWR _0787_
+ sky130_fd_sc_hd__a22o_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ po_0.muxf_0.rf_w_data\[2\] _1151_ _1460_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__mux2_1
XFILLER_85_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2233_ _0714_ _0715_ _0722_ _0712_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__o22ai_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2164_ po_0._1_\[6\] _1526_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__and2b_1
XFILLER_80_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2095_ _1542_ _0601_ _1536_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__a21o_1
XFILLER_65_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2997_ _1269_ _1278_ _1290_ _1264_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__nand4_1
X_1948_ _0000_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__buf_4
X_1879_ po_0.regf_0.rf\[12\]\[12\] po_0.regf_0.rf\[13\]\[12\] po_0.regf_0.rf\[14\]\[12\]
+ po_0.regf_0.rf\[15\]\[12\] _1578_ _1579_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux4_1
X_3618_ net116 _0266_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_3549_ net173 _0201_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfxtp_1
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2920_ _1557_ net73 _1225_ _1223_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__a2bb2o_1
X_2851_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1802_ po_0.regf_0.rf\[4\]\[3\] po_0.regf_0.rf\[5\]\[3\] po_0.regf_0.rf\[6\]\[3\]
+ po_0.regf_0.rf\[7\]\[3\] _1578_ _1579_ VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__mux4_1
X_2782_ _1106_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
X_1733_ uc_0._21_\[6\] VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__clkbuf_2
XFILLER_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3403_ net115 _0059_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_1664_ _1500_ _1502_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__or2_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ net154 _0022_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ uc_0._21_\[8\] _1124_ _1442_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__mux2_1
XFILLER_85_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2216_ net40 VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ po_0.regf_0.rf\[2\]\[14\] _0895_ _1397_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__mux2_1
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2147_ _0646_ VGND VGND VPWR VPWR po_0.alu_0._10_\[5\] sky130_fd_sc_hd__clkbuf_1
X_2078_ po_0.regf_0.rf\[4\]\[15\] po_0.regf_0.rf\[5\]\[15\] po_0.regf_0.rf\[6\]\[15\]
+ po_0.regf_0.rf\[7\]\[15\] _0451_ _0452_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__mux4_1
XFILLER_26_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3050_ po_0.regf_0.rf\[4\]\[13\] _0882_ _1318_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__mux2_1
X_2001_ _0511_ _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__and2b_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2903_ uc_0._21_\[6\] net73 VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__nand2_1
X_2834_ _1123_ _1133_ _1144_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__a21o_1
X_2765_ po_0.regf_0.rf\[11\]\[13\] _0978_ _1081_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__mux2_1
X_2696_ _0896_ po_0.regf_0.rf\[13\]\[14\] _1042_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__mux2_1
X_1716_ _1541_ _1542_ _1518_ _1543_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__or4b_1
X_1647_ _1489_ _1493_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__or2_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _1559_ net58 _1472_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__mux2_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _0738_ _1438_ _1443_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__a21bo_1
XFILLER_73_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3179_ _1397_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__buf_2
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2550_ _0882_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__clkbuf_2
X_2481_ _0778_ po_0.regf_0.rf\[7\]\[3\] _0931_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__mux2_1
XFILLER_68_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3102_ _1363_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__clkbuf_1
X_3033_ po_0.regf_0.rf\[4\]\[5\] _0796_ _1319_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__mux2_1
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2817_ uc_0._01_ _1128_ _1129_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__nor3_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2748_ po_0.regf_0.rf\[11\]\[5\] _0961_ _1082_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__mux2_1
X_2679_ _1042_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__buf_2
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1981_ po_0.regf_0.rf\[12\]\[4\] po_0.regf_0.rf\[13\]\[4\] po_0.regf_0.rf\[14\]\[4\]
+ po_0.regf_0.rf\[15\]\[4\] _0444_ _0445_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__mux4_1
X_3651_ net166 _0299_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_2602_ po_0.regf_0.rf\[15\]\[3\] _0957_ _1004_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__mux2_1
X_3582_ net171 _0234_ VGND VGND VPWR VPWR uc_0._21_\[10\] sky130_fd_sc_hd__dfxtp_1
X_2533_ po_0.regf_0.rf\[9\]\[7\] _0966_ _0964_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__mux2_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2464_ po_0.regf_0.rf\[6\]\[13\] _0883_ _0908_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__mux2_1
X_2395_ _0729_ po_0.alu_0._11_\[12\] _0747_ net84 _0871_ VGND VGND VPWR VPWR _0872_
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3016_ net66 _1290_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__or2b_1
XFILLER_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout131 net132 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout120 net121 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout142 net153 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
Xfanout153 net191 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout164 net168 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
Xfanout186 net188 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
Xfanout175 net176 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2180_ _0668_ _0670_ _0675_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__a21bo_1
XFILLER_65_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1964_ po_0.regf_0.rf\[8\]\[2\] po_0.regf_0.rf\[9\]\[2\] po_0.regf_0.rf\[10\]\[2\]
+ po_0.regf_0.rf\[11\]\[2\] _0488_ _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__mux4_1
X_3703_ po_0.alu_0._10_\[0\] _1624_ VGND VGND VPWR VPWR po_0.alu_0._11_\[0\] sky130_fd_sc_hd__ebufn_1
X_1895_ po_0.regf_0.rf\[12\]\[14\] po_0.regf_0.rf\[13\]\[14\] po_0.regf_0.rf\[14\]\[14\]
+ po_0.regf_0.rf\[15\]\[14\] _0361_ _0362_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__mux4_1
X_3634_ net117 _0282_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_3565_ net115 _0217_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3496_ net140 _0148_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2516_ _0767_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__clkbuf_2
X_2447_ po_0.regf_0.rf\[6\]\[5\] _0797_ _0909_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__mux2_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2378_ _1522_ po_0._1_\[10\] _0855_ _0679_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__a22oi_2
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1680_ _1499_ _1492_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__or2_1
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3350_ po_0.regf_0._5_\[6\] net91 VGND VGND VPWR VPWR po_0._1_\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ _0729_ po_0.alu_0._11_\[4\] _0747_ _0629_ _0785_ VGND VGND VPWR VPWR _0786_
+ sky130_fd_sc_hd__a221o_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _1462_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__clkbuf_1
X_2232_ po_0._1_\[14\] _0707_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__and2b_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2163_ _0658_ _0659_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__and2_1
XFILLER_65_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2094_ _0601_ _1542_ _1539_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__a21bo_1
X_2996_ _1269_ _1278_ _1264_ net95 VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__a31o_1
X_1947_ po_0.regf_0.rf\[0\]\[1\] po_0.regf_0.rf\[1\]\[1\] po_0.regf_0.rf\[2\]\[1\]
+ po_0.regf_0.rf\[3\]\[1\] _0472_ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__mux4_1
X_1878_ _1585_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__and2b_1
X_3617_ net121 _0265_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_3548_ net173 _0200_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfxtp_2
X_3479_ net133 _0131_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2850_ net70 VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1801_ _1571_ _1619_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__and2b_1
X_2781_ po_0.regf_0.rf\[10\]\[4\] _0959_ _1101_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__mux2_1
X_1732_ _1556_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
X_1663_ _1503_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__clkbuf_1
X_3402_ net158 _0058_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ net134 _0021_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _1451_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__clkbuf_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _0699_ _0703_ _0706_ VGND VGND VPWR VPWR po_0.alu_0._10_\[13\] sky130_fd_sc_hd__a21oi_1
XFILLER_66_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3195_ _1413_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2146_ _0644_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__or2_1
X_2077_ po_0.regf_0.rf\[0\]\[15\] po_0.regf_0.rf\[1\]\[15\] po_0.regf_0.rf\[2\]\[15\]
+ po_0.regf_0.rf\[3\]\[15\] _0475_ _0476_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__mux4_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2979_ _1235_ net98 _1263_ _1225_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__nor4_1
XFILLER_69_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2000_ po_0.regf_0.rf\[8\]\[6\] po_0.regf_0.rf\[9\]\[6\] po_0.regf_0.rf\[10\]\[6\]
+ po_0.regf_0.rf\[11\]\[6\] _0512_ _0513_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__mux4_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2902_ _1207_ _1127_ _1208_ _1147_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__a31o_1
X_2833_ net69 VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__clkbuf_2
X_2764_ _1096_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__clkbuf_1
X_1715_ uc_0._21_\[13\] uc_0._21_\[14\] uc_0._21_\[15\] uc_0._21_\[12\] VGND VGND
+ VPWR VPWR _1543_ sky130_fd_sc_hd__a211o_1
X_2695_ _1058_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
X_1646_ _1492_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__clkbuf_2
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3316_ _1480_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__clkbuf_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _1546_ _1440_ _1441_ _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__a211oi_4
X_3178_ _1404_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2129_ po_0._1_\[4\] VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__clkbuf_2
XFILLER_81_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2480_ _0934_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
X_3101_ po_0.regf_0.rf\[3\]\[2\] _0767_ _1360_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__mux2_1
X_3032_ _1324_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2816_ uc_0._02_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__clkbuf_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2747_ _1087_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
X_2678_ _1049_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1980_ _0465_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__and2b_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3650_ net123 _0298_ VGND VGND VPWR VPWR po_0.regf_0.rf\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_2601_ _1007_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
X_3581_ net167 _0233_ VGND VGND VPWR VPWR uc_0._21_\[9\] sky130_fd_sc_hd__dfxtp_1
X_2532_ _0820_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__clkbuf_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2463_ _0923_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
X_2394_ _0692_ _0869_ _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__o21a_1
X_3015_ _1147_ _1312_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__nor2_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout110 net111 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xfanout121 net125 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout132 net133 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
Xfanout143 net147 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
Xfanout154 net157 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
Xfanout165 net168 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout187 net188 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
Xfanout176 net177 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1963_ _0459_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__clkbuf_4
X_3702_ net173 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
X_1894_ po_0.regf_0.rf\[8\]\[14\] po_0.regf_0.rf\[9\]\[14\] po_0.regf_0.rf\[10\]\[14\]
+ po_0.regf_0.rf\[11\]\[14\] _0361_ _0362_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux4_1
X_3633_ net119 _0281_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_3564_ net119 _0216_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_3495_ net143 _0147_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_2515_ _0954_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
X_2446_ _0914_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
X_2377_ _0671_ po_0._1_\[9\] _0846_ _0831_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__o22a_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2300_ _0780_ _0783_ _0784_ _0748_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__o211a_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ po_0.muxf_0.rf_w_data\[1\] _1136_ _1460_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__mux2_1
X_2231_ _0716_ _0717_ _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__nand3b_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2162_ _0658_ _0659_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__nor2_1
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2093_ _1535_ _1541_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__or2_1
XFILLER_80_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2995_ _1286_ _1291_ _1292_ _1293_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__nand4_1
X_1946_ _0459_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__buf_2
X_1877_ po_0.regf_0.rf\[8\]\[12\] po_0.regf_0.rf\[9\]\[12\] po_0.regf_0.rf\[10\]\[12\]
+ po_0.regf_0.rf\[11\]\[12\] _1573_ _1575_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__mux4_1
X_3616_ net156 _0264_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3547_ net172 _0199_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfxtp_1
X_3478_ net139 _0130_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2429_ net7 _0728_ _0901_ _0902_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__a22o_2
XFILLER_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1800_ po_0.regf_0.rf\[0\]\[3\] po_0.regf_0.rf\[1\]\[3\] po_0.regf_0.rf\[2\]\[3\]
+ po_0.regf_0.rf\[3\]\[3\] _1573_ _1575_ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__mux4_1
X_2780_ _1105_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
X_1731_ po_0.regf_0.rq_addr\[1\] _1555_ _1553_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__mux2_1
X_1662_ _1500_ _1502_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__or2_1
X_3401_ net115 _0057_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_3332_ net136 _0020_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ po_0.regf_0.rp_addr\[3\] uc_0._21_\[11\] _0595_ VGND VGND VPWR VPWR _1451_
+ sky130_fd_sc_hd__mux2_1
X_3194_ po_0.regf_0.rf\[2\]\[13\] _0882_ _1397_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__mux2_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _0701_ _0702_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__o21ai_1
X_2145_ _0643_ _0642_ _0639_ _0634_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__a211oi_1
XFILLER_66_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2076_ _0450_ _0588_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__and2b_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2978_ _1258_ _1271_ _1257_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__and3_1
X_1929_ _0442_ _0443_ _0448_ _0454_ _0456_ VGND VGND VPWR VPWR po_0.regf_0._3_\[0\]
+ sky130_fd_sc_hd__a32oi_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2901_ _1161_ _1179_ _1193_ _1175_ _1206_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__a41o_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2832_ _1133_ _1135_ _1143_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__o21a_1
X_2763_ po_0.regf_0.rf\[11\]\[12\] _0976_ _1081_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__mux2_1
X_1714_ uc_0.bc_0._05_\[3\] VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__clkbuf_2
X_2694_ _0883_ po_0.regf_0.rf\[13\]\[13\] _1042_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__mux2_1
X_1645_ _1491_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _1557_ net57 _1472_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__mux2_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3246_ _1552_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__clkbuf_4
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ po_0.regf_0.rf\[2\]\[5\] _0796_ _1398_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__mux2_1
X_2128_ net45 VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__clkbuf_2
XFILLER_81_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2059_ po_0.regf_0.rf\[4\]\[13\] po_0.regf_0.rf\[5\]\[13\] po_0.regf_0.rf\[6\]\[13\]
+ po_0.regf_0.rf\[7\]\[13\] _0439_ _0440_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__mux4_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3100_ _1362_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__clkbuf_1
Xoutput80 net80 VGND VGND VPWR VPWR leds[1] sky130_fd_sc_hd__buf_2
X_3031_ po_0.regf_0.rf\[4\]\[4\] _0788_ _1319_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__mux2_1
XFILLER_51_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2815_ uc_0._00_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__clkbuf_2
XFILLER_31_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2746_ po_0.regf_0.rf\[11\]\[4\] _0959_ _1082_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__mux2_1
X_2677_ _0797_ po_0.regf_0.rf\[13\]\[5\] _1043_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__mux2_1
XFILLER_86_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3229_ po_0.regf_0.rf\[8\]\[13\] _0882_ _1416_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__mux2_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2600_ po_0.regf_0.rf\[15\]\[2\] _0955_ _1004_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__mux2_1
X_3580_ net178 _0232_ VGND VGND VPWR VPWR uc_0._21_\[8\] sky130_fd_sc_hd__dfxtp_1
X_2531_ _0965_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
X_2462_ po_0.regf_0.rf\[6\]\[12\] _0874_ _0908_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__mux2_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2393_ _0869_ _0692_ _0731_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3014_ _1297_ _1310_ _1127_ _1311_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__o211a_1
XFILLER_36_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2729_ _1077_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout111 net114 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
Xfanout100 net102 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout122 net123 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout133 net142 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout144 net147 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
Xfanout155 net157 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout177 net190 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout188 net189 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout166 net168 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1962_ _0457_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__buf_4
X_3701_ net182 uc_0.bc_0._70_\[3\] VGND VGND VPWR VPWR uc_0.bc_0._05_\[3\] sky130_fd_sc_hd__dfxtp_1
X_1893_ _0418_ _0420_ _1596_ _0423_ VGND VGND VPWR VPWR po_0.regf_0._5_\[13\] sky130_fd_sc_hd__o22a_1
X_3632_ net154 _0280_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_3563_ net154 _0215_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3494_ net149 _0146_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_2514_ po_0.regf_0.rf\[9\]\[1\] _0953_ _0951_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__mux2_1
X_2445_ po_0.regf_0.rf\[6\]\[4\] _0789_ _0909_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__mux2_1
X_2376_ _0854_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _0711_ _0705_ _0718_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2161_ po_0._1_\[7\] VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2092_ _0600_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2994_ _1286_ _1291_ _1292_ _1293_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__a22o_1
XFILLER_61_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1945_ _0457_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__clkbuf_4
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1876_ _0403_ _0405_ _1596_ _0408_ VGND VGND VPWR VPWR po_0.regf_0._5_\[11\] sky130_fd_sc_hd__o22a_1
X_3615_ net157 _0263_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3546_ net171 _0198_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfxtp_2
X_3477_ net137 _0129_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2428_ _1491_ po_0.alu_0._11_\[15\] _0859_ net41 _0732_ VGND VGND VPWR VPWR _0902_
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2359_ _0666_ _0831_ _0673_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1730_ uc_0._21_\[5\] VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__clkbuf_2
X_1661_ _1492_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__dlymetal6s2s_1
X_3400_ net119 _0056_ VGND VGND VPWR VPWR po_0.regf_0.rf\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_3331_ net129 _0019_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _1450_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__clkbuf_1
X_3193_ _1412_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__clkbuf_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _0694_ _0697_ _0704_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__o21bai_2
XFILLER_38_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2144_ _0634_ _0639_ _0642_ _0643_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__o211a_1
X_2075_ po_0.regf_0.rf\[8\]\[15\] po_0.regf_0.rf\[9\]\[15\] po_0.regf_0.rf\[10\]\[15\]
+ po_0.regf_0.rf\[11\]\[15\] _0472_ _0473_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__mux4_1
XFILLER_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2977_ net96 VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__clkbuf_2
X_1928_ _0455_ _0447_ _0443_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a21oi_1
X_1859_ _0392_ _0393_ _1613_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__mux2_1
XFILLER_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3529_ net151 _0181_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2900_ _1206_ _1201_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__nand2_1
X_2831_ _1139_ _1121_ _1140_ _1142_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__a31o_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2762_ _1095_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__clkbuf_1
X_1713_ uc_0.bc_0._05_\[2\] VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2693_ _1057_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1644_ _1490_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__clkbuf_2
XFILLER_86_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ _1479_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__clkbuf_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _1520_ uc_0.bc_0._70_\[0\] _1357_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__and3_2
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3176_ _1403_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2127_ _0628_ VGND VGND VPWR VPWR po_0.alu_0._10_\[3\] sky130_fd_sc_hd__clkbuf_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2058_ po_0.regf_0.rf\[0\]\[13\] po_0.regf_0.rf\[1\]\[13\] po_0.regf_0.rf\[2\]\[13\]
+ po_0.regf_0.rf\[3\]\[13\] _0451_ _0452_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__mux4_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput70 net70 VGND VGND VPWR VPWR I_addr[3] sky130_fd_sc_hd__buf_2
Xoutput81 net81 VGND VGND VPWR VPWR leds[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3030_ _1323_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2814_ _1126_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__clkbuf_2
X_2745_ _1086_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
X_2676_ _1048_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3228_ _1431_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__clkbuf_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3159_ _0883_ po_0.regf_0.rf\[0\]\[13\] _1378_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__mux2_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2530_ po_0.regf_0.rf\[9\]\[6\] _0963_ _0964_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__mux2_1
XFILLER_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2461_ _0922_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
X_2392_ _0683_ _0865_ _0866_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__o22ai_4
XFILLER_68_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3013_ _1290_ _1264_ _1283_ net67 VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__a31o_1
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2728_ po_0.regf_0.rf\[12\]\[12\] _0976_ _1062_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__mux2_1
X_2659_ _0883_ po_0.regf_0.rf\[14\]\[13\] _1023_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__mux2_1
Xfanout101 net102 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
Xfanout112 net114 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
Xfanout134 net136 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout145 net147 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
Xfanout123 net124 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
Xfanout156 net157 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout189 net190 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout167 net168 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_1
Xfanout178 net189 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3700_ net182 uc_0.bc_0._70_\[2\] VGND VGND VPWR VPWR uc_0.bc_0._05_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1961_ _0438_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__buf_2
X_1892_ _0421_ _0422_ _1613_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux2_1
X_3631_ net160 _0279_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_3562_ net155 _0214_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_2513_ _0755_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__clkbuf_2
X_3493_ net138 _0145_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_2444_ _0913_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
X_2375_ po_0.regf_0.rf\[5\]\[10\] _0853_ _0810_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__mux2_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ net48 VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2091_ po_0.regf_0.rp_addr\[3\] uc_0._21_\[11\] _0596_ VGND VGND VPWR VPWR _0600_
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2993_ net64 net95 VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__or2_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1944_ _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__buf_2
X_3614_ net137 _0262_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_1875_ _0406_ _0407_ _1613_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux2_1
X_3545_ net171 _0197_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfxtp_2
X_3476_ net132 _0128_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2427_ _0899_ _0900_ _0762_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__nand3_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2358_ _0666_ _0673_ _0831_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__or3_1
XFILLER_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2289_ _0731_ _0771_ _0772_ _0774_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__o31ai_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1660_ _1501_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__clkbuf_1
X_3330_ net136 _0018_ VGND VGND VPWR VPWR po_0.regf_0.rf\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ po_0.regf_0.rp_addr\[2\] uc_0._21_\[10\] _0595_ VGND VGND VPWR VPWR _1450_
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3192_ po_0.regf_0.rf\[2\]\[12\] _0873_ _1397_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__mux2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _0692_ _0701_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__or2_1
XFILLER_78_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2143_ net46 po_0._1_\[5\] VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__or2_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2074_ _0586_ _0530_ _0003_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__a21bo_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2976_ _1119_ _1156_ _1248_ _1269_ _1277_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__o41a_1
X_1927_ po_0.regf_0.rf\[4\]\[0\] po_0.regf_0.rf\[5\]\[0\] po_0.regf_0.rf\[6\]\[0\]
+ po_0.regf_0.rf\[7\]\[0\] _0444_ _0445_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__mux4_1
X_1858_ po_0.regf_0.rf\[12\]\[9\] po_0.regf_0.rf\[13\]\[9\] po_0.regf_0.rf\[14\]\[9\]
+ po_0.regf_0.rf\[15\]\[9\] _1600_ _1601_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__mux4_1
X_1789_ _1572_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__buf_4
XFILLER_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3528_ net150 _0180_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_3459_ net107 _0111_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2830_ _1123_ _1133_ _1130_ _1141_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__o22a_1
X_2761_ po_0.regf_0.rf\[11\]\[11\] _0974_ _1089_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__mux2_1
X_2692_ _0874_ po_0.regf_0.rf\[13\]\[12\] _1042_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__mux2_1
X_1712_ _1523_ _1529_ _1532_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__o21ai_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 _0493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1643_ po_0.alu_0.s1 VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__inv_2
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _1555_ net56 _1472_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__mux2_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _1439_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__inv_2
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3175_ po_0.regf_0.rf\[2\]\[4\] _0788_ _1398_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__mux2_1
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2126_ _0622_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__and2_1
XFILLER_66_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2057_ _0567_ _0569_ _0443_ _0572_ VGND VGND VPWR VPWR po_0.regf_0._3_\[12\] sky130_fd_sc_hd__o22a_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2959_ _1257_ _1260_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__nand2_1
XFILLER_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput60 net60 VGND VGND VPWR VPWR D_wr sky130_fd_sc_hd__buf_2
Xoutput71 net71 VGND VGND VPWR VPWR I_addr[4] sky130_fd_sc_hd__clkbuf_4
Xoutput82 net82 VGND VGND VPWR VPWR leds[3] sky130_fd_sc_hd__buf_2
XFILLER_48_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2813_ uc_0._02_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__clkbuf_2
X_2744_ po_0.regf_0.rf\[11\]\[3\] _0957_ _1082_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__mux2_1
X_2675_ _0789_ po_0.regf_0.rf\[13\]\[4\] _1043_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__mux2_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ po_0.regf_0.rf\[8\]\[12\] _0873_ _1416_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__mux2_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3158_ _1393_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2109_ po_0._1_\[1\] _0610_ _0604_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__o21ai_1
X_3089_ uc_0._21_\[15\] net23 _1343_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__mux2_1
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2460_ po_0.regf_0.rf\[6\]\[11\] _0862_ _0916_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__mux2_1
X_2391_ _0826_ _0782_ _0626_ _0867_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__a31oi_4
XFILLER_68_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3012_ net94 net67 VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__xor2_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2727_ _1076_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
X_2658_ _1038_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
X_2589_ _1000_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
Xfanout102 net106 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
Xfanout113 net114 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout135 net136 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_1
Xfanout146 net147 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout124 net125 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout157 net170 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout168 net169 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout179 net186 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1960_ _0485_ _0447_ _0463_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__a21bo_1
X_1891_ po_0.regf_0.rf\[4\]\[13\] po_0.regf_0.rf\[5\]\[13\] po_0.regf_0.rf\[6\]\[13\]
+ po_0.regf_0.rf\[7\]\[13\] _1561_ _1563_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__mux4_1
X_3630_ net148 _0278_ VGND VGND VPWR VPWR po_0.regf_0.rf\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_3561_ net135 _0213_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_2512_ _0952_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
X_3492_ net132 _0144_ VGND VGND VPWR VPWR po_0.regf_0.rf\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_2443_ po_0.regf_0.rf\[6\]\[3\] _0778_ _0909_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__mux2_1
X_2374_ _0852_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2090_ _0599_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2992_ net96 net95 VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__nand2_1
X_1943_ _0003_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__buf_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3613_ net139 _0261_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1874_ po_0.regf_0.rf\[4\]\[11\] po_0.regf_0.rf\[5\]\[11\] po_0.regf_0.rf\[6\]\[11\]
+ po_0.regf_0.rf\[7\]\[11\] _1561_ _1563_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__mux4_1
X_3544_ net176 _0196_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfxtp_1
X_3475_ net100 _0127_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_2426_ _0714_ _0715_ _0889_ _0708_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__o211ai_1
XFILLER_29_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2357_ _0837_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2288_ _0773_ po_0.alu_0._11_\[3\] _0746_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__a21oi_1
XFILLER_56_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _1449_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__clkbuf_1
X_3191_ _1411_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__clkbuf_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _0701_ _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__and2_1
XFILLER_66_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2142_ _0640_ _0641_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__nand2_1
X_2073_ po_0.regf_0.rf\[12\]\[15\] po_0.regf_0.rf\[13\]\[15\] po_0.regf_0.rf\[14\]\[15\]
+ po_0.regf_0.rf\[15\]\[15\] _0488_ _0489_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__mux4_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2975_ _1272_ _1273_ _1121_ _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__a31o_1
X_1926_ _0450_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__or2b_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1857_ po_0.regf_0.rf\[8\]\[9\] po_0.regf_0.rf\[9\]\[9\] po_0.regf_0.rf\[10\]\[9\]
+ po_0.regf_0.rf\[11\]\[9\] _1609_ _1610_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__mux4_1
X_3527_ net146 _0179_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1788_ _1591_ _1607_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__and2b_1
X_3458_ net112 _0110_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_3389_ net109 _0045_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_2409_ _0884_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2760_ _1094_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__clkbuf_1
X_1711_ uc_0.bc_0._05_\[0\] VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__dlymetal6s2s_1
X_2691_ _1056_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
X_1642_ _1488_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__clkbuf_2
XANTENNA_2 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _1478_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__clkbuf_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _1357_ _1517_ _1520_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__or3b_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _1402_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__clkbuf_1
X_2125_ _0623_ _0624_ _0625_ _0626_ _0615_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__o2111ai_1
XFILLER_54_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2056_ _0570_ _0571_ _0438_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__mux2_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2958_ _1257_ _1260_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__or2_1
XFILLER_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1909_ _0432_ _0434_ _1568_ _0437_ VGND VGND VPWR VPWR po_0.regf_0._5_\[15\] sky130_fd_sc_hd__o22a_1
X_2889_ _1185_ _1192_ _1194_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__nand3b_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput50 net50 VGND VGND VPWR VPWR D_W_data[9] sky130_fd_sc_hd__clkbuf_4
Xoutput61 net61 VGND VGND VPWR VPWR I_addr[0] sky130_fd_sc_hd__buf_2
Xoutput72 net72 VGND VGND VPWR VPWR I_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_48_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2812_ _1123_ _1124_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2743_ _1085_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
X_2674_ _1047_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3226_ _1430_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__clkbuf_1
X_3157_ _0874_ po_0.regf_0.rf\[0\]\[12\] _1378_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__mux2_1
XFILLER_39_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2108_ _0610_ po_0._1_\[1\] VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__nand2_1
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3088_ _1354_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__clkbuf_1
X_2039_ po_0.regf_0.rf\[4\]\[10\] po_0.regf_0.rf\[5\]\[10\] po_0.regf_0.rf\[6\]\[10\]
+ po_0.regf_0.rf\[7\]\[10\] _0451_ _0452_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__mux4_1
XFILLER_52_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2390_ _0829_ _0828_ _0660_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3011_ _1302_ _1309_ _1135_ net94 VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2726_ po_0.regf_0.rf\[12\]\[11\] _0974_ _1070_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__mux2_1
X_2657_ _0874_ po_0.regf_0.rf\[14\]\[12\] _1023_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__mux2_1
X_2588_ po_0.regf_0.rf\[1\]\[13\] _0978_ _0984_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__mux2_1
Xfanout103 net106 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
Xfanout136 net142 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
Xfanout114 net126 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
Xfanout147 net153 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
Xfanout125 net126 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout158 net161 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
Xfanout169 net170 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3209_ _1421_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1890_ po_0.regf_0.rf\[0\]\[13\] po_0.regf_0.rf\[1\]\[13\] po_0.regf_0.rf\[2\]\[13\]
+ po_0.regf_0.rf\[3\]\[13\] _1609_ _1610_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux4_1
X_3560_ net136 _0212_ VGND VGND VPWR VPWR po_0.regf_0.rf\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_2511_ po_0.regf_0.rf\[9\]\[0\] _0949_ _0951_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__mux2_1
X_3491_ net100 _0143_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_2442_ _0912_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2373_ net2 _0823_ _0851_ _0753_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__a22o_2
XFILLER_68_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2709_ po_0.regf_0.rf\[12\]\[3\] _0957_ _1063_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__mux2_1
X_3689_ net180 _0337_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dfxtp_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2991_ net96 _1269_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__or2b_1
X_1942_ _0465_ _0468_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__and2b_1
X_1873_ po_0.regf_0.rf\[0\]\[11\] po_0.regf_0.rf\[1\]\[11\] po_0.regf_0.rf\[2\]\[11\]
+ po_0.regf_0.rf\[3\]\[11\] _1609_ _1610_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__mux4_1
X_3612_ net131 _0260_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_3543_ net176 _0195_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfxtp_1
X_3474_ net103 _0126_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_2425_ _0718_ _0898_ _0716_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__o21bai_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2356_ po_0.regf_0.rf\[5\]\[8\] _0836_ _0810_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__mux2_1
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2287_ po_0.alu_0.s1 VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__clkbuf_2
XFILLER_84_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ po_0._1_\[12\] net84 VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__or2b_1
X_3190_ po_0.regf_0.rf\[2\]\[11\] _0861_ _1405_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__mux2_1
X_2141_ po_0._1_\[5\] VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__clkbuf_2
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2072_ _0579_ _0581_ _0583_ _0585_ VGND VGND VPWR VPWR po_0.regf_0._3_\[14\] sky130_fd_sc_hd__o22a_1
XFILLER_38_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2974_ _1274_ _1275_ _1134_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__o21ai_1
X_1925_ po_0.regf_0.rf\[0\]\[0\] po_0.regf_0.rf\[1\]\[0\] po_0.regf_0.rf\[2\]\[0\]
+ po_0.regf_0.rf\[3\]\[0\] _0451_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__mux4_1
X_1856_ _0390_ _1585_ _1568_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__a21o_1
X_1787_ po_0.regf_0.rf\[8\]\[2\] po_0.regf_0.rf\[9\]\[2\] po_0.regf_0.rf\[10\]\[2\]
+ po_0.regf_0.rf\[11\]\[2\] _1592_ _1593_ VGND VGND VPWR VPWR _1607_ sky130_fd_sc_hd__mux4_1
X_3526_ net150 _0178_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3457_ net127 _0109_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_3388_ net105 _0044_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_2408_ po_0.regf_0.rf\[5\]\[13\] _0883_ _0743_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__mux2_1
X_2339_ _0820_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1710_ _1538_ VGND VGND VPWR VPWR uc_0.bc_0._70_\[1\] sky130_fd_sc_hd__inv_2
X_2690_ _0862_ po_0.regf_0.rf\[13\]\[11\] _1050_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__mux2_1
XFILLER_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1641_ _1487_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__clkbuf_2
XANTENNA_3 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3311_ _1549_ net55 _1472_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__mux2_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ net88 _1358_ _0596_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__a21o_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ po_0.regf_0.rf\[2\]\[3\] _0777_ _1398_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__mux2_1
X_2124_ net44 po_0._1_\[3\] VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__or2_2
X_2055_ po_0.regf_0.rf\[4\]\[12\] po_0.regf_0.rf\[5\]\[12\] po_0.regf_0.rf\[6\]\[12\]
+ po_0.regf_0.rf\[7\]\[12\] _0451_ _0452_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__mux4_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2957_ _1258_ _1241_ _1247_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__o2bb2ai_1
X_1908_ _0435_ _0436_ _1566_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__mux2_1
X_2888_ uc_0._21_\[4\] net71 _1195_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__o21ai_1
X_1839_ po_0.regf_0.rf\[12\]\[7\] po_0.regf_0.rf\[13\]\[7\] po_0.regf_0.rf\[14\]\[7\]
+ po_0.regf_0.rf\[15\]\[7\] _1578_ _1579_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__mux4_1
X_3509_ net146 _0161_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput51 net51 VGND VGND VPWR VPWR D_addr[0] sky130_fd_sc_hd__buf_2
Xoutput40 net40 VGND VGND VPWR VPWR D_W_data[14] sky130_fd_sc_hd__buf_2
Xoutput73 net73 VGND VGND VPWR VPWR I_addr[6] sky130_fd_sc_hd__clkbuf_4
Xoutput62 net62 VGND VGND VPWR VPWR I_addr[10] sky130_fd_sc_hd__buf_2
XFILLER_48_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2811_ uc_0._21_\[0\] VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__clkbuf_2
XFILLER_31_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2742_ po_0.regf_0.rf\[11\]\[2\] _0955_ _1082_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__mux2_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2673_ _0778_ po_0.regf_0.rf\[13\]\[3\] _1043_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__mux2_1
XFILLER_86_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3225_ po_0.regf_0.rf\[8\]\[11\] _0861_ _1424_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__mux2_1
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3156_ _1392_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2107_ net87 VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__inv_2
X_3087_ uc_0._21_\[14\] net22 _1343_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__mux2_1
X_2038_ po_0.regf_0.rf\[0\]\[10\] po_0.regf_0.rf\[1\]\[10\] po_0.regf_0.rf\[2\]\[10\]
+ po_0.regf_0.rf\[3\]\[10\] _0524_ _0525_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__mux4_1
XFILLER_50_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3010_ _1307_ _1308_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__nand2_1
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2725_ _1075_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
X_2656_ _1037_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
Xfanout104 net106 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
X_2587_ _0999_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout137 net141 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
Xfanout115 net117 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
Xfanout126 net191 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout148 net152 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
Xfanout159 net161 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
X_3208_ po_0.regf_0.rf\[8\]\[3\] _0777_ _1417_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__mux2_1
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3139_ _1383_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3490_ net104 _0142_ VGND VGND VPWR VPWR po_0.regf_0.rf\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_2510_ _0950_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__buf_2
X_2441_ po_0.regf_0.rf\[6\]\[2\] _0768_ _0909_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__mux2_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2372_ _0848_ _0762_ _0849_ _0850_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__a31o_1
XFILLER_68_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2708_ _1066_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
X_3688_ net175 _0336_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dfxtp_1
X_2639_ _1028_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2990_ net95 VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1941_ po_0.regf_0.rf\[8\]\[1\] po_0.regf_0.rf\[9\]\[1\] po_0.regf_0.rf\[10\]\[1\]
+ po_0.regf_0.rf\[11\]\[1\] _0466_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__mux4_1
X_1872_ _1603_ _0404_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__and2b_1
X_3611_ net139 _0259_ VGND VGND VPWR VPWR po_0.regf_0.rf\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_3542_ net174 _0194_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfxtp_2
X_3473_ net110 _0125_ VGND VGND VPWR VPWR po_0.regf_0.rf\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_2424_ _0885_ _0887_ _0888_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__a21oi_1
X_2355_ _0835_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__clkbuf_2
XFILLER_84_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2286_ _0619_ _0621_ _0761_ _0770_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__o211a_1
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2140_ net46 VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__clkbuf_2
X_2071_ _0584_ _0447_ _0470_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__a21o_1
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2973_ _1269_ _1264_ _1157_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__o21ai_1
X_1924_ _0001_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__clkbuf_4
X_1855_ po_0.regf_0.rf\[4\]\[9\] po_0.regf_0.rf\[5\]\[9\] po_0.regf_0.rf\[6\]\[9\]
+ po_0.regf_0.rf\[7\]\[9\] _1562_ _1564_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux4_1
X_1786_ _1605_ _1567_ _1589_ VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__a21o_1
X_3525_ net146 _0177_ VGND VGND VPWR VPWR po_0.regf_0.rf\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_3456_ net107 _0108_ VGND VGND VPWR VPWR po_0.regf_0.rf\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_2407_ _0882_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__dlymetal6s2s_1
X_3387_ net115 _0043_ VGND VGND VPWR VPWR po_0.regf_0.rf\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2338_ po_0.muxf_0.rf_w_data\[7\] _0725_ _0727_ net14 _0819_ VGND VGND VPWR VPWR
+ _0820_ sky130_fd_sc_hd__a221o_4
XFILLER_69_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2269_ po_0.regf_0.rf\[5\]\[1\] _0756_ _0744_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__mux2_1
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1640_ po_0.alu_0.s0 VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__clkbuf_2
XANTENNA_4 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3310_ _1477_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__clkbuf_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _1438_ net92 _1553_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__a21o_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3172_ _1401_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2123_ _0620_ _0618_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__nand2_1
XFILLER_66_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2054_ po_0.regf_0.rf\[0\]\[12\] po_0.regf_0.rf\[1\]\[12\] po_0.regf_0.rf\[2\]\[12\]
+ po_0.regf_0.rf\[3\]\[12\] _0524_ _0525_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__mux4_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2956_ _1235_ _1225_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__nor2_1
X_1907_ po_0.regf_0.rf\[4\]\[15\] po_0.regf_0.rf\[5\]\[15\] po_0.regf_0.rf\[6\]\[15\]
+ po_0.regf_0.rf\[7\]\[15\] _1561_ _1563_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__mux4_1
X_2887_ _1192_ _1194_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__nand2_1
X_1838_ _1591_ _0374_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__and2b_1
X_1769_ _1588_ _1567_ _1589_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__a21o_1
X_3508_ net145 _0160_ VGND VGND VPWR VPWR po_0.regf_0.rf\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_3439_ net120 _0091_ VGND VGND VPWR VPWR po_0.regf_0.rf\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput52 net52 VGND VGND VPWR VPWR D_addr[1] sky130_fd_sc_hd__clkbuf_4
Xoutput41 net41 VGND VGND VPWR VPWR D_W_data[15] sky130_fd_sc_hd__buf_2
Xoutput63 net97 VGND VGND VPWR VPWR I_addr[11] sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 VGND VGND VPWR VPWR I_addr[7] sky130_fd_sc_hd__buf_2
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2810_ _1122_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__clkbuf_2
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2741_ _1084_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
X_2672_ _1046_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3224_ _1429_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__clkbuf_1
.ends

