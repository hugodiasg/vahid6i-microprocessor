// This is the unpowered netlist.
module vahid6i (D_rd,
    D_wr,
    I_rd,
    clock,
    led_clock,
    reset,
    D_R_data,
    D_W_data,
    D_addr,
    I_addr,
    I_data,
    leds);
 output D_rd;
 output D_wr;
 output I_rd;
 input clock;
 output led_clock;
 input reset;
 input [15:0] D_R_data;
 output [15:0] D_W_data;
 output [7:0] D_addr;
 output [15:0] I_addr;
 input [15:0] I_data;
 output [3:0] leds;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \po_0._1_[0] ;
 wire \po_0._1_[10] ;
 wire \po_0._1_[11] ;
 wire \po_0._1_[12] ;
 wire \po_0._1_[13] ;
 wire \po_0._1_[14] ;
 wire \po_0._1_[15] ;
 wire \po_0._1_[1] ;
 wire \po_0._1_[2] ;
 wire \po_0._1_[3] ;
 wire \po_0._1_[4] ;
 wire \po_0._1_[5] ;
 wire \po_0._1_[6] ;
 wire \po_0._1_[7] ;
 wire \po_0._1_[8] ;
 wire \po_0._1_[9] ;
 wire \po_0.alu_0._10_[0] ;
 wire \po_0.alu_0._10_[10] ;
 wire \po_0.alu_0._10_[11] ;
 wire \po_0.alu_0._10_[12] ;
 wire \po_0.alu_0._10_[13] ;
 wire \po_0.alu_0._10_[14] ;
 wire \po_0.alu_0._10_[15] ;
 wire \po_0.alu_0._10_[1] ;
 wire \po_0.alu_0._10_[2] ;
 wire \po_0.alu_0._10_[3] ;
 wire \po_0.alu_0._10_[4] ;
 wire \po_0.alu_0._10_[5] ;
 wire \po_0.alu_0._10_[6] ;
 wire \po_0.alu_0._10_[7] ;
 wire \po_0.alu_0._10_[8] ;
 wire \po_0.alu_0._10_[9] ;
 wire \po_0.alu_0._11_[0] ;
 wire \po_0.alu_0._11_[10] ;
 wire \po_0.alu_0._11_[11] ;
 wire \po_0.alu_0._11_[12] ;
 wire \po_0.alu_0._11_[13] ;
 wire \po_0.alu_0._11_[14] ;
 wire \po_0.alu_0._11_[15] ;
 wire \po_0.alu_0._11_[1] ;
 wire \po_0.alu_0._11_[2] ;
 wire \po_0.alu_0._11_[3] ;
 wire \po_0.alu_0._11_[4] ;
 wire \po_0.alu_0._11_[5] ;
 wire \po_0.alu_0._11_[6] ;
 wire \po_0.alu_0._11_[7] ;
 wire \po_0.alu_0._11_[8] ;
 wire \po_0.alu_0._11_[9] ;
 wire \po_0.alu_0.s0 ;
 wire \po_0.alu_0.s1 ;
 wire \po_0.muxf_0.rf_w_data[0] ;
 wire \po_0.muxf_0.rf_w_data[1] ;
 wire \po_0.muxf_0.rf_w_data[2] ;
 wire \po_0.muxf_0.rf_w_data[3] ;
 wire \po_0.muxf_0.rf_w_data[4] ;
 wire \po_0.muxf_0.rf_w_data[5] ;
 wire \po_0.muxf_0.rf_w_data[6] ;
 wire \po_0.muxf_0.rf_w_data[7] ;
 wire \po_0.muxf_0.s0 ;
 wire \po_0.muxf_0.s1 ;
 wire \po_0.regf_0._3_[0] ;
 wire \po_0.regf_0._3_[10] ;
 wire \po_0.regf_0._3_[11] ;
 wire \po_0.regf_0._3_[12] ;
 wire \po_0.regf_0._3_[13] ;
 wire \po_0.regf_0._3_[14] ;
 wire \po_0.regf_0._3_[15] ;
 wire \po_0.regf_0._3_[1] ;
 wire \po_0.regf_0._3_[2] ;
 wire \po_0.regf_0._3_[3] ;
 wire \po_0.regf_0._3_[4] ;
 wire \po_0.regf_0._3_[5] ;
 wire \po_0.regf_0._3_[6] ;
 wire \po_0.regf_0._3_[7] ;
 wire \po_0.regf_0._3_[8] ;
 wire \po_0.regf_0._3_[9] ;
 wire \po_0.regf_0._5_[0] ;
 wire \po_0.regf_0._5_[10] ;
 wire \po_0.regf_0._5_[11] ;
 wire \po_0.regf_0._5_[12] ;
 wire \po_0.regf_0._5_[13] ;
 wire \po_0.regf_0._5_[14] ;
 wire \po_0.regf_0._5_[15] ;
 wire \po_0.regf_0._5_[1] ;
 wire \po_0.regf_0._5_[2] ;
 wire \po_0.regf_0._5_[3] ;
 wire \po_0.regf_0._5_[4] ;
 wire \po_0.regf_0._5_[5] ;
 wire \po_0.regf_0._5_[6] ;
 wire \po_0.regf_0._5_[7] ;
 wire \po_0.regf_0._5_[8] ;
 wire \po_0.regf_0._5_[9] ;
 wire \po_0.regf_0.rf[0][0] ;
 wire \po_0.regf_0.rf[0][10] ;
 wire \po_0.regf_0.rf[0][11] ;
 wire \po_0.regf_0.rf[0][12] ;
 wire \po_0.regf_0.rf[0][13] ;
 wire \po_0.regf_0.rf[0][14] ;
 wire \po_0.regf_0.rf[0][15] ;
 wire \po_0.regf_0.rf[0][1] ;
 wire \po_0.regf_0.rf[0][2] ;
 wire \po_0.regf_0.rf[0][3] ;
 wire \po_0.regf_0.rf[0][4] ;
 wire \po_0.regf_0.rf[0][5] ;
 wire \po_0.regf_0.rf[0][6] ;
 wire \po_0.regf_0.rf[0][7] ;
 wire \po_0.regf_0.rf[0][8] ;
 wire \po_0.regf_0.rf[0][9] ;
 wire \po_0.regf_0.rf[10][0] ;
 wire \po_0.regf_0.rf[10][10] ;
 wire \po_0.regf_0.rf[10][11] ;
 wire \po_0.regf_0.rf[10][12] ;
 wire \po_0.regf_0.rf[10][13] ;
 wire \po_0.regf_0.rf[10][14] ;
 wire \po_0.regf_0.rf[10][15] ;
 wire \po_0.regf_0.rf[10][1] ;
 wire \po_0.regf_0.rf[10][2] ;
 wire \po_0.regf_0.rf[10][3] ;
 wire \po_0.regf_0.rf[10][4] ;
 wire \po_0.regf_0.rf[10][5] ;
 wire \po_0.regf_0.rf[10][6] ;
 wire \po_0.regf_0.rf[10][7] ;
 wire \po_0.regf_0.rf[10][8] ;
 wire \po_0.regf_0.rf[10][9] ;
 wire \po_0.regf_0.rf[11][0] ;
 wire \po_0.regf_0.rf[11][10] ;
 wire \po_0.regf_0.rf[11][11] ;
 wire \po_0.regf_0.rf[11][12] ;
 wire \po_0.regf_0.rf[11][13] ;
 wire \po_0.regf_0.rf[11][14] ;
 wire \po_0.regf_0.rf[11][15] ;
 wire \po_0.regf_0.rf[11][1] ;
 wire \po_0.regf_0.rf[11][2] ;
 wire \po_0.regf_0.rf[11][3] ;
 wire \po_0.regf_0.rf[11][4] ;
 wire \po_0.regf_0.rf[11][5] ;
 wire \po_0.regf_0.rf[11][6] ;
 wire \po_0.regf_0.rf[11][7] ;
 wire \po_0.regf_0.rf[11][8] ;
 wire \po_0.regf_0.rf[11][9] ;
 wire \po_0.regf_0.rf[12][0] ;
 wire \po_0.regf_0.rf[12][10] ;
 wire \po_0.regf_0.rf[12][11] ;
 wire \po_0.regf_0.rf[12][12] ;
 wire \po_0.regf_0.rf[12][13] ;
 wire \po_0.regf_0.rf[12][14] ;
 wire \po_0.regf_0.rf[12][15] ;
 wire \po_0.regf_0.rf[12][1] ;
 wire \po_0.regf_0.rf[12][2] ;
 wire \po_0.regf_0.rf[12][3] ;
 wire \po_0.regf_0.rf[12][4] ;
 wire \po_0.regf_0.rf[12][5] ;
 wire \po_0.regf_0.rf[12][6] ;
 wire \po_0.regf_0.rf[12][7] ;
 wire \po_0.regf_0.rf[12][8] ;
 wire \po_0.regf_0.rf[12][9] ;
 wire \po_0.regf_0.rf[13][0] ;
 wire \po_0.regf_0.rf[13][10] ;
 wire \po_0.regf_0.rf[13][11] ;
 wire \po_0.regf_0.rf[13][12] ;
 wire \po_0.regf_0.rf[13][13] ;
 wire \po_0.regf_0.rf[13][14] ;
 wire \po_0.regf_0.rf[13][15] ;
 wire \po_0.regf_0.rf[13][1] ;
 wire \po_0.regf_0.rf[13][2] ;
 wire \po_0.regf_0.rf[13][3] ;
 wire \po_0.regf_0.rf[13][4] ;
 wire \po_0.regf_0.rf[13][5] ;
 wire \po_0.regf_0.rf[13][6] ;
 wire \po_0.regf_0.rf[13][7] ;
 wire \po_0.regf_0.rf[13][8] ;
 wire \po_0.regf_0.rf[13][9] ;
 wire \po_0.regf_0.rf[14][0] ;
 wire \po_0.regf_0.rf[14][10] ;
 wire \po_0.regf_0.rf[14][11] ;
 wire \po_0.regf_0.rf[14][12] ;
 wire \po_0.regf_0.rf[14][13] ;
 wire \po_0.regf_0.rf[14][14] ;
 wire \po_0.regf_0.rf[14][15] ;
 wire \po_0.regf_0.rf[14][1] ;
 wire \po_0.regf_0.rf[14][2] ;
 wire \po_0.regf_0.rf[14][3] ;
 wire \po_0.regf_0.rf[14][4] ;
 wire \po_0.regf_0.rf[14][5] ;
 wire \po_0.regf_0.rf[14][6] ;
 wire \po_0.regf_0.rf[14][7] ;
 wire \po_0.regf_0.rf[14][8] ;
 wire \po_0.regf_0.rf[14][9] ;
 wire \po_0.regf_0.rf[15][0] ;
 wire \po_0.regf_0.rf[15][10] ;
 wire \po_0.regf_0.rf[15][11] ;
 wire \po_0.regf_0.rf[15][12] ;
 wire \po_0.regf_0.rf[15][13] ;
 wire \po_0.regf_0.rf[15][14] ;
 wire \po_0.regf_0.rf[15][15] ;
 wire \po_0.regf_0.rf[15][1] ;
 wire \po_0.regf_0.rf[15][2] ;
 wire \po_0.regf_0.rf[15][3] ;
 wire \po_0.regf_0.rf[15][4] ;
 wire \po_0.regf_0.rf[15][5] ;
 wire \po_0.regf_0.rf[15][6] ;
 wire \po_0.regf_0.rf[15][7] ;
 wire \po_0.regf_0.rf[15][8] ;
 wire \po_0.regf_0.rf[15][9] ;
 wire \po_0.regf_0.rf[1][0] ;
 wire \po_0.regf_0.rf[1][10] ;
 wire \po_0.regf_0.rf[1][11] ;
 wire \po_0.regf_0.rf[1][12] ;
 wire \po_0.regf_0.rf[1][13] ;
 wire \po_0.regf_0.rf[1][14] ;
 wire \po_0.regf_0.rf[1][15] ;
 wire \po_0.regf_0.rf[1][1] ;
 wire \po_0.regf_0.rf[1][2] ;
 wire \po_0.regf_0.rf[1][3] ;
 wire \po_0.regf_0.rf[1][4] ;
 wire \po_0.regf_0.rf[1][5] ;
 wire \po_0.regf_0.rf[1][6] ;
 wire \po_0.regf_0.rf[1][7] ;
 wire \po_0.regf_0.rf[1][8] ;
 wire \po_0.regf_0.rf[1][9] ;
 wire \po_0.regf_0.rf[2][0] ;
 wire \po_0.regf_0.rf[2][10] ;
 wire \po_0.regf_0.rf[2][11] ;
 wire \po_0.regf_0.rf[2][12] ;
 wire \po_0.regf_0.rf[2][13] ;
 wire \po_0.regf_0.rf[2][14] ;
 wire \po_0.regf_0.rf[2][15] ;
 wire \po_0.regf_0.rf[2][1] ;
 wire \po_0.regf_0.rf[2][2] ;
 wire \po_0.regf_0.rf[2][3] ;
 wire \po_0.regf_0.rf[2][4] ;
 wire \po_0.regf_0.rf[2][5] ;
 wire \po_0.regf_0.rf[2][6] ;
 wire \po_0.regf_0.rf[2][7] ;
 wire \po_0.regf_0.rf[2][8] ;
 wire \po_0.regf_0.rf[2][9] ;
 wire \po_0.regf_0.rf[3][0] ;
 wire \po_0.regf_0.rf[3][10] ;
 wire \po_0.regf_0.rf[3][11] ;
 wire \po_0.regf_0.rf[3][12] ;
 wire \po_0.regf_0.rf[3][13] ;
 wire \po_0.regf_0.rf[3][14] ;
 wire \po_0.regf_0.rf[3][15] ;
 wire \po_0.regf_0.rf[3][1] ;
 wire \po_0.regf_0.rf[3][2] ;
 wire \po_0.regf_0.rf[3][3] ;
 wire \po_0.regf_0.rf[3][4] ;
 wire \po_0.regf_0.rf[3][5] ;
 wire \po_0.regf_0.rf[3][6] ;
 wire \po_0.regf_0.rf[3][7] ;
 wire \po_0.regf_0.rf[3][8] ;
 wire \po_0.regf_0.rf[3][9] ;
 wire \po_0.regf_0.rf[4][0] ;
 wire \po_0.regf_0.rf[4][10] ;
 wire \po_0.regf_0.rf[4][11] ;
 wire \po_0.regf_0.rf[4][12] ;
 wire \po_0.regf_0.rf[4][13] ;
 wire \po_0.regf_0.rf[4][14] ;
 wire \po_0.regf_0.rf[4][15] ;
 wire \po_0.regf_0.rf[4][1] ;
 wire \po_0.regf_0.rf[4][2] ;
 wire \po_0.regf_0.rf[4][3] ;
 wire \po_0.regf_0.rf[4][4] ;
 wire \po_0.regf_0.rf[4][5] ;
 wire \po_0.regf_0.rf[4][6] ;
 wire \po_0.regf_0.rf[4][7] ;
 wire \po_0.regf_0.rf[4][8] ;
 wire \po_0.regf_0.rf[4][9] ;
 wire \po_0.regf_0.rf[5][0] ;
 wire \po_0.regf_0.rf[5][10] ;
 wire \po_0.regf_0.rf[5][11] ;
 wire \po_0.regf_0.rf[5][12] ;
 wire \po_0.regf_0.rf[5][13] ;
 wire \po_0.regf_0.rf[5][14] ;
 wire \po_0.regf_0.rf[5][15] ;
 wire \po_0.regf_0.rf[5][1] ;
 wire \po_0.regf_0.rf[5][2] ;
 wire \po_0.regf_0.rf[5][3] ;
 wire \po_0.regf_0.rf[5][4] ;
 wire \po_0.regf_0.rf[5][5] ;
 wire \po_0.regf_0.rf[5][6] ;
 wire \po_0.regf_0.rf[5][7] ;
 wire \po_0.regf_0.rf[5][8] ;
 wire \po_0.regf_0.rf[5][9] ;
 wire \po_0.regf_0.rf[6][0] ;
 wire \po_0.regf_0.rf[6][10] ;
 wire \po_0.regf_0.rf[6][11] ;
 wire \po_0.regf_0.rf[6][12] ;
 wire \po_0.regf_0.rf[6][13] ;
 wire \po_0.regf_0.rf[6][14] ;
 wire \po_0.regf_0.rf[6][15] ;
 wire \po_0.regf_0.rf[6][1] ;
 wire \po_0.regf_0.rf[6][2] ;
 wire \po_0.regf_0.rf[6][3] ;
 wire \po_0.regf_0.rf[6][4] ;
 wire \po_0.regf_0.rf[6][5] ;
 wire \po_0.regf_0.rf[6][6] ;
 wire \po_0.regf_0.rf[6][7] ;
 wire \po_0.regf_0.rf[6][8] ;
 wire \po_0.regf_0.rf[6][9] ;
 wire \po_0.regf_0.rf[7][0] ;
 wire \po_0.regf_0.rf[7][10] ;
 wire \po_0.regf_0.rf[7][11] ;
 wire \po_0.regf_0.rf[7][12] ;
 wire \po_0.regf_0.rf[7][13] ;
 wire \po_0.regf_0.rf[7][14] ;
 wire \po_0.regf_0.rf[7][15] ;
 wire \po_0.regf_0.rf[7][1] ;
 wire \po_0.regf_0.rf[7][2] ;
 wire \po_0.regf_0.rf[7][3] ;
 wire \po_0.regf_0.rf[7][4] ;
 wire \po_0.regf_0.rf[7][5] ;
 wire \po_0.regf_0.rf[7][6] ;
 wire \po_0.regf_0.rf[7][7] ;
 wire \po_0.regf_0.rf[7][8] ;
 wire \po_0.regf_0.rf[7][9] ;
 wire \po_0.regf_0.rf[8][0] ;
 wire \po_0.regf_0.rf[8][10] ;
 wire \po_0.regf_0.rf[8][11] ;
 wire \po_0.regf_0.rf[8][12] ;
 wire \po_0.regf_0.rf[8][13] ;
 wire \po_0.regf_0.rf[8][14] ;
 wire \po_0.regf_0.rf[8][15] ;
 wire \po_0.regf_0.rf[8][1] ;
 wire \po_0.regf_0.rf[8][2] ;
 wire \po_0.regf_0.rf[8][3] ;
 wire \po_0.regf_0.rf[8][4] ;
 wire \po_0.regf_0.rf[8][5] ;
 wire \po_0.regf_0.rf[8][6] ;
 wire \po_0.regf_0.rf[8][7] ;
 wire \po_0.regf_0.rf[8][8] ;
 wire \po_0.regf_0.rf[8][9] ;
 wire \po_0.regf_0.rf[9][0] ;
 wire \po_0.regf_0.rf[9][10] ;
 wire \po_0.regf_0.rf[9][11] ;
 wire \po_0.regf_0.rf[9][12] ;
 wire \po_0.regf_0.rf[9][13] ;
 wire \po_0.regf_0.rf[9][14] ;
 wire \po_0.regf_0.rf[9][15] ;
 wire \po_0.regf_0.rf[9][1] ;
 wire \po_0.regf_0.rf[9][2] ;
 wire \po_0.regf_0.rf[9][3] ;
 wire \po_0.regf_0.rf[9][4] ;
 wire \po_0.regf_0.rf[9][5] ;
 wire \po_0.regf_0.rf[9][6] ;
 wire \po_0.regf_0.rf[9][7] ;
 wire \po_0.regf_0.rf[9][8] ;
 wire \po_0.regf_0.rf[9][9] ;
 wire \po_0.regf_0.rp_addr[0] ;
 wire \po_0.regf_0.rp_addr[1] ;
 wire \po_0.regf_0.rp_addr[2] ;
 wire \po_0.regf_0.rp_addr[3] ;
 wire \po_0.regf_0.rp_rd ;
 wire \po_0.regf_0.rq_addr[0] ;
 wire \po_0.regf_0.rq_addr[1] ;
 wire \po_0.regf_0.rq_addr[2] ;
 wire \po_0.regf_0.rq_addr[3] ;
 wire \po_0.regf_0.rq_rd ;
 wire \po_0.regf_0.w_addr[0] ;
 wire \po_0.regf_0.w_addr[1] ;
 wire \po_0.regf_0.w_addr[2] ;
 wire \po_0.regf_0.w_addr[3] ;
 wire \po_0.regf_0.w_wr ;
 wire \uc_0._00_ ;
 wire \uc_0._01_ ;
 wire \uc_0._02_ ;
 wire \uc_0._03_ ;
 wire \uc_0._20_[10] ;
 wire \uc_0._20_[11] ;
 wire \uc_0._20_[8] ;
 wire \uc_0._20_[9] ;
 wire \uc_0.bc_0._54_[0] ;
 wire \uc_0.bc_0._54_[1] ;
 wire \uc_0.bc_0._54_[2] ;
 wire \uc_0.bc_0._54_[3] ;
 wire \uc_0.bc_0._55_[0] ;
 wire \uc_0.bc_0._55_[1] ;
 wire \uc_0.bc_0._55_[2] ;
 wire \uc_0.bc_0._55_[3] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0423_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\po_0.regf_0._5_[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net39));
 sky130_fd_sc_hd__fill_1 FILLER_0_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_82 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__clkbuf_2 _1574_ (.A(\po_0.alu_0.s0 ),
    .X(_1401_));
 sky130_fd_sc_hd__clkbuf_2 _1575_ (.A(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__clkbuf_2 _1576_ (.A(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_2 _1577_ (.A(\po_0.alu_0.s1 ),
    .X(_1404_));
 sky130_fd_sc_hd__clkbuf_2 _1578_ (.A(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_2 _1579_ (.A(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1580_ (.A(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__or2b_1 _1581_ (.A(_1403_),
    .B_N(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _1582_ (.A(_1408_),
    .X(_1565_));
 sky130_fd_sc_hd__or2b_1 _1583_ (.A(_1403_),
    .B_N(_1407_),
    .X(_1409_));
 sky130_fd_sc_hd__clkbuf_1 _1584_ (.A(_1409_),
    .X(_1564_));
 sky130_fd_sc_hd__or2b_1 _1585_ (.A(_1403_),
    .B_N(_1407_),
    .X(_1410_));
 sky130_fd_sc_hd__clkbuf_1 _1586_ (.A(_1410_),
    .X(_1563_));
 sky130_fd_sc_hd__or2b_1 _1587_ (.A(_1403_),
    .B_N(_1407_),
    .X(_1411_));
 sky130_fd_sc_hd__clkbuf_1 _1588_ (.A(_1411_),
    .X(_1562_));
 sky130_fd_sc_hd__or2b_1 _1589_ (.A(_1403_),
    .B_N(_1407_),
    .X(_1412_));
 sky130_fd_sc_hd__clkbuf_1 _1590_ (.A(_1412_),
    .X(_1561_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1591_ (.A(_1402_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_2 _1592_ (.A(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _1593_ (.A(_1406_),
    .X(_1415_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1594_ (.A(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__or2b_1 _1595_ (.A(_1414_),
    .B_N(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__clkbuf_1 _1596_ (.A(_1417_),
    .X(_1560_));
 sky130_fd_sc_hd__or2b_1 _1597_ (.A(_1414_),
    .B_N(_1416_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _1598_ (.A(_1418_),
    .X(_1559_));
 sky130_fd_sc_hd__or2b_1 _1599_ (.A(_1414_),
    .B_N(_1416_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_1 _1600_ (.A(_1419_),
    .X(_1558_));
 sky130_fd_sc_hd__or2b_1 _1601_ (.A(_1414_),
    .B_N(_1416_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _1602_ (.A(_1420_),
    .X(_1566_));
 sky130_fd_sc_hd__or2b_1 _1603_ (.A(_1414_),
    .B_N(_1416_),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_1 _1604_ (.A(_1421_),
    .X(_1567_));
 sky130_fd_sc_hd__or2b_1 _1605_ (.A(_1414_),
    .B_N(_1416_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_1 _1606_ (.A(_1422_),
    .X(_1568_));
 sky130_fd_sc_hd__or2b_1 _1607_ (.A(_1413_),
    .B_N(_1415_),
    .X(_1423_));
 sky130_fd_sc_hd__clkbuf_1 _1608_ (.A(_1423_),
    .X(_1569_));
 sky130_fd_sc_hd__or2b_1 _1609_ (.A(_1413_),
    .B_N(_1415_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_1 _1610_ (.A(_1424_),
    .X(_1570_));
 sky130_fd_sc_hd__or2b_1 _1611_ (.A(_1413_),
    .B_N(_1415_),
    .X(_1425_));
 sky130_fd_sc_hd__clkbuf_1 _1612_ (.A(_1425_),
    .X(_1571_));
 sky130_fd_sc_hd__or2b_1 _1613_ (.A(_1413_),
    .B_N(_1415_),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_1 _1614_ (.A(_1426_),
    .X(_1572_));
 sky130_fd_sc_hd__or2b_1 _1615_ (.A(_1413_),
    .B_N(_1415_),
    .X(_1427_));
 sky130_fd_sc_hd__clkbuf_1 _1616_ (.A(_1427_),
    .X(_1573_));
 sky130_fd_sc_hd__or2_1 _1617_ (.A(\po_0._1_[0] ),
    .B(net87),
    .X(_1428_));
 sky130_fd_sc_hd__nand2_1 _1618_ (.A(\po_0._1_[0] ),
    .B(net87),
    .Y(_1429_));
 sky130_fd_sc_hd__and2_1 _1619_ (.A(_1428_),
    .B(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__clkbuf_1 _1620_ (.A(_1430_),
    .X(\po_0.alu_0._10_[0] ));
 sky130_fd_sc_hd__or3b_1 _1621_ (.A(net82),
    .B(net81),
    .C_N(net80),
    .X(_1431_));
 sky130_fd_sc_hd__a311oi_2 _1622_ (.A1(_1431_),
    .A2(\uc_0.bc_0._55_[1] ),
    .A3(\uc_0.bc_0._55_[0] ),
    .B1(\uc_0.bc_0._55_[2] ),
    .C1(\uc_0.bc_0._55_[3] ),
    .Y(_1432_));
 sky130_fd_sc_hd__and4bb_1 _1623_ (.A_N(\uc_0.bc_0._55_[1] ),
    .B_N(\uc_0.bc_0._55_[2] ),
    .C(\uc_0.bc_0._55_[3] ),
    .D(\uc_0.bc_0._55_[0] ),
    .X(_1433_));
 sky130_fd_sc_hd__nor4_1 _1624_ (.A(net39),
    .B(net83),
    .C(net41),
    .D(net40),
    .Y(_1434_));
 sky130_fd_sc_hd__nor4_1 _1625_ (.A(net50),
    .B(net49),
    .C(net84),
    .D(net36),
    .Y(_1435_));
 sky130_fd_sc_hd__nand3_1 _1626_ (.A(_1433_),
    .B(_1434_),
    .C(_1435_),
    .Y(_1436_));
 sky130_fd_sc_hd__or4_2 _1627_ (.A(net87),
    .B(net86),
    .C(net44),
    .D(net43),
    .X(_1437_));
 sky130_fd_sc_hd__or4_2 _1628_ (.A(net46),
    .B(net45),
    .C(net85),
    .D(net47),
    .X(_1438_));
 sky130_fd_sc_hd__nor3_2 _1629_ (.A(_1436_),
    .B(_1437_),
    .C(_1438_),
    .Y(_1439_));
 sky130_fd_sc_hd__clkbuf_2 _1630_ (.A(net34),
    .X(_1440_));
 sky130_fd_sc_hd__o21bai_2 _1631_ (.A1(_1432_),
    .A2(_1439_),
    .B1_N(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__inv_2 _1632_ (.A(_1441_),
    .Y(\uc_0.bc_0._54_[1] ));
 sky130_fd_sc_hd__inv_2 _1633_ (.A(\uc_0.bc_0._55_[0] ),
    .Y(_1442_));
 sky130_fd_sc_hd__a2111o_1 _1634_ (.A1(net80),
    .A2(net81),
    .B1(net82),
    .C1(net79),
    .D1(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__a211oi_1 _1635_ (.A1(_1443_),
    .A2(\uc_0.bc_0._55_[1] ),
    .B1(\uc_0.bc_0._55_[2] ),
    .C1(\uc_0.bc_0._55_[3] ),
    .Y(_1444_));
 sky130_fd_sc_hd__nor2_1 _1636_ (.A(net34),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__o31ai_2 _1637_ (.A1(_1436_),
    .A2(_1437_),
    .A3(_1438_),
    .B1(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__inv_2 _1638_ (.A(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__buf_2 _1639_ (.A(_1447_),
    .X(\uc_0.bc_0._54_[0] ));
 sky130_fd_sc_hd__and4bb_1 _1640_ (.A_N(\uc_0.bc_0._55_[2] ),
    .B_N(\uc_0.bc_0._55_[3] ),
    .C(\uc_0.bc_0._55_[0] ),
    .D(\uc_0.bc_0._55_[1] ),
    .X(_1448_));
 sky130_fd_sc_hd__and4bb_1 _1641_ (.A_N(net80),
    .B_N(net82),
    .C(net81),
    .D(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__o21ba_1 _1642_ (.A1(_1439_),
    .A2(_1449_),
    .B1_N(_1440_),
    .X(_1450_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1643_ (.A(_1450_),
    .X(\uc_0.bc_0._54_[3] ));
 sky130_fd_sc_hd__or3b_1 _1644_ (.A(net82),
    .B(net81),
    .C_N(_1448_),
    .X(_1451_));
 sky130_fd_sc_hd__nor2_1 _1645_ (.A(_1440_),
    .B(_1451_),
    .Y(\uc_0.bc_0._54_[2] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1646_ (.A(_0006_),
    .X(_1452_));
 sky130_fd_sc_hd__clkbuf_2 _1647_ (.A(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__clkbuf_2 _1648_ (.A(_0004_),
    .X(_1454_));
 sky130_fd_sc_hd__clkbuf_4 _1649_ (.A(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1650_ (.A(_0005_),
    .X(_1456_));
 sky130_fd_sc_hd__buf_2 _1651_ (.A(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__mux4_1 _1652_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(\po_0.regf_0.rf[9][0] ),
    .A2(\po_0.regf_0.rf[10][0] ),
    .A3(\po_0.regf_0.rf[11][0] ),
    .S0(_1455_),
    .S1(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__and2b_1 _1653_ (.A_N(_1453_),
    .B(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__clkbuf_4 _1654_ (.A(_0004_),
    .X(_1460_));
 sky130_fd_sc_hd__clkbuf_4 _1655_ (.A(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__buf_2 _1656_ (.A(_0005_),
    .X(_1462_));
 sky130_fd_sc_hd__clkbuf_4 _1657_ (.A(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__mux4_1 _1658_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(\po_0.regf_0.rf[13][0] ),
    .A2(\po_0.regf_0.rf[14][0] ),
    .A3(\po_0.regf_0.rf[15][0] ),
    .S0(_1461_),
    .S1(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__buf_2 _1659_ (.A(_0006_),
    .X(_1465_));
 sky130_fd_sc_hd__buf_2 _1660_ (.A(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__clkbuf_2 _1661_ (.A(_0007_),
    .X(_1467_));
 sky130_fd_sc_hd__buf_2 _1662_ (.A(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__a21bo_1 _1663_ (.A1(_1464_),
    .A2(_1466_),
    .B1_N(_1468_),
    .X(_1469_));
 sky130_fd_sc_hd__buf_2 _1664_ (.A(_1452_),
    .X(_1470_));
 sky130_fd_sc_hd__clkbuf_4 _1665_ (.A(_1454_),
    .X(_1471_));
 sky130_fd_sc_hd__clkbuf_4 _1666_ (.A(_1456_),
    .X(_1472_));
 sky130_fd_sc_hd__mux4_1 _1667_ (.A0(\po_0.regf_0.rf[0][0] ),
    .A1(\po_0.regf_0.rf[1][0] ),
    .A2(\po_0.regf_0.rf[2][0] ),
    .A3(\po_0.regf_0.rf[3][0] ),
    .S0(_1471_),
    .S1(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__and2b_1 _1668_ (.A_N(_1470_),
    .B(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__clkbuf_4 _1669_ (.A(_1460_),
    .X(_1475_));
 sky130_fd_sc_hd__buf_2 _1670_ (.A(_1462_),
    .X(_1476_));
 sky130_fd_sc_hd__mux4_1 _1671_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(\po_0.regf_0.rf[5][0] ),
    .A2(\po_0.regf_0.rf[6][0] ),
    .A3(\po_0.regf_0.rf[7][0] ),
    .S0(_1475_),
    .S1(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__buf_2 _1672_ (.A(_1465_),
    .X(_1478_));
 sky130_fd_sc_hd__buf_2 _1673_ (.A(_1467_),
    .X(_1479_));
 sky130_fd_sc_hd__a21o_1 _1674_ (.A1(_1477_),
    .A2(_1478_),
    .B1(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__o22a_1 _1675_ (.A1(_1459_),
    .A2(_1469_),
    .B1(_1474_),
    .B2(_1480_),
    .X(\po_0.regf_0._5_[0] ));
 sky130_fd_sc_hd__clkbuf_4 _1676_ (.A(_1454_),
    .X(_1481_));
 sky130_fd_sc_hd__buf_2 _1677_ (.A(_1456_),
    .X(_1482_));
 sky130_fd_sc_hd__mux4_1 _1678_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(\po_0.regf_0.rf[13][1] ),
    .A2(\po_0.regf_0.rf[14][1] ),
    .A3(\po_0.regf_0.rf[15][1] ),
    .S0(_1481_),
    .S1(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__buf_2 _1679_ (.A(_1452_),
    .X(_1484_));
 sky130_fd_sc_hd__clkbuf_2 _1680_ (.A(_1467_),
    .X(_1485_));
 sky130_fd_sc_hd__a21bo_1 _1681_ (.A1(_1483_),
    .A2(_1484_),
    .B1_N(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_2 _1682_ (.A(_1452_),
    .X(_1487_));
 sky130_fd_sc_hd__clkbuf_4 _1683_ (.A(_1454_),
    .X(_1488_));
 sky130_fd_sc_hd__buf_2 _1684_ (.A(_1456_),
    .X(_1489_));
 sky130_fd_sc_hd__mux4_1 _1685_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(\po_0.regf_0.rf[9][1] ),
    .A2(\po_0.regf_0.rf[10][1] ),
    .A3(\po_0.regf_0.rf[11][1] ),
    .S0(_1488_),
    .S1(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__and2b_1 _1686_ (.A_N(_1487_),
    .B(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__clkbuf_2 _1687_ (.A(_0007_),
    .X(_1492_));
 sky130_fd_sc_hd__buf_2 _1688_ (.A(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__clkbuf_4 _1689_ (.A(_0004_),
    .X(_1494_));
 sky130_fd_sc_hd__buf_2 _1690_ (.A(_0005_),
    .X(_1495_));
 sky130_fd_sc_hd__mux4_1 _1691_ (.A0(\po_0.regf_0.rf[0][1] ),
    .A1(\po_0.regf_0.rf[1][1] ),
    .A2(\po_0.regf_0.rf[2][1] ),
    .A3(\po_0.regf_0.rf[3][1] ),
    .S0(_1494_),
    .S1(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__clkbuf_4 _1692_ (.A(_0004_),
    .X(_1497_));
 sky130_fd_sc_hd__buf_2 _1693_ (.A(_0005_),
    .X(_1498_));
 sky130_fd_sc_hd__mux4_1 _1694_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(\po_0.regf_0.rf[5][1] ),
    .A2(\po_0.regf_0.rf[6][1] ),
    .A3(\po_0.regf_0.rf[7][1] ),
    .S0(_1497_),
    .S1(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__buf_2 _1695_ (.A(_1452_),
    .X(_1500_));
 sky130_fd_sc_hd__mux2_1 _1696_ (.A0(_1496_),
    .A1(_1499_),
    .S(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__o22a_1 _1697_ (.A1(_1486_),
    .A2(_1491_),
    .B1(_1493_),
    .B2(_1501_),
    .X(\po_0.regf_0._5_[1] ));
 sky130_fd_sc_hd__mux4_1 _1698_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(\po_0.regf_0.rf[13][2] ),
    .A2(\po_0.regf_0.rf[14][2] ),
    .A3(\po_0.regf_0.rf[15][2] ),
    .S0(_1481_),
    .S1(_1482_),
    .X(_1502_));
 sky130_fd_sc_hd__a21bo_1 _1699_ (.A1(_1502_),
    .A2(_1484_),
    .B1_N(_1485_),
    .X(_1503_));
 sky130_fd_sc_hd__mux4_1 _1700_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(\po_0.regf_0.rf[9][2] ),
    .A2(\po_0.regf_0.rf[10][2] ),
    .A3(\po_0.regf_0.rf[11][2] ),
    .S0(_1488_),
    .S1(_1489_),
    .X(_1504_));
 sky130_fd_sc_hd__and2b_1 _1701_ (.A_N(_1487_),
    .B(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__mux4_1 _1702_ (.A0(\po_0.regf_0.rf[0][2] ),
    .A1(\po_0.regf_0.rf[1][2] ),
    .A2(\po_0.regf_0.rf[2][2] ),
    .A3(\po_0.regf_0.rf[3][2] ),
    .S0(_1494_),
    .S1(_1495_),
    .X(_1506_));
 sky130_fd_sc_hd__mux4_1 _1703_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(\po_0.regf_0.rf[5][2] ),
    .A2(\po_0.regf_0.rf[6][2] ),
    .A3(\po_0.regf_0.rf[7][2] ),
    .S0(_1497_),
    .S1(_1498_),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _1704_ (.A0(_1506_),
    .A1(_1507_),
    .S(_1500_),
    .X(_1508_));
 sky130_fd_sc_hd__o22a_1 _1705_ (.A1(_1503_),
    .A2(_1505_),
    .B1(_1493_),
    .B2(_1508_),
    .X(\po_0.regf_0._5_[2] ));
 sky130_fd_sc_hd__mux4_1 _1706_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(\po_0.regf_0.rf[13][3] ),
    .A2(\po_0.regf_0.rf[14][3] ),
    .A3(\po_0.regf_0.rf[15][3] ),
    .S0(_1481_),
    .S1(_1482_),
    .X(_1509_));
 sky130_fd_sc_hd__a21bo_1 _1707_ (.A1(_1509_),
    .A2(_1470_),
    .B1_N(_1485_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_2 _1708_ (.A(_1452_),
    .X(_1511_));
 sky130_fd_sc_hd__clkbuf_4 _1709_ (.A(_1454_),
    .X(_1512_));
 sky130_fd_sc_hd__buf_2 _1710_ (.A(_1456_),
    .X(_1513_));
 sky130_fd_sc_hd__mux4_1 _1711_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(\po_0.regf_0.rf[9][3] ),
    .A2(\po_0.regf_0.rf[10][3] ),
    .A3(\po_0.regf_0.rf[11][3] ),
    .S0(_1512_),
    .S1(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__and2b_1 _1712_ (.A_N(_1511_),
    .B(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__mux4_1 _1713_ (.A0(\po_0.regf_0.rf[0][3] ),
    .A1(\po_0.regf_0.rf[1][3] ),
    .A2(\po_0.regf_0.rf[2][3] ),
    .A3(\po_0.regf_0.rf[3][3] ),
    .S0(_1494_),
    .S1(_1495_),
    .X(_1516_));
 sky130_fd_sc_hd__mux4_1 _1714_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(\po_0.regf_0.rf[5][3] ),
    .A2(\po_0.regf_0.rf[6][3] ),
    .A3(\po_0.regf_0.rf[7][3] ),
    .S0(_1497_),
    .S1(_1498_),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_1 _1715_ (.A0(_1516_),
    .A1(_1517_),
    .S(_1500_),
    .X(_1518_));
 sky130_fd_sc_hd__o22a_1 _1716_ (.A1(_1510_),
    .A2(_1515_),
    .B1(_1493_),
    .B2(_1518_),
    .X(\po_0.regf_0._5_[3] ));
 sky130_fd_sc_hd__mux4_1 _1717_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(\po_0.regf_0.rf[9][4] ),
    .A2(\po_0.regf_0.rf[10][4] ),
    .A3(\po_0.regf_0.rf[11][4] ),
    .S0(_1455_),
    .S1(_1457_),
    .X(_1519_));
 sky130_fd_sc_hd__and2b_1 _1718_ (.A_N(_1453_),
    .B(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__mux4_1 _1719_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(\po_0.regf_0.rf[13][4] ),
    .A2(\po_0.regf_0.rf[14][4] ),
    .A3(\po_0.regf_0.rf[15][4] ),
    .S0(_1461_),
    .S1(_1463_),
    .X(_1521_));
 sky130_fd_sc_hd__a21bo_1 _1720_ (.A1(_1521_),
    .A2(_1466_),
    .B1_N(_1468_),
    .X(_1522_));
 sky130_fd_sc_hd__mux4_1 _1721_ (.A0(\po_0.regf_0.rf[0][4] ),
    .A1(\po_0.regf_0.rf[1][4] ),
    .A2(\po_0.regf_0.rf[2][4] ),
    .A3(\po_0.regf_0.rf[3][4] ),
    .S0(_1488_),
    .S1(_1489_),
    .X(_1523_));
 sky130_fd_sc_hd__and2b_1 _1722_ (.A_N(_1487_),
    .B(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__mux4_1 _1723_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(\po_0.regf_0.rf[5][4] ),
    .A2(\po_0.regf_0.rf[6][4] ),
    .A3(\po_0.regf_0.rf[7][4] ),
    .S0(_1475_),
    .S1(_1476_),
    .X(_1525_));
 sky130_fd_sc_hd__a21o_1 _1724_ (.A1(_1525_),
    .A2(_1478_),
    .B1(_1479_),
    .X(_1526_));
 sky130_fd_sc_hd__o22a_1 _1725_ (.A1(_1520_),
    .A2(_1522_),
    .B1(_1524_),
    .B2(_1526_),
    .X(\po_0.regf_0._5_[4] ));
 sky130_fd_sc_hd__mux4_1 _1726_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(\po_0.regf_0.rf[9][5] ),
    .A2(\po_0.regf_0.rf[10][5] ),
    .A3(\po_0.regf_0.rf[11][5] ),
    .S0(_1455_),
    .S1(_1457_),
    .X(_1527_));
 sky130_fd_sc_hd__and2b_1 _1727_ (.A_N(_1453_),
    .B(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__mux4_1 _1728_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(\po_0.regf_0.rf[13][5] ),
    .A2(\po_0.regf_0.rf[14][5] ),
    .A3(\po_0.regf_0.rf[15][5] ),
    .S0(_1461_),
    .S1(_1463_),
    .X(_1529_));
 sky130_fd_sc_hd__a21bo_1 _1729_ (.A1(_1529_),
    .A2(_1466_),
    .B1_N(_1468_),
    .X(_1530_));
 sky130_fd_sc_hd__mux4_1 _1730_ (.A0(\po_0.regf_0.rf[0][5] ),
    .A1(\po_0.regf_0.rf[1][5] ),
    .A2(\po_0.regf_0.rf[2][5] ),
    .A3(\po_0.regf_0.rf[3][5] ),
    .S0(_1488_),
    .S1(_1489_),
    .X(_1531_));
 sky130_fd_sc_hd__and2b_1 _1731_ (.A_N(_1487_),
    .B(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__mux4_1 _1732_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(\po_0.regf_0.rf[5][5] ),
    .A2(\po_0.regf_0.rf[6][5] ),
    .A3(\po_0.regf_0.rf[7][5] ),
    .S0(_1475_),
    .S1(_1476_),
    .X(_1533_));
 sky130_fd_sc_hd__a21o_1 _1733_ (.A1(_1533_),
    .A2(_1478_),
    .B1(_1479_),
    .X(_1534_));
 sky130_fd_sc_hd__o22a_1 _1734_ (.A1(_1528_),
    .A2(_1530_),
    .B1(_1532_),
    .B2(_1534_),
    .X(\po_0.regf_0._5_[5] ));
 sky130_fd_sc_hd__mux4_1 _1735_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(\po_0.regf_0.rf[13][6] ),
    .A2(\po_0.regf_0.rf[14][6] ),
    .A3(\po_0.regf_0.rf[15][6] ),
    .S0(_1481_),
    .S1(_1482_),
    .X(_1535_));
 sky130_fd_sc_hd__a21bo_1 _1736_ (.A1(_1535_),
    .A2(_1470_),
    .B1_N(_1485_),
    .X(_1536_));
 sky130_fd_sc_hd__mux4_1 _1737_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(\po_0.regf_0.rf[9][6] ),
    .A2(\po_0.regf_0.rf[10][6] ),
    .A3(\po_0.regf_0.rf[11][6] ),
    .S0(_1512_),
    .S1(_1513_),
    .X(_1537_));
 sky130_fd_sc_hd__and2b_1 _1738_ (.A_N(_1511_),
    .B(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__mux4_1 _1739_ (.A0(\po_0.regf_0.rf[0][6] ),
    .A1(\po_0.regf_0.rf[1][6] ),
    .A2(\po_0.regf_0.rf[2][6] ),
    .A3(\po_0.regf_0.rf[3][6] ),
    .S0(_1494_),
    .S1(_1495_),
    .X(_1539_));
 sky130_fd_sc_hd__mux4_1 _1740_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(\po_0.regf_0.rf[5][6] ),
    .A2(\po_0.regf_0.rf[6][6] ),
    .A3(\po_0.regf_0.rf[7][6] ),
    .S0(_1460_),
    .S1(_1462_),
    .X(_1540_));
 sky130_fd_sc_hd__mux2_1 _1741_ (.A0(_1539_),
    .A1(_1540_),
    .S(_1500_),
    .X(_1541_));
 sky130_fd_sc_hd__o22a_1 _1742_ (.A1(_1536_),
    .A2(_1538_),
    .B1(_1493_),
    .B2(_1541_),
    .X(\po_0.regf_0._5_[6] ));
 sky130_fd_sc_hd__clkbuf_4 _1743_ (.A(_1454_),
    .X(_1542_));
 sky130_fd_sc_hd__buf_2 _1744_ (.A(_1456_),
    .X(_1543_));
 sky130_fd_sc_hd__mux4_1 _1745_ (.A0(\po_0.regf_0.rf[4][7] ),
    .A1(\po_0.regf_0.rf[5][7] ),
    .A2(\po_0.regf_0.rf[6][7] ),
    .A3(\po_0.regf_0.rf[7][7] ),
    .S0(_1542_),
    .S1(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__a21o_1 _1746_ (.A1(_1544_),
    .A2(_1484_),
    .B1(_1492_),
    .X(_1545_));
 sky130_fd_sc_hd__mux4_1 _1747_ (.A0(\po_0.regf_0.rf[0][7] ),
    .A1(\po_0.regf_0.rf[1][7] ),
    .A2(\po_0.regf_0.rf[2][7] ),
    .A3(\po_0.regf_0.rf[3][7] ),
    .S0(_1512_),
    .S1(_1513_),
    .X(_1546_));
 sky130_fd_sc_hd__and2b_1 _1748_ (.A_N(_1511_),
    .B(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__mux4_1 _1749_ (.A0(\po_0.regf_0.rf[12][7] ),
    .A1(\po_0.regf_0.rf[13][7] ),
    .A2(\po_0.regf_0.rf[14][7] ),
    .A3(\po_0.regf_0.rf[15][7] ),
    .S0(_1475_),
    .S1(_1476_),
    .X(_1548_));
 sky130_fd_sc_hd__a21bo_1 _1750_ (.A1(_1548_),
    .A2(_1478_),
    .B1_N(_1492_),
    .X(_1549_));
 sky130_fd_sc_hd__clkbuf_2 _1751_ (.A(_1465_),
    .X(_1550_));
 sky130_fd_sc_hd__mux4_1 _1752_ (.A0(\po_0.regf_0.rf[8][7] ),
    .A1(\po_0.regf_0.rf[9][7] ),
    .A2(\po_0.regf_0.rf[10][7] ),
    .A3(\po_0.regf_0.rf[11][7] ),
    .S0(_1471_),
    .S1(_1472_),
    .X(_1551_));
 sky130_fd_sc_hd__and2b_1 _1753_ (.A_N(_1550_),
    .B(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__o22a_1 _1754_ (.A1(_1545_),
    .A2(_1547_),
    .B1(_1549_),
    .B2(_1552_),
    .X(\po_0.regf_0._5_[7] ));
 sky130_fd_sc_hd__mux4_1 _1755_ (.A0(\po_0.regf_0.rf[4][8] ),
    .A1(\po_0.regf_0.rf[5][8] ),
    .A2(\po_0.regf_0.rf[6][8] ),
    .A3(\po_0.regf_0.rf[7][8] ),
    .S0(_1542_),
    .S1(_1543_),
    .X(_1553_));
 sky130_fd_sc_hd__a21o_1 _1756_ (.A1(_1553_),
    .A2(_1484_),
    .B1(_1492_),
    .X(_1554_));
 sky130_fd_sc_hd__mux4_1 _1757_ (.A0(\po_0.regf_0.rf[0][8] ),
    .A1(\po_0.regf_0.rf[1][8] ),
    .A2(\po_0.regf_0.rf[2][8] ),
    .A3(\po_0.regf_0.rf[3][8] ),
    .S0(_1512_),
    .S1(_1513_),
    .X(_1555_));
 sky130_fd_sc_hd__and2b_1 _1758_ (.A_N(_1511_),
    .B(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__mux4_1 _1759_ (.A0(\po_0.regf_0.rf[12][8] ),
    .A1(\po_0.regf_0.rf[13][8] ),
    .A2(\po_0.regf_0.rf[14][8] ),
    .A3(\po_0.regf_0.rf[15][8] ),
    .S0(_1461_),
    .S1(_1463_),
    .X(_1557_));
 sky130_fd_sc_hd__a21bo_1 _1760_ (.A1(_1557_),
    .A2(_1466_),
    .B1_N(_1468_),
    .X(_0338_));
 sky130_fd_sc_hd__mux4_1 _1761_ (.A0(\po_0.regf_0.rf[8][8] ),
    .A1(\po_0.regf_0.rf[9][8] ),
    .A2(\po_0.regf_0.rf[10][8] ),
    .A3(\po_0.regf_0.rf[11][8] ),
    .S0(_1471_),
    .S1(_1472_),
    .X(_0339_));
 sky130_fd_sc_hd__and2b_1 _1762_ (.A_N(_1550_),
    .B(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__o22a_1 _1763_ (.A1(_1554_),
    .A2(_1556_),
    .B1(_0338_),
    .B2(_0340_),
    .X(\po_0.regf_0._5_[8] ));
 sky130_fd_sc_hd__mux4_1 _1764_ (.A0(\po_0.regf_0.rf[4][9] ),
    .A1(\po_0.regf_0.rf[5][9] ),
    .A2(\po_0.regf_0.rf[6][9] ),
    .A3(\po_0.regf_0.rf[7][9] ),
    .S0(_1542_),
    .S1(_1543_),
    .X(_0341_));
 sky130_fd_sc_hd__a21o_1 _1765_ (.A1(_0341_),
    .A2(_1484_),
    .B1(_1492_),
    .X(_0342_));
 sky130_fd_sc_hd__mux4_1 _1766_ (.A0(\po_0.regf_0.rf[0][9] ),
    .A1(\po_0.regf_0.rf[1][9] ),
    .A2(\po_0.regf_0.rf[2][9] ),
    .A3(\po_0.regf_0.rf[3][9] ),
    .S0(_1512_),
    .S1(_1513_),
    .X(_0343_));
 sky130_fd_sc_hd__and2b_1 _1767_ (.A_N(_1511_),
    .B(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__mux4_1 _1768_ (.A0(\po_0.regf_0.rf[12][9] ),
    .A1(\po_0.regf_0.rf[13][9] ),
    .A2(\po_0.regf_0.rf[14][9] ),
    .A3(\po_0.regf_0.rf[15][9] ),
    .S0(_1461_),
    .S1(_1463_),
    .X(_0345_));
 sky130_fd_sc_hd__a21bo_1 _1769_ (.A1(_0345_),
    .A2(_1466_),
    .B1_N(_1468_),
    .X(_0346_));
 sky130_fd_sc_hd__mux4_1 _1770_ (.A0(\po_0.regf_0.rf[8][9] ),
    .A1(\po_0.regf_0.rf[9][9] ),
    .A2(\po_0.regf_0.rf[10][9] ),
    .A3(\po_0.regf_0.rf[11][9] ),
    .S0(_1471_),
    .S1(_1472_),
    .X(_0347_));
 sky130_fd_sc_hd__and2b_1 _1771_ (.A_N(_1550_),
    .B(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__o22a_1 _1772_ (.A1(_0342_),
    .A2(_0344_),
    .B1(_0346_),
    .B2(_0348_),
    .X(\po_0.regf_0._5_[9] ));
 sky130_fd_sc_hd__mux4_1 _1773_ (.A0(\po_0.regf_0.rf[12][10] ),
    .A1(\po_0.regf_0.rf[13][10] ),
    .A2(\po_0.regf_0.rf[14][10] ),
    .A3(\po_0.regf_0.rf[15][10] ),
    .S0(_1481_),
    .S1(_1482_),
    .X(_0349_));
 sky130_fd_sc_hd__a21bo_1 _1774_ (.A1(_0349_),
    .A2(_1470_),
    .B1_N(_1467_),
    .X(_0350_));
 sky130_fd_sc_hd__mux4_1 _1775_ (.A0(\po_0.regf_0.rf[8][10] ),
    .A1(\po_0.regf_0.rf[9][10] ),
    .A2(\po_0.regf_0.rf[10][10] ),
    .A3(\po_0.regf_0.rf[11][10] ),
    .S0(_1512_),
    .S1(_1513_),
    .X(_0351_));
 sky130_fd_sc_hd__and2b_1 _1776_ (.A_N(_1511_),
    .B(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__mux4_1 _1777_ (.A0(\po_0.regf_0.rf[0][10] ),
    .A1(\po_0.regf_0.rf[1][10] ),
    .A2(\po_0.regf_0.rf[2][10] ),
    .A3(\po_0.regf_0.rf[3][10] ),
    .S0(_1497_),
    .S1(_1498_),
    .X(_0353_));
 sky130_fd_sc_hd__mux4_1 _1778_ (.A0(\po_0.regf_0.rf[4][10] ),
    .A1(\po_0.regf_0.rf[5][10] ),
    .A2(\po_0.regf_0.rf[6][10] ),
    .A3(\po_0.regf_0.rf[7][10] ),
    .S0(_1460_),
    .S1(_1462_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _1779_ (.A0(_0353_),
    .A1(_0354_),
    .S(_1465_),
    .X(_0355_));
 sky130_fd_sc_hd__o22a_1 _1780_ (.A1(_0350_),
    .A2(_0352_),
    .B1(_1493_),
    .B2(_0355_),
    .X(\po_0.regf_0._5_[10] ));
 sky130_fd_sc_hd__mux4_1 _1781_ (.A0(\po_0.regf_0.rf[8][11] ),
    .A1(\po_0.regf_0.rf[9][11] ),
    .A2(\po_0.regf_0.rf[10][11] ),
    .A3(\po_0.regf_0.rf[11][11] ),
    .S0(_1494_),
    .S1(_1495_),
    .X(_0356_));
 sky130_fd_sc_hd__and2b_1 _1782_ (.A_N(_1500_),
    .B(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__mux4_1 _1783_ (.A0(\po_0.regf_0.rf[12][11] ),
    .A1(\po_0.regf_0.rf[13][11] ),
    .A2(\po_0.regf_0.rf[14][11] ),
    .A3(\po_0.regf_0.rf[15][11] ),
    .S0(_1542_),
    .S1(_1543_),
    .X(_0358_));
 sky130_fd_sc_hd__a21bo_1 _1784_ (.A1(_0358_),
    .A2(_1550_),
    .B1_N(_1485_),
    .X(_0359_));
 sky130_fd_sc_hd__mux4_1 _1785_ (.A0(\po_0.regf_0.rf[0][11] ),
    .A1(\po_0.regf_0.rf[1][11] ),
    .A2(\po_0.regf_0.rf[2][11] ),
    .A3(\po_0.regf_0.rf[3][11] ),
    .S0(_1488_),
    .S1(_1489_),
    .X(_0360_));
 sky130_fd_sc_hd__and2b_1 _1786_ (.A_N(_1487_),
    .B(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__mux4_1 _1787_ (.A0(\po_0.regf_0.rf[4][11] ),
    .A1(\po_0.regf_0.rf[5][11] ),
    .A2(\po_0.regf_0.rf[6][11] ),
    .A3(\po_0.regf_0.rf[7][11] ),
    .S0(_1475_),
    .S1(_1476_),
    .X(_0362_));
 sky130_fd_sc_hd__a21o_1 _1788_ (.A1(_0362_),
    .A2(_1478_),
    .B1(_1479_),
    .X(_0363_));
 sky130_fd_sc_hd__o22a_1 _1789_ (.A1(_0357_),
    .A2(_0359_),
    .B1(_0361_),
    .B2(_0363_),
    .X(\po_0.regf_0._5_[11] ));
 sky130_fd_sc_hd__mux4_1 _1790_ (.A0(\po_0.regf_0.rf[4][12] ),
    .A1(\po_0.regf_0.rf[5][12] ),
    .A2(\po_0.regf_0.rf[6][12] ),
    .A3(\po_0.regf_0.rf[7][12] ),
    .S0(_1542_),
    .S1(_1543_),
    .X(_0364_));
 sky130_fd_sc_hd__a21o_1 _1791_ (.A1(_0364_),
    .A2(_1484_),
    .B1(_1492_),
    .X(_0365_));
 sky130_fd_sc_hd__mux4_1 _1792_ (.A0(\po_0.regf_0.rf[0][12] ),
    .A1(\po_0.regf_0.rf[1][12] ),
    .A2(\po_0.regf_0.rf[2][12] ),
    .A3(\po_0.regf_0.rf[3][12] ),
    .S0(_1455_),
    .S1(_1457_),
    .X(_0366_));
 sky130_fd_sc_hd__and2b_1 _1793_ (.A_N(_1453_),
    .B(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__mux4_1 _1794_ (.A0(\po_0.regf_0.rf[12][12] ),
    .A1(\po_0.regf_0.rf[13][12] ),
    .A2(\po_0.regf_0.rf[14][12] ),
    .A3(\po_0.regf_0.rf[15][12] ),
    .S0(_1461_),
    .S1(_1463_),
    .X(_0368_));
 sky130_fd_sc_hd__a21bo_1 _1795_ (.A1(_0368_),
    .A2(_1466_),
    .B1_N(_1468_),
    .X(_0369_));
 sky130_fd_sc_hd__mux4_1 _1796_ (.A0(\po_0.regf_0.rf[8][12] ),
    .A1(\po_0.regf_0.rf[9][12] ),
    .A2(\po_0.regf_0.rf[10][12] ),
    .A3(\po_0.regf_0.rf[11][12] ),
    .S0(_1471_),
    .S1(_1472_),
    .X(_0370_));
 sky130_fd_sc_hd__and2b_1 _1797_ (.A_N(_1550_),
    .B(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__o22a_1 _1798_ (.A1(_0365_),
    .A2(_0367_),
    .B1(_0369_),
    .B2(_0371_),
    .X(\po_0.regf_0._5_[12] ));
 sky130_fd_sc_hd__mux4_1 _1799_ (.A0(\po_0.regf_0.rf[8][13] ),
    .A1(\po_0.regf_0.rf[9][13] ),
    .A2(\po_0.regf_0.rf[10][13] ),
    .A3(\po_0.regf_0.rf[11][13] ),
    .S0(_1494_),
    .S1(_1495_),
    .X(_0372_));
 sky130_fd_sc_hd__and2b_1 _1800_ (.A_N(_1500_),
    .B(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__mux4_1 _1801_ (.A0(\po_0.regf_0.rf[12][13] ),
    .A1(\po_0.regf_0.rf[13][13] ),
    .A2(\po_0.regf_0.rf[14][13] ),
    .A3(\po_0.regf_0.rf[15][13] ),
    .S0(_1542_),
    .S1(_1543_),
    .X(_0374_));
 sky130_fd_sc_hd__a21bo_1 _1802_ (.A1(_0374_),
    .A2(_1550_),
    .B1_N(_1485_),
    .X(_0375_));
 sky130_fd_sc_hd__mux4_1 _1803_ (.A0(\po_0.regf_0.rf[0][13] ),
    .A1(\po_0.regf_0.rf[1][13] ),
    .A2(\po_0.regf_0.rf[2][13] ),
    .A3(\po_0.regf_0.rf[3][13] ),
    .S0(_1488_),
    .S1(_1489_),
    .X(_0376_));
 sky130_fd_sc_hd__and2b_1 _1804_ (.A_N(_1487_),
    .B(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__mux4_1 _1805_ (.A0(\po_0.regf_0.rf[4][13] ),
    .A1(\po_0.regf_0.rf[5][13] ),
    .A2(\po_0.regf_0.rf[6][13] ),
    .A3(\po_0.regf_0.rf[7][13] ),
    .S0(_1475_),
    .S1(_1476_),
    .X(_0378_));
 sky130_fd_sc_hd__a21o_1 _1806_ (.A1(_0378_),
    .A2(_1478_),
    .B1(_1479_),
    .X(_0379_));
 sky130_fd_sc_hd__o22a_1 _1807_ (.A1(_0373_),
    .A2(_0375_),
    .B1(_0377_),
    .B2(_0379_),
    .X(\po_0.regf_0._5_[13] ));
 sky130_fd_sc_hd__mux4_1 _1808_ (.A0(\po_0.regf_0.rf[12][14] ),
    .A1(\po_0.regf_0.rf[13][14] ),
    .A2(\po_0.regf_0.rf[14][14] ),
    .A3(\po_0.regf_0.rf[15][14] ),
    .S0(_1481_),
    .S1(_1482_),
    .X(_0380_));
 sky130_fd_sc_hd__a21bo_1 _1809_ (.A1(_0380_),
    .A2(_1470_),
    .B1_N(_1467_),
    .X(_0381_));
 sky130_fd_sc_hd__mux4_1 _1810_ (.A0(\po_0.regf_0.rf[8][14] ),
    .A1(\po_0.regf_0.rf[9][14] ),
    .A2(\po_0.regf_0.rf[10][14] ),
    .A3(\po_0.regf_0.rf[11][14] ),
    .S0(_1455_),
    .S1(_1457_),
    .X(_0382_));
 sky130_fd_sc_hd__and2b_1 _1811_ (.A_N(_1453_),
    .B(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__mux4_1 _1812_ (.A0(\po_0.regf_0.rf[0][14] ),
    .A1(\po_0.regf_0.rf[1][14] ),
    .A2(\po_0.regf_0.rf[2][14] ),
    .A3(\po_0.regf_0.rf[3][14] ),
    .S0(_1497_),
    .S1(_1498_),
    .X(_0384_));
 sky130_fd_sc_hd__mux4_1 _1813_ (.A0(\po_0.regf_0.rf[4][14] ),
    .A1(\po_0.regf_0.rf[5][14] ),
    .A2(\po_0.regf_0.rf[6][14] ),
    .A3(\po_0.regf_0.rf[7][14] ),
    .S0(_1460_),
    .S1(_1462_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _1814_ (.A0(_0384_),
    .A1(_0385_),
    .S(_1465_),
    .X(_0386_));
 sky130_fd_sc_hd__o22a_1 _1815_ (.A1(_0381_),
    .A2(_0383_),
    .B1(_1493_),
    .B2(_0386_),
    .X(\po_0.regf_0._5_[14] ));
 sky130_fd_sc_hd__mux4_1 _1816_ (.A0(\po_0.regf_0.rf[12][15] ),
    .A1(\po_0.regf_0.rf[13][15] ),
    .A2(\po_0.regf_0.rf[14][15] ),
    .A3(\po_0.regf_0.rf[15][15] ),
    .S0(_1471_),
    .S1(_1472_),
    .X(_0387_));
 sky130_fd_sc_hd__a21bo_1 _1817_ (.A1(_0387_),
    .A2(_1470_),
    .B1_N(_1467_),
    .X(_0388_));
 sky130_fd_sc_hd__mux4_1 _1818_ (.A0(\po_0.regf_0.rf[8][15] ),
    .A1(\po_0.regf_0.rf[9][15] ),
    .A2(\po_0.regf_0.rf[10][15] ),
    .A3(\po_0.regf_0.rf[11][15] ),
    .S0(_1455_),
    .S1(_1457_),
    .X(_0389_));
 sky130_fd_sc_hd__and2b_1 _1819_ (.A_N(_1453_),
    .B(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__mux4_1 _1820_ (.A0(\po_0.regf_0.rf[0][15] ),
    .A1(\po_0.regf_0.rf[1][15] ),
    .A2(\po_0.regf_0.rf[2][15] ),
    .A3(\po_0.regf_0.rf[3][15] ),
    .S0(_1497_),
    .S1(_1498_),
    .X(_0391_));
 sky130_fd_sc_hd__mux4_1 _1821_ (.A0(\po_0.regf_0.rf[4][15] ),
    .A1(\po_0.regf_0.rf[5][15] ),
    .A2(\po_0.regf_0.rf[6][15] ),
    .A3(\po_0.regf_0.rf[7][15] ),
    .S0(_1460_),
    .S1(_1462_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _1822_ (.A0(_0391_),
    .A1(_0392_),
    .S(_1465_),
    .X(_0393_));
 sky130_fd_sc_hd__o22a_1 _1823_ (.A1(_0388_),
    .A2(_0390_),
    .B1(_1479_),
    .B2(_0393_),
    .X(\po_0.regf_0._5_[15] ));
 sky130_fd_sc_hd__clkbuf_2 _1824_ (.A(_0000_),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_4 _1825_ (.A(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1826_ (.A(_0001_),
    .X(_0396_));
 sky130_fd_sc_hd__buf_2 _1827_ (.A(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__mux4_1 _1828_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(\po_0.regf_0.rf[13][0] ),
    .A2(\po_0.regf_0.rf[14][0] ),
    .A3(\po_0.regf_0.rf[15][0] ),
    .S0(_0395_),
    .S1(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__buf_2 _1829_ (.A(_0002_),
    .X(_0399_));
 sky130_fd_sc_hd__buf_2 _1830_ (.A(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_2 _1831_ (.A(_0003_),
    .X(_0401_));
 sky130_fd_sc_hd__a21bo_1 _1832_ (.A1(_0398_),
    .A2(_0400_),
    .B1_N(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_2 _1833_ (.A(_0399_),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_4 _1834_ (.A(_0000_),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_4 _1835_ (.A(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__buf_2 _1836_ (.A(_0001_),
    .X(_0406_));
 sky130_fd_sc_hd__buf_2 _1837_ (.A(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__mux4_1 _1838_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(\po_0.regf_0.rf[9][0] ),
    .A2(\po_0.regf_0.rf[10][0] ),
    .A3(\po_0.regf_0.rf[11][0] ),
    .S0(_0405_),
    .S1(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__and2b_1 _1839_ (.A_N(_0403_),
    .B(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__buf_2 _1840_ (.A(_0003_),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_4 _1841_ (.A(_0404_),
    .X(_0411_));
 sky130_fd_sc_hd__buf_2 _1842_ (.A(_0406_),
    .X(_0412_));
 sky130_fd_sc_hd__mux4_1 _1843_ (.A0(\po_0.regf_0.rf[0][0] ),
    .A1(\po_0.regf_0.rf[1][0] ),
    .A2(\po_0.regf_0.rf[2][0] ),
    .A3(\po_0.regf_0.rf[3][0] ),
    .S0(_0411_),
    .S1(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__buf_4 _1844_ (.A(_0404_),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_4 _1845_ (.A(_0406_),
    .X(_0415_));
 sky130_fd_sc_hd__mux4_1 _1846_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(\po_0.regf_0.rf[5][0] ),
    .A2(\po_0.regf_0.rf[6][0] ),
    .A3(\po_0.regf_0.rf[7][0] ),
    .S0(_0414_),
    .S1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_2 _1847_ (.A(_0002_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _1848_ (.A0(_0413_),
    .A1(_0416_),
    .S(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__o22a_1 _1849_ (.A1(_0402_),
    .A2(_0409_),
    .B1(_0410_),
    .B2(_0418_),
    .X(\po_0.regf_0._3_[0] ));
 sky130_fd_sc_hd__clkbuf_4 _1850_ (.A(_0394_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_4 _1851_ (.A(_0396_),
    .X(_0420_));
 sky130_fd_sc_hd__mux4_1 _1852_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(\po_0.regf_0.rf[5][1] ),
    .A2(\po_0.regf_0.rf[6][1] ),
    .A3(\po_0.regf_0.rf[7][1] ),
    .S0(_0419_),
    .S1(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_2 _1853_ (.A(_0002_),
    .X(_0422_));
 sky130_fd_sc_hd__buf_2 _1854_ (.A(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__buf_2 _1855_ (.A(_0003_),
    .X(_0424_));
 sky130_fd_sc_hd__a21o_1 _1856_ (.A1(_0421_),
    .A2(_0423_),
    .B1(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__mux4_1 _1857_ (.A0(\po_0.regf_0.rf[0][1] ),
    .A1(\po_0.regf_0.rf[1][1] ),
    .A2(\po_0.regf_0.rf[2][1] ),
    .A3(\po_0.regf_0.rf[3][1] ),
    .S0(_0405_),
    .S1(_0407_),
    .X(_0426_));
 sky130_fd_sc_hd__and2b_1 _1858_ (.A_N(_0403_),
    .B(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_4 _1859_ (.A(_0394_),
    .X(_0428_));
 sky130_fd_sc_hd__buf_2 _1860_ (.A(_0396_),
    .X(_0429_));
 sky130_fd_sc_hd__mux4_1 _1861_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(\po_0.regf_0.rf[13][1] ),
    .A2(\po_0.regf_0.rf[14][1] ),
    .A3(\po_0.regf_0.rf[15][1] ),
    .S0(_0428_),
    .S1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_2 _1862_ (.A(_0422_),
    .X(_0431_));
 sky130_fd_sc_hd__buf_2 _1863_ (.A(_0003_),
    .X(_0432_));
 sky130_fd_sc_hd__a21bo_1 _1864_ (.A1(_0430_),
    .A2(_0431_),
    .B1_N(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_2 _1865_ (.A(_0422_),
    .X(_0434_));
 sky130_fd_sc_hd__buf_4 _1866_ (.A(_0394_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_4 _1867_ (.A(_0396_),
    .X(_0436_));
 sky130_fd_sc_hd__mux4_1 _1868_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(\po_0.regf_0.rf[9][1] ),
    .A2(\po_0.regf_0.rf[10][1] ),
    .A3(\po_0.regf_0.rf[11][1] ),
    .S0(_0435_),
    .S1(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__and2b_1 _1869_ (.A_N(_0434_),
    .B(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__o22a_1 _1870_ (.A1(_0425_),
    .A2(_0427_),
    .B1(_0433_),
    .B2(_0438_),
    .X(\po_0.regf_0._3_[1] ));
 sky130_fd_sc_hd__mux4_1 _1871_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(\po_0.regf_0.rf[9][2] ),
    .A2(\po_0.regf_0.rf[10][2] ),
    .A3(\po_0.regf_0.rf[11][2] ),
    .S0(_0411_),
    .S1(_0412_),
    .X(_0439_));
 sky130_fd_sc_hd__and2b_1 _1872_ (.A_N(_0417_),
    .B(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_4 _1873_ (.A(_0394_),
    .X(_0441_));
 sky130_fd_sc_hd__buf_2 _1874_ (.A(_0396_),
    .X(_0442_));
 sky130_fd_sc_hd__mux4_1 _1875_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(\po_0.regf_0.rf[13][2] ),
    .A2(\po_0.regf_0.rf[14][2] ),
    .A3(\po_0.regf_0.rf[15][2] ),
    .S0(_0441_),
    .S1(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__buf_2 _1876_ (.A(_0422_),
    .X(_0444_));
 sky130_fd_sc_hd__buf_2 _1877_ (.A(_0003_),
    .X(_0445_));
 sky130_fd_sc_hd__a21bo_1 _1878_ (.A1(_0443_),
    .A2(_0444_),
    .B1_N(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__buf_2 _1879_ (.A(_0399_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_4 _1880_ (.A(_0394_),
    .X(_0448_));
 sky130_fd_sc_hd__buf_2 _1881_ (.A(_0396_),
    .X(_0449_));
 sky130_fd_sc_hd__mux4_1 _1882_ (.A0(\po_0.regf_0.rf[0][2] ),
    .A1(\po_0.regf_0.rf[1][2] ),
    .A2(\po_0.regf_0.rf[2][2] ),
    .A3(\po_0.regf_0.rf[3][2] ),
    .S0(_0448_),
    .S1(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__and2b_1 _1883_ (.A_N(_0447_),
    .B(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__mux4_1 _1884_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(\po_0.regf_0.rf[5][2] ),
    .A2(\po_0.regf_0.rf[6][2] ),
    .A3(\po_0.regf_0.rf[7][2] ),
    .S0(_0428_),
    .S1(_0429_),
    .X(_0452_));
 sky130_fd_sc_hd__a21o_1 _1885_ (.A1(_0452_),
    .A2(_0431_),
    .B1(_0410_),
    .X(_0453_));
 sky130_fd_sc_hd__o22a_1 _1886_ (.A1(_0440_),
    .A2(_0446_),
    .B1(_0451_),
    .B2(_0453_),
    .X(\po_0.regf_0._3_[2] ));
 sky130_fd_sc_hd__mux4_1 _1887_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(\po_0.regf_0.rf[13][3] ),
    .A2(\po_0.regf_0.rf[14][3] ),
    .A3(\po_0.regf_0.rf[15][3] ),
    .S0(_0395_),
    .S1(_0397_),
    .X(_0454_));
 sky130_fd_sc_hd__a21bo_1 _1888_ (.A1(_0454_),
    .A2(_0447_),
    .B1_N(_0401_),
    .X(_0455_));
 sky130_fd_sc_hd__mux4_1 _1889_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(\po_0.regf_0.rf[9][3] ),
    .A2(\po_0.regf_0.rf[10][3] ),
    .A3(\po_0.regf_0.rf[11][3] ),
    .S0(_0405_),
    .S1(_0407_),
    .X(_0456_));
 sky130_fd_sc_hd__and2b_1 _1890_ (.A_N(_0403_),
    .B(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__mux4_1 _1891_ (.A0(\po_0.regf_0.rf[0][3] ),
    .A1(\po_0.regf_0.rf[1][3] ),
    .A2(\po_0.regf_0.rf[2][3] ),
    .A3(\po_0.regf_0.rf[3][3] ),
    .S0(_0411_),
    .S1(_0412_),
    .X(_0458_));
 sky130_fd_sc_hd__mux4_1 _1892_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(\po_0.regf_0.rf[5][3] ),
    .A2(\po_0.regf_0.rf[6][3] ),
    .A3(\po_0.regf_0.rf[7][3] ),
    .S0(_0414_),
    .S1(_0415_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _1893_ (.A0(_0458_),
    .A1(_0459_),
    .S(_0417_),
    .X(_0460_));
 sky130_fd_sc_hd__o22a_1 _1894_ (.A1(_0455_),
    .A2(_0457_),
    .B1(_0410_),
    .B2(_0460_),
    .X(\po_0.regf_0._3_[3] ));
 sky130_fd_sc_hd__mux4_1 _1895_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(\po_0.regf_0.rf[5][4] ),
    .A2(\po_0.regf_0.rf[6][4] ),
    .A3(\po_0.regf_0.rf[7][4] ),
    .S0(_0419_),
    .S1(_0420_),
    .X(_0461_));
 sky130_fd_sc_hd__a21o_1 _1896_ (.A1(_0461_),
    .A2(_0423_),
    .B1(_0424_),
    .X(_0462_));
 sky130_fd_sc_hd__mux4_1 _1897_ (.A0(\po_0.regf_0.rf[0][4] ),
    .A1(\po_0.regf_0.rf[1][4] ),
    .A2(\po_0.regf_0.rf[2][4] ),
    .A3(\po_0.regf_0.rf[3][4] ),
    .S0(_0405_),
    .S1(_0407_),
    .X(_0463_));
 sky130_fd_sc_hd__and2b_1 _1898_ (.A_N(_0403_),
    .B(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__mux4_1 _1899_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(\po_0.regf_0.rf[13][4] ),
    .A2(\po_0.regf_0.rf[14][4] ),
    .A3(\po_0.regf_0.rf[15][4] ),
    .S0(_0428_),
    .S1(_0429_),
    .X(_0465_));
 sky130_fd_sc_hd__a21bo_1 _1900_ (.A1(_0465_),
    .A2(_0431_),
    .B1_N(_0432_),
    .X(_0466_));
 sky130_fd_sc_hd__mux4_1 _1901_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(\po_0.regf_0.rf[9][4] ),
    .A2(\po_0.regf_0.rf[10][4] ),
    .A3(\po_0.regf_0.rf[11][4] ),
    .S0(_0435_),
    .S1(_0436_),
    .X(_0467_));
 sky130_fd_sc_hd__and2b_1 _1902_ (.A_N(_0434_),
    .B(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__o22a_1 _1903_ (.A1(_0462_),
    .A2(_0464_),
    .B1(_0466_),
    .B2(_0468_),
    .X(\po_0.regf_0._3_[4] ));
 sky130_fd_sc_hd__mux4_1 _1904_ (.A0(\po_0.regf_0.rf[0][5] ),
    .A1(\po_0.regf_0.rf[1][5] ),
    .A2(\po_0.regf_0.rf[2][5] ),
    .A3(\po_0.regf_0.rf[3][5] ),
    .S0(_0404_),
    .S1(_0406_),
    .X(_0469_));
 sky130_fd_sc_hd__mux4_1 _1905_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(\po_0.regf_0.rf[5][5] ),
    .A2(\po_0.regf_0.rf[6][5] ),
    .A3(\po_0.regf_0.rf[7][5] ),
    .S0(_0404_),
    .S1(_0406_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _1906_ (.A0(_0469_),
    .A1(_0470_),
    .S(_0399_),
    .X(_0471_));
 sky130_fd_sc_hd__mux4_1 _1907_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(\po_0.regf_0.rf[9][5] ),
    .A2(\po_0.regf_0.rf[10][5] ),
    .A3(\po_0.regf_0.rf[11][5] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_0472_));
 sky130_fd_sc_hd__mux4_1 _1908_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(\po_0.regf_0.rf[13][5] ),
    .A2(\po_0.regf_0.rf[14][5] ),
    .A3(\po_0.regf_0.rf[15][5] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _1909_ (.A0(_0472_),
    .A1(_0473_),
    .S(_0399_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _1910_ (.A0(_0471_),
    .A1(_0474_),
    .S(_0445_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_1 _1911_ (.A(_0475_),
    .X(\po_0.regf_0._3_[5] ));
 sky130_fd_sc_hd__mux4_1 _1912_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(\po_0.regf_0.rf[5][6] ),
    .A2(\po_0.regf_0.rf[6][6] ),
    .A3(\po_0.regf_0.rf[7][6] ),
    .S0(_0419_),
    .S1(_0420_),
    .X(_0476_));
 sky130_fd_sc_hd__a21o_1 _1913_ (.A1(_0476_),
    .A2(_0400_),
    .B1(_0424_),
    .X(_0477_));
 sky130_fd_sc_hd__mux4_1 _1914_ (.A0(\po_0.regf_0.rf[0][6] ),
    .A1(\po_0.regf_0.rf[1][6] ),
    .A2(\po_0.regf_0.rf[2][6] ),
    .A3(\po_0.regf_0.rf[3][6] ),
    .S0(_0405_),
    .S1(_0407_),
    .X(_0478_));
 sky130_fd_sc_hd__and2b_1 _1915_ (.A_N(_0403_),
    .B(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__mux4_1 _1916_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(\po_0.regf_0.rf[13][6] ),
    .A2(\po_0.regf_0.rf[14][6] ),
    .A3(\po_0.regf_0.rf[15][6] ),
    .S0(_0441_),
    .S1(_0442_),
    .X(_0480_));
 sky130_fd_sc_hd__a21bo_1 _1917_ (.A1(_0480_),
    .A2(_0444_),
    .B1_N(_0432_),
    .X(_0481_));
 sky130_fd_sc_hd__mux4_1 _1918_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(\po_0.regf_0.rf[9][6] ),
    .A2(\po_0.regf_0.rf[10][6] ),
    .A3(\po_0.regf_0.rf[11][6] ),
    .S0(_0435_),
    .S1(_0436_),
    .X(_0482_));
 sky130_fd_sc_hd__and2b_1 _1919_ (.A_N(_0434_),
    .B(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__o22a_1 _1920_ (.A1(_0477_),
    .A2(_0479_),
    .B1(_0481_),
    .B2(_0483_),
    .X(\po_0.regf_0._3_[6] ));
 sky130_fd_sc_hd__mux4_1 _1921_ (.A0(\po_0.regf_0.rf[8][7] ),
    .A1(\po_0.regf_0.rf[9][7] ),
    .A2(\po_0.regf_0.rf[10][7] ),
    .A3(\po_0.regf_0.rf[11][7] ),
    .S0(_0411_),
    .S1(_0412_),
    .X(_0484_));
 sky130_fd_sc_hd__and2b_1 _1922_ (.A_N(_0417_),
    .B(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__mux4_1 _1923_ (.A0(\po_0.regf_0.rf[12][7] ),
    .A1(\po_0.regf_0.rf[13][7] ),
    .A2(\po_0.regf_0.rf[14][7] ),
    .A3(\po_0.regf_0.rf[15][7] ),
    .S0(_0419_),
    .S1(_0420_),
    .X(_0486_));
 sky130_fd_sc_hd__a21bo_1 _1924_ (.A1(_0486_),
    .A2(_0434_),
    .B1_N(_0401_),
    .X(_0487_));
 sky130_fd_sc_hd__mux4_1 _1925_ (.A0(\po_0.regf_0.rf[0][7] ),
    .A1(\po_0.regf_0.rf[1][7] ),
    .A2(\po_0.regf_0.rf[2][7] ),
    .A3(\po_0.regf_0.rf[3][7] ),
    .S0(_0448_),
    .S1(_0449_),
    .X(_0488_));
 sky130_fd_sc_hd__and2b_1 _1926_ (.A_N(_0447_),
    .B(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__mux4_1 _1927_ (.A0(\po_0.regf_0.rf[4][7] ),
    .A1(\po_0.regf_0.rf[5][7] ),
    .A2(\po_0.regf_0.rf[6][7] ),
    .A3(\po_0.regf_0.rf[7][7] ),
    .S0(_0428_),
    .S1(_0429_),
    .X(_0490_));
 sky130_fd_sc_hd__a21o_1 _1928_ (.A1(_0490_),
    .A2(_0431_),
    .B1(_0410_),
    .X(_0491_));
 sky130_fd_sc_hd__o22a_1 _1929_ (.A1(_0485_),
    .A2(_0487_),
    .B1(_0489_),
    .B2(_0491_),
    .X(\po_0.regf_0._3_[7] ));
 sky130_fd_sc_hd__mux4_1 _1930_ (.A0(\po_0.regf_0.rf[4][8] ),
    .A1(\po_0.regf_0.rf[5][8] ),
    .A2(\po_0.regf_0.rf[6][8] ),
    .A3(\po_0.regf_0.rf[7][8] ),
    .S0(_0395_),
    .S1(_0397_),
    .X(_0492_));
 sky130_fd_sc_hd__a21o_1 _1931_ (.A1(_0492_),
    .A2(_0400_),
    .B1(_0424_),
    .X(_0493_));
 sky130_fd_sc_hd__clkbuf_2 _1932_ (.A(_0399_),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_4 _1933_ (.A(_0404_),
    .X(_0495_));
 sky130_fd_sc_hd__buf_2 _1934_ (.A(_0406_),
    .X(_0496_));
 sky130_fd_sc_hd__mux4_1 _1935_ (.A0(\po_0.regf_0.rf[0][8] ),
    .A1(\po_0.regf_0.rf[1][8] ),
    .A2(\po_0.regf_0.rf[2][8] ),
    .A3(\po_0.regf_0.rf[3][8] ),
    .S0(_0495_),
    .S1(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__and2b_1 _1936_ (.A_N(_0494_),
    .B(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__mux4_1 _1937_ (.A0(\po_0.regf_0.rf[12][8] ),
    .A1(\po_0.regf_0.rf[13][8] ),
    .A2(\po_0.regf_0.rf[14][8] ),
    .A3(\po_0.regf_0.rf[15][8] ),
    .S0(_0441_),
    .S1(_0442_),
    .X(_0499_));
 sky130_fd_sc_hd__a21bo_1 _1938_ (.A1(_0499_),
    .A2(_0444_),
    .B1_N(_0445_),
    .X(_0500_));
 sky130_fd_sc_hd__mux4_1 _1939_ (.A0(\po_0.regf_0.rf[8][8] ),
    .A1(\po_0.regf_0.rf[9][8] ),
    .A2(\po_0.regf_0.rf[10][8] ),
    .A3(\po_0.regf_0.rf[11][8] ),
    .S0(_0435_),
    .S1(_0436_),
    .X(_0501_));
 sky130_fd_sc_hd__and2b_1 _1940_ (.A_N(_0423_),
    .B(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__o22a_1 _1941_ (.A1(_0493_),
    .A2(_0498_),
    .B1(_0500_),
    .B2(_0502_),
    .X(\po_0.regf_0._3_[8] ));
 sky130_fd_sc_hd__mux4_1 _1942_ (.A0(\po_0.regf_0.rf[12][9] ),
    .A1(\po_0.regf_0.rf[13][9] ),
    .A2(\po_0.regf_0.rf[14][9] ),
    .A3(\po_0.regf_0.rf[15][9] ),
    .S0(_0435_),
    .S1(_0436_),
    .X(_0503_));
 sky130_fd_sc_hd__a21bo_1 _1943_ (.A1(_0503_),
    .A2(_0447_),
    .B1_N(_0401_),
    .X(_0504_));
 sky130_fd_sc_hd__mux4_1 _1944_ (.A0(\po_0.regf_0.rf[8][9] ),
    .A1(\po_0.regf_0.rf[9][9] ),
    .A2(\po_0.regf_0.rf[10][9] ),
    .A3(\po_0.regf_0.rf[11][9] ),
    .S0(_0495_),
    .S1(_0496_),
    .X(_0505_));
 sky130_fd_sc_hd__and2b_1 _1945_ (.A_N(_0494_),
    .B(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__mux4_1 _1946_ (.A0(\po_0.regf_0.rf[0][9] ),
    .A1(\po_0.regf_0.rf[1][9] ),
    .A2(\po_0.regf_0.rf[2][9] ),
    .A3(\po_0.regf_0.rf[3][9] ),
    .S0(_0414_),
    .S1(_0415_),
    .X(_0507_));
 sky130_fd_sc_hd__mux4_1 _1947_ (.A0(\po_0.regf_0.rf[4][9] ),
    .A1(\po_0.regf_0.rf[5][9] ),
    .A2(\po_0.regf_0.rf[6][9] ),
    .A3(\po_0.regf_0.rf[7][9] ),
    .S0(_0414_),
    .S1(_0415_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _1948_ (.A0(_0507_),
    .A1(_0508_),
    .S(_0422_),
    .X(_0509_));
 sky130_fd_sc_hd__o22a_1 _1949_ (.A1(_0504_),
    .A2(_0506_),
    .B1(_0410_),
    .B2(_0509_),
    .X(\po_0.regf_0._3_[9] ));
 sky130_fd_sc_hd__mux4_1 _1950_ (.A0(\po_0.regf_0.rf[4][10] ),
    .A1(\po_0.regf_0.rf[5][10] ),
    .A2(\po_0.regf_0.rf[6][10] ),
    .A3(\po_0.regf_0.rf[7][10] ),
    .S0(_0395_),
    .S1(_0397_),
    .X(_0510_));
 sky130_fd_sc_hd__a21o_1 _1951_ (.A1(_0510_),
    .A2(_0400_),
    .B1(_0432_),
    .X(_0511_));
 sky130_fd_sc_hd__mux4_1 _1952_ (.A0(\po_0.regf_0.rf[0][10] ),
    .A1(\po_0.regf_0.rf[1][10] ),
    .A2(\po_0.regf_0.rf[2][10] ),
    .A3(\po_0.regf_0.rf[3][10] ),
    .S0(_0495_),
    .S1(_0496_),
    .X(_0512_));
 sky130_fd_sc_hd__and2b_1 _1953_ (.A_N(_0494_),
    .B(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__mux4_1 _1954_ (.A0(\po_0.regf_0.rf[12][10] ),
    .A1(\po_0.regf_0.rf[13][10] ),
    .A2(\po_0.regf_0.rf[14][10] ),
    .A3(\po_0.regf_0.rf[15][10] ),
    .S0(_0441_),
    .S1(_0442_),
    .X(_0514_));
 sky130_fd_sc_hd__a21bo_1 _1955_ (.A1(_0514_),
    .A2(_0444_),
    .B1_N(_0445_),
    .X(_0515_));
 sky130_fd_sc_hd__mux4_1 _1956_ (.A0(\po_0.regf_0.rf[8][10] ),
    .A1(\po_0.regf_0.rf[9][10] ),
    .A2(\po_0.regf_0.rf[10][10] ),
    .A3(\po_0.regf_0.rf[11][10] ),
    .S0(_0448_),
    .S1(_0449_),
    .X(_0516_));
 sky130_fd_sc_hd__and2b_1 _1957_ (.A_N(_0423_),
    .B(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__o22a_1 _1958_ (.A1(_0511_),
    .A2(_0513_),
    .B1(_0515_),
    .B2(_0517_),
    .X(\po_0.regf_0._3_[10] ));
 sky130_fd_sc_hd__mux4_1 _1959_ (.A0(\po_0.regf_0.rf[4][11] ),
    .A1(\po_0.regf_0.rf[5][11] ),
    .A2(\po_0.regf_0.rf[6][11] ),
    .A3(\po_0.regf_0.rf[7][11] ),
    .S0(_0395_),
    .S1(_0397_),
    .X(_0518_));
 sky130_fd_sc_hd__a21o_1 _1960_ (.A1(_0518_),
    .A2(_0400_),
    .B1(_0432_),
    .X(_0519_));
 sky130_fd_sc_hd__mux4_1 _1961_ (.A0(\po_0.regf_0.rf[0][11] ),
    .A1(\po_0.regf_0.rf[1][11] ),
    .A2(\po_0.regf_0.rf[2][11] ),
    .A3(\po_0.regf_0.rf[3][11] ),
    .S0(_0495_),
    .S1(_0496_),
    .X(_0520_));
 sky130_fd_sc_hd__and2b_1 _1962_ (.A_N(_0494_),
    .B(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__mux4_1 _1963_ (.A0(\po_0.regf_0.rf[12][11] ),
    .A1(\po_0.regf_0.rf[13][11] ),
    .A2(\po_0.regf_0.rf[14][11] ),
    .A3(\po_0.regf_0.rf[15][11] ),
    .S0(_0441_),
    .S1(_0442_),
    .X(_0522_));
 sky130_fd_sc_hd__a21bo_1 _1964_ (.A1(_0522_),
    .A2(_0444_),
    .B1_N(_0445_),
    .X(_0523_));
 sky130_fd_sc_hd__mux4_1 _1965_ (.A0(\po_0.regf_0.rf[8][11] ),
    .A1(\po_0.regf_0.rf[9][11] ),
    .A2(\po_0.regf_0.rf[10][11] ),
    .A3(\po_0.regf_0.rf[11][11] ),
    .S0(_0448_),
    .S1(_0449_),
    .X(_0524_));
 sky130_fd_sc_hd__and2b_1 _1966_ (.A_N(_0423_),
    .B(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__o22a_1 _1967_ (.A1(_0519_),
    .A2(_0521_),
    .B1(_0523_),
    .B2(_0525_),
    .X(\po_0.regf_0._3_[11] ));
 sky130_fd_sc_hd__mux4_1 _1968_ (.A0(\po_0.regf_0.rf[8][12] ),
    .A1(\po_0.regf_0.rf[9][12] ),
    .A2(\po_0.regf_0.rf[10][12] ),
    .A3(\po_0.regf_0.rf[11][12] ),
    .S0(_0411_),
    .S1(_0412_),
    .X(_0526_));
 sky130_fd_sc_hd__and2b_1 _1969_ (.A_N(_0417_),
    .B(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__mux4_1 _1970_ (.A0(\po_0.regf_0.rf[12][12] ),
    .A1(\po_0.regf_0.rf[13][12] ),
    .A2(\po_0.regf_0.rf[14][12] ),
    .A3(\po_0.regf_0.rf[15][12] ),
    .S0(_0419_),
    .S1(_0420_),
    .X(_0528_));
 sky130_fd_sc_hd__a21bo_1 _1971_ (.A1(_0528_),
    .A2(_0434_),
    .B1_N(_0401_),
    .X(_0529_));
 sky130_fd_sc_hd__mux4_1 _1972_ (.A0(\po_0.regf_0.rf[0][12] ),
    .A1(\po_0.regf_0.rf[1][12] ),
    .A2(\po_0.regf_0.rf[2][12] ),
    .A3(\po_0.regf_0.rf[3][12] ),
    .S0(_0448_),
    .S1(_0449_),
    .X(_0530_));
 sky130_fd_sc_hd__and2b_1 _1973_ (.A_N(_0447_),
    .B(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__mux4_1 _1974_ (.A0(\po_0.regf_0.rf[4][12] ),
    .A1(\po_0.regf_0.rf[5][12] ),
    .A2(\po_0.regf_0.rf[6][12] ),
    .A3(\po_0.regf_0.rf[7][12] ),
    .S0(_0428_),
    .S1(_0429_),
    .X(_0532_));
 sky130_fd_sc_hd__a21o_1 _1975_ (.A1(_0532_),
    .A2(_0431_),
    .B1(_0424_),
    .X(_0533_));
 sky130_fd_sc_hd__o22a_1 _1976_ (.A1(_0527_),
    .A2(_0529_),
    .B1(_0531_),
    .B2(_0533_),
    .X(\po_0.regf_0._3_[12] ));
 sky130_fd_sc_hd__mux4_1 _1977_ (.A0(\po_0.regf_0.rf[4][13] ),
    .A1(\po_0.regf_0.rf[5][13] ),
    .A2(\po_0.regf_0.rf[6][13] ),
    .A3(\po_0.regf_0.rf[7][13] ),
    .S0(_0395_),
    .S1(_0397_),
    .X(_0534_));
 sky130_fd_sc_hd__a21o_1 _1978_ (.A1(_0534_),
    .A2(_0400_),
    .B1(_0432_),
    .X(_0535_));
 sky130_fd_sc_hd__mux4_1 _1979_ (.A0(\po_0.regf_0.rf[0][13] ),
    .A1(\po_0.regf_0.rf[1][13] ),
    .A2(\po_0.regf_0.rf[2][13] ),
    .A3(\po_0.regf_0.rf[3][13] ),
    .S0(_0495_),
    .S1(_0496_),
    .X(_0536_));
 sky130_fd_sc_hd__and2b_1 _1980_ (.A_N(_0494_),
    .B(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__mux4_1 _1981_ (.A0(\po_0.regf_0.rf[12][13] ),
    .A1(\po_0.regf_0.rf[13][13] ),
    .A2(\po_0.regf_0.rf[14][13] ),
    .A3(\po_0.regf_0.rf[15][13] ),
    .S0(_0441_),
    .S1(_0442_),
    .X(_0538_));
 sky130_fd_sc_hd__a21bo_1 _1982_ (.A1(_0538_),
    .A2(_0444_),
    .B1_N(_0445_),
    .X(_0539_));
 sky130_fd_sc_hd__mux4_1 _1983_ (.A0(\po_0.regf_0.rf[8][13] ),
    .A1(\po_0.regf_0.rf[9][13] ),
    .A2(\po_0.regf_0.rf[10][13] ),
    .A3(\po_0.regf_0.rf[11][13] ),
    .S0(_0448_),
    .S1(_0449_),
    .X(_0540_));
 sky130_fd_sc_hd__and2b_1 _1984_ (.A_N(_0423_),
    .B(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__o22a_1 _1985_ (.A1(_0535_),
    .A2(_0537_),
    .B1(_0539_),
    .B2(_0541_),
    .X(\po_0.regf_0._3_[13] ));
 sky130_fd_sc_hd__mux4_1 _1986_ (.A0(\po_0.regf_0.rf[12][14] ),
    .A1(\po_0.regf_0.rf[13][14] ),
    .A2(\po_0.regf_0.rf[14][14] ),
    .A3(\po_0.regf_0.rf[15][14] ),
    .S0(_0435_),
    .S1(_0436_),
    .X(_0542_));
 sky130_fd_sc_hd__a21bo_1 _1987_ (.A1(_0542_),
    .A2(_0447_),
    .B1_N(_0003_),
    .X(_0543_));
 sky130_fd_sc_hd__mux4_1 _1988_ (.A0(\po_0.regf_0.rf[8][14] ),
    .A1(\po_0.regf_0.rf[9][14] ),
    .A2(\po_0.regf_0.rf[10][14] ),
    .A3(\po_0.regf_0.rf[11][14] ),
    .S0(_0495_),
    .S1(_0496_),
    .X(_0544_));
 sky130_fd_sc_hd__and2b_1 _1989_ (.A_N(_0494_),
    .B(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__mux4_1 _1990_ (.A0(\po_0.regf_0.rf[0][14] ),
    .A1(\po_0.regf_0.rf[1][14] ),
    .A2(\po_0.regf_0.rf[2][14] ),
    .A3(\po_0.regf_0.rf[3][14] ),
    .S0(_0414_),
    .S1(_0415_),
    .X(_0546_));
 sky130_fd_sc_hd__mux4_1 _1991_ (.A0(\po_0.regf_0.rf[4][14] ),
    .A1(\po_0.regf_0.rf[5][14] ),
    .A2(\po_0.regf_0.rf[6][14] ),
    .A3(\po_0.regf_0.rf[7][14] ),
    .S0(_0414_),
    .S1(_0415_),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _1992_ (.A0(_0546_),
    .A1(_0547_),
    .S(_0422_),
    .X(_0548_));
 sky130_fd_sc_hd__o22a_1 _1993_ (.A1(_0543_),
    .A2(_0545_),
    .B1(_0410_),
    .B2(_0548_),
    .X(\po_0.regf_0._3_[14] ));
 sky130_fd_sc_hd__mux4_1 _1994_ (.A0(\po_0.regf_0.rf[8][15] ),
    .A1(\po_0.regf_0.rf[9][15] ),
    .A2(\po_0.regf_0.rf[10][15] ),
    .A3(\po_0.regf_0.rf[11][15] ),
    .S0(_0411_),
    .S1(_0412_),
    .X(_0549_));
 sky130_fd_sc_hd__and2b_1 _1995_ (.A_N(_0417_),
    .B(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__mux4_1 _1996_ (.A0(\po_0.regf_0.rf[12][15] ),
    .A1(\po_0.regf_0.rf[13][15] ),
    .A2(\po_0.regf_0.rf[14][15] ),
    .A3(\po_0.regf_0.rf[15][15] ),
    .S0(_0419_),
    .S1(_0420_),
    .X(_0551_));
 sky130_fd_sc_hd__a21bo_1 _1997_ (.A1(_0551_),
    .A2(_0434_),
    .B1_N(_0401_),
    .X(_0552_));
 sky130_fd_sc_hd__mux4_1 _1998_ (.A0(\po_0.regf_0.rf[0][15] ),
    .A1(\po_0.regf_0.rf[1][15] ),
    .A2(\po_0.regf_0.rf[2][15] ),
    .A3(\po_0.regf_0.rf[3][15] ),
    .S0(_0405_),
    .S1(_0407_),
    .X(_0553_));
 sky130_fd_sc_hd__and2b_1 _1999_ (.A_N(_0403_),
    .B(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__mux4_1 _2000_ (.A0(\po_0.regf_0.rf[4][15] ),
    .A1(\po_0.regf_0.rf[5][15] ),
    .A2(\po_0.regf_0.rf[6][15] ),
    .A3(\po_0.regf_0.rf[7][15] ),
    .S0(_0428_),
    .S1(_0429_),
    .X(_0555_));
 sky130_fd_sc_hd__a21o_1 _2001_ (.A1(_0555_),
    .A2(_0431_),
    .B1(_0424_),
    .X(_0556_));
 sky130_fd_sc_hd__o22a_1 _2002_ (.A1(_0550_),
    .A2(_0552_),
    .B1(_0554_),
    .B2(_0556_),
    .X(\po_0.regf_0._3_[15] ));
 sky130_fd_sc_hd__buf_2 _2003_ (.A(\po_0.muxf_0.rf_w_data[4] ),
    .X(_0557_));
 sky130_fd_sc_hd__or3_2 _2004_ (.A(_1441_),
    .B(_1451_),
    .C(_1447_),
    .X(_0558_));
 sky130_fd_sc_hd__clkbuf_2 _2005_ (.A(_1446_),
    .X(_0559_));
 sky130_fd_sc_hd__or2_1 _2006_ (.A(_1439_),
    .B(_1449_),
    .X(_0560_));
 sky130_fd_sc_hd__or4bb_2 _2007_ (.A(_1440_),
    .B(\uc_0.bc_0._54_[1] ),
    .C_N(_0559_),
    .D_N(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__nand2_4 _2008_ (.A(_0558_),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__buf_2 _2009_ (.A(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__buf_2 _2010_ (.A(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _2011_ (.A0(\po_0.regf_0.rq_addr[0] ),
    .A1(_0557_),
    .S(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_1 _2012_ (.A(_0565_),
    .X(_0012_));
 sky130_fd_sc_hd__buf_2 _2013_ (.A(\po_0.muxf_0.rf_w_data[5] ),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _2014_ (.A0(\po_0.regf_0.rq_addr[1] ),
    .A1(_0566_),
    .S(_0564_),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_1 _2015_ (.A(_0567_),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_2 _2016_ (.A(\po_0.muxf_0.rf_w_data[6] ),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _2017_ (.A0(\po_0.regf_0.rq_addr[2] ),
    .A1(_0568_),
    .S(_0564_),
    .X(_0569_));
 sky130_fd_sc_hd__clkbuf_1 _2018_ (.A(_0569_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_4 _2019_ (.A(\po_0.muxf_0.rf_w_data[7] ),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _2020_ (.A0(\po_0.regf_0.rq_addr[3] ),
    .A1(_0570_),
    .S(_0564_),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_1 _2021_ (.A(_0571_),
    .X(_0015_));
 sky130_fd_sc_hd__buf_2 _2022_ (.A(_1441_),
    .X(_0572_));
 sky130_fd_sc_hd__or2_1 _2023_ (.A(\uc_0.bc_0._54_[3] ),
    .B(\uc_0.bc_0._54_[2] ),
    .X(_0573_));
 sky130_fd_sc_hd__a31oi_4 _2024_ (.A1(_0572_),
    .A2(_1447_),
    .A3(_0573_),
    .B1(_0562_),
    .Y(_0574_));
 sky130_fd_sc_hd__buf_2 _2025_ (.A(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _2026_ (.A0(\uc_0._20_[8] ),
    .A1(\po_0.regf_0.rp_addr[0] ),
    .S(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__clkbuf_1 _2027_ (.A(_0576_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _2028_ (.A0(\uc_0._20_[9] ),
    .A1(\po_0.regf_0.rp_addr[1] ),
    .S(_0575_),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_1 _2029_ (.A(_0577_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _2030_ (.A0(\uc_0._20_[10] ),
    .A1(\po_0.regf_0.rp_addr[2] ),
    .S(_0575_),
    .X(_0578_));
 sky130_fd_sc_hd__clkbuf_1 _2031_ (.A(_0578_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _2032_ (.A0(\uc_0._20_[11] ),
    .A1(\po_0.regf_0.rp_addr[3] ),
    .S(_0575_),
    .X(_0579_));
 sky130_fd_sc_hd__clkbuf_1 _2033_ (.A(_0579_),
    .X(_0011_));
 sky130_fd_sc_hd__and2b_1 _2034_ (.A_N(net87),
    .B(\po_0._1_[0] ),
    .X(_0580_));
 sky130_fd_sc_hd__and2_1 _2035_ (.A(net86),
    .B(\po_0._1_[1] ),
    .X(_0581_));
 sky130_fd_sc_hd__nor2_1 _2036_ (.A(net86),
    .B(\po_0._1_[1] ),
    .Y(_0582_));
 sky130_fd_sc_hd__nor2_1 _2037_ (.A(_0581_),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__xor2_1 _2038_ (.A(_0580_),
    .B(_0583_),
    .X(\po_0.alu_0._10_[1] ));
 sky130_fd_sc_hd__inv_2 _2039_ (.A(net86),
    .Y(_0584_));
 sky130_fd_sc_hd__nand2_1 _2040_ (.A(_0584_),
    .B(\po_0._1_[1] ),
    .Y(_0585_));
 sky130_fd_sc_hd__o21ai_1 _2041_ (.A1(\po_0._1_[1] ),
    .A2(_0584_),
    .B1(_0580_),
    .Y(_0586_));
 sky130_fd_sc_hd__and2_1 _2042_ (.A(net43),
    .B(\po_0._1_[2] ),
    .X(_0587_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2043_ (.A(net43),
    .X(_0588_));
 sky130_fd_sc_hd__nor2_1 _2044_ (.A(_0588_),
    .B(\po_0._1_[2] ),
    .Y(_0589_));
 sky130_fd_sc_hd__nor2_1 _2045_ (.A(_0587_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__a21oi_1 _2046_ (.A1(_0585_),
    .A2(_0586_),
    .B1(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__and2b_1 _2047_ (.A_N(_0588_),
    .B(\po_0._1_[2] ),
    .X(_0592_));
 sky130_fd_sc_hd__and2b_1 _2048_ (.A_N(\po_0._1_[2] ),
    .B(_0588_),
    .X(_0593_));
 sky130_fd_sc_hd__o211ai_1 _2049_ (.A1(_0592_),
    .A2(_0593_),
    .B1(_0585_),
    .C1(_0586_),
    .Y(_0594_));
 sky130_fd_sc_hd__or2b_1 _2050_ (.A(_0591_),
    .B_N(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__clkbuf_1 _2051_ (.A(_0595_),
    .X(\po_0.alu_0._10_[2] ));
 sky130_fd_sc_hd__or2b_1 _2052_ (.A(\po_0._1_[2] ),
    .B_N(_0588_),
    .X(_0596_));
 sky130_fd_sc_hd__o211ai_1 _2053_ (.A1(_0587_),
    .A2(_0589_),
    .B1(_0585_),
    .C1(_0586_),
    .Y(_0597_));
 sky130_fd_sc_hd__buf_2 _2054_ (.A(net44),
    .X(_0598_));
 sky130_fd_sc_hd__and2_1 _2055_ (.A(_0598_),
    .B(\po_0._1_[3] ),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_2 _2056_ (.A(_0598_),
    .B(\po_0._1_[3] ),
    .Y(_0600_));
 sky130_fd_sc_hd__o2bb2ai_1 _2057_ (.A1_N(_0596_),
    .A2_N(_0597_),
    .B1(_0599_),
    .B2(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__nor2_1 _2058_ (.A(_0599_),
    .B(_0600_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand3_1 _2059_ (.A(_0596_),
    .B(_0597_),
    .C(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__and2_1 _2060_ (.A(_0601_),
    .B(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__clkbuf_1 _2061_ (.A(_0604_),
    .X(\po_0.alu_0._10_[3] ));
 sky130_fd_sc_hd__clkbuf_2 _2062_ (.A(net45),
    .X(_0605_));
 sky130_fd_sc_hd__and2_1 _2063_ (.A(_0605_),
    .B(\po_0._1_[4] ),
    .X(_0606_));
 sky130_fd_sc_hd__nor2_1 _2064_ (.A(_0605_),
    .B(\po_0._1_[4] ),
    .Y(_0607_));
 sky130_fd_sc_hd__or2b_1 _2065_ (.A(\po_0._1_[3] ),
    .B_N(_0598_),
    .X(_0608_));
 sky130_fd_sc_hd__a2bb2oi_1 _2066_ (.A1_N(_0606_),
    .A2_N(_0607_),
    .B1(_0608_),
    .B2(_0601_),
    .Y(_0609_));
 sky130_fd_sc_hd__nor2_2 _2067_ (.A(_0606_),
    .B(_0607_),
    .Y(_0610_));
 sky130_fd_sc_hd__nand3_1 _2068_ (.A(_0601_),
    .B(_0610_),
    .C(_0608_),
    .Y(_0611_));
 sky130_fd_sc_hd__and2b_1 _2069_ (.A_N(_0609_),
    .B(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__clkbuf_1 _2070_ (.A(_0612_),
    .X(\po_0.alu_0._10_[4] ));
 sky130_fd_sc_hd__clkbuf_2 _2071_ (.A(net46),
    .X(_0613_));
 sky130_fd_sc_hd__nor2_2 _2072_ (.A(_0613_),
    .B(\po_0._1_[5] ),
    .Y(_0614_));
 sky130_fd_sc_hd__and2_1 _2073_ (.A(_0613_),
    .B(\po_0._1_[5] ),
    .X(_0615_));
 sky130_fd_sc_hd__and2b_1 _2074_ (.A_N(\po_0._1_[4] ),
    .B(_0605_),
    .X(_0616_));
 sky130_fd_sc_hd__o22ai_2 _2075_ (.A1(_0614_),
    .A2(_0615_),
    .B1(_0616_),
    .B2(_0609_),
    .Y(_0617_));
 sky130_fd_sc_hd__or4_1 _2076_ (.A(_0609_),
    .B(_0614_),
    .C(_0615_),
    .D(_0616_),
    .X(_0618_));
 sky130_fd_sc_hd__and2_1 _2077_ (.A(_0617_),
    .B(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__clkbuf_1 _2078_ (.A(_0619_),
    .X(\po_0.alu_0._10_[5] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2079_ (.A(net47),
    .X(_0620_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2080_ (.A(\po_0._1_[6] ),
    .X(_0621_));
 sky130_fd_sc_hd__and2_1 _2081_ (.A(_0620_),
    .B(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__nor2_1 _2082_ (.A(_0620_),
    .B(_0621_),
    .Y(_0623_));
 sky130_fd_sc_hd__or2b_1 _2083_ (.A(\po_0._1_[5] ),
    .B_N(_0613_),
    .X(_0624_));
 sky130_fd_sc_hd__a2bb2oi_1 _2084_ (.A1_N(_0622_),
    .A2_N(_0623_),
    .B1(_0624_),
    .B2(_0617_),
    .Y(_0625_));
 sky130_fd_sc_hd__or2b_1 _2085_ (.A(\po_0._1_[6] ),
    .B_N(net47),
    .X(_0626_));
 sky130_fd_sc_hd__or2b_1 _2086_ (.A(net47),
    .B_N(_0621_),
    .X(_0627_));
 sky130_fd_sc_hd__nand2_2 _2087_ (.A(_0626_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__and3_1 _2088_ (.A(_0617_),
    .B(_0628_),
    .C(_0624_),
    .X(_0629_));
 sky130_fd_sc_hd__nor2_1 _2089_ (.A(_0625_),
    .B(_0629_),
    .Y(\po_0.alu_0._10_[6] ));
 sky130_fd_sc_hd__and2b_1 _2090_ (.A_N(_0621_),
    .B(_0620_),
    .X(_0630_));
 sky130_fd_sc_hd__nor2_1 _2091_ (.A(net85),
    .B(\po_0._1_[7] ),
    .Y(_0631_));
 sky130_fd_sc_hd__and2_1 _2092_ (.A(net85),
    .B(\po_0._1_[7] ),
    .X(_0632_));
 sky130_fd_sc_hd__nor2_1 _2093_ (.A(_0631_),
    .B(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__o21bai_2 _2094_ (.A1(_0630_),
    .A2(_0625_),
    .B1_N(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__or4_1 _2095_ (.A(_0630_),
    .B(_0625_),
    .C(_0631_),
    .D(_0632_),
    .X(_0635_));
 sky130_fd_sc_hd__and2_1 _2096_ (.A(_0634_),
    .B(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__clkbuf_1 _2097_ (.A(_0636_),
    .X(\po_0.alu_0._10_[7] ));
 sky130_fd_sc_hd__clkbuf_2 _2098_ (.A(net49),
    .X(_0637_));
 sky130_fd_sc_hd__nand2_1 _2099_ (.A(_0637_),
    .B(\po_0._1_[8] ),
    .Y(_0638_));
 sky130_fd_sc_hd__or2_1 _2100_ (.A(_0637_),
    .B(\po_0._1_[8] ),
    .X(_0639_));
 sky130_fd_sc_hd__nand2_1 _2101_ (.A(_0638_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__or2b_1 _2102_ (.A(\po_0._1_[7] ),
    .B_N(net85),
    .X(_0641_));
 sky130_fd_sc_hd__nand2_1 _2103_ (.A(_0634_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__xor2_1 _2104_ (.A(_0640_),
    .B(_0642_),
    .X(\po_0.alu_0._10_[8] ));
 sky130_fd_sc_hd__xor2_2 _2105_ (.A(net50),
    .B(\po_0._1_[9] ),
    .X(_0643_));
 sky130_fd_sc_hd__and2b_1 _2106_ (.A_N(\po_0._1_[8] ),
    .B(_0637_),
    .X(_0644_));
 sky130_fd_sc_hd__a21oi_1 _2107_ (.A1(_0640_),
    .A2(_0642_),
    .B1(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__xor2_1 _2108_ (.A(_0643_),
    .B(_0645_),
    .X(\po_0.alu_0._10_[9] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2109_ (.A(net36),
    .X(_0646_));
 sky130_fd_sc_hd__or2b_1 _2110_ (.A(_0646_),
    .B_N(\po_0._1_[10] ),
    .X(_0647_));
 sky130_fd_sc_hd__or2b_1 _2111_ (.A(\po_0._1_[10] ),
    .B_N(_0646_),
    .X(_0648_));
 sky130_fd_sc_hd__nand2_1 _2112_ (.A(_0647_),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__clkbuf_2 _2113_ (.A(net50),
    .X(_0650_));
 sky130_fd_sc_hd__or2b_1 _2114_ (.A(\po_0._1_[9] ),
    .B_N(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__or3b_1 _2115_ (.A(\po_0._1_[8] ),
    .B(_0643_),
    .C_N(_0637_),
    .X(_0652_));
 sky130_fd_sc_hd__xnor2_1 _2116_ (.A(_0650_),
    .B(\po_0._1_[9] ),
    .Y(_0653_));
 sky130_fd_sc_hd__nand3_1 _2117_ (.A(_0640_),
    .B(_0642_),
    .C(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__nand3_1 _2118_ (.A(_0651_),
    .B(_0652_),
    .C(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__xnor2_1 _2119_ (.A(_0649_),
    .B(_0655_),
    .Y(\po_0.alu_0._10_[10] ));
 sky130_fd_sc_hd__nor2_1 _2120_ (.A(net84),
    .B(\po_0._1_[11] ),
    .Y(_0656_));
 sky130_fd_sc_hd__and2_1 _2121_ (.A(net84),
    .B(\po_0._1_[11] ),
    .X(_0657_));
 sky130_fd_sc_hd__nor2_2 _2122_ (.A(_0656_),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__and3_1 _2123_ (.A(_0648_),
    .B(_0651_),
    .C(_0652_),
    .X(_0659_));
 sky130_fd_sc_hd__a21boi_1 _2124_ (.A1(_0654_),
    .A2(_0659_),
    .B1_N(_0647_),
    .Y(_0660_));
 sky130_fd_sc_hd__xnor2_1 _2125_ (.A(_0658_),
    .B(_0660_),
    .Y(\po_0.alu_0._10_[11] ));
 sky130_fd_sc_hd__and2_1 _2126_ (.A(net83),
    .B(\po_0._1_[12] ),
    .X(_0661_));
 sky130_fd_sc_hd__nor2_1 _2127_ (.A(net83),
    .B(\po_0._1_[12] ),
    .Y(_0662_));
 sky130_fd_sc_hd__or2_1 _2128_ (.A(_0661_),
    .B(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2129_ (.A(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__inv_2 _2130_ (.A(\po_0._1_[11] ),
    .Y(_0665_));
 sky130_fd_sc_hd__nor2_1 _2131_ (.A(_0658_),
    .B(_0659_),
    .Y(_0666_));
 sky130_fd_sc_hd__a22o_1 _2132_ (.A1(net84),
    .A2(_0665_),
    .B1(_0666_),
    .B2(_0647_),
    .X(_0667_));
 sky130_fd_sc_hd__and2_1 _2133_ (.A(_0638_),
    .B(_0639_),
    .X(_0668_));
 sky130_fd_sc_hd__or4_1 _2134_ (.A(_0668_),
    .B(_0643_),
    .C(_0649_),
    .D(_0658_),
    .X(_0669_));
 sky130_fd_sc_hd__a21oi_2 _2135_ (.A1(_0634_),
    .A2(_0641_),
    .B1(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__nor2_1 _2136_ (.A(_0667_),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__xnor2_1 _2137_ (.A(_0664_),
    .B(_0671_),
    .Y(\po_0.alu_0._10_[12] ));
 sky130_fd_sc_hd__inv_2 _2138_ (.A(net83),
    .Y(_0672_));
 sky130_fd_sc_hd__nor2_1 _2139_ (.A(net39),
    .B(\po_0._1_[13] ),
    .Y(_0673_));
 sky130_fd_sc_hd__and2_1 _2140_ (.A(net39),
    .B(\po_0._1_[13] ),
    .X(_0674_));
 sky130_fd_sc_hd__nor2_1 _2141_ (.A(_0673_),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__o21ai_1 _2142_ (.A1(_0667_),
    .A2(_0670_),
    .B1(_0664_),
    .Y(_0676_));
 sky130_fd_sc_hd__o211ai_1 _2143_ (.A1(_0672_),
    .A2(\po_0._1_[12] ),
    .B1(_0675_),
    .C1(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__o21ai_1 _2144_ (.A1(_0673_),
    .A2(_0674_),
    .B1(_0664_),
    .Y(_0678_));
 sky130_fd_sc_hd__o21bai_2 _2145_ (.A1(_0667_),
    .A2(_0670_),
    .B1_N(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__o311a_1 _2146_ (.A1(_0672_),
    .A2(\po_0._1_[12] ),
    .A3(_0675_),
    .B1(_0677_),
    .C1(_0679_),
    .X(\po_0.alu_0._10_[13] ));
 sky130_fd_sc_hd__clkbuf_2 _2147_ (.A(net40),
    .X(_0680_));
 sky130_fd_sc_hd__nand2_1 _2148_ (.A(_0680_),
    .B(\po_0._1_[14] ),
    .Y(_0681_));
 sky130_fd_sc_hd__or2_1 _2149_ (.A(_0680_),
    .B(\po_0._1_[14] ),
    .X(_0682_));
 sky130_fd_sc_hd__inv_2 _2150_ (.A(net39),
    .Y(_0683_));
 sky130_fd_sc_hd__or3_1 _2151_ (.A(_0672_),
    .B(\po_0._1_[12] ),
    .C(_0675_),
    .X(_0684_));
 sky130_fd_sc_hd__o21a_1 _2152_ (.A1(_0683_),
    .A2(\po_0._1_[13] ),
    .B1(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__a22oi_1 _2153_ (.A1(_0681_),
    .A2(_0682_),
    .B1(_0679_),
    .B2(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__and4_1 _2154_ (.A(_0679_),
    .B(_0681_),
    .C(_0682_),
    .D(_0685_),
    .X(_0687_));
 sky130_fd_sc_hd__nor2_1 _2155_ (.A(_0686_),
    .B(_0687_),
    .Y(\po_0.alu_0._10_[14] ));
 sky130_fd_sc_hd__inv_2 _2156_ (.A(_0680_),
    .Y(_0688_));
 sky130_fd_sc_hd__and2b_1 _2157_ (.A_N(\po_0._1_[15] ),
    .B(net41),
    .X(_0689_));
 sky130_fd_sc_hd__and2b_1 _2158_ (.A_N(net41),
    .B(\po_0._1_[15] ),
    .X(_0690_));
 sky130_fd_sc_hd__nor2_1 _2159_ (.A(_0689_),
    .B(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__and2_1 _2160_ (.A(_0680_),
    .B(\po_0._1_[14] ),
    .X(_0692_));
 sky130_fd_sc_hd__nor2_1 _2161_ (.A(_0680_),
    .B(\po_0._1_[14] ),
    .Y(_0693_));
 sky130_fd_sc_hd__o2bb2ai_1 _2162_ (.A1_N(_0685_),
    .A2_N(_0679_),
    .B1(_0692_),
    .B2(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__o211ai_1 _2163_ (.A1(_0688_),
    .A2(\po_0._1_[14] ),
    .B1(_0691_),
    .C1(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__nor2_1 _2164_ (.A(\po_0._1_[14] ),
    .B(_0688_),
    .Y(_0696_));
 sky130_fd_sc_hd__o22ai_1 _2165_ (.A1(_0689_),
    .A2(_0690_),
    .B1(_0696_),
    .B2(_0686_),
    .Y(_0697_));
 sky130_fd_sc_hd__nand2_1 _2166_ (.A(_0695_),
    .B(_0697_),
    .Y(\po_0.alu_0._10_[15] ));
 sky130_fd_sc_hd__inv_2 _2167_ (.A(\po_0.muxf_0.s1 ),
    .Y(_0698_));
 sky130_fd_sc_hd__and2_1 _2168_ (.A(_0698_),
    .B(\po_0.muxf_0.s0 ),
    .X(_0699_));
 sky130_fd_sc_hd__buf_2 _2169_ (.A(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__buf_2 _2170_ (.A(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__nor2_1 _2171_ (.A(\po_0.muxf_0.s0 ),
    .B(_0698_),
    .Y(_0702_));
 sky130_fd_sc_hd__buf_2 _2172_ (.A(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__buf_2 _2173_ (.A(\po_0.muxf_0.rf_w_data[0] ),
    .X(_0704_));
 sky130_fd_sc_hd__nor2_2 _2174_ (.A(_1404_),
    .B(_1401_),
    .Y(_0705_));
 sky130_fd_sc_hd__clkbuf_2 _2175_ (.A(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__or2b_1 _2176_ (.A(_1404_),
    .B_N(\po_0.alu_0.s0 ),
    .X(_0707_));
 sky130_fd_sc_hd__buf_2 _2177_ (.A(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _2178_ (.A0(\po_0.alu_0._10_[0] ),
    .A1(\po_0.alu_0._11_[0] ),
    .S(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__or3_1 _2179_ (.A(net87),
    .B(_1404_),
    .C(_1401_),
    .X(_0710_));
 sky130_fd_sc_hd__nor2_1 _2180_ (.A(_0699_),
    .B(_0702_),
    .Y(_0711_));
 sky130_fd_sc_hd__o211a_1 _2181_ (.A1(_0706_),
    .A2(_0709_),
    .B1(_0710_),
    .C1(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__a221o_2 _2182_ (.A1(net1),
    .A2(_0701_),
    .B1(_0703_),
    .B2(_0704_),
    .C1(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2183_ (.A(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2184_ (.A(\po_0.regf_0.w_addr[3] ),
    .X(_0715_));
 sky130_fd_sc_hd__clkbuf_2 _2185_ (.A(\po_0.regf_0.w_wr ),
    .X(_0716_));
 sky130_fd_sc_hd__and2_1 _2186_ (.A(\po_0.regf_0.w_addr[1] ),
    .B(\po_0.regf_0.w_addr[0] ),
    .X(_0717_));
 sky130_fd_sc_hd__clkbuf_2 _2187_ (.A(\po_0.regf_0.w_addr[2] ),
    .X(_0718_));
 sky130_fd_sc_hd__nand4b_4 _2188_ (.A_N(_0715_),
    .B(_0716_),
    .C(_0717_),
    .D(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__buf_2 _2189_ (.A(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _2190_ (.A0(_0714_),
    .A1(\po_0.regf_0.rf[7][0] ),
    .S(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__clkbuf_1 _2191_ (.A(_0721_),
    .X(_0016_));
 sky130_fd_sc_hd__clkbuf_2 _2192_ (.A(\po_0.muxf_0.s0 ),
    .X(_0722_));
 sky130_fd_sc_hd__clkbuf_2 _2193_ (.A(_0698_),
    .X(_0723_));
 sky130_fd_sc_hd__buf_2 _2194_ (.A(\po_0.muxf_0.rf_w_data[1] ),
    .X(_0724_));
 sky130_fd_sc_hd__and2b_1 _2195_ (.A_N(\po_0.alu_0.s1 ),
    .B(\po_0.alu_0.s0 ),
    .X(_0725_));
 sky130_fd_sc_hd__a2bb2o_1 _2196_ (.A1_N(_0581_),
    .A2_N(_0582_),
    .B1(\po_0._1_[0] ),
    .B2(net87),
    .X(_0726_));
 sky130_fd_sc_hd__o311a_1 _2197_ (.A1(_1429_),
    .A2(_0581_),
    .A3(_0582_),
    .B1(_0725_),
    .C1(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__a221o_1 _2198_ (.A1(_1405_),
    .A2(\po_0.alu_0._11_[1] ),
    .B1(_0705_),
    .B2(net86),
    .C1(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__clkbuf_2 _2199_ (.A(_0711_),
    .X(_0729_));
 sky130_fd_sc_hd__a22o_1 _2200_ (.A1(_0724_),
    .A2(_0702_),
    .B1(_0728_),
    .B2(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__a31o_2 _2201_ (.A1(_0722_),
    .A2(_0723_),
    .A3(net8),
    .B1(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2202_ (.A(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _2203_ (.A0(_0732_),
    .A1(\po_0.regf_0.rf[7][1] ),
    .S(_0720_),
    .X(_0733_));
 sky130_fd_sc_hd__clkbuf_1 _2204_ (.A(_0733_),
    .X(_0017_));
 sky130_fd_sc_hd__clkbuf_4 _2205_ (.A(\po_0.muxf_0.rf_w_data[2] ),
    .X(_0734_));
 sky130_fd_sc_hd__nand2_1 _2206_ (.A(net86),
    .B(\po_0._1_[1] ),
    .Y(_0735_));
 sky130_fd_sc_hd__o21ai_2 _2207_ (.A1(_1429_),
    .A2(_0582_),
    .B1(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__a21oi_1 _2208_ (.A1(_0590_),
    .A2(_0736_),
    .B1(_0707_),
    .Y(_0737_));
 sky130_fd_sc_hd__o31a_1 _2209_ (.A1(_0592_),
    .A2(_0593_),
    .A3(_0736_),
    .B1(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__a221o_1 _2210_ (.A1(_1405_),
    .A2(\po_0.alu_0._11_[2] ),
    .B1(_0705_),
    .B2(_0588_),
    .C1(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__a22o_1 _2211_ (.A1(_0734_),
    .A2(_0702_),
    .B1(_0739_),
    .B2(_0729_),
    .X(_0740_));
 sky130_fd_sc_hd__a31o_2 _2212_ (.A1(_0722_),
    .A2(_0723_),
    .A3(net9),
    .B1(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2213_ (.A(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _2214_ (.A0(_0742_),
    .A1(\po_0.regf_0.rf[7][2] ),
    .S(_0720_),
    .X(_0743_));
 sky130_fd_sc_hd__clkbuf_1 _2215_ (.A(_0743_),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_4 _2216_ (.A(\po_0.muxf_0.rf_w_data[3] ),
    .X(_0744_));
 sky130_fd_sc_hd__clkbuf_2 _2217_ (.A(_1405_),
    .X(_0745_));
 sky130_fd_sc_hd__o21a_1 _2218_ (.A1(_0592_),
    .A2(_0593_),
    .B1(_0736_),
    .X(_0746_));
 sky130_fd_sc_hd__or3_1 _2219_ (.A(_0587_),
    .B(_0602_),
    .C(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__o21ai_1 _2220_ (.A1(_0587_),
    .A2(_0746_),
    .B1(_0602_),
    .Y(_0748_));
 sky130_fd_sc_hd__and3_1 _2221_ (.A(_0747_),
    .B(_0725_),
    .C(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__a211o_1 _2222_ (.A1(_1405_),
    .A2(\po_0.alu_0._11_[3] ),
    .B1(_0706_),
    .C1(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__o311a_1 _2223_ (.A1(_0598_),
    .A2(_0745_),
    .A3(_1402_),
    .B1(_0711_),
    .C1(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__a221o_4 _2224_ (.A1(net10),
    .A2(_0700_),
    .B1(_0703_),
    .B2(_0744_),
    .C1(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2225_ (.A(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _2226_ (.A0(_0753_),
    .A1(\po_0.regf_0.rf[7][3] ),
    .S(_0720_),
    .X(_0754_));
 sky130_fd_sc_hd__clkbuf_1 _2227_ (.A(_0754_),
    .X(_0019_));
 sky130_fd_sc_hd__a22o_1 _2228_ (.A1(_0588_),
    .A2(\po_0._1_[2] ),
    .B1(\po_0._1_[3] ),
    .B2(net44),
    .X(_0755_));
 sky130_fd_sc_hd__o22a_1 _2229_ (.A1(_0598_),
    .A2(\po_0._1_[3] ),
    .B1(_0755_),
    .B2(_0746_),
    .X(_0756_));
 sky130_fd_sc_hd__o221ai_4 _2230_ (.A1(_0598_),
    .A2(\po_0._1_[3] ),
    .B1(_0755_),
    .B2(_0746_),
    .C1(_0610_),
    .Y(_0757_));
 sky130_fd_sc_hd__buf_2 _2231_ (.A(_0725_),
    .X(_0758_));
 sky130_fd_sc_hd__o211a_1 _2232_ (.A1(_0610_),
    .A2(_0756_),
    .B1(_0757_),
    .C1(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__a221o_1 _2233_ (.A1(_1405_),
    .A2(\po_0.alu_0._11_[4] ),
    .B1(_0705_),
    .B2(_0605_),
    .C1(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__a22o_1 _2234_ (.A1(_0557_),
    .A2(_0702_),
    .B1(_0760_),
    .B2(_0729_),
    .X(_0761_));
 sky130_fd_sc_hd__a31o_2 _2235_ (.A1(_0722_),
    .A2(_0723_),
    .A3(net11),
    .B1(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2236_ (.A(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__mux2_1 _2237_ (.A0(_0763_),
    .A1(\po_0.regf_0.rf[7][4] ),
    .S(_0720_),
    .X(_0764_));
 sky130_fd_sc_hd__clkbuf_1 _2238_ (.A(_0764_),
    .X(_0020_));
 sky130_fd_sc_hd__nand2_1 _2239_ (.A(_0605_),
    .B(\po_0._1_[4] ),
    .Y(_0765_));
 sky130_fd_sc_hd__or2_1 _2240_ (.A(_0614_),
    .B(_0615_),
    .X(_0766_));
 sky130_fd_sc_hd__a21oi_1 _2241_ (.A1(_0765_),
    .A2(_0757_),
    .B1(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__a31o_1 _2242_ (.A1(_0765_),
    .A2(_0766_),
    .A3(_0757_),
    .B1(_0707_),
    .X(_0768_));
 sky130_fd_sc_hd__nor2_1 _2243_ (.A(_0767_),
    .B(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__a211o_1 _2244_ (.A1(\po_0.alu_0._11_[5] ),
    .A2(_0708_),
    .B1(_0705_),
    .C1(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__o311a_1 _2245_ (.A1(_0613_),
    .A2(_0745_),
    .A3(_1401_),
    .B1(_0711_),
    .C1(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__a221o_4 _2246_ (.A1(net12),
    .A2(_0700_),
    .B1(_0703_),
    .B2(_0566_),
    .C1(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2247_ (.A(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _2248_ (.A0(_0773_),
    .A1(\po_0.regf_0.rf[7][5] ),
    .S(_0720_),
    .X(_0774_));
 sky130_fd_sc_hd__clkbuf_1 _2249_ (.A(_0774_),
    .X(_0021_));
 sky130_fd_sc_hd__clkbuf_2 _2250_ (.A(_1404_),
    .X(_0775_));
 sky130_fd_sc_hd__a22o_1 _2251_ (.A1(_0775_),
    .A2(\po_0.alu_0._11_[6] ),
    .B1(_0706_),
    .B2(_0620_),
    .X(_0776_));
 sky130_fd_sc_hd__a22oi_2 _2252_ (.A1(_0605_),
    .A2(\po_0._1_[4] ),
    .B1(\po_0._1_[5] ),
    .B2(_0613_),
    .Y(_0777_));
 sky130_fd_sc_hd__o2bb2a_1 _2253_ (.A1_N(_0777_),
    .A2_N(_0757_),
    .B1(\po_0._1_[5] ),
    .B2(_0613_),
    .X(_0778_));
 sky130_fd_sc_hd__a21oi_1 _2254_ (.A1(_0778_),
    .A2(_0628_),
    .B1(_1404_),
    .Y(_0779_));
 sky130_fd_sc_hd__o211a_1 _2255_ (.A1(_0778_),
    .A2(_0628_),
    .B1(_1401_),
    .C1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__o21a_1 _2256_ (.A1(_0776_),
    .A2(_0780_),
    .B1(_0729_),
    .X(_0781_));
 sky130_fd_sc_hd__a221o_4 _2257_ (.A1(net13),
    .A2(_0700_),
    .B1(_0703_),
    .B2(_0568_),
    .C1(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2258_ (.A(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__buf_2 _2259_ (.A(_0719_),
    .X(_0784_));
 sky130_fd_sc_hd__mux2_1 _2260_ (.A0(_0783_),
    .A1(\po_0.regf_0.rf[7][6] ),
    .S(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__clkbuf_1 _2261_ (.A(_0785_),
    .X(_0022_));
 sky130_fd_sc_hd__a221o_1 _2262_ (.A1(_0620_),
    .A2(_0621_),
    .B1(_0778_),
    .B2(_0628_),
    .C1(_0633_),
    .X(_0786_));
 sky130_fd_sc_hd__or2_1 _2263_ (.A(_0622_),
    .B(_0623_),
    .X(_0787_));
 sky130_fd_sc_hd__a211oi_1 _2264_ (.A1(_0757_),
    .A2(_0777_),
    .B1(_0614_),
    .C1(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__o21ai_1 _2265_ (.A1(_0622_),
    .A2(_0788_),
    .B1(_0633_),
    .Y(_0789_));
 sky130_fd_sc_hd__a21o_1 _2266_ (.A1(_0775_),
    .A2(\po_0.alu_0._11_[7] ),
    .B1(_0706_),
    .X(_0790_));
 sky130_fd_sc_hd__a31o_1 _2267_ (.A1(_0786_),
    .A2(_0789_),
    .A3(_0758_),
    .B1(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__or3_1 _2268_ (.A(net85),
    .B(_0775_),
    .C(_1401_),
    .X(_0792_));
 sky130_fd_sc_hd__buf_2 _2269_ (.A(_0711_),
    .X(_0793_));
 sky130_fd_sc_hd__a22o_1 _2270_ (.A1(net14),
    .A2(_0700_),
    .B1(_0703_),
    .B2(_0570_),
    .X(_0794_));
 sky130_fd_sc_hd__a31o_2 _2271_ (.A1(_0791_),
    .A2(_0792_),
    .A3(_0793_),
    .B1(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2272_ (.A(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _2273_ (.A0(_0796_),
    .A1(\po_0.regf_0.rf[7][7] ),
    .S(_0784_),
    .X(_0797_));
 sky130_fd_sc_hd__clkbuf_1 _2274_ (.A(_0797_),
    .X(_0023_));
 sky130_fd_sc_hd__nor2_1 _2275_ (.A(_0614_),
    .B(_0615_),
    .Y(_0798_));
 sky130_fd_sc_hd__nand4_2 _2276_ (.A(_0610_),
    .B(_0798_),
    .C(_0628_),
    .D(_0633_),
    .Y(_0799_));
 sky130_fd_sc_hd__a21oi_1 _2277_ (.A1(_0590_),
    .A2(_0736_),
    .B1(_0755_),
    .Y(_0800_));
 sky130_fd_sc_hd__or2_1 _2278_ (.A(net48),
    .B(\po_0._1_[7] ),
    .X(_0801_));
 sky130_fd_sc_hd__nand2_1 _2279_ (.A(_0620_),
    .B(_0621_),
    .Y(_0802_));
 sky130_fd_sc_hd__o31ai_1 _2280_ (.A1(_0614_),
    .A2(_0623_),
    .A3(_0777_),
    .B1(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__a21oi_2 _2281_ (.A1(_0801_),
    .A2(_0803_),
    .B1(_0632_),
    .Y(_0804_));
 sky130_fd_sc_hd__o31ai_4 _2282_ (.A1(_0600_),
    .A2(_0799_),
    .A3(_0800_),
    .B1(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__a21o_1 _2283_ (.A1(_0638_),
    .A2(_0639_),
    .B1(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__nand2_1 _2284_ (.A(_0805_),
    .B(_0668_),
    .Y(_0807_));
 sky130_fd_sc_hd__a22o_1 _2285_ (.A1(_0775_),
    .A2(\po_0.alu_0._11_[8] ),
    .B1(_0706_),
    .B2(_0637_),
    .X(_0808_));
 sky130_fd_sc_hd__a31o_1 _2286_ (.A1(_0806_),
    .A2(_0807_),
    .A3(_0758_),
    .B1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__a22o_2 _2287_ (.A1(net15),
    .A2(_0701_),
    .B1(_0809_),
    .B2(_0793_),
    .X(_0810_));
 sky130_fd_sc_hd__clkbuf_2 _2288_ (.A(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _2289_ (.A0(_0811_),
    .A1(\po_0.regf_0.rf[7][8] ),
    .S(_0784_),
    .X(_0812_));
 sky130_fd_sc_hd__clkbuf_1 _2290_ (.A(_0812_),
    .X(_0024_));
 sky130_fd_sc_hd__a21oi_1 _2291_ (.A1(_0638_),
    .A2(_0807_),
    .B1(_0653_),
    .Y(_0813_));
 sky130_fd_sc_hd__and3_1 _2292_ (.A(_0638_),
    .B(_0653_),
    .C(_0807_),
    .X(_0814_));
 sky130_fd_sc_hd__clkbuf_2 _2293_ (.A(_0705_),
    .X(_0815_));
 sky130_fd_sc_hd__a21oi_1 _2294_ (.A1(_1406_),
    .A2(\po_0.alu_0._11_[9] ),
    .B1(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__o31ai_1 _2295_ (.A1(_0813_),
    .A2(_0708_),
    .A3(_0814_),
    .B1(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__o31a_1 _2296_ (.A1(_0650_),
    .A2(_1406_),
    .A3(_1402_),
    .B1(_0793_),
    .X(_0818_));
 sky130_fd_sc_hd__a32o_4 _2297_ (.A1(_0722_),
    .A2(_0723_),
    .A3(net16),
    .B1(_0817_),
    .B2(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2298_ (.A(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _2299_ (.A0(_0820_),
    .A1(\po_0.regf_0.rf[7][9] ),
    .S(_0784_),
    .X(_0821_));
 sky130_fd_sc_hd__clkbuf_1 _2300_ (.A(_0821_),
    .X(_0025_));
 sky130_fd_sc_hd__a22oi_2 _2301_ (.A1(_0637_),
    .A2(\po_0._1_[8] ),
    .B1(\po_0._1_[9] ),
    .B2(_0650_),
    .Y(_0822_));
 sky130_fd_sc_hd__a2bb2o_1 _2302_ (.A1_N(_0650_),
    .A2_N(\po_0._1_[9] ),
    .B1(_0647_),
    .B2(_0648_),
    .X(_0823_));
 sky130_fd_sc_hd__a21oi_1 _2303_ (.A1(_0807_),
    .A2(_0822_),
    .B1(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__a2bb2o_1 _2304_ (.A1_N(_0650_),
    .A2_N(\po_0._1_[9] ),
    .B1(_0822_),
    .B2(_0807_),
    .X(_0825_));
 sky130_fd_sc_hd__and3_1 _2305_ (.A(_0825_),
    .B(_0648_),
    .C(_0647_),
    .X(_0826_));
 sky130_fd_sc_hd__a22oi_1 _2306_ (.A1(_0745_),
    .A2(\po_0.alu_0._11_[10] ),
    .B1(_0815_),
    .B2(_0646_),
    .Y(_0827_));
 sky130_fd_sc_hd__o31ai_1 _2307_ (.A1(_0824_),
    .A2(_0708_),
    .A3(_0826_),
    .B1(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__a22o_2 _2308_ (.A1(net2),
    .A2(_0701_),
    .B1(_0828_),
    .B2(_0793_),
    .X(_0829_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2309_ (.A(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_1 _2310_ (.A0(_0830_),
    .A1(\po_0.regf_0.rf[7][10] ),
    .S(_0784_),
    .X(_0831_));
 sky130_fd_sc_hd__clkbuf_1 _2311_ (.A(_0831_),
    .X(_0026_));
 sky130_fd_sc_hd__a211o_1 _2312_ (.A1(_0646_),
    .A2(\po_0._1_[10] ),
    .B1(_0658_),
    .C1(_0824_),
    .X(_0832_));
 sky130_fd_sc_hd__and2_1 _2313_ (.A(_0646_),
    .B(\po_0._1_[10] ),
    .X(_0833_));
 sky130_fd_sc_hd__o21ai_1 _2314_ (.A1(_0833_),
    .A2(_0824_),
    .B1(_0658_),
    .Y(_0834_));
 sky130_fd_sc_hd__a21o_1 _2315_ (.A1(_0775_),
    .A2(\po_0.alu_0._11_[11] ),
    .B1(_0706_),
    .X(_0835_));
 sky130_fd_sc_hd__a31o_1 _2316_ (.A1(_0832_),
    .A2(_0758_),
    .A3(_0834_),
    .B1(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__o31a_1 _2317_ (.A1(net84),
    .A2(_1406_),
    .A3(_1402_),
    .B1(_0729_),
    .X(_0837_));
 sky130_fd_sc_hd__a32o_4 _2318_ (.A1(_0722_),
    .A2(_0723_),
    .A3(net3),
    .B1(_0836_),
    .B2(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2319_ (.A(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _2320_ (.A0(_0839_),
    .A1(\po_0.regf_0.rf[7][11] ),
    .S(_0784_),
    .X(_0840_));
 sky130_fd_sc_hd__clkbuf_1 _2321_ (.A(_0840_),
    .X(_0027_));
 sky130_fd_sc_hd__a22o_1 _2322_ (.A1(_0646_),
    .A2(\po_0._1_[10] ),
    .B1(\po_0._1_[11] ),
    .B2(net84),
    .X(_0841_));
 sky130_fd_sc_hd__o21ba_1 _2323_ (.A1(_0822_),
    .A2(_0823_),
    .B1_N(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__and4_1 _2324_ (.A(_0668_),
    .B(_0643_),
    .C(_0649_),
    .D(_0658_),
    .X(_0843_));
 sky130_fd_sc_hd__a2bb2oi_1 _2325_ (.A1_N(_0656_),
    .A2_N(_0842_),
    .B1(_0843_),
    .B2(_0805_),
    .Y(_0844_));
 sky130_fd_sc_hd__a21oi_1 _2326_ (.A1(_0844_),
    .A2(_0664_),
    .B1(_0708_),
    .Y(_0845_));
 sky130_fd_sc_hd__o31a_1 _2327_ (.A1(_0661_),
    .A2(_0662_),
    .A3(_0844_),
    .B1(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__a221o_1 _2328_ (.A1(_0745_),
    .A2(\po_0.alu_0._11_[12] ),
    .B1(_0815_),
    .B2(net83),
    .C1(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__a22o_2 _2329_ (.A1(net4),
    .A2(_0701_),
    .B1(_0847_),
    .B2(_0793_),
    .X(_0848_));
 sky130_fd_sc_hd__clkbuf_2 _2330_ (.A(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _2331_ (.A0(_0849_),
    .A1(\po_0.regf_0.rf[7][12] ),
    .S(_0719_),
    .X(_0850_));
 sky130_fd_sc_hd__clkbuf_1 _2332_ (.A(_0850_),
    .X(_0028_));
 sky130_fd_sc_hd__a211o_1 _2333_ (.A1(_0683_),
    .A2(_0815_),
    .B1(_0703_),
    .C1(_0700_),
    .X(_0851_));
 sky130_fd_sc_hd__nand2_1 _2334_ (.A(net38),
    .B(\po_0._1_[12] ),
    .Y(_0852_));
 sky130_fd_sc_hd__o21ai_1 _2335_ (.A1(_0664_),
    .A2(_0844_),
    .B1(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__o21a_1 _2336_ (.A1(_0675_),
    .A2(_0853_),
    .B1(_0758_),
    .X(_0854_));
 sky130_fd_sc_hd__nand2_1 _2337_ (.A(_0853_),
    .B(_0675_),
    .Y(_0855_));
 sky130_fd_sc_hd__a21o_1 _2338_ (.A1(_1406_),
    .A2(\po_0.alu_0._11_[13] ),
    .B1(_0815_),
    .X(_0856_));
 sky130_fd_sc_hd__a21oi_1 _2339_ (.A1(_0854_),
    .A2(_0855_),
    .B1(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__o2bb2ai_4 _2340_ (.A1_N(net5),
    .A2_N(_0701_),
    .B1(_0851_),
    .B2(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2341_ (.A(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__mux2_1 _2342_ (.A0(_0859_),
    .A1(\po_0.regf_0.rf[7][13] ),
    .S(_0719_),
    .X(_0860_));
 sky130_fd_sc_hd__clkbuf_1 _2343_ (.A(_0860_),
    .X(_0029_));
 sky130_fd_sc_hd__o2bb2ai_1 _2344_ (.A1_N(_0843_),
    .A2_N(_0805_),
    .B1(_0656_),
    .B2(_0842_),
    .Y(_0861_));
 sky130_fd_sc_hd__nor4_1 _2345_ (.A(_0661_),
    .B(_0662_),
    .C(_0673_),
    .D(_0674_),
    .Y(_0862_));
 sky130_fd_sc_hd__nand2_1 _2346_ (.A(_0861_),
    .B(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__o21ba_1 _2347_ (.A1(_0852_),
    .A2(_0673_),
    .B1_N(_0674_),
    .X(_0864_));
 sky130_fd_sc_hd__nand2_1 _2348_ (.A(_0681_),
    .B(_0682_),
    .Y(_0865_));
 sky130_fd_sc_hd__a21oi_1 _2349_ (.A1(_0863_),
    .A2(_0864_),
    .B1(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__a31o_1 _2350_ (.A1(_0865_),
    .A2(_0863_),
    .A3(_0864_),
    .B1(_0708_),
    .X(_0867_));
 sky130_fd_sc_hd__a22oi_1 _2351_ (.A1(_0745_),
    .A2(\po_0.alu_0._11_[14] ),
    .B1(_0815_),
    .B2(_0680_),
    .Y(_0868_));
 sky130_fd_sc_hd__o21ai_1 _2352_ (.A1(_0866_),
    .A2(_0867_),
    .B1(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__a22o_2 _2353_ (.A1(net6),
    .A2(_0701_),
    .B1(_0869_),
    .B2(_0793_),
    .X(_0870_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2354_ (.A(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_1 _2355_ (.A0(_0871_),
    .A1(\po_0.regf_0.rf[7][14] ),
    .S(_0719_),
    .X(_0872_));
 sky130_fd_sc_hd__clkbuf_1 _2356_ (.A(_0872_),
    .X(_0030_));
 sky130_fd_sc_hd__o21ai_1 _2357_ (.A1(_0692_),
    .A2(_0866_),
    .B1(_0691_),
    .Y(_0873_));
 sky130_fd_sc_hd__a21boi_1 _2358_ (.A1(_0861_),
    .A2(_0862_),
    .B1_N(_0864_),
    .Y(_0874_));
 sky130_fd_sc_hd__o221ai_1 _2359_ (.A1(_0689_),
    .A2(_0690_),
    .B1(_0865_),
    .B2(_0874_),
    .C1(_0681_),
    .Y(_0875_));
 sky130_fd_sc_hd__nand3_1 _2360_ (.A(_0873_),
    .B(_0758_),
    .C(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__or2b_1 _2361_ (.A(\po_0.alu_0._11_[15] ),
    .B_N(_0775_),
    .X(_0877_));
 sky130_fd_sc_hd__o311a_1 _2362_ (.A1(net41),
    .A2(_0745_),
    .A3(_1402_),
    .B1(_0877_),
    .C1(_0729_),
    .X(_0878_));
 sky130_fd_sc_hd__a32o_2 _2363_ (.A1(\po_0.muxf_0.s0 ),
    .A2(_0698_),
    .A3(net7),
    .B1(_0876_),
    .B2(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2364_ (.A(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__mux2_1 _2365_ (.A0(_0880_),
    .A1(\po_0.regf_0.rf[7][15] ),
    .S(_0719_),
    .X(_0881_));
 sky130_fd_sc_hd__clkbuf_1 _2366_ (.A(_0881_),
    .X(_0031_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2367_ (.A(\po_0.regf_0.w_addr[3] ),
    .X(_0882_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2368_ (.A(\po_0.regf_0.w_addr[0] ),
    .X(_0883_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2369_ (.A(\po_0.regf_0.w_addr[1] ),
    .X(_0884_));
 sky130_fd_sc_hd__and2b_1 _2370_ (.A_N(_0883_),
    .B(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2371_ (.A(\po_0.regf_0.w_addr[2] ),
    .X(_0886_));
 sky130_fd_sc_hd__and4b_4 _2372_ (.A_N(_0882_),
    .B(_0716_),
    .C(_0885_),
    .D(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__buf_2 _2373_ (.A(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _2374_ (.A0(\po_0.regf_0.rf[6][0] ),
    .A1(_0714_),
    .S(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__clkbuf_1 _2375_ (.A(_0889_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2376_ (.A0(\po_0.regf_0.rf[6][1] ),
    .A1(_0732_),
    .S(_0888_),
    .X(_0890_));
 sky130_fd_sc_hd__clkbuf_1 _2377_ (.A(_0890_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _2378_ (.A0(\po_0.regf_0.rf[6][2] ),
    .A1(_0742_),
    .S(_0888_),
    .X(_0891_));
 sky130_fd_sc_hd__clkbuf_1 _2379_ (.A(_0891_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2380_ (.A0(\po_0.regf_0.rf[6][3] ),
    .A1(_0753_),
    .S(_0888_),
    .X(_0892_));
 sky130_fd_sc_hd__clkbuf_1 _2381_ (.A(_0892_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2382_ (.A0(\po_0.regf_0.rf[6][4] ),
    .A1(_0763_),
    .S(_0888_),
    .X(_0893_));
 sky130_fd_sc_hd__clkbuf_1 _2383_ (.A(_0893_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2384_ (.A0(\po_0.regf_0.rf[6][5] ),
    .A1(_0773_),
    .S(_0888_),
    .X(_0894_));
 sky130_fd_sc_hd__clkbuf_1 _2385_ (.A(_0894_),
    .X(_0037_));
 sky130_fd_sc_hd__buf_2 _2386_ (.A(_0887_),
    .X(_0895_));
 sky130_fd_sc_hd__mux2_1 _2387_ (.A0(\po_0.regf_0.rf[6][6] ),
    .A1(_0783_),
    .S(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__clkbuf_1 _2388_ (.A(_0896_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2389_ (.A0(\po_0.regf_0.rf[6][7] ),
    .A1(_0796_),
    .S(_0895_),
    .X(_0897_));
 sky130_fd_sc_hd__clkbuf_1 _2390_ (.A(_0897_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2391_ (.A0(\po_0.regf_0.rf[6][8] ),
    .A1(_0811_),
    .S(_0895_),
    .X(_0898_));
 sky130_fd_sc_hd__clkbuf_1 _2392_ (.A(_0898_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2393_ (.A0(\po_0.regf_0.rf[6][9] ),
    .A1(_0820_),
    .S(_0895_),
    .X(_0899_));
 sky130_fd_sc_hd__clkbuf_1 _2394_ (.A(_0899_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _2395_ (.A0(\po_0.regf_0.rf[6][10] ),
    .A1(_0830_),
    .S(_0895_),
    .X(_0900_));
 sky130_fd_sc_hd__clkbuf_1 _2396_ (.A(_0900_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _2397_ (.A0(\po_0.regf_0.rf[6][11] ),
    .A1(_0839_),
    .S(_0895_),
    .X(_0901_));
 sky130_fd_sc_hd__clkbuf_1 _2398_ (.A(_0901_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _2399_ (.A0(\po_0.regf_0.rf[6][12] ),
    .A1(_0849_),
    .S(_0887_),
    .X(_0902_));
 sky130_fd_sc_hd__clkbuf_1 _2400_ (.A(_0902_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _2401_ (.A0(\po_0.regf_0.rf[6][13] ),
    .A1(_0859_),
    .S(_0887_),
    .X(_0903_));
 sky130_fd_sc_hd__clkbuf_1 _2402_ (.A(_0903_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(\po_0.regf_0.rf[6][14] ),
    .A1(_0871_),
    .S(_0887_),
    .X(_0904_));
 sky130_fd_sc_hd__clkbuf_1 _2404_ (.A(_0904_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2405_ (.A0(\po_0.regf_0.rf[6][15] ),
    .A1(_0880_),
    .S(_0887_),
    .X(_0905_));
 sky130_fd_sc_hd__clkbuf_1 _2406_ (.A(_0905_),
    .X(_0047_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2407_ (.A(\po_0.regf_0.w_wr ),
    .X(_0906_));
 sky130_fd_sc_hd__and2b_1 _2408_ (.A_N(_0884_),
    .B(_0883_),
    .X(_0907_));
 sky130_fd_sc_hd__and4b_4 _2409_ (.A_N(_0882_),
    .B(_0906_),
    .C(_0907_),
    .D(_0886_),
    .X(_0908_));
 sky130_fd_sc_hd__buf_2 _2410_ (.A(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(\po_0.regf_0.rf[5][0] ),
    .A1(_0714_),
    .S(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__clkbuf_1 _2412_ (.A(_0910_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _2413_ (.A0(\po_0.regf_0.rf[5][1] ),
    .A1(_0732_),
    .S(_0909_),
    .X(_0911_));
 sky130_fd_sc_hd__clkbuf_1 _2414_ (.A(_0911_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _2415_ (.A0(\po_0.regf_0.rf[5][2] ),
    .A1(_0742_),
    .S(_0909_),
    .X(_0912_));
 sky130_fd_sc_hd__clkbuf_1 _2416_ (.A(_0912_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _2417_ (.A0(\po_0.regf_0.rf[5][3] ),
    .A1(_0753_),
    .S(_0909_),
    .X(_0913_));
 sky130_fd_sc_hd__clkbuf_1 _2418_ (.A(_0913_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(\po_0.regf_0.rf[5][4] ),
    .A1(_0763_),
    .S(_0909_),
    .X(_0914_));
 sky130_fd_sc_hd__clkbuf_1 _2420_ (.A(_0914_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _2421_ (.A0(\po_0.regf_0.rf[5][5] ),
    .A1(_0773_),
    .S(_0909_),
    .X(_0915_));
 sky130_fd_sc_hd__clkbuf_1 _2422_ (.A(_0915_),
    .X(_0053_));
 sky130_fd_sc_hd__buf_2 _2423_ (.A(_0908_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _2424_ (.A0(\po_0.regf_0.rf[5][6] ),
    .A1(_0783_),
    .S(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__clkbuf_1 _2425_ (.A(_0917_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2426_ (.A0(\po_0.regf_0.rf[5][7] ),
    .A1(_0796_),
    .S(_0916_),
    .X(_0918_));
 sky130_fd_sc_hd__clkbuf_1 _2427_ (.A(_0918_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2428_ (.A0(\po_0.regf_0.rf[5][8] ),
    .A1(_0811_),
    .S(_0916_),
    .X(_0919_));
 sky130_fd_sc_hd__clkbuf_1 _2429_ (.A(_0919_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2430_ (.A0(\po_0.regf_0.rf[5][9] ),
    .A1(_0820_),
    .S(_0916_),
    .X(_0920_));
 sky130_fd_sc_hd__clkbuf_1 _2431_ (.A(_0920_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2432_ (.A0(\po_0.regf_0.rf[5][10] ),
    .A1(_0830_),
    .S(_0916_),
    .X(_0921_));
 sky130_fd_sc_hd__clkbuf_1 _2433_ (.A(_0921_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _2434_ (.A0(\po_0.regf_0.rf[5][11] ),
    .A1(_0839_),
    .S(_0916_),
    .X(_0922_));
 sky130_fd_sc_hd__clkbuf_1 _2435_ (.A(_0922_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _2436_ (.A0(\po_0.regf_0.rf[5][12] ),
    .A1(_0849_),
    .S(_0908_),
    .X(_0923_));
 sky130_fd_sc_hd__clkbuf_1 _2437_ (.A(_0923_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(\po_0.regf_0.rf[5][13] ),
    .A1(_0859_),
    .S(_0908_),
    .X(_0924_));
 sky130_fd_sc_hd__clkbuf_1 _2439_ (.A(_0924_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2440_ (.A0(\po_0.regf_0.rf[5][14] ),
    .A1(_0871_),
    .S(_0908_),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_1 _2441_ (.A(_0925_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2442_ (.A0(\po_0.regf_0.rf[5][15] ),
    .A1(_0880_),
    .S(_0908_),
    .X(_0926_));
 sky130_fd_sc_hd__clkbuf_1 _2443_ (.A(_0926_),
    .X(_0063_));
 sky130_fd_sc_hd__clkbuf_2 _2444_ (.A(_0713_),
    .X(_0927_));
 sky130_fd_sc_hd__and4b_2 _2445_ (.A_N(_0886_),
    .B(_0715_),
    .C(_0906_),
    .D(_0907_),
    .X(_0928_));
 sky130_fd_sc_hd__buf_2 _2446_ (.A(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__mux2_1 _2447_ (.A0(\po_0.regf_0.rf[9][0] ),
    .A1(_0927_),
    .S(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__clkbuf_1 _2448_ (.A(_0930_),
    .X(_0064_));
 sky130_fd_sc_hd__clkbuf_2 _2449_ (.A(_0731_),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_1 _2450_ (.A0(\po_0.regf_0.rf[9][1] ),
    .A1(_0931_),
    .S(_0929_),
    .X(_0932_));
 sky130_fd_sc_hd__clkbuf_1 _2451_ (.A(_0932_),
    .X(_0065_));
 sky130_fd_sc_hd__clkbuf_2 _2452_ (.A(_0741_),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_1 _2453_ (.A0(\po_0.regf_0.rf[9][2] ),
    .A1(_0933_),
    .S(_0929_),
    .X(_0934_));
 sky130_fd_sc_hd__clkbuf_1 _2454_ (.A(_0934_),
    .X(_0066_));
 sky130_fd_sc_hd__clkbuf_2 _2455_ (.A(_0752_),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_1 _2456_ (.A0(\po_0.regf_0.rf[9][3] ),
    .A1(_0935_),
    .S(_0929_),
    .X(_0936_));
 sky130_fd_sc_hd__clkbuf_1 _2457_ (.A(_0936_),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_2 _2458_ (.A(_0762_),
    .X(_0937_));
 sky130_fd_sc_hd__mux2_1 _2459_ (.A0(\po_0.regf_0.rf[9][4] ),
    .A1(_0937_),
    .S(_0929_),
    .X(_0938_));
 sky130_fd_sc_hd__clkbuf_1 _2460_ (.A(_0938_),
    .X(_0068_));
 sky130_fd_sc_hd__clkbuf_2 _2461_ (.A(_0772_),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_1 _2462_ (.A0(\po_0.regf_0.rf[9][5] ),
    .A1(_0939_),
    .S(_0929_),
    .X(_0940_));
 sky130_fd_sc_hd__clkbuf_1 _2463_ (.A(_0940_),
    .X(_0069_));
 sky130_fd_sc_hd__clkbuf_2 _2464_ (.A(_0782_),
    .X(_0941_));
 sky130_fd_sc_hd__buf_2 _2465_ (.A(_0928_),
    .X(_0942_));
 sky130_fd_sc_hd__mux2_1 _2466_ (.A0(\po_0.regf_0.rf[9][6] ),
    .A1(_0941_),
    .S(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__clkbuf_1 _2467_ (.A(_0943_),
    .X(_0070_));
 sky130_fd_sc_hd__clkbuf_2 _2468_ (.A(_0795_),
    .X(_0944_));
 sky130_fd_sc_hd__mux2_1 _2469_ (.A0(\po_0.regf_0.rf[9][7] ),
    .A1(_0944_),
    .S(_0942_),
    .X(_0945_));
 sky130_fd_sc_hd__clkbuf_1 _2470_ (.A(_0945_),
    .X(_0071_));
 sky130_fd_sc_hd__clkbuf_2 _2471_ (.A(_0810_),
    .X(_0946_));
 sky130_fd_sc_hd__mux2_1 _2472_ (.A0(\po_0.regf_0.rf[9][8] ),
    .A1(_0946_),
    .S(_0942_),
    .X(_0947_));
 sky130_fd_sc_hd__clkbuf_1 _2473_ (.A(_0947_),
    .X(_0072_));
 sky130_fd_sc_hd__clkbuf_2 _2474_ (.A(_0819_),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _2475_ (.A0(\po_0.regf_0.rf[9][9] ),
    .A1(_0948_),
    .S(_0942_),
    .X(_0949_));
 sky130_fd_sc_hd__clkbuf_1 _2476_ (.A(_0949_),
    .X(_0073_));
 sky130_fd_sc_hd__clkbuf_2 _2477_ (.A(_0829_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _2478_ (.A0(\po_0.regf_0.rf[9][10] ),
    .A1(_0950_),
    .S(_0942_),
    .X(_0951_));
 sky130_fd_sc_hd__clkbuf_1 _2479_ (.A(_0951_),
    .X(_0074_));
 sky130_fd_sc_hd__clkbuf_2 _2480_ (.A(_0838_),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_1 _2481_ (.A0(\po_0.regf_0.rf[9][11] ),
    .A1(_0952_),
    .S(_0942_),
    .X(_0953_));
 sky130_fd_sc_hd__clkbuf_1 _2482_ (.A(_0953_),
    .X(_0075_));
 sky130_fd_sc_hd__clkbuf_2 _2483_ (.A(_0848_),
    .X(_0954_));
 sky130_fd_sc_hd__mux2_1 _2484_ (.A0(\po_0.regf_0.rf[9][12] ),
    .A1(_0954_),
    .S(_0928_),
    .X(_0955_));
 sky130_fd_sc_hd__clkbuf_1 _2485_ (.A(_0955_),
    .X(_0076_));
 sky130_fd_sc_hd__clkbuf_2 _2486_ (.A(_0858_),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _2487_ (.A0(\po_0.regf_0.rf[9][13] ),
    .A1(_0956_),
    .S(_0928_),
    .X(_0957_));
 sky130_fd_sc_hd__clkbuf_1 _2488_ (.A(_0957_),
    .X(_0077_));
 sky130_fd_sc_hd__clkbuf_2 _2489_ (.A(_0870_),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _2490_ (.A0(\po_0.regf_0.rf[9][14] ),
    .A1(_0958_),
    .S(_0928_),
    .X(_0959_));
 sky130_fd_sc_hd__clkbuf_1 _2491_ (.A(_0959_),
    .X(_0078_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2492_ (.A(_0879_),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_1 _2493_ (.A0(\po_0.regf_0.rf[9][15] ),
    .A1(_0960_),
    .S(_0928_),
    .X(_0961_));
 sky130_fd_sc_hd__clkbuf_1 _2494_ (.A(_0961_),
    .X(_0079_));
 sky130_fd_sc_hd__and4bb_2 _2495_ (.A_N(_0718_),
    .B_N(\po_0.regf_0.w_addr[3] ),
    .C(_0906_),
    .D(_0907_),
    .X(_0962_));
 sky130_fd_sc_hd__buf_2 _2496_ (.A(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_1 _2497_ (.A0(\po_0.regf_0.rf[1][0] ),
    .A1(_0927_),
    .S(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__clkbuf_1 _2498_ (.A(_0964_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2499_ (.A0(\po_0.regf_0.rf[1][1] ),
    .A1(_0931_),
    .S(_0963_),
    .X(_0965_));
 sky130_fd_sc_hd__clkbuf_1 _2500_ (.A(_0965_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2501_ (.A0(\po_0.regf_0.rf[1][2] ),
    .A1(_0933_),
    .S(_0963_),
    .X(_0966_));
 sky130_fd_sc_hd__clkbuf_1 _2502_ (.A(_0966_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2503_ (.A0(\po_0.regf_0.rf[1][3] ),
    .A1(_0935_),
    .S(_0963_),
    .X(_0967_));
 sky130_fd_sc_hd__clkbuf_1 _2504_ (.A(_0967_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2505_ (.A0(\po_0.regf_0.rf[1][4] ),
    .A1(_0937_),
    .S(_0963_),
    .X(_0968_));
 sky130_fd_sc_hd__clkbuf_1 _2506_ (.A(_0968_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2507_ (.A0(\po_0.regf_0.rf[1][5] ),
    .A1(_0939_),
    .S(_0963_),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_1 _2508_ (.A(_0969_),
    .X(_0085_));
 sky130_fd_sc_hd__buf_2 _2509_ (.A(_0962_),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(\po_0.regf_0.rf[1][6] ),
    .A1(_0941_),
    .S(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__clkbuf_1 _2511_ (.A(_0971_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(\po_0.regf_0.rf[1][7] ),
    .A1(_0944_),
    .S(_0970_),
    .X(_0972_));
 sky130_fd_sc_hd__clkbuf_1 _2513_ (.A(_0972_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2514_ (.A0(\po_0.regf_0.rf[1][8] ),
    .A1(_0946_),
    .S(_0970_),
    .X(_0973_));
 sky130_fd_sc_hd__clkbuf_1 _2515_ (.A(_0973_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2516_ (.A0(\po_0.regf_0.rf[1][9] ),
    .A1(_0948_),
    .S(_0970_),
    .X(_0974_));
 sky130_fd_sc_hd__clkbuf_1 _2517_ (.A(_0974_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2518_ (.A0(\po_0.regf_0.rf[1][10] ),
    .A1(_0950_),
    .S(_0970_),
    .X(_0975_));
 sky130_fd_sc_hd__clkbuf_1 _2519_ (.A(_0975_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(\po_0.regf_0.rf[1][11] ),
    .A1(_0952_),
    .S(_0970_),
    .X(_0976_));
 sky130_fd_sc_hd__clkbuf_1 _2521_ (.A(_0976_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(\po_0.regf_0.rf[1][12] ),
    .A1(_0954_),
    .S(_0962_),
    .X(_0977_));
 sky130_fd_sc_hd__clkbuf_1 _2523_ (.A(_0977_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(\po_0.regf_0.rf[1][13] ),
    .A1(_0956_),
    .S(_0962_),
    .X(_0978_));
 sky130_fd_sc_hd__clkbuf_1 _2525_ (.A(_0978_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(\po_0.regf_0.rf[1][14] ),
    .A1(_0958_),
    .S(_0962_),
    .X(_0979_));
 sky130_fd_sc_hd__clkbuf_1 _2527_ (.A(_0979_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _2528_ (.A0(\po_0.regf_0.rf[1][15] ),
    .A1(_0960_),
    .S(_0962_),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_1 _2529_ (.A(_0980_),
    .X(_0095_));
 sky130_fd_sc_hd__and4_2 _2530_ (.A(_0718_),
    .B(_0715_),
    .C(_0716_),
    .D(_0717_),
    .X(_0981_));
 sky130_fd_sc_hd__buf_2 _2531_ (.A(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _2532_ (.A0(\po_0.regf_0.rf[15][0] ),
    .A1(_0927_),
    .S(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__clkbuf_1 _2533_ (.A(_0983_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _2534_ (.A0(\po_0.regf_0.rf[15][1] ),
    .A1(_0931_),
    .S(_0982_),
    .X(_0984_));
 sky130_fd_sc_hd__clkbuf_1 _2535_ (.A(_0984_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _2536_ (.A0(\po_0.regf_0.rf[15][2] ),
    .A1(_0933_),
    .S(_0982_),
    .X(_0985_));
 sky130_fd_sc_hd__clkbuf_1 _2537_ (.A(_0985_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(\po_0.regf_0.rf[15][3] ),
    .A1(_0935_),
    .S(_0982_),
    .X(_0986_));
 sky130_fd_sc_hd__clkbuf_1 _2539_ (.A(_0986_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _2540_ (.A0(\po_0.regf_0.rf[15][4] ),
    .A1(_0937_),
    .S(_0982_),
    .X(_0987_));
 sky130_fd_sc_hd__clkbuf_1 _2541_ (.A(_0987_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(\po_0.regf_0.rf[15][5] ),
    .A1(_0939_),
    .S(_0982_),
    .X(_0988_));
 sky130_fd_sc_hd__clkbuf_1 _2543_ (.A(_0988_),
    .X(_0101_));
 sky130_fd_sc_hd__buf_2 _2544_ (.A(_0981_),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_1 _2545_ (.A0(\po_0.regf_0.rf[15][6] ),
    .A1(_0941_),
    .S(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__clkbuf_1 _2546_ (.A(_0990_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _2547_ (.A0(\po_0.regf_0.rf[15][7] ),
    .A1(_0944_),
    .S(_0989_),
    .X(_0991_));
 sky130_fd_sc_hd__clkbuf_1 _2548_ (.A(_0991_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _2549_ (.A0(\po_0.regf_0.rf[15][8] ),
    .A1(_0946_),
    .S(_0989_),
    .X(_0992_));
 sky130_fd_sc_hd__clkbuf_1 _2550_ (.A(_0992_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(\po_0.regf_0.rf[15][9] ),
    .A1(_0948_),
    .S(_0989_),
    .X(_0993_));
 sky130_fd_sc_hd__clkbuf_1 _2552_ (.A(_0993_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2553_ (.A0(\po_0.regf_0.rf[15][10] ),
    .A1(_0950_),
    .S(_0989_),
    .X(_0994_));
 sky130_fd_sc_hd__clkbuf_1 _2554_ (.A(_0994_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(\po_0.regf_0.rf[15][11] ),
    .A1(_0952_),
    .S(_0989_),
    .X(_0995_));
 sky130_fd_sc_hd__clkbuf_1 _2556_ (.A(_0995_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(\po_0.regf_0.rf[15][12] ),
    .A1(_0954_),
    .S(_0981_),
    .X(_0996_));
 sky130_fd_sc_hd__clkbuf_1 _2558_ (.A(_0996_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _2559_ (.A0(\po_0.regf_0.rf[15][13] ),
    .A1(_0956_),
    .S(_0981_),
    .X(_0997_));
 sky130_fd_sc_hd__clkbuf_1 _2560_ (.A(_0997_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(\po_0.regf_0.rf[15][14] ),
    .A1(_0958_),
    .S(_0981_),
    .X(_0998_));
 sky130_fd_sc_hd__clkbuf_1 _2562_ (.A(_0998_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _2563_ (.A0(\po_0.regf_0.rf[15][15] ),
    .A1(_0960_),
    .S(_0981_),
    .X(_0999_));
 sky130_fd_sc_hd__clkbuf_1 _2564_ (.A(_0999_),
    .X(_0111_));
 sky130_fd_sc_hd__nand3_1 _2565_ (.A(\po_0.regf_0.w_addr[2] ),
    .B(\po_0.regf_0.w_addr[3] ),
    .C(\po_0.regf_0.w_wr ),
    .Y(_1000_));
 sky130_fd_sc_hd__or3b_4 _2566_ (.A(_0883_),
    .B(_1000_),
    .C_N(_0884_),
    .X(_1001_));
 sky130_fd_sc_hd__buf_2 _2567_ (.A(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_1 _2568_ (.A0(_0714_),
    .A1(\po_0.regf_0.rf[14][0] ),
    .S(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__clkbuf_1 _2569_ (.A(_1003_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _2570_ (.A0(_0732_),
    .A1(\po_0.regf_0.rf[14][1] ),
    .S(_1002_),
    .X(_1004_));
 sky130_fd_sc_hd__clkbuf_1 _2571_ (.A(_1004_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(_0742_),
    .A1(\po_0.regf_0.rf[14][2] ),
    .S(_1002_),
    .X(_1005_));
 sky130_fd_sc_hd__clkbuf_1 _2573_ (.A(_1005_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(_0753_),
    .A1(\po_0.regf_0.rf[14][3] ),
    .S(_1002_),
    .X(_1006_));
 sky130_fd_sc_hd__clkbuf_1 _2575_ (.A(_1006_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(_0763_),
    .A1(\po_0.regf_0.rf[14][4] ),
    .S(_1002_),
    .X(_1007_));
 sky130_fd_sc_hd__clkbuf_1 _2577_ (.A(_1007_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(_0773_),
    .A1(\po_0.regf_0.rf[14][5] ),
    .S(_1002_),
    .X(_1008_));
 sky130_fd_sc_hd__clkbuf_1 _2579_ (.A(_1008_),
    .X(_0117_));
 sky130_fd_sc_hd__buf_2 _2580_ (.A(_1001_),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_1 _2581_ (.A0(_0783_),
    .A1(\po_0.regf_0.rf[14][6] ),
    .S(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__clkbuf_1 _2582_ (.A(_1010_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _2583_ (.A0(_0796_),
    .A1(\po_0.regf_0.rf[14][7] ),
    .S(_1009_),
    .X(_1011_));
 sky130_fd_sc_hd__clkbuf_1 _2584_ (.A(_1011_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _2585_ (.A0(_0811_),
    .A1(\po_0.regf_0.rf[14][8] ),
    .S(_1009_),
    .X(_1012_));
 sky130_fd_sc_hd__clkbuf_1 _2586_ (.A(_1012_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(_0820_),
    .A1(\po_0.regf_0.rf[14][9] ),
    .S(_1009_),
    .X(_1013_));
 sky130_fd_sc_hd__clkbuf_1 _2588_ (.A(_1013_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2589_ (.A0(_0830_),
    .A1(\po_0.regf_0.rf[14][10] ),
    .S(_1009_),
    .X(_1014_));
 sky130_fd_sc_hd__clkbuf_1 _2590_ (.A(_1014_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _2591_ (.A0(_0839_),
    .A1(\po_0.regf_0.rf[14][11] ),
    .S(_1009_),
    .X(_1015_));
 sky130_fd_sc_hd__clkbuf_1 _2592_ (.A(_1015_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _2593_ (.A0(_0849_),
    .A1(\po_0.regf_0.rf[14][12] ),
    .S(_1001_),
    .X(_1016_));
 sky130_fd_sc_hd__clkbuf_1 _2594_ (.A(_1016_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _2595_ (.A0(_0859_),
    .A1(\po_0.regf_0.rf[14][13] ),
    .S(_1001_),
    .X(_1017_));
 sky130_fd_sc_hd__clkbuf_1 _2596_ (.A(_1017_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2597_ (.A0(_0871_),
    .A1(\po_0.regf_0.rf[14][14] ),
    .S(_1001_),
    .X(_1018_));
 sky130_fd_sc_hd__clkbuf_1 _2598_ (.A(_1018_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _2599_ (.A0(_0880_),
    .A1(\po_0.regf_0.rf[14][15] ),
    .S(_1001_),
    .X(_1019_));
 sky130_fd_sc_hd__clkbuf_1 _2600_ (.A(_1019_),
    .X(_0127_));
 sky130_fd_sc_hd__or3b_4 _2601_ (.A(_1000_),
    .B(_0884_),
    .C_N(_0883_),
    .X(_1020_));
 sky130_fd_sc_hd__buf_2 _2602_ (.A(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_1 _2603_ (.A0(_0714_),
    .A1(\po_0.regf_0.rf[13][0] ),
    .S(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__clkbuf_1 _2604_ (.A(_1022_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _2605_ (.A0(_0732_),
    .A1(\po_0.regf_0.rf[13][1] ),
    .S(_1021_),
    .X(_1023_));
 sky130_fd_sc_hd__clkbuf_1 _2606_ (.A(_1023_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _2607_ (.A0(_0742_),
    .A1(\po_0.regf_0.rf[13][2] ),
    .S(_1021_),
    .X(_1024_));
 sky130_fd_sc_hd__clkbuf_1 _2608_ (.A(_1024_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(_0753_),
    .A1(\po_0.regf_0.rf[13][3] ),
    .S(_1021_),
    .X(_1025_));
 sky130_fd_sc_hd__clkbuf_1 _2610_ (.A(_1025_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(_0763_),
    .A1(\po_0.regf_0.rf[13][4] ),
    .S(_1021_),
    .X(_1026_));
 sky130_fd_sc_hd__clkbuf_1 _2612_ (.A(_1026_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2613_ (.A0(_0773_),
    .A1(\po_0.regf_0.rf[13][5] ),
    .S(_1021_),
    .X(_1027_));
 sky130_fd_sc_hd__clkbuf_1 _2614_ (.A(_1027_),
    .X(_0133_));
 sky130_fd_sc_hd__buf_2 _2615_ (.A(_1020_),
    .X(_1028_));
 sky130_fd_sc_hd__mux2_1 _2616_ (.A0(_0783_),
    .A1(\po_0.regf_0.rf[13][6] ),
    .S(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__clkbuf_1 _2617_ (.A(_1029_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _2618_ (.A0(_0796_),
    .A1(\po_0.regf_0.rf[13][7] ),
    .S(_1028_),
    .X(_1030_));
 sky130_fd_sc_hd__clkbuf_1 _2619_ (.A(_1030_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _2620_ (.A0(_0811_),
    .A1(\po_0.regf_0.rf[13][8] ),
    .S(_1028_),
    .X(_1031_));
 sky130_fd_sc_hd__clkbuf_1 _2621_ (.A(_1031_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _2622_ (.A0(_0820_),
    .A1(\po_0.regf_0.rf[13][9] ),
    .S(_1028_),
    .X(_1032_));
 sky130_fd_sc_hd__clkbuf_1 _2623_ (.A(_1032_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _2624_ (.A0(_0830_),
    .A1(\po_0.regf_0.rf[13][10] ),
    .S(_1028_),
    .X(_1033_));
 sky130_fd_sc_hd__clkbuf_1 _2625_ (.A(_1033_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _2626_ (.A0(_0839_),
    .A1(\po_0.regf_0.rf[13][11] ),
    .S(_1028_),
    .X(_1034_));
 sky130_fd_sc_hd__clkbuf_1 _2627_ (.A(_1034_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _2628_ (.A0(_0849_),
    .A1(\po_0.regf_0.rf[13][12] ),
    .S(_1020_),
    .X(_1035_));
 sky130_fd_sc_hd__clkbuf_1 _2629_ (.A(_1035_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _2630_ (.A0(_0859_),
    .A1(\po_0.regf_0.rf[13][13] ),
    .S(_1020_),
    .X(_1036_));
 sky130_fd_sc_hd__clkbuf_1 _2631_ (.A(_1036_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(_0871_),
    .A1(\po_0.regf_0.rf[13][14] ),
    .S(_1020_),
    .X(_1037_));
 sky130_fd_sc_hd__clkbuf_1 _2633_ (.A(_1037_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(_0880_),
    .A1(\po_0.regf_0.rf[13][15] ),
    .S(_1020_),
    .X(_1038_));
 sky130_fd_sc_hd__clkbuf_1 _2635_ (.A(_1038_),
    .X(_0143_));
 sky130_fd_sc_hd__nor2_1 _2636_ (.A(_0884_),
    .B(_0883_),
    .Y(_1039_));
 sky130_fd_sc_hd__and4_2 _2637_ (.A(_0718_),
    .B(_0715_),
    .C(_0716_),
    .D(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__buf_2 _2638_ (.A(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__mux2_1 _2639_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(_0927_),
    .S(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__clkbuf_1 _2640_ (.A(_1042_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2641_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(_0931_),
    .S(_1041_),
    .X(_1043_));
 sky130_fd_sc_hd__clkbuf_1 _2642_ (.A(_1043_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2643_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(_0933_),
    .S(_1041_),
    .X(_1044_));
 sky130_fd_sc_hd__clkbuf_1 _2644_ (.A(_1044_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(_0935_),
    .S(_1041_),
    .X(_1045_));
 sky130_fd_sc_hd__clkbuf_1 _2646_ (.A(_1045_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2647_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(_0937_),
    .S(_1041_),
    .X(_1046_));
 sky130_fd_sc_hd__clkbuf_1 _2648_ (.A(_1046_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2649_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(_0939_),
    .S(_1041_),
    .X(_1047_));
 sky130_fd_sc_hd__clkbuf_1 _2650_ (.A(_1047_),
    .X(_0149_));
 sky130_fd_sc_hd__buf_2 _2651_ (.A(_1040_),
    .X(_1048_));
 sky130_fd_sc_hd__mux2_1 _2652_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(_0941_),
    .S(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__clkbuf_1 _2653_ (.A(_1049_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2654_ (.A0(\po_0.regf_0.rf[12][7] ),
    .A1(_0944_),
    .S(_1048_),
    .X(_1050_));
 sky130_fd_sc_hd__clkbuf_1 _2655_ (.A(_1050_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2656_ (.A0(\po_0.regf_0.rf[12][8] ),
    .A1(_0946_),
    .S(_1048_),
    .X(_1051_));
 sky130_fd_sc_hd__clkbuf_1 _2657_ (.A(_1051_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2658_ (.A0(\po_0.regf_0.rf[12][9] ),
    .A1(_0948_),
    .S(_1048_),
    .X(_1052_));
 sky130_fd_sc_hd__clkbuf_1 _2659_ (.A(_1052_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2660_ (.A0(\po_0.regf_0.rf[12][10] ),
    .A1(_0950_),
    .S(_1048_),
    .X(_1053_));
 sky130_fd_sc_hd__clkbuf_1 _2661_ (.A(_1053_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2662_ (.A0(\po_0.regf_0.rf[12][11] ),
    .A1(_0952_),
    .S(_1048_),
    .X(_1054_));
 sky130_fd_sc_hd__clkbuf_1 _2663_ (.A(_1054_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2664_ (.A0(\po_0.regf_0.rf[12][12] ),
    .A1(_0954_),
    .S(_1040_),
    .X(_1055_));
 sky130_fd_sc_hd__clkbuf_1 _2665_ (.A(_1055_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2666_ (.A0(\po_0.regf_0.rf[12][13] ),
    .A1(_0956_),
    .S(_1040_),
    .X(_1056_));
 sky130_fd_sc_hd__clkbuf_1 _2667_ (.A(_1056_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2668_ (.A0(\po_0.regf_0.rf[12][14] ),
    .A1(_0958_),
    .S(_1040_),
    .X(_1057_));
 sky130_fd_sc_hd__clkbuf_1 _2669_ (.A(_1057_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2670_ (.A0(\po_0.regf_0.rf[12][15] ),
    .A1(_0960_),
    .S(_1040_),
    .X(_1058_));
 sky130_fd_sc_hd__clkbuf_1 _2671_ (.A(_1058_),
    .X(_0159_));
 sky130_fd_sc_hd__and4b_2 _2672_ (.A_N(\po_0.regf_0.w_addr[2] ),
    .B(_0715_),
    .C(\po_0.regf_0.w_wr ),
    .D(_0717_),
    .X(_1059_));
 sky130_fd_sc_hd__buf_2 _2673_ (.A(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__mux2_1 _2674_ (.A0(\po_0.regf_0.rf[11][0] ),
    .A1(_0927_),
    .S(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__clkbuf_1 _2675_ (.A(_1061_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2676_ (.A0(\po_0.regf_0.rf[11][1] ),
    .A1(_0931_),
    .S(_1060_),
    .X(_1062_));
 sky130_fd_sc_hd__clkbuf_1 _2677_ (.A(_1062_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2678_ (.A0(\po_0.regf_0.rf[11][2] ),
    .A1(_0933_),
    .S(_1060_),
    .X(_1063_));
 sky130_fd_sc_hd__clkbuf_1 _2679_ (.A(_1063_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2680_ (.A0(\po_0.regf_0.rf[11][3] ),
    .A1(_0935_),
    .S(_1060_),
    .X(_1064_));
 sky130_fd_sc_hd__clkbuf_1 _2681_ (.A(_1064_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2682_ (.A0(\po_0.regf_0.rf[11][4] ),
    .A1(_0937_),
    .S(_1060_),
    .X(_1065_));
 sky130_fd_sc_hd__clkbuf_1 _2683_ (.A(_1065_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2684_ (.A0(\po_0.regf_0.rf[11][5] ),
    .A1(_0939_),
    .S(_1060_),
    .X(_1066_));
 sky130_fd_sc_hd__clkbuf_1 _2685_ (.A(_1066_),
    .X(_0165_));
 sky130_fd_sc_hd__buf_2 _2686_ (.A(_1059_),
    .X(_1067_));
 sky130_fd_sc_hd__mux2_1 _2687_ (.A0(\po_0.regf_0.rf[11][6] ),
    .A1(_0941_),
    .S(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__clkbuf_1 _2688_ (.A(_1068_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2689_ (.A0(\po_0.regf_0.rf[11][7] ),
    .A1(_0944_),
    .S(_1067_),
    .X(_1069_));
 sky130_fd_sc_hd__clkbuf_1 _2690_ (.A(_1069_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2691_ (.A0(\po_0.regf_0.rf[11][8] ),
    .A1(_0946_),
    .S(_1067_),
    .X(_1070_));
 sky130_fd_sc_hd__clkbuf_1 _2692_ (.A(_1070_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2693_ (.A0(\po_0.regf_0.rf[11][9] ),
    .A1(_0948_),
    .S(_1067_),
    .X(_1071_));
 sky130_fd_sc_hd__clkbuf_1 _2694_ (.A(_1071_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _2695_ (.A0(\po_0.regf_0.rf[11][10] ),
    .A1(_0950_),
    .S(_1067_),
    .X(_1072_));
 sky130_fd_sc_hd__clkbuf_1 _2696_ (.A(_1072_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2697_ (.A0(\po_0.regf_0.rf[11][11] ),
    .A1(_0952_),
    .S(_1067_),
    .X(_1073_));
 sky130_fd_sc_hd__clkbuf_1 _2698_ (.A(_1073_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _2699_ (.A0(\po_0.regf_0.rf[11][12] ),
    .A1(_0954_),
    .S(_1059_),
    .X(_1074_));
 sky130_fd_sc_hd__clkbuf_1 _2700_ (.A(_1074_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2701_ (.A0(\po_0.regf_0.rf[11][13] ),
    .A1(_0956_),
    .S(_1059_),
    .X(_1075_));
 sky130_fd_sc_hd__clkbuf_1 _2702_ (.A(_1075_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2703_ (.A0(\po_0.regf_0.rf[11][14] ),
    .A1(_0958_),
    .S(_1059_),
    .X(_1076_));
 sky130_fd_sc_hd__clkbuf_1 _2704_ (.A(_1076_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _2705_ (.A0(\po_0.regf_0.rf[11][15] ),
    .A1(_0960_),
    .S(_1059_),
    .X(_1077_));
 sky130_fd_sc_hd__clkbuf_1 _2706_ (.A(_1077_),
    .X(_0175_));
 sky130_fd_sc_hd__and4b_2 _2707_ (.A_N(\po_0.regf_0.w_addr[2] ),
    .B(_0882_),
    .C(\po_0.regf_0.w_wr ),
    .D(_0885_),
    .X(_1078_));
 sky130_fd_sc_hd__buf_2 _2708_ (.A(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__mux2_1 _2709_ (.A0(\po_0.regf_0.rf[10][0] ),
    .A1(_0927_),
    .S(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__clkbuf_1 _2710_ (.A(_1080_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2711_ (.A0(\po_0.regf_0.rf[10][1] ),
    .A1(_0931_),
    .S(_1079_),
    .X(_1081_));
 sky130_fd_sc_hd__clkbuf_1 _2712_ (.A(_1081_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2713_ (.A0(\po_0.regf_0.rf[10][2] ),
    .A1(_0933_),
    .S(_1079_),
    .X(_1082_));
 sky130_fd_sc_hd__clkbuf_1 _2714_ (.A(_1082_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2715_ (.A0(\po_0.regf_0.rf[10][3] ),
    .A1(_0935_),
    .S(_1079_),
    .X(_1083_));
 sky130_fd_sc_hd__clkbuf_1 _2716_ (.A(_1083_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _2717_ (.A0(\po_0.regf_0.rf[10][4] ),
    .A1(_0937_),
    .S(_1079_),
    .X(_1084_));
 sky130_fd_sc_hd__clkbuf_1 _2718_ (.A(_1084_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2719_ (.A0(\po_0.regf_0.rf[10][5] ),
    .A1(_0939_),
    .S(_1079_),
    .X(_1085_));
 sky130_fd_sc_hd__clkbuf_1 _2720_ (.A(_1085_),
    .X(_0181_));
 sky130_fd_sc_hd__buf_2 _2721_ (.A(_1078_),
    .X(_1086_));
 sky130_fd_sc_hd__mux2_1 _2722_ (.A0(\po_0.regf_0.rf[10][6] ),
    .A1(_0941_),
    .S(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__clkbuf_1 _2723_ (.A(_1087_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2724_ (.A0(\po_0.regf_0.rf[10][7] ),
    .A1(_0944_),
    .S(_1086_),
    .X(_1088_));
 sky130_fd_sc_hd__clkbuf_1 _2725_ (.A(_1088_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2726_ (.A0(\po_0.regf_0.rf[10][8] ),
    .A1(_0946_),
    .S(_1086_),
    .X(_1089_));
 sky130_fd_sc_hd__clkbuf_1 _2727_ (.A(_1089_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _2728_ (.A0(\po_0.regf_0.rf[10][9] ),
    .A1(_0948_),
    .S(_1086_),
    .X(_1090_));
 sky130_fd_sc_hd__clkbuf_1 _2729_ (.A(_1090_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _2730_ (.A0(\po_0.regf_0.rf[10][10] ),
    .A1(_0950_),
    .S(_1086_),
    .X(_1091_));
 sky130_fd_sc_hd__clkbuf_1 _2731_ (.A(_1091_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2732_ (.A0(\po_0.regf_0.rf[10][11] ),
    .A1(_0952_),
    .S(_1086_),
    .X(_1092_));
 sky130_fd_sc_hd__clkbuf_1 _2733_ (.A(_1092_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _2734_ (.A0(\po_0.regf_0.rf[10][12] ),
    .A1(_0954_),
    .S(_1078_),
    .X(_1093_));
 sky130_fd_sc_hd__clkbuf_1 _2735_ (.A(_1093_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _2736_ (.A0(\po_0.regf_0.rf[10][13] ),
    .A1(_0956_),
    .S(_1078_),
    .X(_1094_));
 sky130_fd_sc_hd__clkbuf_1 _2737_ (.A(_1094_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _2738_ (.A0(\po_0.regf_0.rf[10][14] ),
    .A1(_0958_),
    .S(_1078_),
    .X(_1095_));
 sky130_fd_sc_hd__clkbuf_1 _2739_ (.A(_1095_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _2740_ (.A0(\po_0.regf_0.rf[10][15] ),
    .A1(_0960_),
    .S(_1078_),
    .X(_1096_));
 sky130_fd_sc_hd__clkbuf_1 _2741_ (.A(_1096_),
    .X(_0191_));
 sky130_fd_sc_hd__or4bb_4 _2742_ (.A(_0718_),
    .B(_0882_),
    .C_N(_0716_),
    .D_N(_1039_),
    .X(_1097_));
 sky130_fd_sc_hd__buf_2 _2743_ (.A(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__mux2_1 _2744_ (.A0(_0714_),
    .A1(\po_0.regf_0.rf[0][0] ),
    .S(_1098_),
    .X(_1099_));
 sky130_fd_sc_hd__clkbuf_1 _2745_ (.A(_1099_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _2746_ (.A0(_0732_),
    .A1(\po_0.regf_0.rf[0][1] ),
    .S(_1098_),
    .X(_1100_));
 sky130_fd_sc_hd__clkbuf_1 _2747_ (.A(_1100_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(_0742_),
    .A1(\po_0.regf_0.rf[0][2] ),
    .S(_1098_),
    .X(_1101_));
 sky130_fd_sc_hd__clkbuf_1 _2749_ (.A(_1101_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _2750_ (.A0(_0753_),
    .A1(\po_0.regf_0.rf[0][3] ),
    .S(_1098_),
    .X(_1102_));
 sky130_fd_sc_hd__clkbuf_1 _2751_ (.A(_1102_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _2752_ (.A0(_0763_),
    .A1(\po_0.regf_0.rf[0][4] ),
    .S(_1098_),
    .X(_1103_));
 sky130_fd_sc_hd__clkbuf_1 _2753_ (.A(_1103_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _2754_ (.A0(_0773_),
    .A1(\po_0.regf_0.rf[0][5] ),
    .S(_1098_),
    .X(_1104_));
 sky130_fd_sc_hd__clkbuf_1 _2755_ (.A(_1104_),
    .X(_0197_));
 sky130_fd_sc_hd__buf_2 _2756_ (.A(_1097_),
    .X(_1105_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(_0783_),
    .A1(\po_0.regf_0.rf[0][6] ),
    .S(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__clkbuf_1 _2758_ (.A(_1106_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2759_ (.A0(_0796_),
    .A1(\po_0.regf_0.rf[0][7] ),
    .S(_1105_),
    .X(_1107_));
 sky130_fd_sc_hd__clkbuf_1 _2760_ (.A(_1107_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _2761_ (.A0(_0811_),
    .A1(\po_0.regf_0.rf[0][8] ),
    .S(_1105_),
    .X(_1108_));
 sky130_fd_sc_hd__clkbuf_1 _2762_ (.A(_1108_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2763_ (.A0(_0820_),
    .A1(\po_0.regf_0.rf[0][9] ),
    .S(_1105_),
    .X(_1109_));
 sky130_fd_sc_hd__clkbuf_1 _2764_ (.A(_1109_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2765_ (.A0(_0830_),
    .A1(\po_0.regf_0.rf[0][10] ),
    .S(_1105_),
    .X(_1110_));
 sky130_fd_sc_hd__clkbuf_1 _2766_ (.A(_1110_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _2767_ (.A0(_0839_),
    .A1(\po_0.regf_0.rf[0][11] ),
    .S(_1105_),
    .X(_1111_));
 sky130_fd_sc_hd__clkbuf_1 _2768_ (.A(_1111_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _2769_ (.A0(_0849_),
    .A1(\po_0.regf_0.rf[0][12] ),
    .S(_1097_),
    .X(_1112_));
 sky130_fd_sc_hd__clkbuf_1 _2770_ (.A(_1112_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _2771_ (.A0(_0859_),
    .A1(\po_0.regf_0.rf[0][13] ),
    .S(_1097_),
    .X(_1113_));
 sky130_fd_sc_hd__clkbuf_1 _2772_ (.A(_1113_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _2773_ (.A0(_0871_),
    .A1(\po_0.regf_0.rf[0][14] ),
    .S(_1097_),
    .X(_1114_));
 sky130_fd_sc_hd__clkbuf_1 _2774_ (.A(_1114_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _2775_ (.A0(_0880_),
    .A1(\po_0.regf_0.rf[0][15] ),
    .S(_1097_),
    .X(_1115_));
 sky130_fd_sc_hd__clkbuf_1 _2776_ (.A(_1115_),
    .X(_0207_));
 sky130_fd_sc_hd__and4b_2 _2777_ (.A_N(\po_0.regf_0.w_addr[2] ),
    .B(_0882_),
    .C(\po_0.regf_0.w_wr ),
    .D(_1039_),
    .X(_1116_));
 sky130_fd_sc_hd__buf_2 _2778_ (.A(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__mux2_1 _2779_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(_0713_),
    .S(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__clkbuf_1 _2780_ (.A(_1118_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _2781_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(_0731_),
    .S(_1117_),
    .X(_1119_));
 sky130_fd_sc_hd__clkbuf_1 _2782_ (.A(_1119_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _2783_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(_0741_),
    .S(_1117_),
    .X(_1120_));
 sky130_fd_sc_hd__clkbuf_1 _2784_ (.A(_1120_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _2785_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(_0752_),
    .S(_1117_),
    .X(_1121_));
 sky130_fd_sc_hd__clkbuf_1 _2786_ (.A(_1121_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _2787_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(_0762_),
    .S(_1117_),
    .X(_1122_));
 sky130_fd_sc_hd__clkbuf_1 _2788_ (.A(_1122_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _2789_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(_0772_),
    .S(_1117_),
    .X(_1123_));
 sky130_fd_sc_hd__clkbuf_1 _2790_ (.A(_1123_),
    .X(_0213_));
 sky130_fd_sc_hd__buf_2 _2791_ (.A(_1116_),
    .X(_1124_));
 sky130_fd_sc_hd__mux2_1 _2792_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(_0782_),
    .S(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__clkbuf_1 _2793_ (.A(_1125_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _2794_ (.A0(\po_0.regf_0.rf[8][7] ),
    .A1(_0795_),
    .S(_1124_),
    .X(_1126_));
 sky130_fd_sc_hd__clkbuf_1 _2795_ (.A(_1126_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _2796_ (.A0(\po_0.regf_0.rf[8][8] ),
    .A1(_0810_),
    .S(_1124_),
    .X(_1127_));
 sky130_fd_sc_hd__clkbuf_1 _2797_ (.A(_1127_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _2798_ (.A0(\po_0.regf_0.rf[8][9] ),
    .A1(_0819_),
    .S(_1124_),
    .X(_1128_));
 sky130_fd_sc_hd__clkbuf_1 _2799_ (.A(_1128_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2800_ (.A0(\po_0.regf_0.rf[8][10] ),
    .A1(_0829_),
    .S(_1124_),
    .X(_1129_));
 sky130_fd_sc_hd__clkbuf_1 _2801_ (.A(_1129_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(\po_0.regf_0.rf[8][11] ),
    .A1(_0838_),
    .S(_1124_),
    .X(_1130_));
 sky130_fd_sc_hd__clkbuf_1 _2803_ (.A(_1130_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _2804_ (.A0(\po_0.regf_0.rf[8][12] ),
    .A1(_0848_),
    .S(_1116_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_1 _2805_ (.A(_1131_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _2806_ (.A0(\po_0.regf_0.rf[8][13] ),
    .A1(_0858_),
    .S(_1116_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _2807_ (.A(_1132_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _2808_ (.A0(\po_0.regf_0.rf[8][14] ),
    .A1(_0870_),
    .S(_1116_),
    .X(_1133_));
 sky130_fd_sc_hd__clkbuf_1 _2809_ (.A(_1133_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _2810_ (.A0(\po_0.regf_0.rf[8][15] ),
    .A1(_0879_),
    .S(_1116_),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _2811_ (.A(_1134_),
    .X(_0223_));
 sky130_fd_sc_hd__buf_2 _2812_ (.A(\uc_0._01_ ),
    .X(_1135_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2813_ (.A(net61),
    .X(_1136_));
 sky130_fd_sc_hd__nand2_1 _2814_ (.A(_1136_),
    .B(\po_0.muxf_0.rf_w_data[0] ),
    .Y(_1137_));
 sky130_fd_sc_hd__clkbuf_2 _2815_ (.A(_1136_),
    .X(_1138_));
 sky130_fd_sc_hd__clkbuf_2 _2816_ (.A(\uc_0._00_ ),
    .X(_1139_));
 sky130_fd_sc_hd__clkbuf_2 _2817_ (.A(\uc_0._02_ ),
    .X(_1140_));
 sky130_fd_sc_hd__nor2_1 _2818_ (.A(_1139_),
    .B(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__clkbuf_2 _2819_ (.A(_1141_),
    .X(_1142_));
 sky130_fd_sc_hd__o21a_1 _2820_ (.A1(_1138_),
    .A2(_0704_),
    .B1(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2821_ (.A(_1140_),
    .X(_1144_));
 sky130_fd_sc_hd__clkbuf_2 _2822_ (.A(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__or2_1 _2823_ (.A(\uc_0._00_ ),
    .B(\uc_0._02_ ),
    .X(_1146_));
 sky130_fd_sc_hd__nor2_1 _2824_ (.A(\uc_0._01_ ),
    .B(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__buf_2 _2825_ (.A(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__mux2_1 _2826_ (.A0(_1145_),
    .A1(_1148_),
    .S(_1138_),
    .X(_1149_));
 sky130_fd_sc_hd__a31o_1 _2827_ (.A1(_1135_),
    .A2(_1137_),
    .A3(_1143_),
    .B1(_1149_),
    .X(_0224_));
 sky130_fd_sc_hd__nor2_2 _2828_ (.A(net68),
    .B(\po_0.muxf_0.rf_w_data[1] ),
    .Y(_1150_));
 sky130_fd_sc_hd__clkbuf_2 _2829_ (.A(net68),
    .X(_1151_));
 sky130_fd_sc_hd__and2_1 _2830_ (.A(_1151_),
    .B(\po_0.muxf_0.rf_w_data[1] ),
    .X(_1152_));
 sky130_fd_sc_hd__or3_1 _2831_ (.A(_1150_),
    .B(_1137_),
    .C(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__a2bb2o_1 _2832_ (.A1_N(_1152_),
    .A2_N(_1150_),
    .B1(_1136_),
    .B2(_0704_),
    .X(_1154_));
 sky130_fd_sc_hd__clkbuf_2 _2833_ (.A(_1151_),
    .X(_1155_));
 sky130_fd_sc_hd__o21ai_1 _2834_ (.A1(_1138_),
    .A2(_1155_),
    .B1(_1140_),
    .Y(_1156_));
 sky130_fd_sc_hd__a21oi_1 _2835_ (.A1(_1138_),
    .A2(_1155_),
    .B1(_1156_),
    .Y(_1157_));
 sky130_fd_sc_hd__a31o_1 _2836_ (.A1(_1153_),
    .A2(_1142_),
    .A3(_1154_),
    .B1(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__mux2_1 _2837_ (.A0(_1158_),
    .A1(_1155_),
    .S(_1148_),
    .X(_1159_));
 sky130_fd_sc_hd__clkbuf_1 _2838_ (.A(_1159_),
    .X(_0225_));
 sky130_fd_sc_hd__nand2_2 _2839_ (.A(net69),
    .B(_0734_),
    .Y(_1160_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2840_ (.A(net69),
    .X(_1161_));
 sky130_fd_sc_hd__or2_1 _2841_ (.A(_1161_),
    .B(_0734_),
    .X(_1162_));
 sky130_fd_sc_hd__o211a_1 _2842_ (.A1(_1151_),
    .A2(_0724_),
    .B1(_1136_),
    .C1(\po_0.muxf_0.rf_w_data[0] ),
    .X(_1163_));
 sky130_fd_sc_hd__a221o_1 _2843_ (.A1(_1155_),
    .A2(_0724_),
    .B1(_1160_),
    .B2(_1162_),
    .C1(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__o211ai_1 _2844_ (.A1(_1152_),
    .A2(_1163_),
    .B1(_1160_),
    .C1(_1162_),
    .Y(_1165_));
 sky130_fd_sc_hd__and3_1 _2845_ (.A(_1136_),
    .B(_1151_),
    .C(_1161_),
    .X(_1166_));
 sky130_fd_sc_hd__a21o_1 _2846_ (.A1(_1136_),
    .A2(_1151_),
    .B1(_1161_),
    .X(_1167_));
 sky130_fd_sc_hd__and3b_1 _2847_ (.A_N(_1166_),
    .B(_1167_),
    .C(_1140_),
    .X(_1168_));
 sky130_fd_sc_hd__a31o_1 _2848_ (.A1(_1164_),
    .A2(_1141_),
    .A3(_1165_),
    .B1(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__mux2_1 _2849_ (.A0(_1169_),
    .A1(_1161_),
    .S(_1148_),
    .X(_1170_));
 sky130_fd_sc_hd__clkbuf_1 _2850_ (.A(_1170_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_2 _2851_ (.A(_1140_),
    .X(_1171_));
 sky130_fd_sc_hd__clkbuf_2 _2852_ (.A(net99),
    .X(_1172_));
 sky130_fd_sc_hd__a31o_1 _2853_ (.A1(_1138_),
    .A2(_1155_),
    .A3(_1161_),
    .B1(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__nand2_1 _2854_ (.A(net99),
    .B(_1166_),
    .Y(_1174_));
 sky130_fd_sc_hd__or2_1 _2855_ (.A(net99),
    .B(_0744_),
    .X(_1175_));
 sky130_fd_sc_hd__nand2_1 _2856_ (.A(net99),
    .B(\po_0.muxf_0.rf_w_data[3] ),
    .Y(_1176_));
 sky130_fd_sc_hd__nor2_1 _2857_ (.A(net69),
    .B(\po_0.muxf_0.rf_w_data[2] ),
    .Y(_1177_));
 sky130_fd_sc_hd__a22oi_4 _2858_ (.A1(net61),
    .A2(\po_0.muxf_0.rf_w_data[0] ),
    .B1(_1151_),
    .B2(\po_0.muxf_0.rf_w_data[1] ),
    .Y(_1178_));
 sky130_fd_sc_hd__o31a_1 _2859_ (.A1(_1150_),
    .A2(_1177_),
    .A3(_1178_),
    .B1(_1160_),
    .X(_1179_));
 sky130_fd_sc_hd__a21oi_1 _2860_ (.A1(_1175_),
    .A2(_1176_),
    .B1(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__and3_1 _2861_ (.A(_1175_),
    .B(_1176_),
    .C(_1179_),
    .X(_1181_));
 sky130_fd_sc_hd__or2_1 _2862_ (.A(_1180_),
    .B(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__a32o_1 _2863_ (.A1(_1171_),
    .A2(_1173_),
    .A3(_1174_),
    .B1(_1182_),
    .B2(_1142_),
    .X(_1183_));
 sky130_fd_sc_hd__mux2_1 _2864_ (.A0(_1183_),
    .A1(_1172_),
    .S(_1148_),
    .X(_1184_));
 sky130_fd_sc_hd__clkbuf_1 _2865_ (.A(_1184_),
    .X(_0227_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2866_ (.A(net71),
    .X(_1185_));
 sky130_fd_sc_hd__clkbuf_2 _2867_ (.A(_1146_),
    .X(_1186_));
 sky130_fd_sc_hd__clkbuf_2 _2868_ (.A(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__nor2_1 _2869_ (.A(_1185_),
    .B(_0557_),
    .Y(_1188_));
 sky130_fd_sc_hd__inv_2 _2870_ (.A(net71),
    .Y(_1189_));
 sky130_fd_sc_hd__inv_2 _2871_ (.A(\po_0.muxf_0.rf_w_data[4] ),
    .Y(_1190_));
 sky130_fd_sc_hd__nor2_1 _2872_ (.A(_1189_),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__o311ai_4 _2873_ (.A1(_1150_),
    .A2(_1177_),
    .A3(_1178_),
    .B1(_1176_),
    .C1(_1160_),
    .Y(_1192_));
 sky130_fd_sc_hd__o21ai_1 _2874_ (.A1(_1172_),
    .A2(_0744_),
    .B1(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__or3_1 _2875_ (.A(_1188_),
    .B(_1191_),
    .C(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__a2bb2o_1 _2876_ (.A1_N(_1188_),
    .A2_N(_1191_),
    .B1(_1192_),
    .B2(_1175_),
    .X(_1195_));
 sky130_fd_sc_hd__or2_1 _2877_ (.A(_1189_),
    .B(_1174_),
    .X(_1196_));
 sky130_fd_sc_hd__a41o_1 _2878_ (.A1(_1138_),
    .A2(_1155_),
    .A3(_1161_),
    .A4(_1172_),
    .B1(_1185_),
    .X(_1197_));
 sky130_fd_sc_hd__a31o_1 _2879_ (.A1(_1196_),
    .A2(_1197_),
    .A3(_1171_),
    .B1(_1147_),
    .X(_1198_));
 sky130_fd_sc_hd__a31o_1 _2880_ (.A1(_1194_),
    .A2(_1142_),
    .A3(_1195_),
    .B1(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__o31a_1 _2881_ (.A1(_1135_),
    .A2(_1185_),
    .A3(_1187_),
    .B1(_1199_),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_2 _2882_ (.A(net72),
    .X(_1200_));
 sky130_fd_sc_hd__o221ai_4 _2883_ (.A1(net70),
    .A2(\po_0.muxf_0.rf_w_data[3] ),
    .B1(net71),
    .B2(\po_0.muxf_0.rf_w_data[4] ),
    .C1(_1192_),
    .Y(_1201_));
 sky130_fd_sc_hd__o21ai_1 _2884_ (.A1(_1189_),
    .A2(_1190_),
    .B1(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__nand2_1 _2885_ (.A(net72),
    .B(\po_0.muxf_0.rf_w_data[5] ),
    .Y(_1203_));
 sky130_fd_sc_hd__or2_1 _2886_ (.A(_1200_),
    .B(_0566_),
    .X(_1204_));
 sky130_fd_sc_hd__a311oi_1 _2887_ (.A1(_1202_),
    .A2(_1203_),
    .A3(_1204_),
    .B1(_1139_),
    .C1(_1171_),
    .Y(_1205_));
 sky130_fd_sc_hd__a21o_1 _2888_ (.A1(_1204_),
    .A2(_1203_),
    .B1(_1202_),
    .X(_1206_));
 sky130_fd_sc_hd__clkbuf_2 _2889_ (.A(_1147_),
    .X(_1207_));
 sky130_fd_sc_hd__and4_1 _2890_ (.A(net99),
    .B(_1185_),
    .C(_1200_),
    .D(_1166_),
    .X(_1208_));
 sky130_fd_sc_hd__clkbuf_2 _2891_ (.A(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__a31o_1 _2892_ (.A1(_1172_),
    .A2(_1185_),
    .A3(_1166_),
    .B1(_1200_),
    .X(_1210_));
 sky130_fd_sc_hd__and3b_1 _2893_ (.A_N(_1209_),
    .B(_1210_),
    .C(_1144_),
    .X(_1211_));
 sky130_fd_sc_hd__a211o_1 _2894_ (.A1(_1205_),
    .A2(_1206_),
    .B1(_1207_),
    .C1(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__o31a_1 _2895_ (.A1(_1135_),
    .A2(_1200_),
    .A3(_1187_),
    .B1(_1212_),
    .X(_0229_));
 sky130_fd_sc_hd__clkbuf_2 _2896_ (.A(net98),
    .X(_1213_));
 sky130_fd_sc_hd__or3_1 _2897_ (.A(\uc_0._01_ ),
    .B(_1139_),
    .C(_1144_),
    .X(_1214_));
 sky130_fd_sc_hd__clkbuf_2 _2898_ (.A(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__nand2_1 _2899_ (.A(_1213_),
    .B(_1209_),
    .Y(_1216_));
 sky130_fd_sc_hd__a41o_1 _2900_ (.A1(_1172_),
    .A2(_1185_),
    .A3(_1200_),
    .A4(_1166_),
    .B1(_1213_),
    .X(_1217_));
 sky130_fd_sc_hd__a31o_1 _2901_ (.A1(_1216_),
    .A2(_1145_),
    .A3(_1217_),
    .B1(_1207_),
    .X(_1218_));
 sky130_fd_sc_hd__nand2_1 _2902_ (.A(net98),
    .B(\po_0.muxf_0.rf_w_data[6] ),
    .Y(_1219_));
 sky130_fd_sc_hd__or2_1 _2903_ (.A(net98),
    .B(\po_0.muxf_0.rf_w_data[6] ),
    .X(_1220_));
 sky130_fd_sc_hd__o211ai_2 _2904_ (.A1(_1189_),
    .A2(_1190_),
    .B1(_1203_),
    .C1(_1201_),
    .Y(_1221_));
 sky130_fd_sc_hd__a22o_1 _2905_ (.A1(_1219_),
    .A2(_1220_),
    .B1(_1221_),
    .B2(_1204_),
    .X(_1222_));
 sky130_fd_sc_hd__o2111ai_2 _2906_ (.A1(_1200_),
    .A2(\po_0.muxf_0.rf_w_data[5] ),
    .B1(_1219_),
    .C1(_1220_),
    .D1(_1221_),
    .Y(_1223_));
 sky130_fd_sc_hd__and3_1 _2907_ (.A(_1222_),
    .B(_1142_),
    .C(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__o22a_1 _2908_ (.A1(_1213_),
    .A2(_1215_),
    .B1(_1218_),
    .B2(_1224_),
    .X(_0230_));
 sky130_fd_sc_hd__clkbuf_2 _2909_ (.A(net74),
    .X(_1225_));
 sky130_fd_sc_hd__or2_2 _2910_ (.A(_1225_),
    .B(_0570_),
    .X(_1226_));
 sky130_fd_sc_hd__nand2_1 _2911_ (.A(net74),
    .B(\po_0.muxf_0.rf_w_data[7] ),
    .Y(_1227_));
 sky130_fd_sc_hd__and2_1 _2912_ (.A(_1219_),
    .B(_1220_),
    .X(_1228_));
 sky130_fd_sc_hd__a32o_1 _2913_ (.A1(_1204_),
    .A2(_1221_),
    .A3(_1228_),
    .B1(net98),
    .B2(_0568_),
    .X(_1229_));
 sky130_fd_sc_hd__a21oi_1 _2914_ (.A1(_1226_),
    .A2(_1227_),
    .B1(_1229_),
    .Y(_1230_));
 sky130_fd_sc_hd__a31o_1 _2915_ (.A1(_1229_),
    .A2(_1226_),
    .A3(_1227_),
    .B1(_1186_),
    .X(_1231_));
 sky130_fd_sc_hd__a21oi_1 _2916_ (.A1(_1213_),
    .A2(_1209_),
    .B1(_1225_),
    .Y(_1232_));
 sky130_fd_sc_hd__and3_1 _2917_ (.A(net98),
    .B(net74),
    .C(_1208_),
    .X(_1233_));
 sky130_fd_sc_hd__clkbuf_2 _2918_ (.A(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__or3b_1 _2919_ (.A(_1232_),
    .B(_1234_),
    .C_N(_1171_),
    .X(_1235_));
 sky130_fd_sc_hd__o211ai_1 _2920_ (.A1(_1230_),
    .A2(_1231_),
    .B1(_1235_),
    .C1(_1215_),
    .Y(_1236_));
 sky130_fd_sc_hd__o31a_1 _2921_ (.A1(_1135_),
    .A2(_1225_),
    .A3(_1187_),
    .B1(_1236_),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_2 _2922_ (.A(net97),
    .X(_1237_));
 sky130_fd_sc_hd__nand2_1 _2923_ (.A(_1237_),
    .B(_1234_),
    .Y(_1238_));
 sky130_fd_sc_hd__a31o_1 _2924_ (.A1(_1213_),
    .A2(_1225_),
    .A3(_1209_),
    .B1(_1237_),
    .X(_1239_));
 sky130_fd_sc_hd__a31o_1 _2925_ (.A1(_1238_),
    .A2(_1145_),
    .A3(_1239_),
    .B1(_1207_),
    .X(_1240_));
 sky130_fd_sc_hd__nand3_2 _2926_ (.A(_1219_),
    .B(_1223_),
    .C(_1227_),
    .Y(_1241_));
 sky130_fd_sc_hd__o21a_1 _2927_ (.A1(net74),
    .A2(\po_0.muxf_0.rf_w_data[7] ),
    .B1(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__clkbuf_2 _2928_ (.A(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__a31o_1 _2929_ (.A1(_1241_),
    .A2(_1237_),
    .A3(_1226_),
    .B1(_1186_),
    .X(_1244_));
 sky130_fd_sc_hd__o21ba_1 _2930_ (.A1(_1237_),
    .A2(_1243_),
    .B1_N(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__o22a_1 _2931_ (.A1(_1237_),
    .A2(_1215_),
    .B1(_1240_),
    .B2(_1245_),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_2 _2932_ (.A(net76),
    .X(_1246_));
 sky130_fd_sc_hd__a41o_1 _2933_ (.A1(net73),
    .A2(_1225_),
    .A3(net97),
    .A4(_1209_),
    .B1(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__clkbuf_2 _2934_ (.A(net97),
    .X(_1248_));
 sky130_fd_sc_hd__clkbuf_2 _2935_ (.A(_1246_),
    .X(_1249_));
 sky130_fd_sc_hd__nand3_1 _2936_ (.A(_1248_),
    .B(_1249_),
    .C(_1234_),
    .Y(_1250_));
 sky130_fd_sc_hd__a311oi_1 _2937_ (.A1(_1248_),
    .A2(_1246_),
    .A3(_1242_),
    .B1(_1144_),
    .C1(_1139_),
    .Y(_1251_));
 sky130_fd_sc_hd__a31o_1 _2938_ (.A1(_1241_),
    .A2(net97),
    .A3(_1226_),
    .B1(_1246_),
    .X(_1252_));
 sky130_fd_sc_hd__a32o_1 _2939_ (.A1(_1171_),
    .A2(_1247_),
    .A3(_1250_),
    .B1(_1251_),
    .B2(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__mux2_1 _2940_ (.A0(_1253_),
    .A1(_1249_),
    .S(_1148_),
    .X(_1254_));
 sky130_fd_sc_hd__clkbuf_1 _2941_ (.A(_1254_),
    .X(_0233_));
 sky130_fd_sc_hd__a31o_1 _2942_ (.A1(net97),
    .A2(_1246_),
    .A3(_1233_),
    .B1(net62),
    .X(_1255_));
 sky130_fd_sc_hd__clkbuf_2 _2943_ (.A(net62),
    .X(_1256_));
 sky130_fd_sc_hd__nand4_1 _2944_ (.A(_1248_),
    .B(_1249_),
    .C(_1256_),
    .D(_1233_),
    .Y(_1257_));
 sky130_fd_sc_hd__a41oi_1 _2945_ (.A1(_1248_),
    .A2(_1249_),
    .A3(_1256_),
    .A4(_1243_),
    .B1(_1186_),
    .Y(_1258_));
 sky130_fd_sc_hd__a31o_1 _2946_ (.A1(_1248_),
    .A2(_1246_),
    .A3(_1242_),
    .B1(_1256_),
    .X(_1259_));
 sky130_fd_sc_hd__a32o_1 _2947_ (.A1(_1144_),
    .A2(_1255_),
    .A3(_1257_),
    .B1(_1258_),
    .B2(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__mux2_1 _2948_ (.A0(_1260_),
    .A1(_1256_),
    .S(_1148_),
    .X(_1261_));
 sky130_fd_sc_hd__clkbuf_1 _2949_ (.A(_1261_),
    .X(_0234_));
 sky130_fd_sc_hd__a41o_1 _2950_ (.A1(_1248_),
    .A2(_1249_),
    .A3(_1256_),
    .A4(_1234_),
    .B1(net63),
    .X(_1262_));
 sky130_fd_sc_hd__and4_1 _2951_ (.A(net97),
    .B(net76),
    .C(net62),
    .D(net63),
    .X(_1263_));
 sky130_fd_sc_hd__clkbuf_2 _2952_ (.A(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__nand2_1 _2953_ (.A(_1234_),
    .B(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__a31o_1 _2954_ (.A1(_1262_),
    .A2(_1265_),
    .A3(_1145_),
    .B1(_1207_),
    .X(_1266_));
 sky130_fd_sc_hd__a41oi_1 _2955_ (.A1(_1237_),
    .A2(_1249_),
    .A3(_1256_),
    .A4(_1243_),
    .B1(net63),
    .Y(_1267_));
 sky130_fd_sc_hd__a311oi_1 _2956_ (.A1(_1226_),
    .A2(_1241_),
    .A3(_1264_),
    .B1(_1187_),
    .C1(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hd__o22a_1 _2957_ (.A1(net63),
    .A2(_1215_),
    .B1(_1266_),
    .B2(_1268_),
    .X(_0235_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2958_ (.A(net64),
    .X(_1269_));
 sky130_fd_sc_hd__nand3_1 _2959_ (.A(_1269_),
    .B(_1234_),
    .C(_1264_),
    .Y(_1270_));
 sky130_fd_sc_hd__a41o_1 _2960_ (.A1(_1213_),
    .A2(_1225_),
    .A3(_1209_),
    .A4(_1263_),
    .B1(_1269_),
    .X(_1271_));
 sky130_fd_sc_hd__a31o_1 _2961_ (.A1(_1270_),
    .A2(_1145_),
    .A3(_1271_),
    .B1(_1207_),
    .X(_1272_));
 sky130_fd_sc_hd__a21oi_1 _2962_ (.A1(_1243_),
    .A2(_1264_),
    .B1(_1269_),
    .Y(_1273_));
 sky130_fd_sc_hd__a311oi_1 _2963_ (.A1(_1269_),
    .A2(_1243_),
    .A3(_1264_),
    .B1(_1187_),
    .C1(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__o22a_1 _2964_ (.A1(_1269_),
    .A2(_1215_),
    .B1(_1272_),
    .B2(_1274_),
    .X(_0236_));
 sky130_fd_sc_hd__a31oi_1 _2965_ (.A1(_1269_),
    .A2(_1243_),
    .A3(_1264_),
    .B1(net65),
    .Y(_1275_));
 sky130_fd_sc_hd__and4_1 _2966_ (.A(net64),
    .B(net65),
    .C(_1242_),
    .D(_1263_),
    .X(_1276_));
 sky130_fd_sc_hd__and4_1 _2967_ (.A(net64),
    .B(net65),
    .C(_1233_),
    .D(_1263_),
    .X(_1277_));
 sky130_fd_sc_hd__a31o_1 _2968_ (.A1(net64),
    .A2(_1233_),
    .A3(_1263_),
    .B1(net65),
    .X(_1278_));
 sky130_fd_sc_hd__nand3b_1 _2969_ (.A_N(_1277_),
    .B(_1171_),
    .C(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__o311a_1 _2970_ (.A1(_1275_),
    .A2(_1186_),
    .A3(_1276_),
    .B1(_1279_),
    .C1(_1214_),
    .X(_1280_));
 sky130_fd_sc_hd__o21ba_1 _2971_ (.A1(net65),
    .A2(_1215_),
    .B1_N(_1280_),
    .X(_0237_));
 sky130_fd_sc_hd__o21ba_1 _2972_ (.A1(\uc_0._01_ ),
    .A2(_1139_),
    .B1_N(_1144_),
    .X(_1281_));
 sky130_fd_sc_hd__and3_1 _2973_ (.A(_1140_),
    .B(net96),
    .C(_1277_),
    .X(_1282_));
 sky130_fd_sc_hd__nor2_1 _2974_ (.A(_1281_),
    .B(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__o31a_1 _2975_ (.A1(net96),
    .A2(_1147_),
    .A3(_1277_),
    .B1(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__a21oi_1 _2976_ (.A1(net96),
    .A2(_1276_),
    .B1(_1186_),
    .Y(_1285_));
 sky130_fd_sc_hd__o21a_1 _2977_ (.A1(net96),
    .A2(_1276_),
    .B1(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__o32a_1 _2978_ (.A1(_1135_),
    .A2(_1187_),
    .A3(net96),
    .B1(_1284_),
    .B2(_1286_),
    .X(_0238_));
 sky130_fd_sc_hd__a31oi_1 _2979_ (.A1(net66),
    .A2(_1142_),
    .A3(_1276_),
    .B1(_1282_),
    .Y(_1287_));
 sky130_fd_sc_hd__o21ai_1 _2980_ (.A1(_1285_),
    .A2(_1283_),
    .B1(net67),
    .Y(_1288_));
 sky130_fd_sc_hd__o31ai_1 _2981_ (.A1(net67),
    .A2(_1207_),
    .A3(_1287_),
    .B1(_1288_),
    .Y(_0239_));
 sky130_fd_sc_hd__buf_2 _2982_ (.A(\uc_0._03_ ),
    .X(_1289_));
 sky130_fd_sc_hd__mux2_1 _2983_ (.A0(_0704_),
    .A1(net17),
    .S(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _2984_ (.A(_1290_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(_0724_),
    .A1(net24),
    .S(_1289_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _2986_ (.A(_1291_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _2987_ (.A0(_0734_),
    .A1(net25),
    .S(_1289_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _2988_ (.A(_1292_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(_0744_),
    .A1(net26),
    .S(_1289_),
    .X(_1293_));
 sky130_fd_sc_hd__clkbuf_1 _2990_ (.A(_1293_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _2991_ (.A0(_0557_),
    .A1(net27),
    .S(_1289_),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _2992_ (.A(_1294_),
    .X(_0244_));
 sky130_fd_sc_hd__clkbuf_4 _2993_ (.A(\uc_0._03_ ),
    .X(_1295_));
 sky130_fd_sc_hd__buf_2 _2994_ (.A(_1295_),
    .X(_1296_));
 sky130_fd_sc_hd__mux2_1 _2995_ (.A0(_0566_),
    .A1(net28),
    .S(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_1 _2996_ (.A(_1297_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(_0568_),
    .A1(net29),
    .S(_1296_),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_1 _2998_ (.A(_1298_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _2999_ (.A0(_0570_),
    .A1(net30),
    .S(_1296_),
    .X(_1299_));
 sky130_fd_sc_hd__clkbuf_1 _3000_ (.A(_1299_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _3001_ (.A0(\uc_0._20_[8] ),
    .A1(net31),
    .S(_1296_),
    .X(_1300_));
 sky130_fd_sc_hd__clkbuf_1 _3002_ (.A(_1300_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _3003_ (.A0(\uc_0._20_[9] ),
    .A1(net32),
    .S(_1296_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_1 _3004_ (.A(_1301_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _3005_ (.A0(\uc_0._20_[10] ),
    .A1(net18),
    .S(_1296_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _3006_ (.A(_1302_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _3007_ (.A0(\uc_0._20_[11] ),
    .A1(net19),
    .S(_1295_),
    .X(_1303_));
 sky130_fd_sc_hd__clkbuf_1 _3008_ (.A(_1303_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(net79),
    .A1(net20),
    .S(_1295_),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_1 _3010_ (.A(_1304_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _3011_ (.A0(net80),
    .A1(net21),
    .S(_1295_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_1 _3012_ (.A(_1305_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _3013_ (.A0(net81),
    .A1(net22),
    .S(_1295_),
    .X(_1306_));
 sky130_fd_sc_hd__clkbuf_1 _3014_ (.A(_1306_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _3015_ (.A0(net82),
    .A1(net23),
    .S(_1295_),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_1 _3016_ (.A(_1307_),
    .X(_0255_));
 sky130_fd_sc_hd__nor4_1 _3017_ (.A(_0559_),
    .B(\uc_0.bc_0._54_[3] ),
    .C(\uc_0.bc_0._54_[2] ),
    .D(\uc_0.bc_0._54_[1] ),
    .Y(_1308_));
 sky130_fd_sc_hd__nor4_1 _3018_ (.A(_0572_),
    .B(\uc_0.bc_0._54_[0] ),
    .C(\uc_0.bc_0._54_[3] ),
    .D(\uc_0.bc_0._54_[2] ),
    .Y(_1309_));
 sky130_fd_sc_hd__nor2_1 _3019_ (.A(_1308_),
    .B(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__buf_2 _3020_ (.A(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__o21a_1 _3021_ (.A1(_1440_),
    .A2(_1139_),
    .B1(_1311_),
    .X(_0256_));
 sky130_fd_sc_hd__and4b_4 _3022_ (.A_N(_0882_),
    .B(_0906_),
    .C(_1039_),
    .D(_0886_),
    .X(_1312_));
 sky130_fd_sc_hd__buf_2 _3023_ (.A(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__mux2_1 _3024_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(_0713_),
    .S(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__clkbuf_1 _3025_ (.A(_1314_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _3026_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(_0731_),
    .S(_1313_),
    .X(_1315_));
 sky130_fd_sc_hd__clkbuf_1 _3027_ (.A(_1315_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _3028_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(_0741_),
    .S(_1313_),
    .X(_1316_));
 sky130_fd_sc_hd__clkbuf_1 _3029_ (.A(_1316_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _3030_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(_0752_),
    .S(_1313_),
    .X(_1317_));
 sky130_fd_sc_hd__clkbuf_1 _3031_ (.A(_1317_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _3032_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(_0762_),
    .S(_1313_),
    .X(_1318_));
 sky130_fd_sc_hd__clkbuf_1 _3033_ (.A(_1318_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _3034_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(_0772_),
    .S(_1313_),
    .X(_1319_));
 sky130_fd_sc_hd__clkbuf_1 _3035_ (.A(_1319_),
    .X(_0262_));
 sky130_fd_sc_hd__buf_2 _3036_ (.A(_1312_),
    .X(_1320_));
 sky130_fd_sc_hd__mux2_1 _3037_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(_0782_),
    .S(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__clkbuf_1 _3038_ (.A(_1321_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _3039_ (.A0(\po_0.regf_0.rf[4][7] ),
    .A1(_0795_),
    .S(_1320_),
    .X(_1322_));
 sky130_fd_sc_hd__clkbuf_1 _3040_ (.A(_1322_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _3041_ (.A0(\po_0.regf_0.rf[4][8] ),
    .A1(_0810_),
    .S(_1320_),
    .X(_1323_));
 sky130_fd_sc_hd__clkbuf_1 _3042_ (.A(_1323_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _3043_ (.A0(\po_0.regf_0.rf[4][9] ),
    .A1(_0819_),
    .S(_1320_),
    .X(_1324_));
 sky130_fd_sc_hd__clkbuf_1 _3044_ (.A(_1324_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _3045_ (.A0(\po_0.regf_0.rf[4][10] ),
    .A1(_0829_),
    .S(_1320_),
    .X(_1325_));
 sky130_fd_sc_hd__clkbuf_1 _3046_ (.A(_1325_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _3047_ (.A0(\po_0.regf_0.rf[4][11] ),
    .A1(_0838_),
    .S(_1320_),
    .X(_1326_));
 sky130_fd_sc_hd__clkbuf_1 _3048_ (.A(_1326_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _3049_ (.A0(\po_0.regf_0.rf[4][12] ),
    .A1(_0848_),
    .S(_1312_),
    .X(_1327_));
 sky130_fd_sc_hd__clkbuf_1 _3050_ (.A(_1327_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _3051_ (.A0(\po_0.regf_0.rf[4][13] ),
    .A1(_0858_),
    .S(_1312_),
    .X(_1328_));
 sky130_fd_sc_hd__clkbuf_1 _3052_ (.A(_1328_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _3053_ (.A0(\po_0.regf_0.rf[4][14] ),
    .A1(_0870_),
    .S(_1312_),
    .X(_1329_));
 sky130_fd_sc_hd__clkbuf_1 _3054_ (.A(_1329_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _3055_ (.A0(\po_0.regf_0.rf[4][15] ),
    .A1(_0879_),
    .S(_1312_),
    .X(_1330_));
 sky130_fd_sc_hd__clkbuf_1 _3056_ (.A(_1330_),
    .X(_0272_));
 sky130_fd_sc_hd__and4bb_4 _3057_ (.A_N(_0886_),
    .B_N(\po_0.regf_0.w_addr[3] ),
    .C(_0906_),
    .D(_0717_),
    .X(_1331_));
 sky130_fd_sc_hd__buf_2 _3058_ (.A(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(\po_0.regf_0.rf[3][0] ),
    .A1(_0713_),
    .S(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__clkbuf_1 _3060_ (.A(_1333_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(\po_0.regf_0.rf[3][1] ),
    .A1(_0731_),
    .S(_1332_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_1 _3062_ (.A(_1334_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _3063_ (.A0(\po_0.regf_0.rf[3][2] ),
    .A1(_0741_),
    .S(_1332_),
    .X(_1335_));
 sky130_fd_sc_hd__clkbuf_1 _3064_ (.A(_1335_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _3065_ (.A0(\po_0.regf_0.rf[3][3] ),
    .A1(_0752_),
    .S(_1332_),
    .X(_1336_));
 sky130_fd_sc_hd__clkbuf_1 _3066_ (.A(_1336_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _3067_ (.A0(\po_0.regf_0.rf[3][4] ),
    .A1(_0762_),
    .S(_1332_),
    .X(_1337_));
 sky130_fd_sc_hd__clkbuf_1 _3068_ (.A(_1337_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _3069_ (.A0(\po_0.regf_0.rf[3][5] ),
    .A1(_0772_),
    .S(_1332_),
    .X(_1338_));
 sky130_fd_sc_hd__clkbuf_1 _3070_ (.A(_1338_),
    .X(_0278_));
 sky130_fd_sc_hd__buf_2 _3071_ (.A(_1331_),
    .X(_1339_));
 sky130_fd_sc_hd__mux2_1 _3072_ (.A0(\po_0.regf_0.rf[3][6] ),
    .A1(_0782_),
    .S(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__clkbuf_1 _3073_ (.A(_1340_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _3074_ (.A0(\po_0.regf_0.rf[3][7] ),
    .A1(_0795_),
    .S(_1339_),
    .X(_1341_));
 sky130_fd_sc_hd__clkbuf_1 _3075_ (.A(_1341_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _3076_ (.A0(\po_0.regf_0.rf[3][8] ),
    .A1(_0810_),
    .S(_1339_),
    .X(_1342_));
 sky130_fd_sc_hd__clkbuf_1 _3077_ (.A(_1342_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _3078_ (.A0(\po_0.regf_0.rf[3][9] ),
    .A1(_0819_),
    .S(_1339_),
    .X(_1343_));
 sky130_fd_sc_hd__clkbuf_1 _3079_ (.A(_1343_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _3080_ (.A0(\po_0.regf_0.rf[3][10] ),
    .A1(_0829_),
    .S(_1339_),
    .X(_1344_));
 sky130_fd_sc_hd__clkbuf_1 _3081_ (.A(_1344_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _3082_ (.A0(\po_0.regf_0.rf[3][11] ),
    .A1(_0838_),
    .S(_1339_),
    .X(_1345_));
 sky130_fd_sc_hd__clkbuf_1 _3083_ (.A(_1345_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _3084_ (.A0(\po_0.regf_0.rf[3][12] ),
    .A1(_0848_),
    .S(_1331_),
    .X(_1346_));
 sky130_fd_sc_hd__clkbuf_1 _3085_ (.A(_1346_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _3086_ (.A0(\po_0.regf_0.rf[3][13] ),
    .A1(_0858_),
    .S(_1331_),
    .X(_1347_));
 sky130_fd_sc_hd__clkbuf_1 _3087_ (.A(_1347_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _3088_ (.A0(\po_0.regf_0.rf[3][14] ),
    .A1(_0870_),
    .S(_1331_),
    .X(_1348_));
 sky130_fd_sc_hd__clkbuf_1 _3089_ (.A(_1348_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _3090_ (.A0(\po_0.regf_0.rf[3][15] ),
    .A1(_0879_),
    .S(_1331_),
    .X(_1349_));
 sky130_fd_sc_hd__clkbuf_1 _3091_ (.A(_1349_),
    .X(_0288_));
 sky130_fd_sc_hd__and4bb_4 _3092_ (.A_N(_0886_),
    .B_N(\po_0.regf_0.w_addr[3] ),
    .C(_0906_),
    .D(_0885_),
    .X(_1350_));
 sky130_fd_sc_hd__buf_2 _3093_ (.A(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__mux2_1 _3094_ (.A0(\po_0.regf_0.rf[2][0] ),
    .A1(_0713_),
    .S(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__clkbuf_1 _3095_ (.A(_1352_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _3096_ (.A0(\po_0.regf_0.rf[2][1] ),
    .A1(_0731_),
    .S(_1351_),
    .X(_1353_));
 sky130_fd_sc_hd__clkbuf_1 _3097_ (.A(_1353_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _3098_ (.A0(\po_0.regf_0.rf[2][2] ),
    .A1(_0741_),
    .S(_1351_),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_1 _3099_ (.A(_1354_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _3100_ (.A0(\po_0.regf_0.rf[2][3] ),
    .A1(_0752_),
    .S(_1351_),
    .X(_1355_));
 sky130_fd_sc_hd__clkbuf_1 _3101_ (.A(_1355_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _3102_ (.A0(\po_0.regf_0.rf[2][4] ),
    .A1(_0762_),
    .S(_1351_),
    .X(_1356_));
 sky130_fd_sc_hd__clkbuf_1 _3103_ (.A(_1356_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _3104_ (.A0(\po_0.regf_0.rf[2][5] ),
    .A1(_0772_),
    .S(_1351_),
    .X(_1357_));
 sky130_fd_sc_hd__clkbuf_1 _3105_ (.A(_1357_),
    .X(_0294_));
 sky130_fd_sc_hd__buf_2 _3106_ (.A(_1350_),
    .X(_1358_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(\po_0.regf_0.rf[2][6] ),
    .A1(_0782_),
    .S(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__clkbuf_1 _3108_ (.A(_1359_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _3109_ (.A0(\po_0.regf_0.rf[2][7] ),
    .A1(_0795_),
    .S(_1358_),
    .X(_1360_));
 sky130_fd_sc_hd__clkbuf_1 _3110_ (.A(_1360_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _3111_ (.A0(\po_0.regf_0.rf[2][8] ),
    .A1(_0810_),
    .S(_1358_),
    .X(_1361_));
 sky130_fd_sc_hd__clkbuf_1 _3112_ (.A(_1361_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _3113_ (.A0(\po_0.regf_0.rf[2][9] ),
    .A1(_0819_),
    .S(_1358_),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _3114_ (.A(_1362_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _3115_ (.A0(\po_0.regf_0.rf[2][10] ),
    .A1(_0829_),
    .S(_1358_),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_1 _3116_ (.A(_1363_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _3117_ (.A0(\po_0.regf_0.rf[2][11] ),
    .A1(_0838_),
    .S(_1358_),
    .X(_1364_));
 sky130_fd_sc_hd__clkbuf_1 _3118_ (.A(_1364_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _3119_ (.A0(\po_0.regf_0.rf[2][12] ),
    .A1(_0848_),
    .S(_1350_),
    .X(_1365_));
 sky130_fd_sc_hd__clkbuf_1 _3120_ (.A(_1365_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _3121_ (.A0(\po_0.regf_0.rf[2][13] ),
    .A1(_0858_),
    .S(_1350_),
    .X(_1366_));
 sky130_fd_sc_hd__clkbuf_1 _3122_ (.A(_1366_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _3123_ (.A0(\po_0.regf_0.rf[2][14] ),
    .A1(_0870_),
    .S(_1350_),
    .X(_1367_));
 sky130_fd_sc_hd__clkbuf_1 _3124_ (.A(_1367_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _3125_ (.A0(\po_0.regf_0.rf[2][15] ),
    .A1(_0879_),
    .S(_1350_),
    .X(_1368_));
 sky130_fd_sc_hd__clkbuf_1 _3126_ (.A(_1368_),
    .X(_0304_));
 sky130_fd_sc_hd__a32o_1 _3127_ (.A1(_0572_),
    .A2(_0559_),
    .A3(\uc_0.bc_0._54_[3] ),
    .B1(_0558_),
    .B2(_1407_),
    .X(_0305_));
 sky130_fd_sc_hd__a21bo_1 _3128_ (.A1(_1403_),
    .A2(_0561_),
    .B1_N(_0558_),
    .X(_0306_));
 sky130_fd_sc_hd__a21o_1 _3129_ (.A1(net92),
    .A2(_1311_),
    .B1(_0564_),
    .X(_0307_));
 sky130_fd_sc_hd__a21bo_1 _3130_ (.A1(net88),
    .A2(_1311_),
    .B1_N(_0575_),
    .X(_0308_));
 sky130_fd_sc_hd__or4_2 _3131_ (.A(_1440_),
    .B(_1432_),
    .C(_1439_),
    .D(_1451_),
    .X(_1369_));
 sky130_fd_sc_hd__or3_2 _3132_ (.A(_1441_),
    .B(_0559_),
    .C(_1451_),
    .X(_1370_));
 sky130_fd_sc_hd__and2_1 _3133_ (.A(_0558_),
    .B(_0561_),
    .X(_1371_));
 sky130_fd_sc_hd__o211ai_4 _3134_ (.A1(\uc_0.bc_0._54_[0] ),
    .A2(_1369_),
    .B1(_1370_),
    .C1(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__a21o_1 _3135_ (.A1(_0716_),
    .A2(_1311_),
    .B1(_1372_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _3136_ (.A0(\po_0.regf_0.rq_addr[0] ),
    .A1(_0557_),
    .S(_0563_),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_1 _3137_ (.A(_1373_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _3138_ (.A0(\po_0.regf_0.rq_addr[1] ),
    .A1(_0566_),
    .S(_0563_),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_1 _3139_ (.A(_1374_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _3140_ (.A0(\po_0.regf_0.rq_addr[2] ),
    .A1(_0568_),
    .S(_0563_),
    .X(_1375_));
 sky130_fd_sc_hd__clkbuf_1 _3141_ (.A(_1375_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _3142_ (.A0(\po_0.regf_0.rq_addr[3] ),
    .A1(_0570_),
    .S(_0563_),
    .X(_1376_));
 sky130_fd_sc_hd__clkbuf_1 _3143_ (.A(_1376_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _3144_ (.A0(\uc_0._20_[8] ),
    .A1(\po_0.regf_0.rp_addr[0] ),
    .S(_0575_),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_1 _3145_ (.A(_1377_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _3146_ (.A0(\uc_0._20_[9] ),
    .A1(\po_0.regf_0.rp_addr[1] ),
    .S(_0574_),
    .X(_1378_));
 sky130_fd_sc_hd__clkbuf_1 _3147_ (.A(_1378_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _3148_ (.A0(\uc_0._20_[10] ),
    .A1(\po_0.regf_0.rp_addr[2] ),
    .S(_0574_),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _3149_ (.A(_1379_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _3150_ (.A0(\uc_0._20_[11] ),
    .A1(\po_0.regf_0.rp_addr[3] ),
    .S(_0574_),
    .X(_1380_));
 sky130_fd_sc_hd__clkbuf_1 _3151_ (.A(_1380_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _3152_ (.A0(\uc_0._20_[8] ),
    .A1(_0704_),
    .S(_0563_),
    .X(_1381_));
 sky130_fd_sc_hd__mux2_1 _3153_ (.A0(_0883_),
    .A1(_1381_),
    .S(_1372_),
    .X(_1382_));
 sky130_fd_sc_hd__clkbuf_1 _3154_ (.A(_1382_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _3155_ (.A0(\uc_0._20_[9] ),
    .A1(_0724_),
    .S(_0562_),
    .X(_1383_));
 sky130_fd_sc_hd__mux2_1 _3156_ (.A0(_0884_),
    .A1(_1383_),
    .S(_1372_),
    .X(_1384_));
 sky130_fd_sc_hd__clkbuf_1 _3157_ (.A(_1384_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _3158_ (.A0(\uc_0._20_[10] ),
    .A1(_0734_),
    .S(_0562_),
    .X(_1385_));
 sky130_fd_sc_hd__mux2_1 _3159_ (.A0(_0718_),
    .A1(_1385_),
    .S(_1372_),
    .X(_1386_));
 sky130_fd_sc_hd__clkbuf_1 _3160_ (.A(_1386_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _3161_ (.A0(\uc_0._20_[11] ),
    .A1(_0744_),
    .S(_0562_),
    .X(_1387_));
 sky130_fd_sc_hd__mux2_1 _3162_ (.A0(_0715_),
    .A1(_1387_),
    .S(_1372_),
    .X(_1388_));
 sky130_fd_sc_hd__clkbuf_1 _3163_ (.A(_1388_),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_2 _3164_ (.A(_1369_),
    .X(_1389_));
 sky130_fd_sc_hd__nor2_1 _3165_ (.A(\uc_0.bc_0._54_[0] ),
    .B(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__o211a_1 _3166_ (.A1(_0722_),
    .A2(_1390_),
    .B1(_1370_),
    .C1(_1371_),
    .X(_0322_));
 sky130_fd_sc_hd__a211oi_1 _3167_ (.A1(_0723_),
    .A2(_1370_),
    .B1(_1390_),
    .C1(_0564_),
    .Y(_0323_));
 sky130_fd_sc_hd__a32o_1 _3168_ (.A1(_0572_),
    .A2(\uc_0.bc_0._54_[0] ),
    .A3(\uc_0.bc_0._54_[2] ),
    .B1(_1311_),
    .B2(net60),
    .X(_0324_));
 sky130_fd_sc_hd__a2bb2o_1 _3169_ (.A1_N(_1389_),
    .A2_N(\uc_0.bc_0._54_[0] ),
    .B1(net59),
    .B2(_1311_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _3170_ (.A0(_0704_),
    .A1(net51),
    .S(_1389_),
    .X(_1391_));
 sky130_fd_sc_hd__clkbuf_1 _3171_ (.A(_1391_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _3172_ (.A0(_0724_),
    .A1(net52),
    .S(_1389_),
    .X(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _3173_ (.A(_1392_),
    .X(_0327_));
 sky130_fd_sc_hd__buf_4 _3174_ (.A(_1369_),
    .X(_1393_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(_0734_),
    .A1(net53),
    .S(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _3176_ (.A(_1394_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _3177_ (.A0(_0744_),
    .A1(net54),
    .S(_1393_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_1 _3178_ (.A(_1395_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _3179_ (.A0(_0557_),
    .A1(net55),
    .S(_1393_),
    .X(_1396_));
 sky130_fd_sc_hd__clkbuf_1 _3180_ (.A(_1396_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _3181_ (.A0(_0566_),
    .A1(net56),
    .S(_1393_),
    .X(_1397_));
 sky130_fd_sc_hd__clkbuf_1 _3182_ (.A(_1397_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _3183_ (.A0(_0568_),
    .A1(net57),
    .S(_1393_),
    .X(_1398_));
 sky130_fd_sc_hd__clkbuf_1 _3184_ (.A(_1398_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _3185_ (.A0(_0570_),
    .A1(net58),
    .S(_1393_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_1 _3186_ (.A(_1399_),
    .X(_0333_));
 sky130_fd_sc_hd__o31a_1 _3187_ (.A1(_0572_),
    .A2(_0559_),
    .A3(_0573_),
    .B1(_1389_),
    .X(_1400_));
 sky130_fd_sc_hd__o31a_1 _3188_ (.A1(net77),
    .A2(_1308_),
    .A3(_1309_),
    .B1(_1400_),
    .X(_0334_));
 sky130_fd_sc_hd__o21a_1 _3189_ (.A1(_1289_),
    .A2(_1309_),
    .B1(_1400_),
    .X(_0335_));
 sky130_fd_sc_hd__o221a_1 _3190_ (.A1(_0572_),
    .A2(_0573_),
    .B1(_1308_),
    .B2(_1145_),
    .C1(_1389_),
    .X(_0336_));
 sky130_fd_sc_hd__a32o_1 _3191_ (.A1(\uc_0.bc_0._54_[1] ),
    .A2(_0559_),
    .A3(_0560_),
    .B1(_1310_),
    .B2(_1135_),
    .X(_0337_));
 sky130_fd_sc_hd__dfxtp_1 _3192_ (.CLK(net134),
    .D(_0016_),
    .Q(\po_0.regf_0.rf[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3193_ (.CLK(net134),
    .D(_0017_),
    .Q(\po_0.regf_0.rf[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3194_ (.CLK(net127),
    .D(_0018_),
    .Q(\po_0.regf_0.rf[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3195_ (.CLK(net127),
    .D(_0019_),
    .Q(\po_0.regf_0.rf[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3196_ (.CLK(net135),
    .D(_0020_),
    .Q(\po_0.regf_0.rf[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3197_ (.CLK(net135),
    .D(_0021_),
    .Q(\po_0.regf_0.rf[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3198_ (.CLK(net108),
    .D(_0022_),
    .Q(\po_0.regf_0.rf[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3199_ (.CLK(net108),
    .D(_0023_),
    .Q(\po_0.regf_0.rf[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3200_ (.CLK(net102),
    .D(_0024_),
    .Q(\po_0.regf_0.rf[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3201_ (.CLK(net102),
    .D(_0025_),
    .Q(\po_0.regf_0.rf[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3202_ (.CLK(net100),
    .D(_0026_),
    .Q(\po_0.regf_0.rf[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3203_ (.CLK(net100),
    .D(_0027_),
    .Q(\po_0.regf_0.rf[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3204_ (.CLK(net109),
    .D(_0028_),
    .Q(\po_0.regf_0.rf[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3205_ (.CLK(net113),
    .D(_0029_),
    .Q(\po_0.regf_0.rf[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3206_ (.CLK(net109),
    .D(_0030_),
    .Q(\po_0.regf_0.rf[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3207_ (.CLK(net126),
    .D(_0031_),
    .Q(\po_0.regf_0.rf[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3208_ (.CLK(net134),
    .D(_0032_),
    .Q(\po_0.regf_0.rf[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3209_ (.CLK(net134),
    .D(_0033_),
    .Q(\po_0.regf_0.rf[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3210_ (.CLK(net127),
    .D(_0034_),
    .Q(\po_0.regf_0.rf[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3211_ (.CLK(net127),
    .D(_0035_),
    .Q(\po_0.regf_0.rf[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3212_ (.CLK(net135),
    .D(_0036_),
    .Q(\po_0.regf_0.rf[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3213_ (.CLK(net135),
    .D(_0037_),
    .Q(\po_0.regf_0.rf[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3214_ (.CLK(net111),
    .D(_0038_),
    .Q(\po_0.regf_0.rf[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3215_ (.CLK(net108),
    .D(_0039_),
    .Q(\po_0.regf_0.rf[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3216_ (.CLK(net102),
    .D(_0040_),
    .Q(\po_0.regf_0.rf[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3217_ (.CLK(net102),
    .D(_0041_),
    .Q(\po_0.regf_0.rf[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3218_ (.CLK(net100),
    .D(_0042_),
    .Q(\po_0.regf_0.rf[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3219_ (.CLK(net100),
    .D(_0043_),
    .Q(\po_0.regf_0.rf[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3220_ (.CLK(net109),
    .D(_0044_),
    .Q(\po_0.regf_0.rf[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3221_ (.CLK(net109),
    .D(_0045_),
    .Q(\po_0.regf_0.rf[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3222_ (.CLK(net109),
    .D(_0046_),
    .Q(\po_0.regf_0.rf[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3223_ (.CLK(net126),
    .D(_0047_),
    .Q(\po_0.regf_0.rf[6][15] ));
 sky130_fd_sc_hd__dlxtp_1 _3224_ (.D(\po_0.regf_0._5_[0] ),
    .GATE(net94),
    .Q(\po_0._1_[0] ));
 sky130_fd_sc_hd__dlxtp_1 _3225_ (.D(\po_0.regf_0._5_[1] ),
    .GATE(net94),
    .Q(\po_0._1_[1] ));
 sky130_fd_sc_hd__dlxtp_1 _3226_ (.D(\po_0.regf_0._5_[2] ),
    .GATE(net94),
    .Q(\po_0._1_[2] ));
 sky130_fd_sc_hd__dlxtp_1 _3227_ (.D(\po_0.regf_0._5_[3] ),
    .GATE(net94),
    .Q(\po_0._1_[3] ));
 sky130_fd_sc_hd__dlxtp_1 _3228_ (.D(\po_0.regf_0._5_[4] ),
    .GATE(net94),
    .Q(\po_0._1_[4] ));
 sky130_fd_sc_hd__dlxtp_1 _3229_ (.D(\po_0.regf_0._5_[5] ),
    .GATE(net95),
    .Q(\po_0._1_[5] ));
 sky130_fd_sc_hd__dlxtp_1 _3230_ (.D(\po_0.regf_0._5_[6] ),
    .GATE(net94),
    .Q(\po_0._1_[6] ));
 sky130_fd_sc_hd__dlxtp_1 _3231_ (.D(\po_0.regf_0._5_[7] ),
    .GATE(net92),
    .Q(\po_0._1_[7] ));
 sky130_fd_sc_hd__dlxtp_1 _3232_ (.D(\po_0.regf_0._5_[8] ),
    .GATE(net92),
    .Q(\po_0._1_[8] ));
 sky130_fd_sc_hd__dlxtp_1 _3233_ (.D(\po_0.regf_0._5_[9] ),
    .GATE(net92),
    .Q(\po_0._1_[9] ));
 sky130_fd_sc_hd__dlxtp_1 _3234_ (.D(\po_0.regf_0._5_[10] ),
    .GATE(net92),
    .Q(\po_0._1_[10] ));
 sky130_fd_sc_hd__dlxtp_1 _3235_ (.D(\po_0.regf_0._5_[11] ),
    .GATE(net93),
    .Q(\po_0._1_[11] ));
 sky130_fd_sc_hd__dlxtp_1 _3236_ (.D(\po_0.regf_0._5_[12] ),
    .GATE(net93),
    .Q(\po_0._1_[12] ));
 sky130_fd_sc_hd__dlxtp_1 _3237_ (.D(\po_0.regf_0._5_[13] ),
    .GATE(net92),
    .Q(\po_0._1_[13] ));
 sky130_fd_sc_hd__dlxtp_1 _3238_ (.D(\po_0.regf_0._5_[14] ),
    .GATE(net93),
    .Q(\po_0._1_[14] ));
 sky130_fd_sc_hd__dlxtp_1 _3239_ (.D(\po_0.regf_0._5_[15] ),
    .GATE(net93),
    .Q(\po_0._1_[15] ));
 sky130_fd_sc_hd__dlxtp_1 _3240_ (.D(\po_0.regf_0._3_[0] ),
    .GATE(net89),
    .Q(net35));
 sky130_fd_sc_hd__dlxtp_1 _3241_ (.D(\po_0.regf_0._3_[1] ),
    .GATE(net89),
    .Q(net42));
 sky130_fd_sc_hd__dlxtp_1 _3242_ (.D(\po_0.regf_0._3_[2] ),
    .GATE(net90),
    .Q(net43));
 sky130_fd_sc_hd__dlxtp_1 _3243_ (.D(\po_0.regf_0._3_[3] ),
    .GATE(net90),
    .Q(net44));
 sky130_fd_sc_hd__dlxtp_1 _3244_ (.D(\po_0.regf_0._3_[4] ),
    .GATE(net90),
    .Q(net45));
 sky130_fd_sc_hd__dlxtp_1 _3245_ (.D(\po_0.regf_0._3_[5] ),
    .GATE(net90),
    .Q(net46));
 sky130_fd_sc_hd__dlxtp_1 _3246_ (.D(\po_0.regf_0._3_[6] ),
    .GATE(net89),
    .Q(net47));
 sky130_fd_sc_hd__dlxtp_1 _3247_ (.D(\po_0.regf_0._3_[7] ),
    .GATE(net88),
    .Q(net48));
 sky130_fd_sc_hd__dlxtp_1 _3248_ (.D(\po_0.regf_0._3_[8] ),
    .GATE(net88),
    .Q(net49));
 sky130_fd_sc_hd__dlxtp_1 _3249_ (.D(\po_0.regf_0._3_[9] ),
    .GATE(net88),
    .Q(net50));
 sky130_fd_sc_hd__dlxtp_1 _3250_ (.D(\po_0.regf_0._3_[10] ),
    .GATE(net88),
    .Q(net36));
 sky130_fd_sc_hd__dlxtp_1 _3251_ (.D(\po_0.regf_0._3_[11] ),
    .GATE(net88),
    .Q(net37));
 sky130_fd_sc_hd__dlxtp_1 _3252_ (.D(\po_0.regf_0._3_[12] ),
    .GATE(net89),
    .Q(net38));
 sky130_fd_sc_hd__dlxtp_1 _3253_ (.D(\po_0.regf_0._3_[13] ),
    .GATE(net91),
    .Q(net39));
 sky130_fd_sc_hd__dlxtp_1 _3254_ (.D(\po_0.regf_0._3_[14] ),
    .GATE(net89),
    .Q(net40));
 sky130_fd_sc_hd__dlxtp_1 _3255_ (.D(\po_0.regf_0._3_[15] ),
    .GATE(net89),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _3256_ (.CLK(net134),
    .D(_0048_),
    .Q(\po_0.regf_0.rf[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3257_ (.CLK(net134),
    .D(_0049_),
    .Q(\po_0.regf_0.rf[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3258_ (.CLK(net133),
    .D(_0050_),
    .Q(\po_0.regf_0.rf[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3259_ (.CLK(net133),
    .D(_0051_),
    .Q(\po_0.regf_0.rf[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3260_ (.CLK(net135),
    .D(_0052_),
    .Q(\po_0.regf_0.rf[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3261_ (.CLK(net135),
    .D(_0053_),
    .Q(\po_0.regf_0.rf[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3262_ (.CLK(net108),
    .D(_0054_),
    .Q(\po_0.regf_0.rf[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3263_ (.CLK(net108),
    .D(_0055_),
    .Q(\po_0.regf_0.rf[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3264_ (.CLK(net102),
    .D(_0056_),
    .Q(\po_0.regf_0.rf[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3265_ (.CLK(net102),
    .D(_0057_),
    .Q(\po_0.regf_0.rf[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3266_ (.CLK(net100),
    .D(_0058_),
    .Q(\po_0.regf_0.rf[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3267_ (.CLK(net101),
    .D(_0059_),
    .Q(\po_0.regf_0.rf[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3268_ (.CLK(net109),
    .D(_0060_),
    .Q(\po_0.regf_0.rf[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3269_ (.CLK(net110),
    .D(_0061_),
    .Q(\po_0.regf_0.rf[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3270_ (.CLK(net126),
    .D(_0062_),
    .Q(\po_0.regf_0.rf[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3271_ (.CLK(net126),
    .D(_0063_),
    .Q(\po_0.regf_0.rf[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _3272_ (.CLK(net160),
    .D(_0008_),
    .Q(_0000_));
 sky130_fd_sc_hd__dfxtp_2 _3273_ (.CLK(net171),
    .D(_0009_),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_1 _3274_ (.CLK(net153),
    .D(_0010_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_2 _3275_ (.CLK(net159),
    .D(_0011_),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_1 _3276_ (.CLK(net173),
    .D(_0064_),
    .Q(\po_0.regf_0.rf[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3277_ (.CLK(net174),
    .D(_0065_),
    .Q(\po_0.regf_0.rf[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3278_ (.CLK(net173),
    .D(_0066_),
    .Q(\po_0.regf_0.rf[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3279_ (.CLK(net171),
    .D(_0067_),
    .Q(\po_0.regf_0.rf[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3280_ (.CLK(net146),
    .D(_0068_),
    .Q(\po_0.regf_0.rf[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3281_ (.CLK(net174),
    .D(_0069_),
    .Q(\po_0.regf_0.rf[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3282_ (.CLK(net152),
    .D(_0070_),
    .Q(\po_0.regf_0.rf[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3283_ (.CLK(net158),
    .D(_0071_),
    .Q(\po_0.regf_0.rf[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3284_ (.CLK(net119),
    .D(_0072_),
    .Q(\po_0.regf_0.rf[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3285_ (.CLK(net150),
    .D(_0073_),
    .Q(\po_0.regf_0.rf[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3286_ (.CLK(net152),
    .D(_0074_),
    .Q(\po_0.regf_0.rf[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3287_ (.CLK(net120),
    .D(_0075_),
    .Q(\po_0.regf_0.rf[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3288_ (.CLK(net170),
    .D(_0076_),
    .Q(\po_0.regf_0.rf[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3289_ (.CLK(net157),
    .D(_0077_),
    .Q(\po_0.regf_0.rf[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3290_ (.CLK(net157),
    .D(_0078_),
    .Q(\po_0.regf_0.rf[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3291_ (.CLK(net170),
    .D(_0079_),
    .Q(\po_0.regf_0.rf[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3292_ (.CLK(net147),
    .D(_0080_),
    .Q(\po_0.regf_0.rf[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3293_ (.CLK(net146),
    .D(_0081_),
    .Q(\po_0.regf_0.rf[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3294_ (.CLK(net141),
    .D(_0082_),
    .Q(\po_0.regf_0.rf[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3295_ (.CLK(net142),
    .D(_0083_),
    .Q(\po_0.regf_0.rf[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3296_ (.CLK(net146),
    .D(_0084_),
    .Q(\po_0.regf_0.rf[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3297_ (.CLK(net144),
    .D(_0085_),
    .Q(\po_0.regf_0.rf[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3298_ (.CLK(net122),
    .D(_0086_),
    .Q(\po_0.regf_0.rf[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3299_ (.CLK(net123),
    .D(_0087_),
    .Q(\po_0.regf_0.rf[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3300_ (.CLK(net119),
    .D(_0088_),
    .Q(\po_0.regf_0.rf[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3301_ (.CLK(net116),
    .D(_0089_),
    .Q(\po_0.regf_0.rf[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3302_ (.CLK(net117),
    .D(_0090_),
    .Q(\po_0.regf_0.rf[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3303_ (.CLK(net120),
    .D(_0091_),
    .Q(\po_0.regf_0.rf[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3304_ (.CLK(net141),
    .D(_0092_),
    .Q(\po_0.regf_0.rf[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3305_ (.CLK(net123),
    .D(_0093_),
    .Q(\po_0.regf_0.rf[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3306_ (.CLK(net122),
    .D(_0094_),
    .Q(\po_0.regf_0.rf[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3307_ (.CLK(net141),
    .D(_0095_),
    .Q(\po_0.regf_0.rf[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3308_ (.CLK(net144),
    .D(_0096_),
    .Q(\po_0.regf_0.rf[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3309_ (.CLK(net144),
    .D(_0097_),
    .Q(\po_0.regf_0.rf[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3310_ (.CLK(net140),
    .D(_0098_),
    .Q(\po_0.regf_0.rf[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3311_ (.CLK(net140),
    .D(_0099_),
    .Q(\po_0.regf_0.rf[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3312_ (.CLK(net144),
    .D(_0100_),
    .Q(\po_0.regf_0.rf[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3313_ (.CLK(net145),
    .D(_0101_),
    .Q(\po_0.regf_0.rf[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3314_ (.CLK(net118),
    .D(_0102_),
    .Q(\po_0.regf_0.rf[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3315_ (.CLK(net112),
    .D(_0103_),
    .Q(\po_0.regf_0.rf[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3316_ (.CLK(net103),
    .D(_0104_),
    .Q(\po_0.regf_0.rf[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3317_ (.CLK(net116),
    .D(_0105_),
    .Q(\po_0.regf_0.rf[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3318_ (.CLK(net116),
    .D(_0106_),
    .Q(\po_0.regf_0.rf[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3319_ (.CLK(net105),
    .D(_0107_),
    .Q(\po_0.regf_0.rf[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3320_ (.CLK(net129),
    .D(_0108_),
    .Q(\po_0.regf_0.rf[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3321_ (.CLK(net122),
    .D(_0109_),
    .Q(\po_0.regf_0.rf[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3322_ (.CLK(net122),
    .D(_0110_),
    .Q(\po_0.regf_0.rf[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3323_ (.CLK(net141),
    .D(_0111_),
    .Q(\po_0.regf_0.rf[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3324_ (.CLK(net136),
    .D(_0112_),
    .Q(\po_0.regf_0.rf[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3325_ (.CLK(net136),
    .D(_0113_),
    .Q(\po_0.regf_0.rf[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3326_ (.CLK(net130),
    .D(_0114_),
    .Q(\po_0.regf_0.rf[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3327_ (.CLK(net130),
    .D(_0115_),
    .Q(\po_0.regf_0.rf[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3328_ (.CLK(net137),
    .D(_0116_),
    .Q(\po_0.regf_0.rf[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3329_ (.CLK(net137),
    .D(_0117_),
    .Q(\po_0.regf_0.rf[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3330_ (.CLK(net112),
    .D(_0118_),
    .Q(\po_0.regf_0.rf[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3331_ (.CLK(net112),
    .D(_0119_),
    .Q(\po_0.regf_0.rf[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3332_ (.CLK(net103),
    .D(_0120_),
    .Q(\po_0.regf_0.rf[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3333_ (.CLK(net103),
    .D(_0121_),
    .Q(\po_0.regf_0.rf[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3334_ (.CLK(net103),
    .D(_0122_),
    .Q(\po_0.regf_0.rf[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3335_ (.CLK(net105),
    .D(_0123_),
    .Q(\po_0.regf_0.rf[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3336_ (.CLK(net129),
    .D(_0124_),
    .Q(\po_0.regf_0.rf[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3337_ (.CLK(net113),
    .D(_0125_),
    .Q(\po_0.regf_0.rf[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3338_ (.CLK(net113),
    .D(_0126_),
    .Q(\po_0.regf_0.rf[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3339_ (.CLK(net128),
    .D(_0127_),
    .Q(\po_0.regf_0.rf[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3340_ (.CLK(net138),
    .D(_0128_),
    .Q(\po_0.regf_0.rf[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3341_ (.CLK(net138),
    .D(_0129_),
    .Q(\po_0.regf_0.rf[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3342_ (.CLK(net131),
    .D(_0130_),
    .Q(\po_0.regf_0.rf[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3343_ (.CLK(net131),
    .D(_0131_),
    .Q(\po_0.regf_0.rf[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3344_ (.CLK(net137),
    .D(_0132_),
    .Q(\po_0.regf_0.rf[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3345_ (.CLK(net138),
    .D(_0133_),
    .Q(\po_0.regf_0.rf[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3346_ (.CLK(net112),
    .D(_0134_),
    .Q(\po_0.regf_0.rf[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3347_ (.CLK(net112),
    .D(_0135_),
    .Q(\po_0.regf_0.rf[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3348_ (.CLK(net104),
    .D(_0136_),
    .Q(\po_0.regf_0.rf[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3349_ (.CLK(net103),
    .D(_0137_),
    .Q(\po_0.regf_0.rf[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3350_ (.CLK(net106),
    .D(_0138_),
    .Q(\po_0.regf_0.rf[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3351_ (.CLK(net105),
    .D(_0139_),
    .Q(\po_0.regf_0.rf[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3352_ (.CLK(net128),
    .D(_0140_),
    .Q(\po_0.regf_0.rf[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3353_ (.CLK(net113),
    .D(_0141_),
    .Q(\po_0.regf_0.rf[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3354_ (.CLK(net128),
    .D(_0142_),
    .Q(\po_0.regf_0.rf[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3355_ (.CLK(net128),
    .D(_0143_),
    .Q(\po_0.regf_0.rf[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3356_ (.CLK(net144),
    .D(_0144_),
    .Q(\po_0.regf_0.rf[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3357_ (.CLK(net145),
    .D(_0145_),
    .Q(\po_0.regf_0.rf[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3358_ (.CLK(net131),
    .D(_0146_),
    .Q(\po_0.regf_0.rf[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3359_ (.CLK(net140),
    .D(_0147_),
    .Q(\po_0.regf_0.rf[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3360_ (.CLK(net145),
    .D(_0148_),
    .Q(\po_0.regf_0.rf[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3361_ (.CLK(net145),
    .D(_0149_),
    .Q(\po_0.regf_0.rf[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3362_ (.CLK(net122),
    .D(_0150_),
    .Q(\po_0.regf_0.rf[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3363_ (.CLK(net114),
    .D(_0151_),
    .Q(\po_0.regf_0.rf[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3364_ (.CLK(net104),
    .D(_0152_),
    .Q(\po_0.regf_0.rf[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3365_ (.CLK(net116),
    .D(_0153_),
    .Q(\po_0.regf_0.rf[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3366_ (.CLK(net116),
    .D(_0154_),
    .Q(\po_0.regf_0.rf[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3367_ (.CLK(net106),
    .D(_0155_),
    .Q(\po_0.regf_0.rf[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3368_ (.CLK(net129),
    .D(_0156_),
    .Q(\po_0.regf_0.rf[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3369_ (.CLK(net124),
    .D(_0157_),
    .Q(\po_0.regf_0.rf[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3370_ (.CLK(net140),
    .D(_0158_),
    .Q(\po_0.regf_0.rf[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3371_ (.CLK(net141),
    .D(_0159_),
    .Q(\po_0.regf_0.rf[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3372_ (.CLK(net173),
    .D(_0160_),
    .Q(\po_0.regf_0.rf[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3373_ (.CLK(net174),
    .D(_0161_),
    .Q(\po_0.regf_0.rf[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3374_ (.CLK(net173),
    .D(_0162_),
    .Q(\po_0.regf_0.rf[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3375_ (.CLK(net171),
    .D(_0163_),
    .Q(\po_0.regf_0.rf[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3376_ (.CLK(net148),
    .D(_0164_),
    .Q(\po_0.regf_0.rf[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3377_ (.CLK(net174),
    .D(_0165_),
    .Q(\po_0.regf_0.rf[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3378_ (.CLK(net152),
    .D(_0166_),
    .Q(\po_0.regf_0.rf[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3379_ (.CLK(net158),
    .D(_0167_),
    .Q(\po_0.regf_0.rf[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3380_ (.CLK(net119),
    .D(_0168_),
    .Q(\po_0.regf_0.rf[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3381_ (.CLK(net150),
    .D(_0169_),
    .Q(\po_0.regf_0.rf[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3382_ (.CLK(net150),
    .D(_0170_),
    .Q(\po_0.regf_0.rf[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3383_ (.CLK(net120),
    .D(_0171_),
    .Q(\po_0.regf_0.rf[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3384_ (.CLK(net170),
    .D(_0172_),
    .Q(\po_0.regf_0.rf[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3385_ (.CLK(net157),
    .D(_0173_),
    .Q(\po_0.regf_0.rf[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3386_ (.CLK(net157),
    .D(_0174_),
    .Q(\po_0.regf_0.rf[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3387_ (.CLK(net170),
    .D(_0175_),
    .Q(\po_0.regf_0.rf[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3388_ (.CLK(net173),
    .D(_0176_),
    .Q(\po_0.regf_0.rf[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3389_ (.CLK(net173),
    .D(_0177_),
    .Q(\po_0.regf_0.rf[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3390_ (.CLK(net171),
    .D(_0178_),
    .Q(\po_0.regf_0.rf[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3391_ (.CLK(net171),
    .D(_0179_),
    .Q(\po_0.regf_0.rf[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3392_ (.CLK(net148),
    .D(_0180_),
    .Q(\po_0.regf_0.rf[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3393_ (.CLK(net175),
    .D(_0181_),
    .Q(\po_0.regf_0.rf[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3394_ (.CLK(net152),
    .D(_0182_),
    .Q(\po_0.regf_0.rf[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3395_ (.CLK(net158),
    .D(_0183_),
    .Q(\po_0.regf_0.rf[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3396_ (.CLK(net119),
    .D(_0184_),
    .Q(\po_0.regf_0.rf[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3397_ (.CLK(net150),
    .D(_0185_),
    .Q(\po_0.regf_0.rf[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3398_ (.CLK(net150),
    .D(_0186_),
    .Q(\po_0.regf_0.rf[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3399_ (.CLK(net120),
    .D(_0187_),
    .Q(\po_0.regf_0.rf[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3400_ (.CLK(net170),
    .D(_0188_),
    .Q(\po_0.regf_0.rf[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3401_ (.CLK(net123),
    .D(_0189_),
    .Q(\po_0.regf_0.rf[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3402_ (.CLK(net157),
    .D(_0190_),
    .Q(\po_0.regf_0.rf[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3403_ (.CLK(net170),
    .D(_0191_),
    .Q(\po_0.regf_0.rf[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3404_ (.CLK(net136),
    .D(_0192_),
    .Q(\po_0.regf_0.rf[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3405_ (.CLK(net136),
    .D(_0193_),
    .Q(\po_0.regf_0.rf[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3406_ (.CLK(net130),
    .D(_0194_),
    .Q(\po_0.regf_0.rf[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3407_ (.CLK(net130),
    .D(_0195_),
    .Q(\po_0.regf_0.rf[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3408_ (.CLK(net137),
    .D(_0196_),
    .Q(\po_0.regf_0.rf[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3409_ (.CLK(net138),
    .D(_0197_),
    .Q(\po_0.regf_0.rf[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3410_ (.CLK(net114),
    .D(_0198_),
    .Q(\po_0.regf_0.rf[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3411_ (.CLK(net112),
    .D(_0199_),
    .Q(\po_0.regf_0.rf[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3412_ (.CLK(net104),
    .D(_0200_),
    .Q(\po_0.regf_0.rf[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3413_ (.CLK(net103),
    .D(_0201_),
    .Q(\po_0.regf_0.rf[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3414_ (.CLK(net105),
    .D(_0202_),
    .Q(\po_0.regf_0.rf[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3415_ (.CLK(net105),
    .D(_0203_),
    .Q(\po_0.regf_0.rf[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3416_ (.CLK(net141),
    .D(_0204_),
    .Q(\po_0.regf_0.rf[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3417_ (.CLK(net113),
    .D(_0205_),
    .Q(\po_0.regf_0.rf[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3418_ (.CLK(net128),
    .D(_0206_),
    .Q(\po_0.regf_0.rf[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3419_ (.CLK(net128),
    .D(_0207_),
    .Q(\po_0.regf_0.rf[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3420_ (.CLK(net176),
    .D(_0208_),
    .Q(\po_0.regf_0.rf[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3421_ (.CLK(net174),
    .D(_0209_),
    .Q(\po_0.regf_0.rf[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3422_ (.CLK(net176),
    .D(_0210_),
    .Q(\po_0.regf_0.rf[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3423_ (.CLK(net171),
    .D(_0211_),
    .Q(\po_0.regf_0.rf[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3424_ (.CLK(net174),
    .D(_0212_),
    .Q(\po_0.regf_0.rf[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3425_ (.CLK(net175),
    .D(_0213_),
    .Q(\po_0.regf_0.rf[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3426_ (.CLK(net156),
    .D(_0214_),
    .Q(\po_0.regf_0.rf[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3427_ (.CLK(net158),
    .D(_0215_),
    .Q(\po_0.regf_0.rf[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3428_ (.CLK(net150),
    .D(_0216_),
    .Q(\po_0.regf_0.rf[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3429_ (.CLK(net151),
    .D(_0217_),
    .Q(\po_0.regf_0.rf[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3430_ (.CLK(net151),
    .D(_0218_),
    .Q(\po_0.regf_0.rf[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3431_ (.CLK(net156),
    .D(_0219_),
    .Q(\po_0.regf_0.rf[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3432_ (.CLK(net172),
    .D(_0220_),
    .Q(\po_0.regf_0.rf[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3433_ (.CLK(net157),
    .D(_0221_),
    .Q(\po_0.regf_0.rf[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3434_ (.CLK(net161),
    .D(_0222_),
    .Q(\po_0.regf_0.rf[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3435_ (.CLK(net172),
    .D(_0223_),
    .Q(\po_0.regf_0.rf[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _3436_ (.CLK(net167),
    .D(_0224_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_2 _3437_ (.CLK(net167),
    .D(_0225_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_2 _3438_ (.CLK(net167),
    .D(_0226_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _3439_ (.CLK(net167),
    .D(_0227_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_2 _3440_ (.CLK(net167),
    .D(_0228_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_2 _3441_ (.CLK(net162),
    .D(_0229_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _3442_ (.CLK(net162),
    .D(_0230_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_2 _3443_ (.CLK(net163),
    .D(_0231_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _3444_ (.CLK(net164),
    .D(_0232_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _3445_ (.CLK(net164),
    .D(_0233_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_2 _3446_ (.CLK(net164),
    .D(_0234_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _3447_ (.CLK(net164),
    .D(_0235_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_4 _3448_ (.CLK(net163),
    .D(_0236_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _3449_ (.CLK(net165),
    .D(_0237_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_1 _3450_ (.CLK(net166),
    .D(_0238_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_2 _3451_ (.CLK(net166),
    .D(_0239_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _3452_ (.CLK(net166),
    .D(_0012_),
    .Q(_0004_));
 sky130_fd_sc_hd__dfxtp_1 _3453_ (.CLK(net153),
    .D(_0013_),
    .Q(_0005_));
 sky130_fd_sc_hd__dfxtp_1 _3454_ (.CLK(net153),
    .D(_0014_),
    .Q(_0006_));
 sky130_fd_sc_hd__dfxtp_1 _3455_ (.CLK(net153),
    .D(_0015_),
    .Q(_0007_));
 sky130_fd_sc_hd__dfxtp_1 _3456_ (.CLK(net177),
    .D(_0240_),
    .Q(\po_0.muxf_0.rf_w_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3457_ (.CLK(net177),
    .D(_0241_),
    .Q(\po_0.muxf_0.rf_w_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3458_ (.CLK(net178),
    .D(_0242_),
    .Q(\po_0.muxf_0.rf_w_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3459_ (.CLK(net167),
    .D(_0243_),
    .Q(\po_0.muxf_0.rf_w_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3460_ (.CLK(net177),
    .D(_0244_),
    .Q(\po_0.muxf_0.rf_w_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3461_ (.CLK(net162),
    .D(_0245_),
    .Q(\po_0.muxf_0.rf_w_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3462_ (.CLK(net162),
    .D(_0246_),
    .Q(\po_0.muxf_0.rf_w_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3463_ (.CLK(net162),
    .D(_0247_),
    .Q(\po_0.muxf_0.rf_w_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3464_ (.CLK(net159),
    .D(_0248_),
    .Q(\uc_0._20_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3465_ (.CLK(net160),
    .D(_0249_),
    .Q(\uc_0._20_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3466_ (.CLK(net155),
    .D(_0250_),
    .Q(\uc_0._20_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3467_ (.CLK(net155),
    .D(_0251_),
    .Q(\uc_0._20_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3468_ (.CLK(net164),
    .D(_0252_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_2 _3469_ (.CLK(net179),
    .D(_0253_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_2 _3470_ (.CLK(net151),
    .D(_0254_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_2 _3471_ (.CLK(net168),
    .D(_0255_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _3472_ (.CLK(net168),
    .D(_0256_),
    .Q(\uc_0._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _3473_ (.CLK(net136),
    .D(_0257_),
    .Q(\po_0.regf_0.rf[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3474_ (.CLK(net136),
    .D(_0258_),
    .Q(\po_0.regf_0.rf[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3475_ (.CLK(net130),
    .D(_0259_),
    .Q(\po_0.regf_0.rf[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3476_ (.CLK(net130),
    .D(_0260_),
    .Q(\po_0.regf_0.rf[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3477_ (.CLK(net137),
    .D(_0261_),
    .Q(\po_0.regf_0.rf[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3478_ (.CLK(net137),
    .D(_0262_),
    .Q(\po_0.regf_0.rf[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3479_ (.CLK(net111),
    .D(_0263_),
    .Q(\po_0.regf_0.rf[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3480_ (.CLK(net110),
    .D(_0264_),
    .Q(\po_0.regf_0.rf[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3481_ (.CLK(net101),
    .D(_0265_),
    .Q(\po_0.regf_0.rf[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3482_ (.CLK(net105),
    .D(_0266_),
    .Q(\po_0.regf_0.rf[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3483_ (.CLK(net101),
    .D(_0267_),
    .Q(\po_0.regf_0.rf[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3484_ (.CLK(net101),
    .D(_0268_),
    .Q(\po_0.regf_0.rf[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3485_ (.CLK(net110),
    .D(_0269_),
    .Q(\po_0.regf_0.rf[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3486_ (.CLK(net113),
    .D(_0270_),
    .Q(\po_0.regf_0.rf[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3487_ (.CLK(net126),
    .D(_0271_),
    .Q(\po_0.regf_0.rf[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3488_ (.CLK(net127),
    .D(_0272_),
    .Q(\po_0.regf_0.rf[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3489_ (.CLK(net147),
    .D(_0273_),
    .Q(\po_0.regf_0.rf[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3490_ (.CLK(net147),
    .D(_0274_),
    .Q(\po_0.regf_0.rf[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3491_ (.CLK(net142),
    .D(_0275_),
    .Q(\po_0.regf_0.rf[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3492_ (.CLK(net142),
    .D(_0276_),
    .Q(\po_0.regf_0.rf[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3493_ (.CLK(net146),
    .D(_0277_),
    .Q(\po_0.regf_0.rf[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3494_ (.CLK(net146),
    .D(_0278_),
    .Q(\po_0.regf_0.rf[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3495_ (.CLK(net118),
    .D(_0279_),
    .Q(\po_0.regf_0.rf[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3496_ (.CLK(net123),
    .D(_0280_),
    .Q(\po_0.regf_0.rf[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3497_ (.CLK(net119),
    .D(_0281_),
    .Q(\po_0.regf_0.rf[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3498_ (.CLK(net117),
    .D(_0282_),
    .Q(\po_0.regf_0.rf[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3499_ (.CLK(net118),
    .D(_0283_),
    .Q(\po_0.regf_0.rf[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3500_ (.CLK(net120),
    .D(_0284_),
    .Q(\po_0.regf_0.rf[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3501_ (.CLK(net123),
    .D(_0285_),
    .Q(\po_0.regf_0.rf[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3502_ (.CLK(net124),
    .D(_0286_),
    .Q(\po_0.regf_0.rf[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3503_ (.CLK(net114),
    .D(_0287_),
    .Q(\po_0.regf_0.rf[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3504_ (.CLK(net140),
    .D(_0288_),
    .Q(\po_0.regf_0.rf[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3505_ (.CLK(net147),
    .D(_0289_),
    .Q(\po_0.regf_0.rf[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3506_ (.CLK(net144),
    .D(_0290_),
    .Q(\po_0.regf_0.rf[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3507_ (.CLK(net143),
    .D(_0291_),
    .Q(\po_0.regf_0.rf[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3508_ (.CLK(net142),
    .D(_0292_),
    .Q(\po_0.regf_0.rf[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3509_ (.CLK(net147),
    .D(_0293_),
    .Q(\po_0.regf_0.rf[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3510_ (.CLK(net146),
    .D(_0294_),
    .Q(\po_0.regf_0.rf[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3511_ (.CLK(net122),
    .D(_0295_),
    .Q(\po_0.regf_0.rf[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3512_ (.CLK(net123),
    .D(_0296_),
    .Q(\po_0.regf_0.rf[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3513_ (.CLK(net119),
    .D(_0297_),
    .Q(\po_0.regf_0.rf[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3514_ (.CLK(net117),
    .D(_0298_),
    .Q(\po_0.regf_0.rf[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3515_ (.CLK(net116),
    .D(_0299_),
    .Q(\po_0.regf_0.rf[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3516_ (.CLK(net120),
    .D(_0300_),
    .Q(\po_0.regf_0.rf[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3517_ (.CLK(net124),
    .D(_0301_),
    .Q(\po_0.regf_0.rf[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3518_ (.CLK(net124),
    .D(_0302_),
    .Q(\po_0.regf_0.rf[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3519_ (.CLK(net114),
    .D(_0303_),
    .Q(\po_0.regf_0.rf[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3520_ (.CLK(net140),
    .D(_0304_),
    .Q(\po_0.regf_0.rf[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3521_ (.CLK(net179),
    .D(_0305_),
    .Q(\po_0.alu_0.s1 ));
 sky130_fd_sc_hd__dfxtp_1 _3522_ (.CLK(net180),
    .D(_0306_),
    .Q(\po_0.alu_0.s0 ));
 sky130_fd_sc_hd__dfxtp_1 _3523_ (.CLK(net166),
    .D(_0307_),
    .Q(\po_0.regf_0.rq_rd ));
 sky130_fd_sc_hd__dfxtp_1 _3524_ (.CLK(net160),
    .D(_0308_),
    .Q(\po_0.regf_0.rp_rd ));
 sky130_fd_sc_hd__dfxtp_1 _3525_ (.CLK(net159),
    .D(_0309_),
    .Q(\po_0.regf_0.w_wr ));
 sky130_fd_sc_hd__dfxtp_1 _3526_ (.CLK(net166),
    .D(_0310_),
    .Q(\po_0.regf_0.rq_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3527_ (.CLK(net162),
    .D(_0311_),
    .Q(\po_0.regf_0.rq_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3528_ (.CLK(net154),
    .D(_0312_),
    .Q(\po_0.regf_0.rq_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3529_ (.CLK(net154),
    .D(_0313_),
    .Q(\po_0.regf_0.rq_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3530_ (.CLK(net160),
    .D(_0314_),
    .Q(\po_0.regf_0.rp_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3531_ (.CLK(net160),
    .D(_0315_),
    .Q(\po_0.regf_0.rp_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3532_ (.CLK(net154),
    .D(_0316_),
    .Q(\po_0.regf_0.rp_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3533_ (.CLK(net153),
    .D(_0317_),
    .Q(\po_0.regf_0.rp_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3534_ (.CLK(net159),
    .D(_0318_),
    .Q(\po_0.regf_0.w_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3535_ (.CLK(net159),
    .D(_0319_),
    .Q(\po_0.regf_0.w_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3536_ (.CLK(net158),
    .D(_0320_),
    .Q(\po_0.regf_0.w_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3537_ (.CLK(net159),
    .D(_0321_),
    .Q(\po_0.regf_0.w_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3538_ (.CLK(net180),
    .D(_0322_),
    .Q(\po_0.muxf_0.s0 ));
 sky130_fd_sc_hd__dfxtp_1 _3539_ (.CLK(net180),
    .D(_0323_),
    .Q(\po_0.muxf_0.s1 ));
 sky130_fd_sc_hd__dfxtp_1 _3540_ (.CLK(net179),
    .D(_0324_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _3541_ (.CLK(net180),
    .D(_0325_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_2 _3542_ (.CLK(net166),
    .D(_0326_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _3543_ (.CLK(net178),
    .D(_0327_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _3544_ (.CLK(net108),
    .D(_0328_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _3545_ (.CLK(net126),
    .D(_0329_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _3546_ (.CLK(net180),
    .D(_0330_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _3547_ (.CLK(net168),
    .D(_0331_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _3548_ (.CLK(net153),
    .D(_0332_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _3549_ (.CLK(net100),
    .D(_0333_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _3550_ (.CLK(net178),
    .D(_0334_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _3551_ (.CLK(net178),
    .D(_0335_),
    .Q(\uc_0._03_ ));
 sky130_fd_sc_hd__dfxtp_1 _3552_ (.CLK(net177),
    .D(_0336_),
    .Q(\uc_0._02_ ));
 sky130_fd_sc_hd__dfxtp_1 _3553_ (.CLK(net177),
    .D(_0337_),
    .Q(\uc_0._01_ ));
 sky130_fd_sc_hd__dfxtp_1 _3554_ (.CLK(net179),
    .D(\uc_0.bc_0._54_[0] ),
    .Q(\uc_0.bc_0._55_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3555_ (.CLK(net177),
    .D(\uc_0.bc_0._54_[1] ),
    .Q(\uc_0.bc_0._55_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3556_ (.CLK(net181),
    .D(\uc_0.bc_0._54_[2] ),
    .Q(\uc_0.bc_0._55_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3557_ (.CLK(net181),
    .D(\uc_0.bc_0._54_[3] ),
    .Q(\uc_0.bc_0._55_[3] ));
 sky130_fd_sc_hd__clkbuf_1 _3558_ (.A(net164),
    .X(net78));
 sky130_fd_sc_hd__ebufn_1 _3559_ (.A(\po_0.alu_0._10_[0] ),
    .TE_B(_1558_),
    .Z(\po_0.alu_0._11_[0] ));
 sky130_fd_sc_hd__ebufn_1 _3560_ (.A(\po_0.alu_0._10_[1] ),
    .TE_B(_1559_),
    .Z(\po_0.alu_0._11_[1] ));
 sky130_fd_sc_hd__ebufn_1 _3561_ (.A(\po_0.alu_0._10_[2] ),
    .TE_B(_1560_),
    .Z(\po_0.alu_0._11_[2] ));
 sky130_fd_sc_hd__ebufn_1 _3562_ (.A(\po_0.alu_0._10_[3] ),
    .TE_B(_1561_),
    .Z(\po_0.alu_0._11_[3] ));
 sky130_fd_sc_hd__ebufn_1 _3563_ (.A(\po_0.alu_0._10_[4] ),
    .TE_B(_1562_),
    .Z(\po_0.alu_0._11_[4] ));
 sky130_fd_sc_hd__ebufn_1 _3564_ (.A(\po_0.alu_0._10_[5] ),
    .TE_B(_1563_),
    .Z(\po_0.alu_0._11_[5] ));
 sky130_fd_sc_hd__ebufn_1 _3565_ (.A(\po_0.alu_0._10_[6] ),
    .TE_B(_1564_),
    .Z(\po_0.alu_0._11_[6] ));
 sky130_fd_sc_hd__ebufn_1 _3566_ (.A(\po_0.alu_0._10_[7] ),
    .TE_B(_1565_),
    .Z(\po_0.alu_0._11_[7] ));
 sky130_fd_sc_hd__ebufn_1 _3567_ (.A(\po_0.alu_0._10_[8] ),
    .TE_B(_1566_),
    .Z(\po_0.alu_0._11_[8] ));
 sky130_fd_sc_hd__ebufn_1 _3568_ (.A(\po_0.alu_0._10_[9] ),
    .TE_B(_1567_),
    .Z(\po_0.alu_0._11_[9] ));
 sky130_fd_sc_hd__ebufn_1 _3569_ (.A(\po_0.alu_0._10_[10] ),
    .TE_B(_1568_),
    .Z(\po_0.alu_0._11_[10] ));
 sky130_fd_sc_hd__ebufn_1 _3570_ (.A(\po_0.alu_0._10_[11] ),
    .TE_B(_1569_),
    .Z(\po_0.alu_0._11_[11] ));
 sky130_fd_sc_hd__ebufn_1 _3571_ (.A(\po_0.alu_0._10_[12] ),
    .TE_B(_1570_),
    .Z(\po_0.alu_0._11_[12] ));
 sky130_fd_sc_hd__ebufn_1 _3572_ (.A(\po_0.alu_0._10_[13] ),
    .TE_B(_1571_),
    .Z(\po_0.alu_0._11_[13] ));
 sky130_fd_sc_hd__ebufn_1 _3573_ (.A(\po_0.alu_0._10_[14] ),
    .TE_B(_1572_),
    .Z(\po_0.alu_0._11_[14] ));
 sky130_fd_sc_hd__ebufn_1 _3574_ (.A(\po_0.alu_0._10_[15] ),
    .TE_B(_1573_),
    .Z(\po_0.alu_0._11_[15] ));
 sky130_fd_sc_hd__clkbuf_2 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout101 (.A(net107),
    .X(net101));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout102 (.A(net107),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 fanout103 (.A(net106),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 fanout104 (.A(net106),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 fanout107 (.A(net115),
    .X(net107));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout108 (.A(net111),
    .X(net108));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout109 (.A(net111),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 fanout111 (.A(net115),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 fanout112 (.A(net114),
    .X(net112));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout115 (.A(net125),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 fanout116 (.A(net118),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 fanout118 (.A(net121),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout119 (.A(net121),
    .X(net119));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 fanout121 (.A(net125),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 fanout122 (.A(net124),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(net183),
    .X(net125));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout127 (.A(net133),
    .X(net127));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout128 (.A(net132),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 fanout129 (.A(net132),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 fanout130 (.A(net132),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 fanout133 (.A(net149),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 fanout134 (.A(net139),
    .X(net134));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout135 (.A(net139),
    .X(net135));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout136 (.A(net138),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 fanout139 (.A(net149),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 fanout140 (.A(net143),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 fanout141 (.A(net143),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout143 (.A(net149),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 fanout144 (.A(net148),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 fanout145 (.A(net148),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 fanout149 (.A(net183),
    .X(net149));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout150 (.A(net152),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 fanout151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout152 (.A(net156),
    .X(net152));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout153 (.A(net155),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout156 (.A(net169),
    .X(net156));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 fanout158 (.A(net161),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 fanout161 (.A(net169),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 fanout163 (.A(net165),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 fanout165 (.A(net169),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 fanout166 (.A(net168),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 fanout169 (.A(net183),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 fanout170 (.A(net172),
    .X(net170));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout172 (.A(net182),
    .X(net172));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout173 (.A(net176),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout176 (.A(net182),
    .X(net176));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout177 (.A(net179),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__buf_2 fanout183 (.A(net33),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(net38),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 fanout84 (.A(net37),
    .X(net84));
 sky130_fd_sc_hd__buf_2 fanout85 (.A(net48),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 fanout86 (.A(net42),
    .X(net86));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout87 (.A(net35),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 fanout88 (.A(net91),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 fanout89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(\po_0.regf_0.rp_rd ),
    .X(net91));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 fanout93 (.A(net95),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 fanout95 (.A(\po_0.regf_0.rq_rd ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(net66),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 fanout97 (.A(net75),
    .X(net97));
 sky130_fd_sc_hd__buf_2 fanout98 (.A(net73),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 fanout99 (.A(net70),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(D_R_data[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(D_R_data[3]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(D_R_data[4]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(D_R_data[5]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(D_R_data[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(D_R_data[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(D_R_data[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(D_R_data[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(I_data[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(I_data[10]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(I_data[11]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(D_R_data[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(I_data[12]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(I_data[13]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(I_data[14]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(I_data[15]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(I_data[1]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(I_data[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(I_data[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(I_data[4]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(I_data[5]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(I_data[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(D_R_data[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(I_data[7]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(I_data[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(I_data[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(clock),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(reset),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(D_R_data[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(D_R_data[13]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(D_R_data[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(D_R_data[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(D_R_data[1]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(D_R_data[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(D_W_data[0]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(D_W_data[10]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(D_W_data[11]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net83),
    .X(D_W_data[12]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(D_W_data[13]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(D_W_data[14]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(D_W_data[15]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(D_W_data[1]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(D_W_data[2]));
 sky130_fd_sc_hd__clkbuf_4 output44 (.A(net44),
    .X(D_W_data[3]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(D_W_data[4]));
 sky130_fd_sc_hd__clkbuf_4 output46 (.A(net46),
    .X(D_W_data[5]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(D_W_data[6]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net85),
    .X(D_W_data[7]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(D_W_data[8]));
 sky130_fd_sc_hd__clkbuf_4 output50 (.A(net50),
    .X(D_W_data[9]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(D_addr[0]));
 sky130_fd_sc_hd__clkbuf_4 output52 (.A(net52),
    .X(D_addr[1]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(D_addr[2]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(D_addr[3]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(D_addr[4]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(D_addr[5]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(D_addr[6]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(D_addr[7]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(D_rd));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(D_wr));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(I_addr[0]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(I_addr[10]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(I_addr[11]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(I_addr[12]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(I_addr[13]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net96),
    .X(I_addr[14]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(I_addr[15]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(I_addr[1]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(I_addr[2]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net99),
    .X(I_addr[3]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(I_addr[4]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(I_addr[5]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net98),
    .X(I_addr[6]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(I_addr[7]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(I_addr[8]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(I_addr[9]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(I_rd));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net78),
    .X(led_clock));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(leds[0]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(leds[1]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(leds[2]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(leds[3]));
endmodule

