magic
tech sky130A
timestamp 0
<< properties >>
string FIXED_BBOX 0 0 0 0
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5931692
string GDS_FILE /openlane/designs/vahid6i/runs/RUN_2023.03.28_22.13.51/results/signoff/vahid6i.magic.gds
string GDS_START 804134
<< end >>

