// This is the unpowered netlist.
module vahid6i (D_rd,
    D_wr,
    I_rd,
    clock,
    led_clock,
    reset,
    D_R_data,
    D_W_data,
    D_addr,
    I_addr,
    I_data,
    leds);
 output D_rd;
 output D_wr;
 output I_rd;
 input clock;
 output led_clock;
 input reset;
 input [15:0] D_R_data;
 output [15:0] D_W_data;
 output [7:0] D_addr;
 output [15:0] I_addr;
 input [15:0] I_data;
 output [3:0] leds;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \po_0._1_[0] ;
 wire \po_0._1_[10] ;
 wire \po_0._1_[11] ;
 wire \po_0._1_[12] ;
 wire \po_0._1_[13] ;
 wire \po_0._1_[14] ;
 wire \po_0._1_[15] ;
 wire \po_0._1_[1] ;
 wire \po_0._1_[2] ;
 wire \po_0._1_[3] ;
 wire \po_0._1_[4] ;
 wire \po_0._1_[5] ;
 wire \po_0._1_[6] ;
 wire \po_0._1_[7] ;
 wire \po_0._1_[8] ;
 wire \po_0._1_[9] ;
 wire \po_0.alu_0._10_[0] ;
 wire \po_0.alu_0._10_[10] ;
 wire \po_0.alu_0._10_[11] ;
 wire \po_0.alu_0._10_[12] ;
 wire \po_0.alu_0._10_[13] ;
 wire \po_0.alu_0._10_[14] ;
 wire \po_0.alu_0._10_[15] ;
 wire \po_0.alu_0._10_[1] ;
 wire \po_0.alu_0._10_[2] ;
 wire \po_0.alu_0._10_[3] ;
 wire \po_0.alu_0._10_[4] ;
 wire \po_0.alu_0._10_[5] ;
 wire \po_0.alu_0._10_[6] ;
 wire \po_0.alu_0._10_[7] ;
 wire \po_0.alu_0._10_[8] ;
 wire \po_0.alu_0._10_[9] ;
 wire \po_0.alu_0._11_[0] ;
 wire \po_0.alu_0._11_[10] ;
 wire \po_0.alu_0._11_[11] ;
 wire \po_0.alu_0._11_[12] ;
 wire \po_0.alu_0._11_[13] ;
 wire \po_0.alu_0._11_[14] ;
 wire \po_0.alu_0._11_[15] ;
 wire \po_0.alu_0._11_[1] ;
 wire \po_0.alu_0._11_[2] ;
 wire \po_0.alu_0._11_[3] ;
 wire \po_0.alu_0._11_[4] ;
 wire \po_0.alu_0._11_[5] ;
 wire \po_0.alu_0._11_[6] ;
 wire \po_0.alu_0._11_[7] ;
 wire \po_0.alu_0._11_[8] ;
 wire \po_0.alu_0._11_[9] ;
 wire \po_0.alu_0.s0 ;
 wire \po_0.alu_0.s1 ;
 wire \po_0.muxf_0.rf_w_data[0] ;
 wire \po_0.muxf_0.rf_w_data[1] ;
 wire \po_0.muxf_0.rf_w_data[2] ;
 wire \po_0.muxf_0.rf_w_data[3] ;
 wire \po_0.muxf_0.rf_w_data[4] ;
 wire \po_0.muxf_0.rf_w_data[5] ;
 wire \po_0.muxf_0.rf_w_data[6] ;
 wire \po_0.muxf_0.rf_w_data[7] ;
 wire \po_0.muxf_0.s0 ;
 wire \po_0.muxf_0.s1 ;
 wire \po_0.regf_0._3_[0] ;
 wire \po_0.regf_0._3_[10] ;
 wire \po_0.regf_0._3_[11] ;
 wire \po_0.regf_0._3_[12] ;
 wire \po_0.regf_0._3_[13] ;
 wire \po_0.regf_0._3_[14] ;
 wire \po_0.regf_0._3_[15] ;
 wire \po_0.regf_0._3_[1] ;
 wire \po_0.regf_0._3_[2] ;
 wire \po_0.regf_0._3_[3] ;
 wire \po_0.regf_0._3_[4] ;
 wire \po_0.regf_0._3_[5] ;
 wire \po_0.regf_0._3_[6] ;
 wire \po_0.regf_0._3_[7] ;
 wire \po_0.regf_0._3_[8] ;
 wire \po_0.regf_0._3_[9] ;
 wire \po_0.regf_0._5_[0] ;
 wire \po_0.regf_0._5_[10] ;
 wire \po_0.regf_0._5_[11] ;
 wire \po_0.regf_0._5_[12] ;
 wire \po_0.regf_0._5_[13] ;
 wire \po_0.regf_0._5_[14] ;
 wire \po_0.regf_0._5_[15] ;
 wire \po_0.regf_0._5_[1] ;
 wire \po_0.regf_0._5_[2] ;
 wire \po_0.regf_0._5_[3] ;
 wire \po_0.regf_0._5_[4] ;
 wire \po_0.regf_0._5_[5] ;
 wire \po_0.regf_0._5_[6] ;
 wire \po_0.regf_0._5_[7] ;
 wire \po_0.regf_0._5_[8] ;
 wire \po_0.regf_0._5_[9] ;
 wire \po_0.regf_0.rf[0][0] ;
 wire \po_0.regf_0.rf[0][10] ;
 wire \po_0.regf_0.rf[0][11] ;
 wire \po_0.regf_0.rf[0][12] ;
 wire \po_0.regf_0.rf[0][13] ;
 wire \po_0.regf_0.rf[0][14] ;
 wire \po_0.regf_0.rf[0][15] ;
 wire \po_0.regf_0.rf[0][1] ;
 wire \po_0.regf_0.rf[0][2] ;
 wire \po_0.regf_0.rf[0][3] ;
 wire \po_0.regf_0.rf[0][4] ;
 wire \po_0.regf_0.rf[0][5] ;
 wire \po_0.regf_0.rf[0][6] ;
 wire \po_0.regf_0.rf[0][7] ;
 wire \po_0.regf_0.rf[0][8] ;
 wire \po_0.regf_0.rf[0][9] ;
 wire \po_0.regf_0.rf[10][0] ;
 wire \po_0.regf_0.rf[10][10] ;
 wire \po_0.regf_0.rf[10][11] ;
 wire \po_0.regf_0.rf[10][12] ;
 wire \po_0.regf_0.rf[10][13] ;
 wire \po_0.regf_0.rf[10][14] ;
 wire \po_0.regf_0.rf[10][15] ;
 wire \po_0.regf_0.rf[10][1] ;
 wire \po_0.regf_0.rf[10][2] ;
 wire \po_0.regf_0.rf[10][3] ;
 wire \po_0.regf_0.rf[10][4] ;
 wire \po_0.regf_0.rf[10][5] ;
 wire \po_0.regf_0.rf[10][6] ;
 wire \po_0.regf_0.rf[10][7] ;
 wire \po_0.regf_0.rf[10][8] ;
 wire \po_0.regf_0.rf[10][9] ;
 wire \po_0.regf_0.rf[11][0] ;
 wire \po_0.regf_0.rf[11][10] ;
 wire \po_0.regf_0.rf[11][11] ;
 wire \po_0.regf_0.rf[11][12] ;
 wire \po_0.regf_0.rf[11][13] ;
 wire \po_0.regf_0.rf[11][14] ;
 wire \po_0.regf_0.rf[11][15] ;
 wire \po_0.regf_0.rf[11][1] ;
 wire \po_0.regf_0.rf[11][2] ;
 wire \po_0.regf_0.rf[11][3] ;
 wire \po_0.regf_0.rf[11][4] ;
 wire \po_0.regf_0.rf[11][5] ;
 wire \po_0.regf_0.rf[11][6] ;
 wire \po_0.regf_0.rf[11][7] ;
 wire \po_0.regf_0.rf[11][8] ;
 wire \po_0.regf_0.rf[11][9] ;
 wire \po_0.regf_0.rf[12][0] ;
 wire \po_0.regf_0.rf[12][10] ;
 wire \po_0.regf_0.rf[12][11] ;
 wire \po_0.regf_0.rf[12][12] ;
 wire \po_0.regf_0.rf[12][13] ;
 wire \po_0.regf_0.rf[12][14] ;
 wire \po_0.regf_0.rf[12][15] ;
 wire \po_0.regf_0.rf[12][1] ;
 wire \po_0.regf_0.rf[12][2] ;
 wire \po_0.regf_0.rf[12][3] ;
 wire \po_0.regf_0.rf[12][4] ;
 wire \po_0.regf_0.rf[12][5] ;
 wire \po_0.regf_0.rf[12][6] ;
 wire \po_0.regf_0.rf[12][7] ;
 wire \po_0.regf_0.rf[12][8] ;
 wire \po_0.regf_0.rf[12][9] ;
 wire \po_0.regf_0.rf[13][0] ;
 wire \po_0.regf_0.rf[13][10] ;
 wire \po_0.regf_0.rf[13][11] ;
 wire \po_0.regf_0.rf[13][12] ;
 wire \po_0.regf_0.rf[13][13] ;
 wire \po_0.regf_0.rf[13][14] ;
 wire \po_0.regf_0.rf[13][15] ;
 wire \po_0.regf_0.rf[13][1] ;
 wire \po_0.regf_0.rf[13][2] ;
 wire \po_0.regf_0.rf[13][3] ;
 wire \po_0.regf_0.rf[13][4] ;
 wire \po_0.regf_0.rf[13][5] ;
 wire \po_0.regf_0.rf[13][6] ;
 wire \po_0.regf_0.rf[13][7] ;
 wire \po_0.regf_0.rf[13][8] ;
 wire \po_0.regf_0.rf[13][9] ;
 wire \po_0.regf_0.rf[14][0] ;
 wire \po_0.regf_0.rf[14][10] ;
 wire \po_0.regf_0.rf[14][11] ;
 wire \po_0.regf_0.rf[14][12] ;
 wire \po_0.regf_0.rf[14][13] ;
 wire \po_0.regf_0.rf[14][14] ;
 wire \po_0.regf_0.rf[14][15] ;
 wire \po_0.regf_0.rf[14][1] ;
 wire \po_0.regf_0.rf[14][2] ;
 wire \po_0.regf_0.rf[14][3] ;
 wire \po_0.regf_0.rf[14][4] ;
 wire \po_0.regf_0.rf[14][5] ;
 wire \po_0.regf_0.rf[14][6] ;
 wire \po_0.regf_0.rf[14][7] ;
 wire \po_0.regf_0.rf[14][8] ;
 wire \po_0.regf_0.rf[14][9] ;
 wire \po_0.regf_0.rf[15][0] ;
 wire \po_0.regf_0.rf[15][10] ;
 wire \po_0.regf_0.rf[15][11] ;
 wire \po_0.regf_0.rf[15][12] ;
 wire \po_0.regf_0.rf[15][13] ;
 wire \po_0.regf_0.rf[15][14] ;
 wire \po_0.regf_0.rf[15][15] ;
 wire \po_0.regf_0.rf[15][1] ;
 wire \po_0.regf_0.rf[15][2] ;
 wire \po_0.regf_0.rf[15][3] ;
 wire \po_0.regf_0.rf[15][4] ;
 wire \po_0.regf_0.rf[15][5] ;
 wire \po_0.regf_0.rf[15][6] ;
 wire \po_0.regf_0.rf[15][7] ;
 wire \po_0.regf_0.rf[15][8] ;
 wire \po_0.regf_0.rf[15][9] ;
 wire \po_0.regf_0.rf[1][0] ;
 wire \po_0.regf_0.rf[1][10] ;
 wire \po_0.regf_0.rf[1][11] ;
 wire \po_0.regf_0.rf[1][12] ;
 wire \po_0.regf_0.rf[1][13] ;
 wire \po_0.regf_0.rf[1][14] ;
 wire \po_0.regf_0.rf[1][15] ;
 wire \po_0.regf_0.rf[1][1] ;
 wire \po_0.regf_0.rf[1][2] ;
 wire \po_0.regf_0.rf[1][3] ;
 wire \po_0.regf_0.rf[1][4] ;
 wire \po_0.regf_0.rf[1][5] ;
 wire \po_0.regf_0.rf[1][6] ;
 wire \po_0.regf_0.rf[1][7] ;
 wire \po_0.regf_0.rf[1][8] ;
 wire \po_0.regf_0.rf[1][9] ;
 wire \po_0.regf_0.rf[2][0] ;
 wire \po_0.regf_0.rf[2][10] ;
 wire \po_0.regf_0.rf[2][11] ;
 wire \po_0.regf_0.rf[2][12] ;
 wire \po_0.regf_0.rf[2][13] ;
 wire \po_0.regf_0.rf[2][14] ;
 wire \po_0.regf_0.rf[2][15] ;
 wire \po_0.regf_0.rf[2][1] ;
 wire \po_0.regf_0.rf[2][2] ;
 wire \po_0.regf_0.rf[2][3] ;
 wire \po_0.regf_0.rf[2][4] ;
 wire \po_0.regf_0.rf[2][5] ;
 wire \po_0.regf_0.rf[2][6] ;
 wire \po_0.regf_0.rf[2][7] ;
 wire \po_0.regf_0.rf[2][8] ;
 wire \po_0.regf_0.rf[2][9] ;
 wire \po_0.regf_0.rf[3][0] ;
 wire \po_0.regf_0.rf[3][10] ;
 wire \po_0.regf_0.rf[3][11] ;
 wire \po_0.regf_0.rf[3][12] ;
 wire \po_0.regf_0.rf[3][13] ;
 wire \po_0.regf_0.rf[3][14] ;
 wire \po_0.regf_0.rf[3][15] ;
 wire \po_0.regf_0.rf[3][1] ;
 wire \po_0.regf_0.rf[3][2] ;
 wire \po_0.regf_0.rf[3][3] ;
 wire \po_0.regf_0.rf[3][4] ;
 wire \po_0.regf_0.rf[3][5] ;
 wire \po_0.regf_0.rf[3][6] ;
 wire \po_0.regf_0.rf[3][7] ;
 wire \po_0.regf_0.rf[3][8] ;
 wire \po_0.regf_0.rf[3][9] ;
 wire \po_0.regf_0.rf[4][0] ;
 wire \po_0.regf_0.rf[4][10] ;
 wire \po_0.regf_0.rf[4][11] ;
 wire \po_0.regf_0.rf[4][12] ;
 wire \po_0.regf_0.rf[4][13] ;
 wire \po_0.regf_0.rf[4][14] ;
 wire \po_0.regf_0.rf[4][15] ;
 wire \po_0.regf_0.rf[4][1] ;
 wire \po_0.regf_0.rf[4][2] ;
 wire \po_0.regf_0.rf[4][3] ;
 wire \po_0.regf_0.rf[4][4] ;
 wire \po_0.regf_0.rf[4][5] ;
 wire \po_0.regf_0.rf[4][6] ;
 wire \po_0.regf_0.rf[4][7] ;
 wire \po_0.regf_0.rf[4][8] ;
 wire \po_0.regf_0.rf[4][9] ;
 wire \po_0.regf_0.rf[5][0] ;
 wire \po_0.regf_0.rf[5][10] ;
 wire \po_0.regf_0.rf[5][11] ;
 wire \po_0.regf_0.rf[5][12] ;
 wire \po_0.regf_0.rf[5][13] ;
 wire \po_0.regf_0.rf[5][14] ;
 wire \po_0.regf_0.rf[5][15] ;
 wire \po_0.regf_0.rf[5][1] ;
 wire \po_0.regf_0.rf[5][2] ;
 wire \po_0.regf_0.rf[5][3] ;
 wire \po_0.regf_0.rf[5][4] ;
 wire \po_0.regf_0.rf[5][5] ;
 wire \po_0.regf_0.rf[5][6] ;
 wire \po_0.regf_0.rf[5][7] ;
 wire \po_0.regf_0.rf[5][8] ;
 wire \po_0.regf_0.rf[5][9] ;
 wire \po_0.regf_0.rf[6][0] ;
 wire \po_0.regf_0.rf[6][10] ;
 wire \po_0.regf_0.rf[6][11] ;
 wire \po_0.regf_0.rf[6][12] ;
 wire \po_0.regf_0.rf[6][13] ;
 wire \po_0.regf_0.rf[6][14] ;
 wire \po_0.regf_0.rf[6][15] ;
 wire \po_0.regf_0.rf[6][1] ;
 wire \po_0.regf_0.rf[6][2] ;
 wire \po_0.regf_0.rf[6][3] ;
 wire \po_0.regf_0.rf[6][4] ;
 wire \po_0.regf_0.rf[6][5] ;
 wire \po_0.regf_0.rf[6][6] ;
 wire \po_0.regf_0.rf[6][7] ;
 wire \po_0.regf_0.rf[6][8] ;
 wire \po_0.regf_0.rf[6][9] ;
 wire \po_0.regf_0.rf[7][0] ;
 wire \po_0.regf_0.rf[7][10] ;
 wire \po_0.regf_0.rf[7][11] ;
 wire \po_0.regf_0.rf[7][12] ;
 wire \po_0.regf_0.rf[7][13] ;
 wire \po_0.regf_0.rf[7][14] ;
 wire \po_0.regf_0.rf[7][15] ;
 wire \po_0.regf_0.rf[7][1] ;
 wire \po_0.regf_0.rf[7][2] ;
 wire \po_0.regf_0.rf[7][3] ;
 wire \po_0.regf_0.rf[7][4] ;
 wire \po_0.regf_0.rf[7][5] ;
 wire \po_0.regf_0.rf[7][6] ;
 wire \po_0.regf_0.rf[7][7] ;
 wire \po_0.regf_0.rf[7][8] ;
 wire \po_0.regf_0.rf[7][9] ;
 wire \po_0.regf_0.rf[8][0] ;
 wire \po_0.regf_0.rf[8][10] ;
 wire \po_0.regf_0.rf[8][11] ;
 wire \po_0.regf_0.rf[8][12] ;
 wire \po_0.regf_0.rf[8][13] ;
 wire \po_0.regf_0.rf[8][14] ;
 wire \po_0.regf_0.rf[8][15] ;
 wire \po_0.regf_0.rf[8][1] ;
 wire \po_0.regf_0.rf[8][2] ;
 wire \po_0.regf_0.rf[8][3] ;
 wire \po_0.regf_0.rf[8][4] ;
 wire \po_0.regf_0.rf[8][5] ;
 wire \po_0.regf_0.rf[8][6] ;
 wire \po_0.regf_0.rf[8][7] ;
 wire \po_0.regf_0.rf[8][8] ;
 wire \po_0.regf_0.rf[8][9] ;
 wire \po_0.regf_0.rf[9][0] ;
 wire \po_0.regf_0.rf[9][10] ;
 wire \po_0.regf_0.rf[9][11] ;
 wire \po_0.regf_0.rf[9][12] ;
 wire \po_0.regf_0.rf[9][13] ;
 wire \po_0.regf_0.rf[9][14] ;
 wire \po_0.regf_0.rf[9][15] ;
 wire \po_0.regf_0.rf[9][1] ;
 wire \po_0.regf_0.rf[9][2] ;
 wire \po_0.regf_0.rf[9][3] ;
 wire \po_0.regf_0.rf[9][4] ;
 wire \po_0.regf_0.rf[9][5] ;
 wire \po_0.regf_0.rf[9][6] ;
 wire \po_0.regf_0.rf[9][7] ;
 wire \po_0.regf_0.rf[9][8] ;
 wire \po_0.regf_0.rf[9][9] ;
 wire \po_0.regf_0.rp_addr[0] ;
 wire \po_0.regf_0.rp_addr[1] ;
 wire \po_0.regf_0.rp_addr[2] ;
 wire \po_0.regf_0.rp_addr[3] ;
 wire \po_0.regf_0.rp_rd ;
 wire \po_0.regf_0.rq_addr[0] ;
 wire \po_0.regf_0.rq_addr[1] ;
 wire \po_0.regf_0.rq_addr[2] ;
 wire \po_0.regf_0.rq_addr[3] ;
 wire \po_0.regf_0.rq_rd ;
 wire \po_0.regf_0.w_addr[0] ;
 wire \po_0.regf_0.w_addr[1] ;
 wire \po_0.regf_0.w_addr[2] ;
 wire \po_0.regf_0.w_addr[3] ;
 wire \po_0.regf_0.w_wr ;
 wire \uc_0._00_ ;
 wire \uc_0._01_ ;
 wire \uc_0._02_ ;
 wire \uc_0._03_ ;
 wire \uc_0._21_[0] ;
 wire \uc_0._21_[10] ;
 wire \uc_0._21_[11] ;
 wire \uc_0._21_[12] ;
 wire \uc_0._21_[13] ;
 wire \uc_0._21_[14] ;
 wire \uc_0._21_[15] ;
 wire \uc_0._21_[1] ;
 wire \uc_0._21_[2] ;
 wire \uc_0._21_[3] ;
 wire \uc_0._21_[4] ;
 wire \uc_0._21_[5] ;
 wire \uc_0._21_[6] ;
 wire \uc_0._21_[7] ;
 wire \uc_0._21_[8] ;
 wire \uc_0._21_[9] ;
 wire \uc_0.bc_0._05_[0] ;
 wire \uc_0.bc_0._05_[1] ;
 wire \uc_0.bc_0._05_[2] ;
 wire \uc_0.bc_0._05_[3] ;
 wire \uc_0.bc_0._70_[0] ;
 wire \uc_0.bc_0._70_[1] ;
 wire \uc_0.bc_0._70_[2] ;
 wire \uc_0.bc_0._70_[3] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net96));
 sky130_fd_sc_hd__decap_8 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_94 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__clkbuf_2 _1640_ (.A(\po_0.alu_0.s0 ),
    .X(_1487_));
 sky130_fd_sc_hd__clkbuf_2 _1641_ (.A(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__clkbuf_2 _1642_ (.A(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__inv_2 _1643_ (.A(\po_0.alu_0.s1 ),
    .Y(_1490_));
 sky130_fd_sc_hd__clkbuf_2 _1644_ (.A(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1645_ (.A(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__clkbuf_2 _1646_ (.A(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__or2_1 _1647_ (.A(_1489_),
    .B(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__clkbuf_1 _1648_ (.A(_1494_),
    .X(_1631_));
 sky130_fd_sc_hd__or2_1 _1649_ (.A(_1489_),
    .B(_1493_),
    .X(_1495_));
 sky130_fd_sc_hd__clkbuf_1 _1650_ (.A(_1495_),
    .X(_1630_));
 sky130_fd_sc_hd__or2_1 _1651_ (.A(_1489_),
    .B(_1493_),
    .X(_1496_));
 sky130_fd_sc_hd__clkbuf_1 _1652_ (.A(_1496_),
    .X(_1629_));
 sky130_fd_sc_hd__or2_1 _1653_ (.A(_1489_),
    .B(_1493_),
    .X(_1497_));
 sky130_fd_sc_hd__clkbuf_1 _1654_ (.A(_1497_),
    .X(_1628_));
 sky130_fd_sc_hd__or2_1 _1655_ (.A(_1489_),
    .B(_1493_),
    .X(_1498_));
 sky130_fd_sc_hd__clkbuf_1 _1656_ (.A(_1498_),
    .X(_1627_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1657_ (.A(_1488_),
    .X(_1499_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1658_ (.A(_1499_),
    .X(_1500_));
 sky130_fd_sc_hd__or2_1 _1659_ (.A(_1500_),
    .B(_1493_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _1660_ (.A(_1501_),
    .X(_1626_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1661_ (.A(_1492_),
    .X(_1502_));
 sky130_fd_sc_hd__or2_1 _1662_ (.A(_1500_),
    .B(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__clkbuf_1 _1663_ (.A(_1503_),
    .X(_1625_));
 sky130_fd_sc_hd__or2_1 _1664_ (.A(_1500_),
    .B(_1502_),
    .X(_1504_));
 sky130_fd_sc_hd__clkbuf_1 _1665_ (.A(_1504_),
    .X(_1624_));
 sky130_fd_sc_hd__or2_1 _1666_ (.A(_1500_),
    .B(_1502_),
    .X(_1505_));
 sky130_fd_sc_hd__clkbuf_1 _1667_ (.A(_1505_),
    .X(_1632_));
 sky130_fd_sc_hd__or2_1 _1668_ (.A(_1500_),
    .B(_1502_),
    .X(_1506_));
 sky130_fd_sc_hd__clkbuf_1 _1669_ (.A(_1506_),
    .X(_1633_));
 sky130_fd_sc_hd__or2_1 _1670_ (.A(_1500_),
    .B(_1502_),
    .X(_1507_));
 sky130_fd_sc_hd__clkbuf_1 _1671_ (.A(_1507_),
    .X(_1634_));
 sky130_fd_sc_hd__or2_1 _1672_ (.A(_1499_),
    .B(_1502_),
    .X(_1508_));
 sky130_fd_sc_hd__clkbuf_1 _1673_ (.A(_1508_),
    .X(_1635_));
 sky130_fd_sc_hd__or2_1 _1674_ (.A(_1499_),
    .B(_1492_),
    .X(_1509_));
 sky130_fd_sc_hd__clkbuf_1 _1675_ (.A(_1509_),
    .X(_1636_));
 sky130_fd_sc_hd__or2_1 _1676_ (.A(_1499_),
    .B(_1492_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_1 _1677_ (.A(_1510_),
    .X(_1637_));
 sky130_fd_sc_hd__or2_1 _1678_ (.A(_1499_),
    .B(_1492_),
    .X(_1511_));
 sky130_fd_sc_hd__clkbuf_1 _1679_ (.A(_1511_),
    .X(_1638_));
 sky130_fd_sc_hd__or2_1 _1680_ (.A(_1499_),
    .B(_1492_),
    .X(_1512_));
 sky130_fd_sc_hd__clkbuf_1 _1681_ (.A(_1512_),
    .X(_1639_));
 sky130_fd_sc_hd__clkbuf_2 _1682_ (.A(net35),
    .X(_1513_));
 sky130_fd_sc_hd__or2_1 _1683_ (.A(\po_0._1_[0] ),
    .B(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__nand2_1 _1684_ (.A(\po_0._1_[0] ),
    .B(net35),
    .Y(_1515_));
 sky130_fd_sc_hd__and2_1 _1685_ (.A(_1514_),
    .B(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__clkbuf_1 _1686_ (.A(_1516_),
    .X(\po_0.alu_0._10_[0] ));
 sky130_fd_sc_hd__clkbuf_2 _1687_ (.A(net34),
    .X(_1517_));
 sky130_fd_sc_hd__nand2_1 _1688_ (.A(\uc_0.bc_0._05_[0] ),
    .B(\uc_0.bc_0._05_[1] ),
    .Y(_1518_));
 sky130_fd_sc_hd__nor2_1 _1689_ (.A(\uc_0.bc_0._05_[2] ),
    .B(\uc_0.bc_0._05_[3] ),
    .Y(_1519_));
 sky130_fd_sc_hd__nor4b_2 _1690_ (.A(\uc_0._21_[15] ),
    .B(\uc_0._21_[14] ),
    .C(_1518_),
    .D_N(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__and2b_1 _1691_ (.A_N(_1517_),
    .B(_1520_),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_2 _1692_ (.A(_1521_),
    .X(\uc_0.bc_0._70_[2] ));
 sky130_fd_sc_hd__clkbuf_2 _1693_ (.A(net36),
    .X(_1522_));
 sky130_fd_sc_hd__or4_1 _1694_ (.A(net50),
    .B(net86),
    .C(net85),
    .D(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__clkbuf_2 _1695_ (.A(net43),
    .X(_1524_));
 sky130_fd_sc_hd__nor4_1 _1696_ (.A(_1513_),
    .B(net87),
    .C(net44),
    .D(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__clkbuf_2 _1697_ (.A(net47),
    .X(_1526_));
 sky130_fd_sc_hd__nor4_1 _1698_ (.A(net46),
    .B(net45),
    .C(net48),
    .D(_1526_),
    .Y(_1527_));
 sky130_fd_sc_hd__nor4_1 _1699_ (.A(net83),
    .B(net84),
    .C(net41),
    .D(net40),
    .Y(_1528_));
 sky130_fd_sc_hd__nand3_2 _1700_ (.A(_1525_),
    .B(_1527_),
    .C(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__nor2_1 _1701_ (.A(_1523_),
    .B(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__nor2_1 _1702_ (.A(\uc_0.bc_0._05_[1] ),
    .B(\uc_0.bc_0._05_[2] ),
    .Y(_1531_));
 sky130_fd_sc_hd__and3_1 _1703_ (.A(\uc_0.bc_0._05_[0] ),
    .B(\uc_0.bc_0._05_[3] ),
    .C(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__nand2_1 _1704_ (.A(_1530_),
    .B(_1532_),
    .Y(_1533_));
 sky130_fd_sc_hd__nand2_1 _1705_ (.A(\uc_0._21_[13] ),
    .B(_1520_),
    .Y(_1534_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1706_ (.A(\uc_0.bc_0._05_[1] ),
    .X(_1535_));
 sky130_fd_sc_hd__xor2_1 _1707_ (.A(\uc_0.bc_0._05_[0] ),
    .B(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__nand2_1 _1708_ (.A(_1536_),
    .B(_1519_),
    .Y(_1537_));
 sky130_fd_sc_hd__a31o_1 _1709_ (.A1(_1533_),
    .A2(_1534_),
    .A3(_1537_),
    .B1(net34),
    .X(_1538_));
 sky130_fd_sc_hd__inv_2 _1710_ (.A(_1538_),
    .Y(\uc_0.bc_0._70_[1] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1711_ (.A(\uc_0.bc_0._05_[0] ),
    .X(_1539_));
 sky130_fd_sc_hd__o21ai_1 _1712_ (.A1(_1523_),
    .A2(_1529_),
    .B1(_1532_),
    .Y(_1540_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1713_ (.A(\uc_0.bc_0._05_[2] ),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_2 _1714_ (.A(\uc_0.bc_0._05_[3] ),
    .X(_1542_));
 sky130_fd_sc_hd__a211o_1 _1715_ (.A1(\uc_0._21_[13] ),
    .A2(\uc_0._21_[14] ),
    .B1(\uc_0._21_[15] ),
    .C1(\uc_0._21_[12] ),
    .X(_1543_));
 sky130_fd_sc_hd__or4b_1 _1716_ (.A(_1541_),
    .B(_1542_),
    .C(_1518_),
    .D_N(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__o2111a_1 _1717_ (.A1(_1519_),
    .A2(_1531_),
    .B1(_1539_),
    .C1(_1540_),
    .D1(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_2 _1718_ (.A(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__nor2_1 _1719_ (.A(_1517_),
    .B(_1546_),
    .Y(\uc_0.bc_0._70_[0] ));
 sky130_fd_sc_hd__or3b_1 _1720_ (.A(\uc_0._21_[13] ),
    .B(\uc_0._21_[15] ),
    .C_N(\uc_0._21_[14] ),
    .X(_1547_));
 sky130_fd_sc_hd__o41a_1 _1721_ (.A1(_1541_),
    .A2(_1542_),
    .A3(_1518_),
    .A4(_1547_),
    .B1(_1533_),
    .X(_1548_));
 sky130_fd_sc_hd__nor2_1 _1722_ (.A(_1517_),
    .B(_1548_),
    .Y(\uc_0.bc_0._70_[3] ));
 sky130_fd_sc_hd__clkbuf_2 _1723_ (.A(\uc_0._21_[4] ),
    .X(_1549_));
 sky130_fd_sc_hd__o211ai_2 _1724_ (.A1(_1517_),
    .A2(_1545_),
    .B1(_1538_),
    .C1(\uc_0.bc_0._70_[3] ),
    .Y(_1550_));
 sky130_fd_sc_hd__nand3_1 _1725_ (.A(_1521_),
    .B(\uc_0.bc_0._70_[1] ),
    .C(_1546_),
    .Y(_1551_));
 sky130_fd_sc_hd__nand2_2 _1726_ (.A(_1550_),
    .B(_1551_),
    .Y(_1552_));
 sky130_fd_sc_hd__buf_2 _1727_ (.A(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__mux2_1 _1728_ (.A0(\po_0.regf_0.rq_addr[0] ),
    .A1(_1549_),
    .S(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__clkbuf_1 _1729_ (.A(_1554_),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_2 _1730_ (.A(\uc_0._21_[5] ),
    .X(_1555_));
 sky130_fd_sc_hd__mux2_1 _1731_ (.A0(\po_0.regf_0.rq_addr[1] ),
    .A1(_1555_),
    .S(_1553_),
    .X(_1556_));
 sky130_fd_sc_hd__clkbuf_1 _1732_ (.A(_1556_),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_2 _1733_ (.A(\uc_0._21_[6] ),
    .X(_1557_));
 sky130_fd_sc_hd__mux2_1 _1734_ (.A0(\po_0.regf_0.rq_addr[2] ),
    .A1(_1557_),
    .S(_1553_),
    .X(_1558_));
 sky130_fd_sc_hd__clkbuf_1 _1735_ (.A(_1558_),
    .X(_0014_));
 sky130_fd_sc_hd__buf_2 _1736_ (.A(\uc_0._21_[7] ),
    .X(_1559_));
 sky130_fd_sc_hd__mux2_1 _1737_ (.A0(\po_0.regf_0.rq_addr[3] ),
    .A1(_1559_),
    .S(_1553_),
    .X(_1560_));
 sky130_fd_sc_hd__clkbuf_1 _1738_ (.A(_1560_),
    .X(_0015_));
 sky130_fd_sc_hd__clkbuf_4 _1739_ (.A(_0004_),
    .X(_1561_));
 sky130_fd_sc_hd__clkbuf_4 _1740_ (.A(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__buf_2 _1741_ (.A(_0005_),
    .X(_1563_));
 sky130_fd_sc_hd__clkbuf_4 _1742_ (.A(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__mux4_1 _1743_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(\po_0.regf_0.rf[5][0] ),
    .A2(\po_0.regf_0.rf[6][0] ),
    .A3(\po_0.regf_0.rf[7][0] ),
    .S0(_1562_),
    .S1(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__clkbuf_2 _1744_ (.A(_0006_),
    .X(_1566_));
 sky130_fd_sc_hd__buf_2 _1745_ (.A(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__buf_2 _1746_ (.A(_0007_),
    .X(_1568_));
 sky130_fd_sc_hd__a21o_1 _1747_ (.A1(_1565_),
    .A2(_1567_),
    .B1(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__buf_2 _1748_ (.A(_0006_),
    .X(_1570_));
 sky130_fd_sc_hd__clkbuf_2 _1749_ (.A(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__clkbuf_2 _1750_ (.A(_0004_),
    .X(_1572_));
 sky130_fd_sc_hd__clkbuf_4 _1751_ (.A(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__clkbuf_2 _1752_ (.A(_0005_),
    .X(_1574_));
 sky130_fd_sc_hd__buf_2 _1753_ (.A(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__mux4_1 _1754_ (.A0(\po_0.regf_0.rf[0][0] ),
    .A1(\po_0.regf_0.rf[1][0] ),
    .A2(\po_0.regf_0.rf[2][0] ),
    .A3(\po_0.regf_0.rf[3][0] ),
    .S0(_1573_),
    .S1(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__and2b_1 _1755_ (.A_N(_1571_),
    .B(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__buf_4 _1756_ (.A(_1561_),
    .X(_1578_));
 sky130_fd_sc_hd__clkbuf_4 _1757_ (.A(_1563_),
    .X(_1579_));
 sky130_fd_sc_hd__mux4_1 _1758_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(\po_0.regf_0.rf[13][0] ),
    .A2(\po_0.regf_0.rf[14][0] ),
    .A3(\po_0.regf_0.rf[15][0] ),
    .S0(_1578_),
    .S1(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__buf_2 _1759_ (.A(_1566_),
    .X(_1581_));
 sky130_fd_sc_hd__clkinv_2 _1760_ (.A(_0007_),
    .Y(_1582_));
 sky130_fd_sc_hd__clkbuf_2 _1761_ (.A(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__a21o_1 _1762_ (.A1(_1580_),
    .A2(_1581_),
    .B1(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__clkbuf_2 _1763_ (.A(_1566_),
    .X(_1585_));
 sky130_fd_sc_hd__mux4_1 _1764_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(\po_0.regf_0.rf[9][0] ),
    .A2(\po_0.regf_0.rf[10][0] ),
    .A3(\po_0.regf_0.rf[11][0] ),
    .S0(_1573_),
    .S1(_1575_),
    .X(_1586_));
 sky130_fd_sc_hd__and2b_1 _1765_ (.A_N(_1585_),
    .B(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__o22a_1 _1766_ (.A1(_1569_),
    .A2(_1577_),
    .B1(_1584_),
    .B2(_1587_),
    .X(\po_0.regf_0._5_[0] ));
 sky130_fd_sc_hd__mux4_1 _1767_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(\po_0.regf_0.rf[13][1] ),
    .A2(\po_0.regf_0.rf[14][1] ),
    .A3(\po_0.regf_0.rf[15][1] ),
    .S0(_1562_),
    .S1(_1564_),
    .X(_1588_));
 sky130_fd_sc_hd__buf_2 _1768_ (.A(_1582_),
    .X(_1589_));
 sky130_fd_sc_hd__a21o_1 _1769_ (.A1(_1588_),
    .A2(_1567_),
    .B1(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__clkbuf_2 _1770_ (.A(_1566_),
    .X(_1591_));
 sky130_fd_sc_hd__clkbuf_4 _1771_ (.A(_1572_),
    .X(_1592_));
 sky130_fd_sc_hd__clkbuf_4 _1772_ (.A(_1574_),
    .X(_1593_));
 sky130_fd_sc_hd__mux4_1 _1773_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(\po_0.regf_0.rf[9][1] ),
    .A2(\po_0.regf_0.rf[10][1] ),
    .A3(\po_0.regf_0.rf[11][1] ),
    .S0(_1592_),
    .S1(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__and2b_1 _1774_ (.A_N(_1591_),
    .B(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__buf_2 _1775_ (.A(_1568_),
    .X(_1596_));
 sky130_fd_sc_hd__buf_4 _1776_ (.A(_1572_),
    .X(_1597_));
 sky130_fd_sc_hd__clkbuf_4 _1777_ (.A(_1574_),
    .X(_1598_));
 sky130_fd_sc_hd__mux4_1 _1778_ (.A0(\po_0.regf_0.rf[0][1] ),
    .A1(\po_0.regf_0.rf[1][1] ),
    .A2(\po_0.regf_0.rf[2][1] ),
    .A3(\po_0.regf_0.rf[3][1] ),
    .S0(_1597_),
    .S1(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__clkbuf_4 _1779_ (.A(_1572_),
    .X(_1600_));
 sky130_fd_sc_hd__buf_2 _1780_ (.A(_1574_),
    .X(_1601_));
 sky130_fd_sc_hd__mux4_1 _1781_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(\po_0.regf_0.rf[5][1] ),
    .A2(\po_0.regf_0.rf[6][1] ),
    .A3(\po_0.regf_0.rf[7][1] ),
    .S0(_1600_),
    .S1(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__buf_2 _1782_ (.A(_0006_),
    .X(_1603_));
 sky130_fd_sc_hd__mux2_1 _1783_ (.A0(_1599_),
    .A1(_1602_),
    .S(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__o22a_1 _1784_ (.A1(_1590_),
    .A2(_1595_),
    .B1(_1596_),
    .B2(_1604_),
    .X(\po_0.regf_0._5_[1] ));
 sky130_fd_sc_hd__mux4_1 _1785_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(\po_0.regf_0.rf[13][2] ),
    .A2(\po_0.regf_0.rf[14][2] ),
    .A3(\po_0.regf_0.rf[15][2] ),
    .S0(_1562_),
    .S1(_1564_),
    .X(_1605_));
 sky130_fd_sc_hd__a21o_1 _1786_ (.A1(_1605_),
    .A2(_1567_),
    .B1(_1589_),
    .X(_1606_));
 sky130_fd_sc_hd__mux4_1 _1787_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(\po_0.regf_0.rf[9][2] ),
    .A2(\po_0.regf_0.rf[10][2] ),
    .A3(\po_0.regf_0.rf[11][2] ),
    .S0(_1592_),
    .S1(_1593_),
    .X(_1607_));
 sky130_fd_sc_hd__and2b_1 _1788_ (.A_N(_1591_),
    .B(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__buf_4 _1789_ (.A(_1572_),
    .X(_1609_));
 sky130_fd_sc_hd__clkbuf_4 _1790_ (.A(_1574_),
    .X(_1610_));
 sky130_fd_sc_hd__mux4_1 _1791_ (.A0(\po_0.regf_0.rf[0][2] ),
    .A1(\po_0.regf_0.rf[1][2] ),
    .A2(\po_0.regf_0.rf[2][2] ),
    .A3(\po_0.regf_0.rf[3][2] ),
    .S0(_1609_),
    .S1(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__mux4_1 _1792_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(\po_0.regf_0.rf[5][2] ),
    .A2(\po_0.regf_0.rf[6][2] ),
    .A3(\po_0.regf_0.rf[7][2] ),
    .S0(_1600_),
    .S1(_1601_),
    .X(_1612_));
 sky130_fd_sc_hd__clkbuf_4 _1793_ (.A(_0006_),
    .X(_1613_));
 sky130_fd_sc_hd__mux2_1 _1794_ (.A0(_1611_),
    .A1(_1612_),
    .S(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__o22a_1 _1795_ (.A1(_1606_),
    .A2(_1608_),
    .B1(_1596_),
    .B2(_1614_),
    .X(\po_0.regf_0._5_[2] ));
 sky130_fd_sc_hd__mux4_1 _1796_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(\po_0.regf_0.rf[9][3] ),
    .A2(\po_0.regf_0.rf[10][3] ),
    .A3(\po_0.regf_0.rf[11][3] ),
    .S0(_1597_),
    .S1(_1598_),
    .X(_1615_));
 sky130_fd_sc_hd__and2b_1 _1797_ (.A_N(_1603_),
    .B(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__mux4_1 _1798_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(\po_0.regf_0.rf[13][3] ),
    .A2(\po_0.regf_0.rf[14][3] ),
    .A3(\po_0.regf_0.rf[15][3] ),
    .S0(_1562_),
    .S1(_1564_),
    .X(_1617_));
 sky130_fd_sc_hd__a21o_1 _1799_ (.A1(_1617_),
    .A2(_1585_),
    .B1(_1583_),
    .X(_1618_));
 sky130_fd_sc_hd__mux4_1 _1800_ (.A0(\po_0.regf_0.rf[0][3] ),
    .A1(\po_0.regf_0.rf[1][3] ),
    .A2(\po_0.regf_0.rf[2][3] ),
    .A3(\po_0.regf_0.rf[3][3] ),
    .S0(_1573_),
    .S1(_1575_),
    .X(_1619_));
 sky130_fd_sc_hd__and2b_1 _1801_ (.A_N(_1571_),
    .B(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__mux4_1 _1802_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(\po_0.regf_0.rf[5][3] ),
    .A2(\po_0.regf_0.rf[6][3] ),
    .A3(\po_0.regf_0.rf[7][3] ),
    .S0(_1578_),
    .S1(_1579_),
    .X(_1621_));
 sky130_fd_sc_hd__a21o_1 _1803_ (.A1(_1621_),
    .A2(_1581_),
    .B1(_1568_),
    .X(_1622_));
 sky130_fd_sc_hd__o22a_1 _1804_ (.A1(_1616_),
    .A2(_1618_),
    .B1(_1620_),
    .B2(_1622_),
    .X(\po_0.regf_0._5_[3] ));
 sky130_fd_sc_hd__mux4_1 _1805_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(\po_0.regf_0.rf[13][4] ),
    .A2(\po_0.regf_0.rf[14][4] ),
    .A3(\po_0.regf_0.rf[15][4] ),
    .S0(_1562_),
    .S1(_1564_),
    .X(_1623_));
 sky130_fd_sc_hd__a21o_1 _1806_ (.A1(_1623_),
    .A2(_1567_),
    .B1(_1589_),
    .X(_0346_));
 sky130_fd_sc_hd__mux4_1 _1807_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(\po_0.regf_0.rf[9][4] ),
    .A2(\po_0.regf_0.rf[10][4] ),
    .A3(\po_0.regf_0.rf[11][4] ),
    .S0(_1592_),
    .S1(_1593_),
    .X(_0347_));
 sky130_fd_sc_hd__and2b_1 _1808_ (.A_N(_1591_),
    .B(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__mux4_1 _1809_ (.A0(\po_0.regf_0.rf[0][4] ),
    .A1(\po_0.regf_0.rf[1][4] ),
    .A2(\po_0.regf_0.rf[2][4] ),
    .A3(\po_0.regf_0.rf[3][4] ),
    .S0(_1609_),
    .S1(_1610_),
    .X(_0349_));
 sky130_fd_sc_hd__mux4_1 _1810_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(\po_0.regf_0.rf[5][4] ),
    .A2(\po_0.regf_0.rf[6][4] ),
    .A3(\po_0.regf_0.rf[7][4] ),
    .S0(_1600_),
    .S1(_1601_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _1811_ (.A0(_0349_),
    .A1(_0350_),
    .S(_1613_),
    .X(_0351_));
 sky130_fd_sc_hd__o22a_1 _1812_ (.A1(_0346_),
    .A2(_0348_),
    .B1(_1596_),
    .B2(_0351_),
    .X(\po_0.regf_0._5_[4] ));
 sky130_fd_sc_hd__buf_4 _1813_ (.A(_1561_),
    .X(_0352_));
 sky130_fd_sc_hd__buf_4 _1814_ (.A(_1563_),
    .X(_0353_));
 sky130_fd_sc_hd__mux4_1 _1815_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(\po_0.regf_0.rf[13][5] ),
    .A2(\po_0.regf_0.rf[14][5] ),
    .A3(\po_0.regf_0.rf[15][5] ),
    .S0(_0352_),
    .S1(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__a21o_1 _1816_ (.A1(_0354_),
    .A2(_1567_),
    .B1(_1589_),
    .X(_0355_));
 sky130_fd_sc_hd__mux4_1 _1817_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(\po_0.regf_0.rf[9][5] ),
    .A2(\po_0.regf_0.rf[10][5] ),
    .A3(\po_0.regf_0.rf[11][5] ),
    .S0(_1592_),
    .S1(_1593_),
    .X(_0356_));
 sky130_fd_sc_hd__and2b_1 _1818_ (.A_N(_1591_),
    .B(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__mux4_1 _1819_ (.A0(\po_0.regf_0.rf[0][5] ),
    .A1(\po_0.regf_0.rf[1][5] ),
    .A2(\po_0.regf_0.rf[2][5] ),
    .A3(\po_0.regf_0.rf[3][5] ),
    .S0(_1609_),
    .S1(_1610_),
    .X(_0358_));
 sky130_fd_sc_hd__mux4_1 _1820_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(\po_0.regf_0.rf[5][5] ),
    .A2(\po_0.regf_0.rf[6][5] ),
    .A3(\po_0.regf_0.rf[7][5] ),
    .S0(_1600_),
    .S1(_1601_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _1821_ (.A0(_0358_),
    .A1(_0359_),
    .S(_1613_),
    .X(_0360_));
 sky130_fd_sc_hd__o22a_1 _1822_ (.A1(_0355_),
    .A2(_0357_),
    .B1(_1596_),
    .B2(_0360_),
    .X(\po_0.regf_0._5_[5] ));
 sky130_fd_sc_hd__clkbuf_4 _1823_ (.A(_0004_),
    .X(_0361_));
 sky130_fd_sc_hd__buf_2 _1824_ (.A(_0005_),
    .X(_0362_));
 sky130_fd_sc_hd__mux4_1 _1825_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(\po_0.regf_0.rf[9][6] ),
    .A2(\po_0.regf_0.rf[10][6] ),
    .A3(\po_0.regf_0.rf[11][6] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__mux4_1 _1826_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(\po_0.regf_0.rf[13][6] ),
    .A2(\po_0.regf_0.rf[14][6] ),
    .A3(\po_0.regf_0.rf[15][6] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _1827_ (.A0(_0363_),
    .A1(_0364_),
    .S(_1570_),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_4 _1828_ (.A(_0004_),
    .X(_0366_));
 sky130_fd_sc_hd__buf_2 _1829_ (.A(_0005_),
    .X(_0367_));
 sky130_fd_sc_hd__mux4_1 _1830_ (.A0(\po_0.regf_0.rf[0][6] ),
    .A1(\po_0.regf_0.rf[1][6] ),
    .A2(\po_0.regf_0.rf[2][6] ),
    .A3(\po_0.regf_0.rf[3][6] ),
    .S0(_0366_),
    .S1(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__mux4_1 _1831_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(\po_0.regf_0.rf[5][6] ),
    .A2(\po_0.regf_0.rf[6][6] ),
    .A3(\po_0.regf_0.rf[7][6] ),
    .S0(_0366_),
    .S1(_0367_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _1832_ (.A0(_0368_),
    .A1(_0369_),
    .S(_1570_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _1833_ (.A0(_0365_),
    .A1(_0370_),
    .S(_1582_),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_1 _1834_ (.A(_0371_),
    .X(\po_0.regf_0._5_[6] ));
 sky130_fd_sc_hd__mux4_1 _1835_ (.A0(\po_0.regf_0.rf[4][7] ),
    .A1(\po_0.regf_0.rf[5][7] ),
    .A2(\po_0.regf_0.rf[6][7] ),
    .A3(\po_0.regf_0.rf[7][7] ),
    .S0(_0352_),
    .S1(_0353_),
    .X(_0372_));
 sky130_fd_sc_hd__a21o_1 _1836_ (.A1(_0372_),
    .A2(_1567_),
    .B1(_0007_),
    .X(_0373_));
 sky130_fd_sc_hd__mux4_1 _1837_ (.A0(\po_0.regf_0.rf[0][7] ),
    .A1(\po_0.regf_0.rf[1][7] ),
    .A2(\po_0.regf_0.rf[2][7] ),
    .A3(\po_0.regf_0.rf[3][7] ),
    .S0(_1592_),
    .S1(_1593_),
    .X(_0374_));
 sky130_fd_sc_hd__and2b_1 _1838_ (.A_N(_1591_),
    .B(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__mux4_1 _1839_ (.A0(\po_0.regf_0.rf[12][7] ),
    .A1(\po_0.regf_0.rf[13][7] ),
    .A2(\po_0.regf_0.rf[14][7] ),
    .A3(\po_0.regf_0.rf[15][7] ),
    .S0(_1578_),
    .S1(_1579_),
    .X(_0376_));
 sky130_fd_sc_hd__a21o_1 _1840_ (.A1(_0376_),
    .A2(_1581_),
    .B1(_1583_),
    .X(_0377_));
 sky130_fd_sc_hd__mux4_1 _1841_ (.A0(\po_0.regf_0.rf[8][7] ),
    .A1(\po_0.regf_0.rf[9][7] ),
    .A2(\po_0.regf_0.rf[10][7] ),
    .A3(\po_0.regf_0.rf[11][7] ),
    .S0(_1573_),
    .S1(_1575_),
    .X(_0378_));
 sky130_fd_sc_hd__and2b_1 _1842_ (.A_N(_1585_),
    .B(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__o22a_1 _1843_ (.A1(_0373_),
    .A2(_0375_),
    .B1(_0377_),
    .B2(_0379_),
    .X(\po_0.regf_0._5_[7] ));
 sky130_fd_sc_hd__mux4_1 _1844_ (.A0(\po_0.regf_0.rf[4][8] ),
    .A1(\po_0.regf_0.rf[5][8] ),
    .A2(\po_0.regf_0.rf[6][8] ),
    .A3(\po_0.regf_0.rf[7][8] ),
    .S0(_0352_),
    .S1(_0353_),
    .X(_0380_));
 sky130_fd_sc_hd__a21o_1 _1845_ (.A1(_0380_),
    .A2(_1571_),
    .B1(_0007_),
    .X(_0381_));
 sky130_fd_sc_hd__mux4_1 _1846_ (.A0(\po_0.regf_0.rf[0][8] ),
    .A1(\po_0.regf_0.rf[1][8] ),
    .A2(\po_0.regf_0.rf[2][8] ),
    .A3(\po_0.regf_0.rf[3][8] ),
    .S0(_1592_),
    .S1(_1593_),
    .X(_0382_));
 sky130_fd_sc_hd__and2b_1 _1847_ (.A_N(_1591_),
    .B(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__mux4_1 _1848_ (.A0(\po_0.regf_0.rf[12][8] ),
    .A1(\po_0.regf_0.rf[13][8] ),
    .A2(\po_0.regf_0.rf[14][8] ),
    .A3(\po_0.regf_0.rf[15][8] ),
    .S0(_1578_),
    .S1(_1579_),
    .X(_0384_));
 sky130_fd_sc_hd__a21o_1 _1849_ (.A1(_0384_),
    .A2(_1581_),
    .B1(_1583_),
    .X(_0385_));
 sky130_fd_sc_hd__mux4_1 _1850_ (.A0(\po_0.regf_0.rf[8][8] ),
    .A1(\po_0.regf_0.rf[9][8] ),
    .A2(\po_0.regf_0.rf[10][8] ),
    .A3(\po_0.regf_0.rf[11][8] ),
    .S0(_1573_),
    .S1(_1575_),
    .X(_0386_));
 sky130_fd_sc_hd__and2b_1 _1851_ (.A_N(_1585_),
    .B(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__o22a_1 _1852_ (.A1(_0381_),
    .A2(_0383_),
    .B1(_0385_),
    .B2(_0387_),
    .X(\po_0.regf_0._5_[8] ));
 sky130_fd_sc_hd__mux4_1 _1853_ (.A0(\po_0.regf_0.rf[0][9] ),
    .A1(\po_0.regf_0.rf[1][9] ),
    .A2(\po_0.regf_0.rf[2][9] ),
    .A3(\po_0.regf_0.rf[3][9] ),
    .S0(_1597_),
    .S1(_1598_),
    .X(_0388_));
 sky130_fd_sc_hd__and2b_1 _1854_ (.A_N(_1603_),
    .B(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__mux4_1 _1855_ (.A0(\po_0.regf_0.rf[4][9] ),
    .A1(\po_0.regf_0.rf[5][9] ),
    .A2(\po_0.regf_0.rf[6][9] ),
    .A3(\po_0.regf_0.rf[7][9] ),
    .S0(_1562_),
    .S1(_1564_),
    .X(_0390_));
 sky130_fd_sc_hd__a21o_1 _1856_ (.A1(_0390_),
    .A2(_1585_),
    .B1(_1568_),
    .X(_0391_));
 sky130_fd_sc_hd__mux4_1 _1857_ (.A0(\po_0.regf_0.rf[8][9] ),
    .A1(\po_0.regf_0.rf[9][9] ),
    .A2(\po_0.regf_0.rf[10][9] ),
    .A3(\po_0.regf_0.rf[11][9] ),
    .S0(_1609_),
    .S1(_1610_),
    .X(_0392_));
 sky130_fd_sc_hd__mux4_1 _1858_ (.A0(\po_0.regf_0.rf[12][9] ),
    .A1(\po_0.regf_0.rf[13][9] ),
    .A2(\po_0.regf_0.rf[14][9] ),
    .A3(\po_0.regf_0.rf[15][9] ),
    .S0(_1600_),
    .S1(_1601_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _1859_ (.A0(_0392_),
    .A1(_0393_),
    .S(_1613_),
    .X(_0394_));
 sky130_fd_sc_hd__o22a_1 _1860_ (.A1(_0389_),
    .A2(_0391_),
    .B1(_1583_),
    .B2(_0394_),
    .X(\po_0.regf_0._5_[9] ));
 sky130_fd_sc_hd__mux4_1 _1861_ (.A0(\po_0.regf_0.rf[8][10] ),
    .A1(\po_0.regf_0.rf[9][10] ),
    .A2(\po_0.regf_0.rf[10][10] ),
    .A3(\po_0.regf_0.rf[11][10] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0395_));
 sky130_fd_sc_hd__mux4_1 _1862_ (.A0(\po_0.regf_0.rf[12][10] ),
    .A1(\po_0.regf_0.rf[13][10] ),
    .A2(\po_0.regf_0.rf[14][10] ),
    .A3(\po_0.regf_0.rf[15][10] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _1863_ (.A0(_0395_),
    .A1(_0396_),
    .S(_1570_),
    .X(_0397_));
 sky130_fd_sc_hd__mux4_1 _1864_ (.A0(\po_0.regf_0.rf[0][10] ),
    .A1(\po_0.regf_0.rf[1][10] ),
    .A2(\po_0.regf_0.rf[2][10] ),
    .A3(\po_0.regf_0.rf[3][10] ),
    .S0(_0366_),
    .S1(_0367_),
    .X(_0398_));
 sky130_fd_sc_hd__mux4_1 _1865_ (.A0(\po_0.regf_0.rf[4][10] ),
    .A1(\po_0.regf_0.rf[5][10] ),
    .A2(\po_0.regf_0.rf[6][10] ),
    .A3(\po_0.regf_0.rf[7][10] ),
    .S0(_0366_),
    .S1(_0367_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _1866_ (.A0(_0398_),
    .A1(_0399_),
    .S(_1570_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _1867_ (.A0(_0397_),
    .A1(_0400_),
    .S(_1582_),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _1868_ (.A(_0401_),
    .X(\po_0.regf_0._5_[10] ));
 sky130_fd_sc_hd__mux4_1 _1869_ (.A0(\po_0.regf_0.rf[12][11] ),
    .A1(\po_0.regf_0.rf[13][11] ),
    .A2(\po_0.regf_0.rf[14][11] ),
    .A3(\po_0.regf_0.rf[15][11] ),
    .S0(_0352_),
    .S1(_0353_),
    .X(_0402_));
 sky130_fd_sc_hd__a21o_1 _1870_ (.A1(_0402_),
    .A2(_1571_),
    .B1(_1589_),
    .X(_0403_));
 sky130_fd_sc_hd__mux4_1 _1871_ (.A0(\po_0.regf_0.rf[8][11] ),
    .A1(\po_0.regf_0.rf[9][11] ),
    .A2(\po_0.regf_0.rf[10][11] ),
    .A3(\po_0.regf_0.rf[11][11] ),
    .S0(_1597_),
    .S1(_1598_),
    .X(_0404_));
 sky130_fd_sc_hd__and2b_1 _1872_ (.A_N(_1603_),
    .B(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__mux4_1 _1873_ (.A0(\po_0.regf_0.rf[0][11] ),
    .A1(\po_0.regf_0.rf[1][11] ),
    .A2(\po_0.regf_0.rf[2][11] ),
    .A3(\po_0.regf_0.rf[3][11] ),
    .S0(_1609_),
    .S1(_1610_),
    .X(_0406_));
 sky130_fd_sc_hd__mux4_1 _1874_ (.A0(\po_0.regf_0.rf[4][11] ),
    .A1(\po_0.regf_0.rf[5][11] ),
    .A2(\po_0.regf_0.rf[6][11] ),
    .A3(\po_0.regf_0.rf[7][11] ),
    .S0(_1561_),
    .S1(_1563_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _1875_ (.A0(_0406_),
    .A1(_0407_),
    .S(_1613_),
    .X(_0408_));
 sky130_fd_sc_hd__o22a_1 _1876_ (.A1(_0403_),
    .A2(_0405_),
    .B1(_1596_),
    .B2(_0408_),
    .X(\po_0.regf_0._5_[11] ));
 sky130_fd_sc_hd__mux4_1 _1877_ (.A0(\po_0.regf_0.rf[8][12] ),
    .A1(\po_0.regf_0.rf[9][12] ),
    .A2(\po_0.regf_0.rf[10][12] ),
    .A3(\po_0.regf_0.rf[11][12] ),
    .S0(_1573_),
    .S1(_1575_),
    .X(_0409_));
 sky130_fd_sc_hd__and2b_1 _1878_ (.A_N(_1585_),
    .B(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__mux4_1 _1879_ (.A0(\po_0.regf_0.rf[12][12] ),
    .A1(\po_0.regf_0.rf[13][12] ),
    .A2(\po_0.regf_0.rf[14][12] ),
    .A3(\po_0.regf_0.rf[15][12] ),
    .S0(_1578_),
    .S1(_1579_),
    .X(_0411_));
 sky130_fd_sc_hd__a21o_1 _1880_ (.A1(_0411_),
    .A2(_1581_),
    .B1(_1583_),
    .X(_0412_));
 sky130_fd_sc_hd__mux4_1 _1881_ (.A0(\po_0.regf_0.rf[4][12] ),
    .A1(\po_0.regf_0.rf[5][12] ),
    .A2(\po_0.regf_0.rf[6][12] ),
    .A3(\po_0.regf_0.rf[7][12] ),
    .S0(_1578_),
    .S1(_1579_),
    .X(_0413_));
 sky130_fd_sc_hd__mux4_1 _1882_ (.A0(\po_0.regf_0.rf[0][12] ),
    .A1(\po_0.regf_0.rf[1][12] ),
    .A2(\po_0.regf_0.rf[2][12] ),
    .A3(\po_0.regf_0.rf[3][12] ),
    .S0(_1572_),
    .S1(_1574_),
    .X(_0414_));
 sky130_fd_sc_hd__and2b_1 _1883_ (.A_N(_1566_),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__a211o_1 _1884_ (.A1(_0413_),
    .A2(_1581_),
    .B1(_1568_),
    .C1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__o21a_1 _1885_ (.A1(_0410_),
    .A2(_0412_),
    .B1(_0416_),
    .X(\po_0.regf_0._5_[12] ));
 sky130_fd_sc_hd__mux4_1 _1886_ (.A0(\po_0.regf_0.rf[12][13] ),
    .A1(\po_0.regf_0.rf[13][13] ),
    .A2(\po_0.regf_0.rf[14][13] ),
    .A3(\po_0.regf_0.rf[15][13] ),
    .S0(_0352_),
    .S1(_0353_),
    .X(_0417_));
 sky130_fd_sc_hd__a21o_1 _1887_ (.A1(_0417_),
    .A2(_1571_),
    .B1(_1589_),
    .X(_0418_));
 sky130_fd_sc_hd__mux4_1 _1888_ (.A0(\po_0.regf_0.rf[8][13] ),
    .A1(\po_0.regf_0.rf[9][13] ),
    .A2(\po_0.regf_0.rf[10][13] ),
    .A3(\po_0.regf_0.rf[11][13] ),
    .S0(_1597_),
    .S1(_1598_),
    .X(_0419_));
 sky130_fd_sc_hd__and2b_1 _1889_ (.A_N(_1603_),
    .B(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__mux4_1 _1890_ (.A0(\po_0.regf_0.rf[0][13] ),
    .A1(\po_0.regf_0.rf[1][13] ),
    .A2(\po_0.regf_0.rf[2][13] ),
    .A3(\po_0.regf_0.rf[3][13] ),
    .S0(_1609_),
    .S1(_1610_),
    .X(_0421_));
 sky130_fd_sc_hd__mux4_1 _1891_ (.A0(\po_0.regf_0.rf[4][13] ),
    .A1(\po_0.regf_0.rf[5][13] ),
    .A2(\po_0.regf_0.rf[6][13] ),
    .A3(\po_0.regf_0.rf[7][13] ),
    .S0(_1561_),
    .S1(_1563_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _1892_ (.A0(_0421_),
    .A1(_0422_),
    .S(_1613_),
    .X(_0423_));
 sky130_fd_sc_hd__o22a_1 _1893_ (.A1(_0418_),
    .A2(_0420_),
    .B1(_1596_),
    .B2(_0423_),
    .X(\po_0.regf_0._5_[13] ));
 sky130_fd_sc_hd__mux4_1 _1894_ (.A0(\po_0.regf_0.rf[8][14] ),
    .A1(\po_0.regf_0.rf[9][14] ),
    .A2(\po_0.regf_0.rf[10][14] ),
    .A3(\po_0.regf_0.rf[11][14] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0424_));
 sky130_fd_sc_hd__mux4_1 _1895_ (.A0(\po_0.regf_0.rf[12][14] ),
    .A1(\po_0.regf_0.rf[13][14] ),
    .A2(\po_0.regf_0.rf[14][14] ),
    .A3(\po_0.regf_0.rf[15][14] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _1896_ (.A0(_0424_),
    .A1(_0425_),
    .S(_1570_),
    .X(_0426_));
 sky130_fd_sc_hd__mux4_1 _1897_ (.A0(\po_0.regf_0.rf[0][14] ),
    .A1(\po_0.regf_0.rf[1][14] ),
    .A2(\po_0.regf_0.rf[2][14] ),
    .A3(\po_0.regf_0.rf[3][14] ),
    .S0(_0366_),
    .S1(_0367_),
    .X(_0427_));
 sky130_fd_sc_hd__mux4_1 _1898_ (.A0(\po_0.regf_0.rf[4][14] ),
    .A1(\po_0.regf_0.rf[5][14] ),
    .A2(\po_0.regf_0.rf[6][14] ),
    .A3(\po_0.regf_0.rf[7][14] ),
    .S0(_0366_),
    .S1(_0367_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _1899_ (.A0(_0427_),
    .A1(_0428_),
    .S(_0006_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _1900_ (.A0(_0426_),
    .A1(_0429_),
    .S(_1582_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _1901_ (.A(_0430_),
    .X(\po_0.regf_0._5_[14] ));
 sky130_fd_sc_hd__mux4_1 _1902_ (.A0(\po_0.regf_0.rf[12][15] ),
    .A1(\po_0.regf_0.rf[13][15] ),
    .A2(\po_0.regf_0.rf[14][15] ),
    .A3(\po_0.regf_0.rf[15][15] ),
    .S0(_0352_),
    .S1(_0353_),
    .X(_0431_));
 sky130_fd_sc_hd__a21o_1 _1903_ (.A1(_0431_),
    .A2(_1571_),
    .B1(_1582_),
    .X(_0432_));
 sky130_fd_sc_hd__mux4_1 _1904_ (.A0(\po_0.regf_0.rf[8][15] ),
    .A1(\po_0.regf_0.rf[9][15] ),
    .A2(\po_0.regf_0.rf[10][15] ),
    .A3(\po_0.regf_0.rf[11][15] ),
    .S0(_1597_),
    .S1(_1598_),
    .X(_0433_));
 sky130_fd_sc_hd__and2b_1 _1905_ (.A_N(_1603_),
    .B(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__mux4_1 _1906_ (.A0(\po_0.regf_0.rf[0][15] ),
    .A1(\po_0.regf_0.rf[1][15] ),
    .A2(\po_0.regf_0.rf[2][15] ),
    .A3(\po_0.regf_0.rf[3][15] ),
    .S0(_1600_),
    .S1(_1601_),
    .X(_0435_));
 sky130_fd_sc_hd__mux4_1 _1907_ (.A0(\po_0.regf_0.rf[4][15] ),
    .A1(\po_0.regf_0.rf[5][15] ),
    .A2(\po_0.regf_0.rf[6][15] ),
    .A3(\po_0.regf_0.rf[7][15] ),
    .S0(_1561_),
    .S1(_1563_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _1908_ (.A0(_0435_),
    .A1(_0436_),
    .S(_1566_),
    .X(_0437_));
 sky130_fd_sc_hd__o22a_1 _1909_ (.A1(_0432_),
    .A2(_0434_),
    .B1(_1568_),
    .B2(_0437_),
    .X(\po_0.regf_0._5_[15] ));
 sky130_fd_sc_hd__buf_2 _1910_ (.A(_0002_),
    .X(_0438_));
 sky130_fd_sc_hd__buf_2 _1911_ (.A(_0000_),
    .X(_0439_));
 sky130_fd_sc_hd__buf_2 _1912_ (.A(_0001_),
    .X(_0440_));
 sky130_fd_sc_hd__mux4_1 _1913_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(\po_0.regf_0.rf[9][0] ),
    .A2(\po_0.regf_0.rf[10][0] ),
    .A3(\po_0.regf_0.rf[11][0] ),
    .S0(_0439_),
    .S1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__or2b_1 _1914_ (.A(_0438_),
    .B_N(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__buf_2 _1915_ (.A(_0003_),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_4 _1916_ (.A(_0439_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_4 _1917_ (.A(_0440_),
    .X(_0445_));
 sky130_fd_sc_hd__mux4_1 _1918_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(\po_0.regf_0.rf[13][0] ),
    .A2(\po_0.regf_0.rf[14][0] ),
    .A3(\po_0.regf_0.rf[15][0] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__buf_2 _1919_ (.A(_0438_),
    .X(_0447_));
 sky130_fd_sc_hd__nand2_1 _1920_ (.A(_0446_),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1921_ (.A(_0002_),
    .X(_0449_));
 sky130_fd_sc_hd__buf_2 _1922_ (.A(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__buf_4 _1923_ (.A(_0000_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_4 _1924_ (.A(_0001_),
    .X(_0452_));
 sky130_fd_sc_hd__mux4_1 _1925_ (.A0(\po_0.regf_0.rf[0][0] ),
    .A1(\po_0.regf_0.rf[1][0] ),
    .A2(\po_0.regf_0.rf[2][0] ),
    .A3(\po_0.regf_0.rf[3][0] ),
    .S0(_0451_),
    .S1(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__or2b_1 _1926_ (.A(_0450_),
    .B_N(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__mux4_1 _1927_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(\po_0.regf_0.rf[5][0] ),
    .A2(\po_0.regf_0.rf[6][0] ),
    .A3(\po_0.regf_0.rf[7][0] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0455_));
 sky130_fd_sc_hd__a21oi_1 _1928_ (.A1(_0455_),
    .A2(_0447_),
    .B1(_0443_),
    .Y(_0456_));
 sky130_fd_sc_hd__a32oi_4 _1929_ (.A1(_0442_),
    .A2(_0443_),
    .A3(_0448_),
    .B1(_0454_),
    .B2(_0456_),
    .Y(\po_0.regf_0._3_[0] ));
 sky130_fd_sc_hd__clkbuf_2 _1930_ (.A(_0000_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_4 _1931_ (.A(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_2 _1932_ (.A(_0001_),
    .X(_0459_));
 sky130_fd_sc_hd__buf_2 _1933_ (.A(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__mux4_1 _1934_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(\po_0.regf_0.rf[13][1] ),
    .A2(\po_0.regf_0.rf[14][1] ),
    .A3(\po_0.regf_0.rf[15][1] ),
    .S0(_0458_),
    .S1(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__buf_2 _1935_ (.A(_0449_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_2 _1936_ (.A(_0003_),
    .X(_0463_));
 sky130_fd_sc_hd__a21bo_1 _1937_ (.A1(_0461_),
    .A2(_0462_),
    .B1_N(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__clkbuf_2 _1938_ (.A(_0449_),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_4 _1939_ (.A(_0457_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_4 _1940_ (.A(_0459_),
    .X(_0467_));
 sky130_fd_sc_hd__mux4_1 _1941_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(\po_0.regf_0.rf[9][1] ),
    .A2(\po_0.regf_0.rf[10][1] ),
    .A3(\po_0.regf_0.rf[11][1] ),
    .S0(_0466_),
    .S1(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__and2b_1 _1942_ (.A_N(_0465_),
    .B(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__buf_2 _1943_ (.A(_0003_),
    .X(_0470_));
 sky130_fd_sc_hd__buf_2 _1944_ (.A(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_4 _1945_ (.A(_0457_),
    .X(_0472_));
 sky130_fd_sc_hd__buf_2 _1946_ (.A(_0459_),
    .X(_0473_));
 sky130_fd_sc_hd__mux4_1 _1947_ (.A0(\po_0.regf_0.rf[0][1] ),
    .A1(\po_0.regf_0.rf[1][1] ),
    .A2(\po_0.regf_0.rf[2][1] ),
    .A3(\po_0.regf_0.rf[3][1] ),
    .S0(_0472_),
    .S1(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__buf_4 _1948_ (.A(_0000_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_4 _1949_ (.A(_0001_),
    .X(_0476_));
 sky130_fd_sc_hd__mux4_1 _1950_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(\po_0.regf_0.rf[5][1] ),
    .A2(\po_0.regf_0.rf[6][1] ),
    .A3(\po_0.regf_0.rf[7][1] ),
    .S0(_0475_),
    .S1(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _1951_ (.A0(_0474_),
    .A1(_0477_),
    .S(_0450_),
    .X(_0478_));
 sky130_fd_sc_hd__o22a_1 _1952_ (.A1(_0464_),
    .A2(_0469_),
    .B1(_0471_),
    .B2(_0478_),
    .X(\po_0.regf_0._3_[1] ));
 sky130_fd_sc_hd__clkbuf_4 _1953_ (.A(_0439_),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_4 _1954_ (.A(_0440_),
    .X(_0480_));
 sky130_fd_sc_hd__mux4_1 _1955_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(\po_0.regf_0.rf[5][2] ),
    .A2(\po_0.regf_0.rf[6][2] ),
    .A3(\po_0.regf_0.rf[7][2] ),
    .S0(_0479_),
    .S1(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__a21o_1 _1956_ (.A1(_0481_),
    .A2(_0462_),
    .B1(_0470_),
    .X(_0482_));
 sky130_fd_sc_hd__mux4_1 _1957_ (.A0(\po_0.regf_0.rf[0][2] ),
    .A1(\po_0.regf_0.rf[1][2] ),
    .A2(\po_0.regf_0.rf[2][2] ),
    .A3(\po_0.regf_0.rf[3][2] ),
    .S0(_0466_),
    .S1(_0467_),
    .X(_0483_));
 sky130_fd_sc_hd__and2b_1 _1958_ (.A_N(_0465_),
    .B(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__mux4_1 _1959_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(\po_0.regf_0.rf[13][2] ),
    .A2(\po_0.regf_0.rf[14][2] ),
    .A3(\po_0.regf_0.rf[15][2] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0485_));
 sky130_fd_sc_hd__a21bo_1 _1960_ (.A1(_0485_),
    .A2(_0447_),
    .B1_N(_0463_),
    .X(_0486_));
 sky130_fd_sc_hd__buf_2 _1961_ (.A(_0438_),
    .X(_0487_));
 sky130_fd_sc_hd__buf_4 _1962_ (.A(_0457_),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_4 _1963_ (.A(_0459_),
    .X(_0489_));
 sky130_fd_sc_hd__mux4_1 _1964_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(\po_0.regf_0.rf[9][2] ),
    .A2(\po_0.regf_0.rf[10][2] ),
    .A3(\po_0.regf_0.rf[11][2] ),
    .S0(_0488_),
    .S1(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__and2b_1 _1965_ (.A_N(_0487_),
    .B(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__o22a_1 _1966_ (.A1(_0482_),
    .A2(_0484_),
    .B1(_0486_),
    .B2(_0491_),
    .X(\po_0.regf_0._3_[2] ));
 sky130_fd_sc_hd__mux4_1 _1967_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(\po_0.regf_0.rf[13][3] ),
    .A2(\po_0.regf_0.rf[14][3] ),
    .A3(\po_0.regf_0.rf[15][3] ),
    .S0(_0458_),
    .S1(_0460_),
    .X(_0492_));
 sky130_fd_sc_hd__buf_2 _1968_ (.A(_0003_),
    .X(_0493_));
 sky130_fd_sc_hd__a21bo_1 _1969_ (.A1(_0492_),
    .A2(_0462_),
    .B1_N(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__mux4_1 _1970_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(\po_0.regf_0.rf[9][3] ),
    .A2(\po_0.regf_0.rf[10][3] ),
    .A3(\po_0.regf_0.rf[11][3] ),
    .S0(_0466_),
    .S1(_0467_),
    .X(_0495_));
 sky130_fd_sc_hd__and2b_1 _1971_ (.A_N(_0465_),
    .B(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__mux4_1 _1972_ (.A0(\po_0.regf_0.rf[0][3] ),
    .A1(\po_0.regf_0.rf[1][3] ),
    .A2(\po_0.regf_0.rf[2][3] ),
    .A3(\po_0.regf_0.rf[3][3] ),
    .S0(_0472_),
    .S1(_0473_),
    .X(_0497_));
 sky130_fd_sc_hd__mux4_1 _1973_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(\po_0.regf_0.rf[5][3] ),
    .A2(\po_0.regf_0.rf[6][3] ),
    .A3(\po_0.regf_0.rf[7][3] ),
    .S0(_0475_),
    .S1(_0476_),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_4 _1974_ (.A(_0449_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _1975_ (.A0(_0497_),
    .A1(_0498_),
    .S(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__o22a_1 _1976_ (.A1(_0494_),
    .A2(_0496_),
    .B1(_0471_),
    .B2(_0500_),
    .X(\po_0.regf_0._3_[3] ));
 sky130_fd_sc_hd__mux4_1 _1977_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(\po_0.regf_0.rf[5][4] ),
    .A2(\po_0.regf_0.rf[6][4] ),
    .A3(\po_0.regf_0.rf[7][4] ),
    .S0(_0479_),
    .S1(_0480_),
    .X(_0501_));
 sky130_fd_sc_hd__a21o_1 _1978_ (.A1(_0501_),
    .A2(_0462_),
    .B1(_0470_),
    .X(_0502_));
 sky130_fd_sc_hd__mux4_1 _1979_ (.A0(\po_0.regf_0.rf[0][4] ),
    .A1(\po_0.regf_0.rf[1][4] ),
    .A2(\po_0.regf_0.rf[2][4] ),
    .A3(\po_0.regf_0.rf[3][4] ),
    .S0(_0466_),
    .S1(_0467_),
    .X(_0503_));
 sky130_fd_sc_hd__and2b_1 _1980_ (.A_N(_0465_),
    .B(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__mux4_1 _1981_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(\po_0.regf_0.rf[13][4] ),
    .A2(\po_0.regf_0.rf[14][4] ),
    .A3(\po_0.regf_0.rf[15][4] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0505_));
 sky130_fd_sc_hd__a21bo_1 _1982_ (.A1(_0505_),
    .A2(_0447_),
    .B1_N(_0463_),
    .X(_0506_));
 sky130_fd_sc_hd__mux4_1 _1983_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(\po_0.regf_0.rf[9][4] ),
    .A2(\po_0.regf_0.rf[10][4] ),
    .A3(\po_0.regf_0.rf[11][4] ),
    .S0(_0488_),
    .S1(_0489_),
    .X(_0507_));
 sky130_fd_sc_hd__and2b_1 _1984_ (.A_N(_0487_),
    .B(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__o22a_1 _1985_ (.A1(_0502_),
    .A2(_0504_),
    .B1(_0506_),
    .B2(_0508_),
    .X(\po_0.regf_0._3_[4] ));
 sky130_fd_sc_hd__mux4_1 _1986_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(\po_0.regf_0.rf[5][5] ),
    .A2(\po_0.regf_0.rf[6][5] ),
    .A3(\po_0.regf_0.rf[7][5] ),
    .S0(_0479_),
    .S1(_0480_),
    .X(_0509_));
 sky130_fd_sc_hd__a21o_1 _1987_ (.A1(_0509_),
    .A2(_0462_),
    .B1(_0470_),
    .X(_0510_));
 sky130_fd_sc_hd__buf_2 _1988_ (.A(_0449_),
    .X(_0511_));
 sky130_fd_sc_hd__clkbuf_4 _1989_ (.A(_0457_),
    .X(_0512_));
 sky130_fd_sc_hd__buf_2 _1990_ (.A(_0459_),
    .X(_0513_));
 sky130_fd_sc_hd__mux4_1 _1991_ (.A0(\po_0.regf_0.rf[0][5] ),
    .A1(\po_0.regf_0.rf[1][5] ),
    .A2(\po_0.regf_0.rf[2][5] ),
    .A3(\po_0.regf_0.rf[3][5] ),
    .S0(_0512_),
    .S1(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__and2b_1 _1992_ (.A_N(_0511_),
    .B(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__mux4_1 _1993_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(\po_0.regf_0.rf[13][5] ),
    .A2(\po_0.regf_0.rf[14][5] ),
    .A3(\po_0.regf_0.rf[15][5] ),
    .S0(_0479_),
    .S1(_0480_),
    .X(_0516_));
 sky130_fd_sc_hd__a21bo_1 _1994_ (.A1(_0516_),
    .A2(_0487_),
    .B1_N(_0463_),
    .X(_0517_));
 sky130_fd_sc_hd__mux4_1 _1995_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(\po_0.regf_0.rf[9][5] ),
    .A2(\po_0.regf_0.rf[10][5] ),
    .A3(\po_0.regf_0.rf[11][5] ),
    .S0(_0488_),
    .S1(_0489_),
    .X(_0518_));
 sky130_fd_sc_hd__and2b_1 _1996_ (.A_N(_0487_),
    .B(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__o22a_1 _1997_ (.A1(_0510_),
    .A2(_0515_),
    .B1(_0517_),
    .B2(_0519_),
    .X(\po_0.regf_0._3_[5] ));
 sky130_fd_sc_hd__mux4_1 _1998_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(\po_0.regf_0.rf[13][6] ),
    .A2(\po_0.regf_0.rf[14][6] ),
    .A3(\po_0.regf_0.rf[15][6] ),
    .S0(_0458_),
    .S1(_0460_),
    .X(_0520_));
 sky130_fd_sc_hd__a21bo_1 _1999_ (.A1(_0520_),
    .A2(_0462_),
    .B1_N(_0493_),
    .X(_0521_));
 sky130_fd_sc_hd__mux4_1 _2000_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(\po_0.regf_0.rf[9][6] ),
    .A2(\po_0.regf_0.rf[10][6] ),
    .A3(\po_0.regf_0.rf[11][6] ),
    .S0(_0512_),
    .S1(_0513_),
    .X(_0522_));
 sky130_fd_sc_hd__and2b_1 _2001_ (.A_N(_0511_),
    .B(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_4 _2002_ (.A(_0457_),
    .X(_0524_));
 sky130_fd_sc_hd__buf_2 _2003_ (.A(_0459_),
    .X(_0525_));
 sky130_fd_sc_hd__mux4_1 _2004_ (.A0(\po_0.regf_0.rf[0][6] ),
    .A1(\po_0.regf_0.rf[1][6] ),
    .A2(\po_0.regf_0.rf[2][6] ),
    .A3(\po_0.regf_0.rf[3][6] ),
    .S0(_0524_),
    .S1(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__mux4_1 _2005_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(\po_0.regf_0.rf[5][6] ),
    .A2(\po_0.regf_0.rf[6][6] ),
    .A3(\po_0.regf_0.rf[7][6] ),
    .S0(_0475_),
    .S1(_0476_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _2006_ (.A0(_0526_),
    .A1(_0527_),
    .S(_0499_),
    .X(_0528_));
 sky130_fd_sc_hd__o22a_1 _2007_ (.A1(_0521_),
    .A2(_0523_),
    .B1(_0471_),
    .B2(_0528_),
    .X(\po_0.regf_0._3_[6] ));
 sky130_fd_sc_hd__mux4_1 _2008_ (.A0(\po_0.regf_0.rf[12][7] ),
    .A1(\po_0.regf_0.rf[13][7] ),
    .A2(\po_0.regf_0.rf[14][7] ),
    .A3(\po_0.regf_0.rf[15][7] ),
    .S0(_0458_),
    .S1(_0460_),
    .X(_0529_));
 sky130_fd_sc_hd__buf_2 _2009_ (.A(_0449_),
    .X(_0530_));
 sky130_fd_sc_hd__a21bo_1 _2010_ (.A1(_0529_),
    .A2(_0530_),
    .B1_N(_0493_),
    .X(_0531_));
 sky130_fd_sc_hd__mux4_1 _2011_ (.A0(\po_0.regf_0.rf[8][7] ),
    .A1(\po_0.regf_0.rf[9][7] ),
    .A2(\po_0.regf_0.rf[10][7] ),
    .A3(\po_0.regf_0.rf[11][7] ),
    .S0(_0512_),
    .S1(_0513_),
    .X(_0532_));
 sky130_fd_sc_hd__and2b_1 _2012_ (.A_N(_0511_),
    .B(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__mux4_1 _2013_ (.A0(\po_0.regf_0.rf[0][7] ),
    .A1(\po_0.regf_0.rf[1][7] ),
    .A2(\po_0.regf_0.rf[2][7] ),
    .A3(\po_0.regf_0.rf[3][7] ),
    .S0(_0524_),
    .S1(_0525_),
    .X(_0534_));
 sky130_fd_sc_hd__mux4_1 _2014_ (.A0(\po_0.regf_0.rf[4][7] ),
    .A1(\po_0.regf_0.rf[5][7] ),
    .A2(\po_0.regf_0.rf[6][7] ),
    .A3(\po_0.regf_0.rf[7][7] ),
    .S0(_0475_),
    .S1(_0476_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _2015_ (.A0(_0534_),
    .A1(_0535_),
    .S(_0499_),
    .X(_0536_));
 sky130_fd_sc_hd__o22a_1 _2016_ (.A1(_0531_),
    .A2(_0533_),
    .B1(_0471_),
    .B2(_0536_),
    .X(\po_0.regf_0._3_[7] ));
 sky130_fd_sc_hd__mux4_1 _2017_ (.A0(\po_0.regf_0.rf[12][8] ),
    .A1(\po_0.regf_0.rf[13][8] ),
    .A2(\po_0.regf_0.rf[14][8] ),
    .A3(\po_0.regf_0.rf[15][8] ),
    .S0(_0458_),
    .S1(_0460_),
    .X(_0537_));
 sky130_fd_sc_hd__a21bo_1 _2018_ (.A1(_0537_),
    .A2(_0530_),
    .B1_N(_0493_),
    .X(_0538_));
 sky130_fd_sc_hd__mux4_1 _2019_ (.A0(\po_0.regf_0.rf[8][8] ),
    .A1(\po_0.regf_0.rf[9][8] ),
    .A2(\po_0.regf_0.rf[10][8] ),
    .A3(\po_0.regf_0.rf[11][8] ),
    .S0(_0512_),
    .S1(_0513_),
    .X(_0539_));
 sky130_fd_sc_hd__and2b_1 _2020_ (.A_N(_0511_),
    .B(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__mux4_1 _2021_ (.A0(\po_0.regf_0.rf[0][8] ),
    .A1(\po_0.regf_0.rf[1][8] ),
    .A2(\po_0.regf_0.rf[2][8] ),
    .A3(\po_0.regf_0.rf[3][8] ),
    .S0(_0524_),
    .S1(_0525_),
    .X(_0541_));
 sky130_fd_sc_hd__mux4_1 _2022_ (.A0(\po_0.regf_0.rf[4][8] ),
    .A1(\po_0.regf_0.rf[5][8] ),
    .A2(\po_0.regf_0.rf[6][8] ),
    .A3(\po_0.regf_0.rf[7][8] ),
    .S0(_0475_),
    .S1(_0476_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _2023_ (.A0(_0541_),
    .A1(_0542_),
    .S(_0499_),
    .X(_0543_));
 sky130_fd_sc_hd__o22a_1 _2024_ (.A1(_0538_),
    .A2(_0540_),
    .B1(_0471_),
    .B2(_0543_),
    .X(\po_0.regf_0._3_[8] ));
 sky130_fd_sc_hd__mux4_1 _2025_ (.A0(\po_0.regf_0.rf[8][9] ),
    .A1(\po_0.regf_0.rf[9][9] ),
    .A2(\po_0.regf_0.rf[10][9] ),
    .A3(\po_0.regf_0.rf[11][9] ),
    .S0(_0472_),
    .S1(_0473_),
    .X(_0544_));
 sky130_fd_sc_hd__and2b_1 _2026_ (.A_N(_0450_),
    .B(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__mux4_1 _2027_ (.A0(\po_0.regf_0.rf[12][9] ),
    .A1(\po_0.regf_0.rf[13][9] ),
    .A2(\po_0.regf_0.rf[14][9] ),
    .A3(\po_0.regf_0.rf[15][9] ),
    .S0(_0479_),
    .S1(_0480_),
    .X(_0546_));
 sky130_fd_sc_hd__a21bo_1 _2028_ (.A1(_0546_),
    .A2(_0487_),
    .B1_N(_0463_),
    .X(_0547_));
 sky130_fd_sc_hd__mux4_1 _2029_ (.A0(\po_0.regf_0.rf[0][9] ),
    .A1(\po_0.regf_0.rf[1][9] ),
    .A2(\po_0.regf_0.rf[2][9] ),
    .A3(\po_0.regf_0.rf[3][9] ),
    .S0(_0466_),
    .S1(_0467_),
    .X(_0548_));
 sky130_fd_sc_hd__and2b_1 _2030_ (.A_N(_0465_),
    .B(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__mux4_1 _2031_ (.A0(\po_0.regf_0.rf[4][9] ),
    .A1(\po_0.regf_0.rf[5][9] ),
    .A2(\po_0.regf_0.rf[6][9] ),
    .A3(\po_0.regf_0.rf[7][9] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0550_));
 sky130_fd_sc_hd__a21o_1 _2032_ (.A1(_0550_),
    .A2(_0447_),
    .B1(_0443_),
    .X(_0551_));
 sky130_fd_sc_hd__o22a_1 _2033_ (.A1(_0545_),
    .A2(_0547_),
    .B1(_0549_),
    .B2(_0551_),
    .X(\po_0.regf_0._3_[9] ));
 sky130_fd_sc_hd__mux4_1 _2034_ (.A0(\po_0.regf_0.rf[12][10] ),
    .A1(\po_0.regf_0.rf[13][10] ),
    .A2(\po_0.regf_0.rf[14][10] ),
    .A3(\po_0.regf_0.rf[15][10] ),
    .S0(_0458_),
    .S1(_0460_),
    .X(_0552_));
 sky130_fd_sc_hd__a21bo_1 _2035_ (.A1(_0552_),
    .A2(_0530_),
    .B1_N(_0493_),
    .X(_0553_));
 sky130_fd_sc_hd__mux4_1 _2036_ (.A0(\po_0.regf_0.rf[8][10] ),
    .A1(\po_0.regf_0.rf[9][10] ),
    .A2(\po_0.regf_0.rf[10][10] ),
    .A3(\po_0.regf_0.rf[11][10] ),
    .S0(_0512_),
    .S1(_0513_),
    .X(_0554_));
 sky130_fd_sc_hd__and2b_1 _2037_ (.A_N(_0511_),
    .B(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__mux4_1 _2038_ (.A0(\po_0.regf_0.rf[0][10] ),
    .A1(\po_0.regf_0.rf[1][10] ),
    .A2(\po_0.regf_0.rf[2][10] ),
    .A3(\po_0.regf_0.rf[3][10] ),
    .S0(_0524_),
    .S1(_0525_),
    .X(_0556_));
 sky130_fd_sc_hd__mux4_1 _2039_ (.A0(\po_0.regf_0.rf[4][10] ),
    .A1(\po_0.regf_0.rf[5][10] ),
    .A2(\po_0.regf_0.rf[6][10] ),
    .A3(\po_0.regf_0.rf[7][10] ),
    .S0(_0451_),
    .S1(_0452_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _2040_ (.A0(_0556_),
    .A1(_0557_),
    .S(_0499_),
    .X(_0558_));
 sky130_fd_sc_hd__o22a_1 _2041_ (.A1(_0553_),
    .A2(_0555_),
    .B1(_0471_),
    .B2(_0558_),
    .X(\po_0.regf_0._3_[10] ));
 sky130_fd_sc_hd__mux4_1 _2042_ (.A0(\po_0.regf_0.rf[12][11] ),
    .A1(\po_0.regf_0.rf[13][11] ),
    .A2(\po_0.regf_0.rf[14][11] ),
    .A3(\po_0.regf_0.rf[15][11] ),
    .S0(_0488_),
    .S1(_0489_),
    .X(_0559_));
 sky130_fd_sc_hd__a21bo_1 _2043_ (.A1(_0559_),
    .A2(_0530_),
    .B1_N(_0493_),
    .X(_0560_));
 sky130_fd_sc_hd__mux4_1 _2044_ (.A0(\po_0.regf_0.rf[8][11] ),
    .A1(\po_0.regf_0.rf[9][11] ),
    .A2(\po_0.regf_0.rf[10][11] ),
    .A3(\po_0.regf_0.rf[11][11] ),
    .S0(_0512_),
    .S1(_0513_),
    .X(_0561_));
 sky130_fd_sc_hd__and2b_1 _2045_ (.A_N(_0511_),
    .B(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__mux4_1 _2046_ (.A0(\po_0.regf_0.rf[0][11] ),
    .A1(\po_0.regf_0.rf[1][11] ),
    .A2(\po_0.regf_0.rf[2][11] ),
    .A3(\po_0.regf_0.rf[3][11] ),
    .S0(_0524_),
    .S1(_0525_),
    .X(_0563_));
 sky130_fd_sc_hd__mux4_1 _2047_ (.A0(\po_0.regf_0.rf[4][11] ),
    .A1(\po_0.regf_0.rf[5][11] ),
    .A2(\po_0.regf_0.rf[6][11] ),
    .A3(\po_0.regf_0.rf[7][11] ),
    .S0(_0451_),
    .S1(_0452_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _2048_ (.A0(_0563_),
    .A1(_0564_),
    .S(_0499_),
    .X(_0565_));
 sky130_fd_sc_hd__o22a_1 _2049_ (.A1(_0560_),
    .A2(_0562_),
    .B1(_0443_),
    .B2(_0565_),
    .X(\po_0.regf_0._3_[11] ));
 sky130_fd_sc_hd__mux4_1 _2050_ (.A0(\po_0.regf_0.rf[12][12] ),
    .A1(\po_0.regf_0.rf[13][12] ),
    .A2(\po_0.regf_0.rf[14][12] ),
    .A3(\po_0.regf_0.rf[15][12] ),
    .S0(_0488_),
    .S1(_0489_),
    .X(_0566_));
 sky130_fd_sc_hd__a21bo_1 _2051_ (.A1(_0566_),
    .A2(_0530_),
    .B1_N(_0003_),
    .X(_0567_));
 sky130_fd_sc_hd__mux4_1 _2052_ (.A0(\po_0.regf_0.rf[8][12] ),
    .A1(\po_0.regf_0.rf[9][12] ),
    .A2(\po_0.regf_0.rf[10][12] ),
    .A3(\po_0.regf_0.rf[11][12] ),
    .S0(_0472_),
    .S1(_0473_),
    .X(_0568_));
 sky130_fd_sc_hd__and2b_1 _2053_ (.A_N(_0450_),
    .B(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__mux4_1 _2054_ (.A0(\po_0.regf_0.rf[0][12] ),
    .A1(\po_0.regf_0.rf[1][12] ),
    .A2(\po_0.regf_0.rf[2][12] ),
    .A3(\po_0.regf_0.rf[3][12] ),
    .S0(_0524_),
    .S1(_0525_),
    .X(_0570_));
 sky130_fd_sc_hd__mux4_1 _2055_ (.A0(\po_0.regf_0.rf[4][12] ),
    .A1(\po_0.regf_0.rf[5][12] ),
    .A2(\po_0.regf_0.rf[6][12] ),
    .A3(\po_0.regf_0.rf[7][12] ),
    .S0(_0451_),
    .S1(_0452_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _2056_ (.A0(_0570_),
    .A1(_0571_),
    .S(_0438_),
    .X(_0572_));
 sky130_fd_sc_hd__o22a_1 _2057_ (.A1(_0567_),
    .A2(_0569_),
    .B1(_0443_),
    .B2(_0572_),
    .X(\po_0.regf_0._3_[12] ));
 sky130_fd_sc_hd__mux4_1 _2058_ (.A0(\po_0.regf_0.rf[0][13] ),
    .A1(\po_0.regf_0.rf[1][13] ),
    .A2(\po_0.regf_0.rf[2][13] ),
    .A3(\po_0.regf_0.rf[3][13] ),
    .S0(_0451_),
    .S1(_0452_),
    .X(_0573_));
 sky130_fd_sc_hd__mux4_1 _2059_ (.A0(\po_0.regf_0.rf[4][13] ),
    .A1(\po_0.regf_0.rf[5][13] ),
    .A2(\po_0.regf_0.rf[6][13] ),
    .A3(\po_0.regf_0.rf[7][13] ),
    .S0(_0439_),
    .S1(_0440_),
    .X(_0574_));
 sky130_fd_sc_hd__mux4_1 _2060_ (.A0(\po_0.regf_0.rf[8][13] ),
    .A1(\po_0.regf_0.rf[9][13] ),
    .A2(\po_0.regf_0.rf[10][13] ),
    .A3(\po_0.regf_0.rf[11][13] ),
    .S0(_0439_),
    .S1(_0440_),
    .X(_0575_));
 sky130_fd_sc_hd__mux4_1 _2061_ (.A0(\po_0.regf_0.rf[12][13] ),
    .A1(\po_0.regf_0.rf[13][13] ),
    .A2(\po_0.regf_0.rf[14][13] ),
    .A3(\po_0.regf_0.rf[15][13] ),
    .S0(_0439_),
    .S1(_0440_),
    .X(_0576_));
 sky130_fd_sc_hd__mux4_1 _2062_ (.A0(_0573_),
    .A1(_0574_),
    .A2(_0575_),
    .A3(_0576_),
    .S0(_0438_),
    .S1(_0470_),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_1 _2063_ (.A(_0577_),
    .X(\po_0.regf_0._3_[13] ));
 sky130_fd_sc_hd__mux4_1 _2064_ (.A0(\po_0.regf_0.rf[8][14] ),
    .A1(\po_0.regf_0.rf[9][14] ),
    .A2(\po_0.regf_0.rf[10][14] ),
    .A3(\po_0.regf_0.rf[11][14] ),
    .S0(_0472_),
    .S1(_0473_),
    .X(_0578_));
 sky130_fd_sc_hd__and2b_1 _2065_ (.A_N(_0450_),
    .B(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__mux4_1 _2066_ (.A0(\po_0.regf_0.rf[12][14] ),
    .A1(\po_0.regf_0.rf[13][14] ),
    .A2(\po_0.regf_0.rf[14][14] ),
    .A3(\po_0.regf_0.rf[15][14] ),
    .S0(_0479_),
    .S1(_0480_),
    .X(_0580_));
 sky130_fd_sc_hd__a21bo_1 _2067_ (.A1(_0580_),
    .A2(_0487_),
    .B1_N(_0463_),
    .X(_0581_));
 sky130_fd_sc_hd__mux4_1 _2068_ (.A0(\po_0.regf_0.rf[0][14] ),
    .A1(\po_0.regf_0.rf[1][14] ),
    .A2(\po_0.regf_0.rf[2][14] ),
    .A3(\po_0.regf_0.rf[3][14] ),
    .S0(_0466_),
    .S1(_0467_),
    .X(_0582_));
 sky130_fd_sc_hd__and2b_1 _2069_ (.A_N(_0465_),
    .B(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__mux4_1 _2070_ (.A0(\po_0.regf_0.rf[4][14] ),
    .A1(\po_0.regf_0.rf[5][14] ),
    .A2(\po_0.regf_0.rf[6][14] ),
    .A3(\po_0.regf_0.rf[7][14] ),
    .S0(_0444_),
    .S1(_0445_),
    .X(_0584_));
 sky130_fd_sc_hd__a21o_1 _2071_ (.A1(_0584_),
    .A2(_0447_),
    .B1(_0470_),
    .X(_0585_));
 sky130_fd_sc_hd__o22a_1 _2072_ (.A1(_0579_),
    .A2(_0581_),
    .B1(_0583_),
    .B2(_0585_),
    .X(\po_0.regf_0._3_[14] ));
 sky130_fd_sc_hd__mux4_1 _2073_ (.A0(\po_0.regf_0.rf[12][15] ),
    .A1(\po_0.regf_0.rf[13][15] ),
    .A2(\po_0.regf_0.rf[14][15] ),
    .A3(\po_0.regf_0.rf[15][15] ),
    .S0(_0488_),
    .S1(_0489_),
    .X(_0586_));
 sky130_fd_sc_hd__a21bo_1 _2074_ (.A1(_0586_),
    .A2(_0530_),
    .B1_N(_0003_),
    .X(_0587_));
 sky130_fd_sc_hd__mux4_1 _2075_ (.A0(\po_0.regf_0.rf[8][15] ),
    .A1(\po_0.regf_0.rf[9][15] ),
    .A2(\po_0.regf_0.rf[10][15] ),
    .A3(\po_0.regf_0.rf[11][15] ),
    .S0(_0472_),
    .S1(_0473_),
    .X(_0588_));
 sky130_fd_sc_hd__and2b_1 _2076_ (.A_N(_0450_),
    .B(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__mux4_1 _2077_ (.A0(\po_0.regf_0.rf[0][15] ),
    .A1(\po_0.regf_0.rf[1][15] ),
    .A2(\po_0.regf_0.rf[2][15] ),
    .A3(\po_0.regf_0.rf[3][15] ),
    .S0(_0475_),
    .S1(_0476_),
    .X(_0590_));
 sky130_fd_sc_hd__mux4_1 _2078_ (.A0(\po_0.regf_0.rf[4][15] ),
    .A1(\po_0.regf_0.rf[5][15] ),
    .A2(\po_0.regf_0.rf[6][15] ),
    .A3(\po_0.regf_0.rf[7][15] ),
    .S0(_0451_),
    .S1(_0452_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _2079_ (.A0(_0590_),
    .A1(_0591_),
    .S(_0438_),
    .X(_0592_));
 sky130_fd_sc_hd__o22a_1 _2080_ (.A1(_0587_),
    .A2(_0589_),
    .B1(_0443_),
    .B2(_0592_),
    .X(\po_0.regf_0._3_[15] ));
 sky130_fd_sc_hd__and3_1 _2081_ (.A(_1533_),
    .B(_1534_),
    .C(_1537_),
    .X(_0593_));
 sky130_fd_sc_hd__or2_1 _2082_ (.A(\uc_0.bc_0._70_[2] ),
    .B(\uc_0.bc_0._70_[3] ),
    .X(_0594_));
 sky130_fd_sc_hd__a31o_2 _2083_ (.A1(_0593_),
    .A2(\uc_0.bc_0._70_[0] ),
    .A3(_0594_),
    .B1(_1552_),
    .X(_0595_));
 sky130_fd_sc_hd__buf_2 _2084_ (.A(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _2085_ (.A0(\po_0.regf_0.rp_addr[0] ),
    .A1(\uc_0._21_[8] ),
    .S(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__clkbuf_1 _2086_ (.A(_0597_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _2087_ (.A0(\po_0.regf_0.rp_addr[1] ),
    .A1(\uc_0._21_[9] ),
    .S(_0596_),
    .X(_0598_));
 sky130_fd_sc_hd__clkbuf_1 _2088_ (.A(_0598_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _2089_ (.A0(\po_0.regf_0.rp_addr[2] ),
    .A1(\uc_0._21_[10] ),
    .S(_0596_),
    .X(_0599_));
 sky130_fd_sc_hd__clkbuf_1 _2090_ (.A(_0599_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _2091_ (.A0(\po_0.regf_0.rp_addr[3] ),
    .A1(\uc_0._21_[11] ),
    .S(_0596_),
    .X(_0600_));
 sky130_fd_sc_hd__clkbuf_1 _2092_ (.A(_0600_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _2093_ (.A(_1535_),
    .B(_1541_),
    .X(_0601_));
 sky130_fd_sc_hd__a21bo_1 _2094_ (.A1(_0601_),
    .A2(_1542_),
    .B1_N(_1539_),
    .X(net79));
 sky130_fd_sc_hd__a21o_1 _2095_ (.A1(_1542_),
    .A2(_0601_),
    .B1(_1536_),
    .X(net80));
 sky130_fd_sc_hd__and4b_1 _2096_ (.A_N(_1542_),
    .B(_1541_),
    .C(_1535_),
    .D(_1539_),
    .X(_0602_));
 sky130_fd_sc_hd__a21oi_1 _2097_ (.A1(_1539_),
    .A2(_1535_),
    .B1(_1541_),
    .Y(_0603_));
 sky130_fd_sc_hd__nor2_2 _2098_ (.A(_0602_),
    .B(_0603_),
    .Y(net81));
 sky130_fd_sc_hd__a31o_1 _2099_ (.A1(_1539_),
    .A2(_1535_),
    .A3(_1541_),
    .B1(_1542_),
    .X(net82));
 sky130_fd_sc_hd__and2b_1 _2100_ (.A_N(_1513_),
    .B(\po_0._1_[0] ),
    .X(_0604_));
 sky130_fd_sc_hd__and2_1 _2101_ (.A(net87),
    .B(\po_0._1_[1] ),
    .X(_0605_));
 sky130_fd_sc_hd__nor2_1 _2102_ (.A(net87),
    .B(\po_0._1_[1] ),
    .Y(_0606_));
 sky130_fd_sc_hd__nor2_1 _2103_ (.A(_0605_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__xor2_1 _2104_ (.A(_0604_),
    .B(_0607_),
    .X(\po_0.alu_0._10_[1] ));
 sky130_fd_sc_hd__and2_1 _2105_ (.A(_1524_),
    .B(\po_0._1_[2] ),
    .X(_0608_));
 sky130_fd_sc_hd__nor2_1 _2106_ (.A(_1524_),
    .B(\po_0._1_[2] ),
    .Y(_0609_));
 sky130_fd_sc_hd__inv_2 _2107_ (.A(net87),
    .Y(_0610_));
 sky130_fd_sc_hd__nand2_1 _2108_ (.A(_0610_),
    .B(\po_0._1_[1] ),
    .Y(_0611_));
 sky130_fd_sc_hd__o21ai_1 _2109_ (.A1(\po_0._1_[1] ),
    .A2(_0610_),
    .B1(_0604_),
    .Y(_0612_));
 sky130_fd_sc_hd__o211ai_1 _2110_ (.A1(_0608_),
    .A2(_0609_),
    .B1(_0611_),
    .C1(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__or2b_1 _2111_ (.A(net43),
    .B_N(\po_0._1_[2] ),
    .X(_0614_));
 sky130_fd_sc_hd__or2b_1 _2112_ (.A(\po_0._1_[2] ),
    .B_N(net43),
    .X(_0615_));
 sky130_fd_sc_hd__a22o_1 _2113_ (.A1(_0614_),
    .A2(_0615_),
    .B1(_0611_),
    .B2(_0612_),
    .X(_0616_));
 sky130_fd_sc_hd__and2_1 _2114_ (.A(_0613_),
    .B(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__clkbuf_1 _2115_ (.A(_0617_),
    .X(\po_0.alu_0._10_[2] ));
 sky130_fd_sc_hd__clkbuf_2 _2116_ (.A(\po_0._1_[3] ),
    .X(_0618_));
 sky130_fd_sc_hd__and2_1 _2117_ (.A(net44),
    .B(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__clkbuf_2 _2118_ (.A(net44),
    .X(_0620_));
 sky130_fd_sc_hd__nor2_1 _2119_ (.A(_0620_),
    .B(_0618_),
    .Y(_0621_));
 sky130_fd_sc_hd__o2bb2ai_1 _2120_ (.A1_N(_0615_),
    .A2_N(_0613_),
    .B1(_0619_),
    .B2(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__nand2_1 _2121_ (.A(_0614_),
    .B(_0615_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand2_1 _2122_ (.A(_0611_),
    .B(_0612_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _2123_ (.A(_0620_),
    .B(_0618_),
    .Y(_0625_));
 sky130_fd_sc_hd__or2_2 _2124_ (.A(net44),
    .B(\po_0._1_[3] ),
    .X(_0626_));
 sky130_fd_sc_hd__o2111ai_1 _2125_ (.A1(_0623_),
    .A2(_0624_),
    .B1(_0625_),
    .C1(_0626_),
    .D1(_0615_),
    .Y(_0627_));
 sky130_fd_sc_hd__and2_1 _2126_ (.A(_0622_),
    .B(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__clkbuf_1 _2127_ (.A(_0628_),
    .X(\po_0.alu_0._10_[3] ));
 sky130_fd_sc_hd__clkbuf_2 _2128_ (.A(net45),
    .X(_0629_));
 sky130_fd_sc_hd__clkbuf_2 _2129_ (.A(\po_0._1_[4] ),
    .X(_0630_));
 sky130_fd_sc_hd__and2_1 _2130_ (.A(_0629_),
    .B(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__nor2_1 _2131_ (.A(_0629_),
    .B(_0630_),
    .Y(_0632_));
 sky130_fd_sc_hd__or2b_1 _2132_ (.A(_0618_),
    .B_N(_0620_),
    .X(_0633_));
 sky130_fd_sc_hd__a2bb2oi_2 _2133_ (.A1_N(_0631_),
    .A2_N(_0632_),
    .B1(_0633_),
    .B2(_0622_),
    .Y(_0634_));
 sky130_fd_sc_hd__nand2_2 _2134_ (.A(_0629_),
    .B(_0630_),
    .Y(_0635_));
 sky130_fd_sc_hd__or2_1 _2135_ (.A(net45),
    .B(\po_0._1_[4] ),
    .X(_0636_));
 sky130_fd_sc_hd__nand4_1 _2136_ (.A(_0622_),
    .B(_0635_),
    .C(_0636_),
    .D(_0633_),
    .Y(_0637_));
 sky130_fd_sc_hd__and2b_1 _2137_ (.A_N(_0634_),
    .B(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__clkbuf_1 _2138_ (.A(_0638_),
    .X(\po_0.alu_0._10_[4] ));
 sky130_fd_sc_hd__and2b_1 _2139_ (.A_N(_0630_),
    .B(_0629_),
    .X(_0639_));
 sky130_fd_sc_hd__clkbuf_2 _2140_ (.A(net46),
    .X(_0640_));
 sky130_fd_sc_hd__clkbuf_2 _2141_ (.A(\po_0._1_[5] ),
    .X(_0641_));
 sky130_fd_sc_hd__nand2_1 _2142_ (.A(_0640_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__or2_2 _2143_ (.A(net46),
    .B(\po_0._1_[5] ),
    .X(_0643_));
 sky130_fd_sc_hd__o211a_1 _2144_ (.A1(_0634_),
    .A2(_0639_),
    .B1(_0642_),
    .C1(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__a211oi_1 _2145_ (.A1(_0643_),
    .A2(_0642_),
    .B1(_0639_),
    .C1(_0634_),
    .Y(_0645_));
 sky130_fd_sc_hd__or2_1 _2146_ (.A(_0644_),
    .B(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__clkbuf_1 _2147_ (.A(_0646_),
    .X(\po_0.alu_0._10_[5] ));
 sky130_fd_sc_hd__and2_1 _2148_ (.A(_1526_),
    .B(\po_0._1_[6] ),
    .X(_0647_));
 sky130_fd_sc_hd__nor2_1 _2149_ (.A(_1526_),
    .B(\po_0._1_[6] ),
    .Y(_0648_));
 sky130_fd_sc_hd__or2b_1 _2150_ (.A(_0641_),
    .B_N(_0640_),
    .X(_0649_));
 sky130_fd_sc_hd__nor2_1 _2151_ (.A(_0640_),
    .B(_0641_),
    .Y(_0650_));
 sky130_fd_sc_hd__and2_1 _2152_ (.A(_0640_),
    .B(_0641_),
    .X(_0651_));
 sky130_fd_sc_hd__o22ai_1 _2153_ (.A1(_0650_),
    .A2(_0651_),
    .B1(_0639_),
    .B2(_0634_),
    .Y(_0652_));
 sky130_fd_sc_hd__a2bb2oi_1 _2154_ (.A1_N(_0647_),
    .A2_N(_0648_),
    .B1(_0649_),
    .B2(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__nand2_1 _2155_ (.A(_1526_),
    .B(\po_0._1_[6] ),
    .Y(_0654_));
 sky130_fd_sc_hd__or2_1 _2156_ (.A(net47),
    .B(\po_0._1_[6] ),
    .X(_0655_));
 sky130_fd_sc_hd__nand4_1 _2157_ (.A(_0652_),
    .B(_0654_),
    .C(_0655_),
    .D(_0649_),
    .Y(_0656_));
 sky130_fd_sc_hd__and2b_1 _2158_ (.A_N(_0653_),
    .B(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__clkbuf_1 _2159_ (.A(_0657_),
    .X(\po_0.alu_0._10_[6] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2160_ (.A(net48),
    .X(_0658_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2161_ (.A(\po_0._1_[7] ),
    .X(_0659_));
 sky130_fd_sc_hd__nor2_1 _2162_ (.A(_0658_),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__and2_1 _2163_ (.A(_0658_),
    .B(_0659_),
    .X(_0661_));
 sky130_fd_sc_hd__and2b_1 _2164_ (.A_N(\po_0._1_[6] ),
    .B(_1526_),
    .X(_0662_));
 sky130_fd_sc_hd__o22ai_2 _2165_ (.A1(_0660_),
    .A2(_0661_),
    .B1(_0662_),
    .B2(_0653_),
    .Y(_0663_));
 sky130_fd_sc_hd__or4_1 _2166_ (.A(_0653_),
    .B(_0660_),
    .C(_0661_),
    .D(_0662_),
    .X(_0664_));
 sky130_fd_sc_hd__and2_1 _2167_ (.A(_0663_),
    .B(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__clkbuf_1 _2168_ (.A(_0665_),
    .X(\po_0.alu_0._10_[7] ));
 sky130_fd_sc_hd__and2_1 _2169_ (.A(net86),
    .B(\po_0._1_[8] ),
    .X(_0666_));
 sky130_fd_sc_hd__nor2_1 _2170_ (.A(net86),
    .B(\po_0._1_[8] ),
    .Y(_0667_));
 sky130_fd_sc_hd__or2_2 _2171_ (.A(_0666_),
    .B(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__or2b_1 _2172_ (.A(_0659_),
    .B_N(_0658_),
    .X(_0669_));
 sky130_fd_sc_hd__nand2_1 _2173_ (.A(_0663_),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__xor2_1 _2174_ (.A(_0668_),
    .B(_0670_),
    .X(\po_0.alu_0._10_[8] ));
 sky130_fd_sc_hd__clkbuf_2 _2175_ (.A(net50),
    .X(_0671_));
 sky130_fd_sc_hd__xor2_1 _2176_ (.A(_0671_),
    .B(\po_0._1_[9] ),
    .X(_0672_));
 sky130_fd_sc_hd__clkbuf_2 _2177_ (.A(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__inv_2 _2178_ (.A(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__or2b_1 _2179_ (.A(\po_0._1_[8] ),
    .B_N(net86),
    .X(_0675_));
 sky130_fd_sc_hd__a21bo_1 _2180_ (.A1(_0668_),
    .A2(_0670_),
    .B1_N(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__xor2_1 _2181_ (.A(_0674_),
    .B(_0676_),
    .X(\po_0.alu_0._10_[9] ));
 sky130_fd_sc_hd__or2b_1 _2182_ (.A(\po_0._1_[10] ),
    .B_N(_1522_),
    .X(_0677_));
 sky130_fd_sc_hd__or2b_1 _2183_ (.A(net36),
    .B_N(\po_0._1_[10] ),
    .X(_0678_));
 sky130_fd_sc_hd__nand2_2 _2184_ (.A(_0677_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__or2b_1 _2185_ (.A(\po_0._1_[9] ),
    .B_N(_0671_),
    .X(_0680_));
 sky130_fd_sc_hd__o211ai_1 _2186_ (.A1(_0666_),
    .A2(_0667_),
    .B1(_0670_),
    .C1(_0674_),
    .Y(_0681_));
 sky130_fd_sc_hd__o211a_1 _2187_ (.A1(_0673_),
    .A2(_0675_),
    .B1(_0680_),
    .C1(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__xor2_1 _2188_ (.A(_0679_),
    .B(_0682_),
    .X(\po_0.alu_0._10_[10] ));
 sky130_fd_sc_hd__nor2_2 _2189_ (.A(net85),
    .B(\po_0._1_[11] ),
    .Y(_0683_));
 sky130_fd_sc_hd__and2_1 _2190_ (.A(net85),
    .B(\po_0._1_[11] ),
    .X(_0684_));
 sky130_fd_sc_hd__nor2_2 _2191_ (.A(_0683_),
    .B(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__o211a_1 _2192_ (.A1(_0675_),
    .A2(_0673_),
    .B1(_0680_),
    .C1(_0677_),
    .X(_0686_));
 sky130_fd_sc_hd__and2b_1 _2193_ (.A_N(_1522_),
    .B(\po_0._1_[10] ),
    .X(_0687_));
 sky130_fd_sc_hd__a21oi_1 _2194_ (.A1(_0681_),
    .A2(_0686_),
    .B1(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__xnor2_1 _2195_ (.A(_0685_),
    .B(_0688_),
    .Y(\po_0.alu_0._10_[11] ));
 sky130_fd_sc_hd__and2_1 _2196_ (.A(net84),
    .B(\po_0._1_[12] ),
    .X(_0689_));
 sky130_fd_sc_hd__nor2_1 _2197_ (.A(net84),
    .B(\po_0._1_[12] ),
    .Y(_0690_));
 sky130_fd_sc_hd__nor2_1 _2198_ (.A(_0689_),
    .B(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__clkbuf_2 _2199_ (.A(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__inv_2 _2200_ (.A(net85),
    .Y(_0693_));
 sky130_fd_sc_hd__o32ai_2 _2201_ (.A1(_0687_),
    .A2(_0685_),
    .A3(_0686_),
    .B1(\po_0._1_[11] ),
    .B2(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__nor2_1 _2202_ (.A(_0666_),
    .B(_0667_),
    .Y(_0695_));
 sky130_fd_sc_hd__or4_1 _2203_ (.A(_0695_),
    .B(_0673_),
    .C(_0679_),
    .D(_0685_),
    .X(_0696_));
 sky130_fd_sc_hd__a21oi_1 _2204_ (.A1(_0663_),
    .A2(_0669_),
    .B1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__or2_1 _2205_ (.A(_0694_),
    .B(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__xnor2_1 _2206_ (.A(_0692_),
    .B(_0698_),
    .Y(\po_0.alu_0._10_[12] ));
 sky130_fd_sc_hd__o21ai_1 _2207_ (.A1(_0689_),
    .A2(_0690_),
    .B1(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__xor2_1 _2208_ (.A(net83),
    .B(\po_0._1_[13] ),
    .X(_0700_));
 sky130_fd_sc_hd__clkbuf_2 _2209_ (.A(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__or2b_1 _2210_ (.A(\po_0._1_[12] ),
    .B_N(net84),
    .X(_0702_));
 sky130_fd_sc_hd__and2_1 _2211_ (.A(_0701_),
    .B(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__or2_1 _2212_ (.A(_0692_),
    .B(_0701_),
    .X(_0704_));
 sky130_fd_sc_hd__o21bai_2 _2213_ (.A1(_0694_),
    .A2(_0697_),
    .B1_N(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__o21ai_1 _2214_ (.A1(_0701_),
    .A2(_0702_),
    .B1(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__a21oi_1 _2215_ (.A1(_0699_),
    .A2(_0703_),
    .B1(_0706_),
    .Y(\po_0.alu_0._10_[13] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2216_ (.A(net40),
    .X(_0707_));
 sky130_fd_sc_hd__nand2_1 _2217_ (.A(_0707_),
    .B(\po_0._1_[14] ),
    .Y(_0708_));
 sky130_fd_sc_hd__or2_1 _2218_ (.A(net40),
    .B(\po_0._1_[14] ),
    .X(_0709_));
 sky130_fd_sc_hd__or2b_1 _2219_ (.A(\po_0._1_[13] ),
    .B_N(net83),
    .X(_0710_));
 sky130_fd_sc_hd__o21a_1 _2220_ (.A1(_0702_),
    .A2(_0701_),
    .B1(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__a22oi_1 _2221_ (.A1(_0708_),
    .A2(_0709_),
    .B1(_0705_),
    .B2(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__and4_1 _2222_ (.A(_0705_),
    .B(_0708_),
    .C(_0709_),
    .D(_0711_),
    .X(_0713_));
 sky130_fd_sc_hd__nor2_1 _2223_ (.A(_0712_),
    .B(_0713_),
    .Y(\po_0.alu_0._10_[14] ));
 sky130_fd_sc_hd__and2b_1 _2224_ (.A_N(\po_0._1_[15] ),
    .B(net41),
    .X(_0714_));
 sky130_fd_sc_hd__and2b_1 _2225_ (.A_N(net41),
    .B(\po_0._1_[15] ),
    .X(_0715_));
 sky130_fd_sc_hd__or2_1 _2226_ (.A(_0714_),
    .B(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__or2b_1 _2227_ (.A(\po_0._1_[14] ),
    .B_N(_0707_),
    .X(_0717_));
 sky130_fd_sc_hd__and2_1 _2228_ (.A(_0707_),
    .B(\po_0._1_[14] ),
    .X(_0718_));
 sky130_fd_sc_hd__nor2_1 _2229_ (.A(_0707_),
    .B(\po_0._1_[14] ),
    .Y(_0719_));
 sky130_fd_sc_hd__o2bb2ai_1 _2230_ (.A1_N(_0711_),
    .A2_N(_0705_),
    .B1(_0718_),
    .B2(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__nand3b_1 _2231_ (.A_N(_0716_),
    .B(_0717_),
    .C(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__and2b_1 _2232_ (.A_N(\po_0._1_[14] ),
    .B(_0707_),
    .X(_0722_));
 sky130_fd_sc_hd__o22ai_1 _2233_ (.A1(_0714_),
    .A2(_0715_),
    .B1(_0722_),
    .B2(_0712_),
    .Y(_0723_));
 sky130_fd_sc_hd__nand2_1 _2234_ (.A(_0721_),
    .B(_0723_),
    .Y(\po_0.alu_0._10_[15] ));
 sky130_fd_sc_hd__and2b_1 _2235_ (.A_N(\po_0.muxf_0.s0 ),
    .B(\po_0.muxf_0.s1 ),
    .X(_0724_));
 sky130_fd_sc_hd__buf_2 _2236_ (.A(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__and2b_1 _2237_ (.A_N(\po_0.muxf_0.s1 ),
    .B(\po_0.muxf_0.s0 ),
    .X(_0726_));
 sky130_fd_sc_hd__clkbuf_2 _2238_ (.A(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__buf_2 _2239_ (.A(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__buf_2 _2240_ (.A(\po_0.alu_0.s1 ),
    .X(_0729_));
 sky130_fd_sc_hd__nand2_1 _2241_ (.A(_1490_),
    .B(\po_0.alu_0.s0 ),
    .Y(_0730_));
 sky130_fd_sc_hd__buf_2 _2242_ (.A(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__nor2_2 _2243_ (.A(_0724_),
    .B(_0726_),
    .Y(_0732_));
 sky130_fd_sc_hd__o221a_1 _2244_ (.A1(_1491_),
    .A2(\po_0.alu_0._11_[0] ),
    .B1(_0731_),
    .B2(\po_0.alu_0._10_[0] ),
    .C1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__o31a_1 _2245_ (.A1(_1513_),
    .A2(_0729_),
    .A3(_1488_),
    .B1(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__a221o_2 _2246_ (.A1(\po_0.muxf_0.rf_w_data[0] ),
    .A2(_0725_),
    .B1(_0728_),
    .B2(net1),
    .C1(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2247_ (.A(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2248_ (.A(\po_0.regf_0.w_addr[3] ),
    .X(_0737_));
 sky130_fd_sc_hd__clkbuf_2 _2249_ (.A(\po_0.regf_0.w_wr ),
    .X(_0738_));
 sky130_fd_sc_hd__clkbuf_2 _2250_ (.A(\po_0.regf_0.w_addr[1] ),
    .X(_0739_));
 sky130_fd_sc_hd__clkbuf_2 _2251_ (.A(\po_0.regf_0.w_addr[0] ),
    .X(_0740_));
 sky130_fd_sc_hd__and2b_1 _2252_ (.A_N(_0739_),
    .B(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2253_ (.A(\po_0.regf_0.w_addr[2] ),
    .X(_0742_));
 sky130_fd_sc_hd__and4b_4 _2254_ (.A_N(_0737_),
    .B(_0738_),
    .C(_0741_),
    .D(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__buf_2 _2255_ (.A(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_1 _2256_ (.A0(\po_0.regf_0.rf[5][0] ),
    .A1(_0736_),
    .S(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__clkbuf_1 _2257_ (.A(_0745_),
    .X(_0016_));
 sky130_fd_sc_hd__nor2_2 _2258_ (.A(\po_0.alu_0.s1 ),
    .B(_1487_),
    .Y(_0746_));
 sky130_fd_sc_hd__clkbuf_2 _2259_ (.A(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__and2_2 _2260_ (.A(_1490_),
    .B(_1487_),
    .X(_0748_));
 sky130_fd_sc_hd__a2bb2o_1 _2261_ (.A1_N(_0605_),
    .A2_N(_0606_),
    .B1(\po_0._1_[0] ),
    .B2(_1513_),
    .X(_0749_));
 sky130_fd_sc_hd__o311a_1 _2262_ (.A1(_1515_),
    .A2(_0605_),
    .A3(_0606_),
    .B1(_0748_),
    .C1(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__a221o_1 _2263_ (.A1(_0729_),
    .A2(\po_0.alu_0._11_[1] ),
    .B1(_0747_),
    .B2(net87),
    .C1(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__clkbuf_2 _2264_ (.A(_0732_),
    .X(_0752_));
 sky130_fd_sc_hd__clkbuf_2 _2265_ (.A(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__a22o_1 _2266_ (.A1(\po_0.muxf_0.rf_w_data[1] ),
    .A2(_0725_),
    .B1(_0727_),
    .B2(net8),
    .X(_0754_));
 sky130_fd_sc_hd__a21o_2 _2267_ (.A1(_0751_),
    .A2(_0753_),
    .B1(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2268_ (.A(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_1 _2269_ (.A0(\po_0.regf_0.rf[5][1] ),
    .A1(_0756_),
    .S(_0744_),
    .X(_0757_));
 sky130_fd_sc_hd__clkbuf_1 _2270_ (.A(_0757_),
    .X(_0017_));
 sky130_fd_sc_hd__a311o_1 _2271_ (.A1(\po_0._1_[0] ),
    .A2(_1513_),
    .A3(_0607_),
    .B1(_0623_),
    .C1(_0605_),
    .X(_0758_));
 sky130_fd_sc_hd__nand2_1 _2272_ (.A(net87),
    .B(\po_0._1_[1] ),
    .Y(_0759_));
 sky130_fd_sc_hd__o21ai_1 _2273_ (.A1(_1515_),
    .A2(_0606_),
    .B1(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__or3b_1 _2274_ (.A(_0608_),
    .B(_0609_),
    .C_N(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__buf_2 _2275_ (.A(_0748_),
    .X(_0762_));
 sky130_fd_sc_hd__clkbuf_2 _2276_ (.A(\po_0.alu_0.s1 ),
    .X(_0763_));
 sky130_fd_sc_hd__a22o_1 _2277_ (.A1(_0763_),
    .A2(\po_0.alu_0._11_[2] ),
    .B1(_0747_),
    .B2(_1524_),
    .X(_0764_));
 sky130_fd_sc_hd__a31o_1 _2278_ (.A1(_0758_),
    .A2(_0761_),
    .A3(_0762_),
    .B1(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__a22o_1 _2279_ (.A1(\po_0.muxf_0.rf_w_data[2] ),
    .A2(_0724_),
    .B1(_0727_),
    .B2(net9),
    .X(_0766_));
 sky130_fd_sc_hd__a21o_2 _2280_ (.A1(_0765_),
    .A2(_0753_),
    .B1(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__clkbuf_2 _2281_ (.A(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__mux2_1 _2282_ (.A0(\po_0.regf_0.rf[5][2] ),
    .A1(_0768_),
    .S(_0744_),
    .X(_0769_));
 sky130_fd_sc_hd__clkbuf_1 _2283_ (.A(_0769_),
    .X(_0018_));
 sky130_fd_sc_hd__nand2_1 _2284_ (.A(_1524_),
    .B(\po_0._1_[2] ),
    .Y(_0770_));
 sky130_fd_sc_hd__a211oi_1 _2285_ (.A1(_0770_),
    .A2(_0761_),
    .B1(_0621_),
    .C1(_0619_),
    .Y(_0771_));
 sky130_fd_sc_hd__o211a_1 _2286_ (.A1(_0619_),
    .A2(_0621_),
    .B1(_0761_),
    .C1(_0770_),
    .X(_0772_));
 sky130_fd_sc_hd__clkbuf_2 _2287_ (.A(\po_0.alu_0.s1 ),
    .X(_0773_));
 sky130_fd_sc_hd__a21oi_1 _2288_ (.A1(_0773_),
    .A2(\po_0.alu_0._11_[3] ),
    .B1(_0746_),
    .Y(_0774_));
 sky130_fd_sc_hd__o31ai_1 _2289_ (.A1(_0731_),
    .A2(_0771_),
    .A3(_0772_),
    .B1(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__o311a_1 _2290_ (.A1(_0620_),
    .A2(_0729_),
    .A3(_1488_),
    .B1(_0732_),
    .C1(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__a221o_2 _2291_ (.A1(\po_0.muxf_0.rf_w_data[3] ),
    .A2(_0725_),
    .B1(_0728_),
    .B2(net10),
    .C1(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2292_ (.A(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_1 _2293_ (.A0(\po_0.regf_0.rf[5][3] ),
    .A1(_0778_),
    .S(_0744_),
    .X(_0779_));
 sky130_fd_sc_hd__clkbuf_1 _2294_ (.A(_0779_),
    .X(_0019_));
 sky130_fd_sc_hd__nor2_1 _2295_ (.A(_0631_),
    .B(_0632_),
    .Y(_0780_));
 sky130_fd_sc_hd__a22o_1 _2296_ (.A1(_1524_),
    .A2(\po_0._1_[2] ),
    .B1(\po_0._1_[3] ),
    .B2(net44),
    .X(_0781_));
 sky130_fd_sc_hd__a21o_2 _2297_ (.A1(_0623_),
    .A2(_0760_),
    .B1(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__o21a_1 _2298_ (.A1(_0620_),
    .A2(_0618_),
    .B1(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__o2111ai_4 _2299_ (.A1(_0620_),
    .A2(_0618_),
    .B1(_0635_),
    .C1(_0636_),
    .D1(_0782_),
    .Y(_0784_));
 sky130_fd_sc_hd__o211a_1 _2300_ (.A1(_0780_),
    .A2(_0783_),
    .B1(_0784_),
    .C1(_0748_),
    .X(_0785_));
 sky130_fd_sc_hd__a221o_1 _2301_ (.A1(_0729_),
    .A2(\po_0.alu_0._11_[4] ),
    .B1(_0747_),
    .B2(_0629_),
    .C1(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__a22o_1 _2302_ (.A1(\po_0.muxf_0.rf_w_data[4] ),
    .A2(_0724_),
    .B1(_0727_),
    .B2(net11),
    .X(_0787_));
 sky130_fd_sc_hd__a21o_2 _2303_ (.A1(_0786_),
    .A2(_0753_),
    .B1(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__clkbuf_2 _2304_ (.A(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__mux2_1 _2305_ (.A0(\po_0.regf_0.rf[5][4] ),
    .A1(_0789_),
    .S(_0744_),
    .X(_0790_));
 sky130_fd_sc_hd__clkbuf_1 _2306_ (.A(_0790_),
    .X(_0020_));
 sky130_fd_sc_hd__a211o_1 _2307_ (.A1(_0635_),
    .A2(_0784_),
    .B1(_0651_),
    .C1(_0650_),
    .X(_0791_));
 sky130_fd_sc_hd__a221o_1 _2308_ (.A1(_0643_),
    .A2(_0642_),
    .B1(_0783_),
    .B2(_0780_),
    .C1(_0631_),
    .X(_0792_));
 sky130_fd_sc_hd__o21a_1 _2309_ (.A1(_1491_),
    .A2(\po_0.alu_0._11_[5] ),
    .B1(_0731_),
    .X(_0793_));
 sky130_fd_sc_hd__a31o_1 _2310_ (.A1(_0791_),
    .A2(_0748_),
    .A3(_0792_),
    .B1(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__o311a_1 _2311_ (.A1(_0640_),
    .A2(_0763_),
    .A3(_1488_),
    .B1(_0732_),
    .C1(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__a221o_4 _2312_ (.A1(\po_0.muxf_0.rf_w_data[5] ),
    .A2(_0725_),
    .B1(_0728_),
    .B2(net12),
    .C1(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2313_ (.A(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_1 _2314_ (.A0(\po_0.regf_0.rf[5][5] ),
    .A1(_0797_),
    .S(_0744_),
    .X(_0798_));
 sky130_fd_sc_hd__clkbuf_1 _2315_ (.A(_0798_),
    .X(_0021_));
 sky130_fd_sc_hd__a22o_1 _2316_ (.A1(_0773_),
    .A2(\po_0.alu_0._11_[6] ),
    .B1(_0746_),
    .B2(_1526_),
    .X(_0799_));
 sky130_fd_sc_hd__a21oi_1 _2317_ (.A1(_0629_),
    .A2(_0630_),
    .B1(_0651_),
    .Y(_0800_));
 sky130_fd_sc_hd__or3_1 _2318_ (.A(_0650_),
    .B(_0647_),
    .C(_0648_),
    .X(_0801_));
 sky130_fd_sc_hd__a21oi_1 _2319_ (.A1(_0784_),
    .A2(_0800_),
    .B1(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__a22o_1 _2320_ (.A1(net45),
    .A2(_0630_),
    .B1(_0641_),
    .B2(net46),
    .X(_0803_));
 sky130_fd_sc_hd__a31o_1 _2321_ (.A1(_0626_),
    .A2(_0782_),
    .A3(_0780_),
    .B1(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__a22o_1 _2322_ (.A1(_0654_),
    .A2(_0655_),
    .B1(_0804_),
    .B2(_0643_),
    .X(_0805_));
 sky130_fd_sc_hd__and3b_1 _2323_ (.A_N(_0802_),
    .B(_0748_),
    .C(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__o21a_1 _2324_ (.A1(_0799_),
    .A2(_0806_),
    .B1(_0752_),
    .X(_0807_));
 sky130_fd_sc_hd__a221o_2 _2325_ (.A1(\po_0.muxf_0.rf_w_data[6] ),
    .A2(_0725_),
    .B1(_0728_),
    .B2(net13),
    .C1(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2326_ (.A(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__buf_2 _2327_ (.A(_0743_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _2328_ (.A0(\po_0.regf_0.rf[5][6] ),
    .A1(_0809_),
    .S(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__clkbuf_1 _2329_ (.A(_0811_),
    .X(_0022_));
 sky130_fd_sc_hd__nor2_1 _2330_ (.A(_0660_),
    .B(_0661_),
    .Y(_0812_));
 sky130_fd_sc_hd__o31ai_1 _2331_ (.A1(_0647_),
    .A2(_0812_),
    .A3(_0802_),
    .B1(_0748_),
    .Y(_0813_));
 sky130_fd_sc_hd__nand2_1 _2332_ (.A(net48),
    .B(_0659_),
    .Y(_0814_));
 sky130_fd_sc_hd__or2_1 _2333_ (.A(net48),
    .B(\po_0._1_[7] ),
    .X(_0815_));
 sky130_fd_sc_hd__o211a_1 _2334_ (.A1(_0647_),
    .A2(_0802_),
    .B1(_0814_),
    .C1(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__o21ai_1 _2335_ (.A1(_1491_),
    .A2(\po_0.alu_0._11_[7] ),
    .B1(_0731_),
    .Y(_0817_));
 sky130_fd_sc_hd__o21ai_1 _2336_ (.A1(_0813_),
    .A2(_0816_),
    .B1(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__o311a_1 _2337_ (.A1(_0658_),
    .A2(_0763_),
    .A3(_1488_),
    .B1(_0732_),
    .C1(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__a221o_4 _2338_ (.A1(\po_0.muxf_0.rf_w_data[7] ),
    .A2(_0725_),
    .B1(_0727_),
    .B2(net14),
    .C1(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2339_ (.A(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__mux2_1 _2340_ (.A0(\po_0.regf_0.rf[5][7] ),
    .A1(_0821_),
    .S(_0810_),
    .X(_0822_));
 sky130_fd_sc_hd__clkbuf_1 _2341_ (.A(_0822_),
    .X(_0023_));
 sky130_fd_sc_hd__clkbuf_2 _2342_ (.A(_0727_),
    .X(_0823_));
 sky130_fd_sc_hd__nand4_1 _2343_ (.A(_0654_),
    .B(_0655_),
    .C(_0815_),
    .D(_0814_),
    .Y(_0824_));
 sky130_fd_sc_hd__nand4_1 _2344_ (.A(_0635_),
    .B(_0636_),
    .C(_0643_),
    .D(_0642_),
    .Y(_0825_));
 sky130_fd_sc_hd__nor2_1 _2345_ (.A(_0824_),
    .B(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__nand3_1 _2346_ (.A(_0826_),
    .B(_0782_),
    .C(_0626_),
    .Y(_0827_));
 sky130_fd_sc_hd__a21oi_1 _2347_ (.A1(_0658_),
    .A2(_0659_),
    .B1(_0647_),
    .Y(_0828_));
 sky130_fd_sc_hd__o2111ai_2 _2348_ (.A1(_0640_),
    .A2(_0641_),
    .B1(_0654_),
    .C1(_0655_),
    .D1(_0803_),
    .Y(_0829_));
 sky130_fd_sc_hd__a2bb2o_1 _2349_ (.A1_N(_0658_),
    .A2_N(_0659_),
    .B1(_0828_),
    .B2(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__a21oi_2 _2350_ (.A1(_0827_),
    .A2(_0830_),
    .B1(_0668_),
    .Y(_0831_));
 sky130_fd_sc_hd__a31o_1 _2351_ (.A1(_0668_),
    .A2(_0827_),
    .A3(_0830_),
    .B1(_0730_),
    .X(_0832_));
 sky130_fd_sc_hd__a2bb2o_1 _2352_ (.A1_N(_0831_),
    .A2_N(_0832_),
    .B1(_0763_),
    .B2(\po_0.alu_0._11_[8] ),
    .X(_0833_));
 sky130_fd_sc_hd__a21o_1 _2353_ (.A1(net86),
    .A2(_0747_),
    .B1(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__a22o_2 _2354_ (.A1(net15),
    .A2(_0823_),
    .B1(_0834_),
    .B2(_0753_),
    .X(_0835_));
 sky130_fd_sc_hd__clkbuf_2 _2355_ (.A(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_1 _2356_ (.A0(\po_0.regf_0.rf[5][8] ),
    .A1(_0836_),
    .S(_0810_),
    .X(_0837_));
 sky130_fd_sc_hd__clkbuf_1 _2357_ (.A(_0837_),
    .X(_0024_));
 sky130_fd_sc_hd__or3_1 _2358_ (.A(_0666_),
    .B(_0673_),
    .C(_0831_),
    .X(_0838_));
 sky130_fd_sc_hd__o21ai_1 _2359_ (.A1(_0666_),
    .A2(_0831_),
    .B1(_0673_),
    .Y(_0839_));
 sky130_fd_sc_hd__a21o_1 _2360_ (.A1(_0773_),
    .A2(\po_0.alu_0._11_[9] ),
    .B1(_0747_),
    .X(_0840_));
 sky130_fd_sc_hd__a31o_1 _2361_ (.A1(_0838_),
    .A2(_0839_),
    .A3(_0762_),
    .B1(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__or3_1 _2362_ (.A(_0671_),
    .B(_0763_),
    .C(_1487_),
    .X(_0842_));
 sky130_fd_sc_hd__a32o_2 _2363_ (.A1(_0841_),
    .A2(_0842_),
    .A3(_0752_),
    .B1(_0823_),
    .B2(net16),
    .X(_0843_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2364_ (.A(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_1 _2365_ (.A0(\po_0.regf_0.rf[5][9] ),
    .A1(_0844_),
    .S(_0810_),
    .X(_0845_));
 sky130_fd_sc_hd__clkbuf_1 _2366_ (.A(_0845_),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_1 _2367_ (.A1(net49),
    .A2(\po_0._1_[8] ),
    .B1(\po_0._1_[9] ),
    .B2(net50),
    .X(_0846_));
 sky130_fd_sc_hd__o22ai_1 _2368_ (.A1(_0671_),
    .A2(\po_0._1_[9] ),
    .B1(_0846_),
    .B2(_0831_),
    .Y(_0847_));
 sky130_fd_sc_hd__a21o_1 _2369_ (.A1(_0677_),
    .A2(_0678_),
    .B1(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__nand3_1 _2370_ (.A(_0847_),
    .B(_0678_),
    .C(_0677_),
    .Y(_0849_));
 sky130_fd_sc_hd__a22o_1 _2371_ (.A1(_0773_),
    .A2(\po_0.alu_0._11_[10] ),
    .B1(_0746_),
    .B2(_1522_),
    .X(_0850_));
 sky130_fd_sc_hd__a31o_1 _2372_ (.A1(_0848_),
    .A2(_0762_),
    .A3(_0849_),
    .B1(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__a22o_2 _2373_ (.A1(net2),
    .A2(_0823_),
    .B1(_0851_),
    .B2(_0753_),
    .X(_0852_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2374_ (.A(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_1 _2375_ (.A0(\po_0.regf_0.rf[5][10] ),
    .A1(_0853_),
    .S(_0810_),
    .X(_0854_));
 sky130_fd_sc_hd__clkbuf_1 _2376_ (.A(_0854_),
    .X(_0026_));
 sky130_fd_sc_hd__o22a_1 _2377_ (.A1(_0671_),
    .A2(\po_0._1_[9] ),
    .B1(_0846_),
    .B2(_0831_),
    .X(_0855_));
 sky130_fd_sc_hd__a22oi_2 _2378_ (.A1(_1522_),
    .A2(\po_0._1_[10] ),
    .B1(_0855_),
    .B2(_0679_),
    .Y(_0856_));
 sky130_fd_sc_hd__a21oi_1 _2379_ (.A1(_0685_),
    .A2(_0856_),
    .B1(_0731_),
    .Y(_0857_));
 sky130_fd_sc_hd__o21ai_1 _2380_ (.A1(_0685_),
    .A2(_0856_),
    .B1(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__or2_1 _2381_ (.A(\po_0.alu_0.s1 ),
    .B(_1487_),
    .X(_0859_));
 sky130_fd_sc_hd__o221a_1 _2382_ (.A1(_1491_),
    .A2(\po_0.alu_0._11_[11] ),
    .B1(_0859_),
    .B2(net85),
    .C1(_0752_),
    .X(_0860_));
 sky130_fd_sc_hd__a22o_2 _2383_ (.A1(net3),
    .A2(_0823_),
    .B1(_0858_),
    .B2(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__clkbuf_2 _2384_ (.A(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__mux2_1 _2385_ (.A0(\po_0.regf_0.rf[5][11] ),
    .A1(_0862_),
    .S(_0810_),
    .X(_0863_));
 sky130_fd_sc_hd__clkbuf_1 _2386_ (.A(_0863_),
    .X(_0027_));
 sky130_fd_sc_hd__o211a_1 _2387_ (.A1(_0671_),
    .A2(\po_0._1_[9] ),
    .B1(_0846_),
    .C1(_0679_),
    .X(_0864_));
 sky130_fd_sc_hd__a221oi_4 _2388_ (.A1(_1522_),
    .A2(\po_0._1_[10] ),
    .B1(\po_0._1_[11] ),
    .B2(net85),
    .C1(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__nand4_2 _2389_ (.A(_0695_),
    .B(_0672_),
    .C(_0679_),
    .D(_0685_),
    .Y(_0866_));
 sky130_fd_sc_hd__a21oi_1 _2390_ (.A1(_0829_),
    .A2(_0828_),
    .B1(_0660_),
    .Y(_0867_));
 sky130_fd_sc_hd__a31oi_4 _2391_ (.A1(_0826_),
    .A2(_0782_),
    .A3(_0626_),
    .B1(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__o22ai_4 _2392_ (.A1(_0683_),
    .A2(_0865_),
    .B1(_0866_),
    .B2(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__a21oi_1 _2393_ (.A1(_0869_),
    .A2(_0692_),
    .B1(_0731_),
    .Y(_0870_));
 sky130_fd_sc_hd__o21a_1 _2394_ (.A1(_0692_),
    .A2(_0869_),
    .B1(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__a221o_1 _2395_ (.A1(_0729_),
    .A2(\po_0.alu_0._11_[12] ),
    .B1(_0747_),
    .B2(net84),
    .C1(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__a22o_2 _2396_ (.A1(net4),
    .A2(_0823_),
    .B1(_0872_),
    .B2(_0753_),
    .X(_0873_));
 sky130_fd_sc_hd__clkbuf_2 _2397_ (.A(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__mux2_1 _2398_ (.A0(\po_0.regf_0.rf[5][12] ),
    .A1(_0874_),
    .S(_0743_),
    .X(_0875_));
 sky130_fd_sc_hd__clkbuf_1 _2399_ (.A(_0875_),
    .X(_0028_));
 sky130_fd_sc_hd__a21o_1 _2400_ (.A1(_0869_),
    .A2(_0692_),
    .B1(_0689_),
    .X(_0876_));
 sky130_fd_sc_hd__nand2_1 _2401_ (.A(_0876_),
    .B(_0701_),
    .Y(_0877_));
 sky130_fd_sc_hd__a211o_1 _2402_ (.A1(_0869_),
    .A2(_0692_),
    .B1(_0689_),
    .C1(_0701_),
    .X(_0878_));
 sky130_fd_sc_hd__a21o_1 _2403_ (.A1(_0773_),
    .A2(\po_0.alu_0._11_[13] ),
    .B1(_0746_),
    .X(_0879_));
 sky130_fd_sc_hd__a31o_1 _2404_ (.A1(_0877_),
    .A2(_0878_),
    .A3(_0762_),
    .B1(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__or3_1 _2405_ (.A(net83),
    .B(_0763_),
    .C(_1487_),
    .X(_0881_));
 sky130_fd_sc_hd__a32o_2 _2406_ (.A1(_0880_),
    .A2(_0752_),
    .A3(_0881_),
    .B1(_0823_),
    .B2(net5),
    .X(_0882_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2407_ (.A(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _2408_ (.A0(\po_0.regf_0.rf[5][13] ),
    .A1(_0883_),
    .S(_0743_),
    .X(_0884_));
 sky130_fd_sc_hd__clkbuf_1 _2409_ (.A(_0884_),
    .X(_0029_));
 sky130_fd_sc_hd__nand3_1 _2410_ (.A(_0869_),
    .B(_0700_),
    .C(_0691_),
    .Y(_0885_));
 sky130_fd_sc_hd__o211a_1 _2411_ (.A1(net83),
    .A2(\po_0._1_[13] ),
    .B1(\po_0._1_[12] ),
    .C1(net38),
    .X(_0886_));
 sky130_fd_sc_hd__a21oi_1 _2412_ (.A1(net83),
    .A2(\po_0._1_[13] ),
    .B1(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__nand2_1 _2413_ (.A(_0708_),
    .B(_0709_),
    .Y(_0888_));
 sky130_fd_sc_hd__a21o_1 _2414_ (.A1(_0885_),
    .A2(_0887_),
    .B1(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__or3b_1 _2415_ (.A(_0689_),
    .B(_0690_),
    .C_N(_0700_),
    .X(_0890_));
 sky130_fd_sc_hd__o22a_1 _2416_ (.A1(_0683_),
    .A2(_0865_),
    .B1(_0866_),
    .B2(_0868_),
    .X(_0891_));
 sky130_fd_sc_hd__o211ai_1 _2417_ (.A1(_0890_),
    .A2(_0891_),
    .B1(_0888_),
    .C1(_0887_),
    .Y(_0892_));
 sky130_fd_sc_hd__a22o_1 _2418_ (.A1(_0773_),
    .A2(\po_0.alu_0._11_[14] ),
    .B1(_0746_),
    .B2(_0707_),
    .X(_0893_));
 sky130_fd_sc_hd__a31o_1 _2419_ (.A1(_0889_),
    .A2(_0892_),
    .A3(_0762_),
    .B1(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__a22o_2 _2420_ (.A1(net6),
    .A2(_0728_),
    .B1(_0894_),
    .B2(_0752_),
    .X(_0895_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2421_ (.A(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_1 _2422_ (.A0(\po_0.regf_0.rf[5][14] ),
    .A1(_0896_),
    .S(_0743_),
    .X(_0897_));
 sky130_fd_sc_hd__clkbuf_1 _2423_ (.A(_0897_),
    .X(_0030_));
 sky130_fd_sc_hd__a21oi_1 _2424_ (.A1(_0885_),
    .A2(_0887_),
    .B1(_0888_),
    .Y(_0898_));
 sky130_fd_sc_hd__o21bai_1 _2425_ (.A1(_0718_),
    .A2(_0898_),
    .B1_N(_0716_),
    .Y(_0899_));
 sky130_fd_sc_hd__o211ai_1 _2426_ (.A1(_0714_),
    .A2(_0715_),
    .B1(_0889_),
    .C1(_0708_),
    .Y(_0900_));
 sky130_fd_sc_hd__nand3_1 _2427_ (.A(_0899_),
    .B(_0900_),
    .C(_0762_),
    .Y(_0901_));
 sky130_fd_sc_hd__o221a_1 _2428_ (.A1(_1491_),
    .A2(\po_0.alu_0._11_[15] ),
    .B1(_0859_),
    .B2(net41),
    .C1(_0732_),
    .X(_0902_));
 sky130_fd_sc_hd__a22o_2 _2429_ (.A1(net7),
    .A2(_0728_),
    .B1(_0901_),
    .B2(_0902_),
    .X(_0903_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2430_ (.A(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _2431_ (.A0(\po_0.regf_0.rf[5][15] ),
    .A1(_0904_),
    .S(_0743_),
    .X(_0905_));
 sky130_fd_sc_hd__clkbuf_1 _2432_ (.A(_0905_),
    .X(_0031_));
 sky130_fd_sc_hd__clkbuf_2 _2433_ (.A(\po_0.regf_0.w_wr ),
    .X(_0906_));
 sky130_fd_sc_hd__and2b_1 _2434_ (.A_N(_0740_),
    .B(_0739_),
    .X(_0907_));
 sky130_fd_sc_hd__and4b_4 _2435_ (.A_N(_0737_),
    .B(_0906_),
    .C(_0907_),
    .D(_0742_),
    .X(_0908_));
 sky130_fd_sc_hd__buf_2 _2436_ (.A(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _2437_ (.A0(\po_0.regf_0.rf[6][0] ),
    .A1(_0736_),
    .S(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__clkbuf_1 _2438_ (.A(_0910_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2439_ (.A0(\po_0.regf_0.rf[6][1] ),
    .A1(_0756_),
    .S(_0909_),
    .X(_0911_));
 sky130_fd_sc_hd__clkbuf_1 _2440_ (.A(_0911_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _2441_ (.A0(\po_0.regf_0.rf[6][2] ),
    .A1(_0768_),
    .S(_0909_),
    .X(_0912_));
 sky130_fd_sc_hd__clkbuf_1 _2442_ (.A(_0912_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2443_ (.A0(\po_0.regf_0.rf[6][3] ),
    .A1(_0778_),
    .S(_0909_),
    .X(_0913_));
 sky130_fd_sc_hd__clkbuf_1 _2444_ (.A(_0913_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2445_ (.A0(\po_0.regf_0.rf[6][4] ),
    .A1(_0789_),
    .S(_0909_),
    .X(_0914_));
 sky130_fd_sc_hd__clkbuf_1 _2446_ (.A(_0914_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2447_ (.A0(\po_0.regf_0.rf[6][5] ),
    .A1(_0797_),
    .S(_0909_),
    .X(_0915_));
 sky130_fd_sc_hd__clkbuf_1 _2448_ (.A(_0915_),
    .X(_0037_));
 sky130_fd_sc_hd__buf_2 _2449_ (.A(_0908_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _2450_ (.A0(\po_0.regf_0.rf[6][6] ),
    .A1(_0809_),
    .S(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__clkbuf_1 _2451_ (.A(_0917_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2452_ (.A0(\po_0.regf_0.rf[6][7] ),
    .A1(_0821_),
    .S(_0916_),
    .X(_0918_));
 sky130_fd_sc_hd__clkbuf_1 _2453_ (.A(_0918_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2454_ (.A0(\po_0.regf_0.rf[6][8] ),
    .A1(_0836_),
    .S(_0916_),
    .X(_0919_));
 sky130_fd_sc_hd__clkbuf_1 _2455_ (.A(_0919_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2456_ (.A0(\po_0.regf_0.rf[6][9] ),
    .A1(_0844_),
    .S(_0916_),
    .X(_0920_));
 sky130_fd_sc_hd__clkbuf_1 _2457_ (.A(_0920_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _2458_ (.A0(\po_0.regf_0.rf[6][10] ),
    .A1(_0853_),
    .S(_0916_),
    .X(_0921_));
 sky130_fd_sc_hd__clkbuf_1 _2459_ (.A(_0921_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _2460_ (.A0(\po_0.regf_0.rf[6][11] ),
    .A1(_0862_),
    .S(_0916_),
    .X(_0922_));
 sky130_fd_sc_hd__clkbuf_1 _2461_ (.A(_0922_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _2462_ (.A0(\po_0.regf_0.rf[6][12] ),
    .A1(_0874_),
    .S(_0908_),
    .X(_0923_));
 sky130_fd_sc_hd__clkbuf_1 _2463_ (.A(_0923_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _2464_ (.A0(\po_0.regf_0.rf[6][13] ),
    .A1(_0883_),
    .S(_0908_),
    .X(_0924_));
 sky130_fd_sc_hd__clkbuf_1 _2465_ (.A(_0924_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2466_ (.A0(\po_0.regf_0.rf[6][14] ),
    .A1(_0896_),
    .S(_0908_),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_1 _2467_ (.A(_0925_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2468_ (.A0(\po_0.regf_0.rf[6][15] ),
    .A1(_0904_),
    .S(_0908_),
    .X(_0926_));
 sky130_fd_sc_hd__clkbuf_1 _2469_ (.A(_0926_),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_2 _2470_ (.A(\po_0.regf_0.w_addr[3] ),
    .X(_0927_));
 sky130_fd_sc_hd__and2_2 _2471_ (.A(\po_0.regf_0.w_addr[0] ),
    .B(\po_0.regf_0.w_addr[1] ),
    .X(_0928_));
 sky130_fd_sc_hd__clkbuf_2 _2472_ (.A(\po_0.regf_0.w_addr[2] ),
    .X(_0929_));
 sky130_fd_sc_hd__nand4b_4 _2473_ (.A_N(_0927_),
    .B(_0738_),
    .C(_0928_),
    .D(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__buf_2 _2474_ (.A(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_1 _2475_ (.A0(_0736_),
    .A1(\po_0.regf_0.rf[7][0] ),
    .S(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__clkbuf_1 _2476_ (.A(_0932_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _2477_ (.A0(_0756_),
    .A1(\po_0.regf_0.rf[7][1] ),
    .S(_0931_),
    .X(_0933_));
 sky130_fd_sc_hd__clkbuf_1 _2478_ (.A(_0933_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _2479_ (.A0(_0768_),
    .A1(\po_0.regf_0.rf[7][2] ),
    .S(_0931_),
    .X(_0934_));
 sky130_fd_sc_hd__clkbuf_1 _2480_ (.A(_0934_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _2481_ (.A0(_0778_),
    .A1(\po_0.regf_0.rf[7][3] ),
    .S(_0931_),
    .X(_0935_));
 sky130_fd_sc_hd__clkbuf_1 _2482_ (.A(_0935_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _2483_ (.A0(_0789_),
    .A1(\po_0.regf_0.rf[7][4] ),
    .S(_0931_),
    .X(_0936_));
 sky130_fd_sc_hd__clkbuf_1 _2484_ (.A(_0936_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _2485_ (.A0(_0797_),
    .A1(\po_0.regf_0.rf[7][5] ),
    .S(_0931_),
    .X(_0937_));
 sky130_fd_sc_hd__clkbuf_1 _2486_ (.A(_0937_),
    .X(_0053_));
 sky130_fd_sc_hd__buf_2 _2487_ (.A(_0930_),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_1 _2488_ (.A0(_0809_),
    .A1(\po_0.regf_0.rf[7][6] ),
    .S(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__clkbuf_1 _2489_ (.A(_0939_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2490_ (.A0(_0821_),
    .A1(\po_0.regf_0.rf[7][7] ),
    .S(_0938_),
    .X(_0940_));
 sky130_fd_sc_hd__clkbuf_1 _2491_ (.A(_0940_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2492_ (.A0(_0836_),
    .A1(\po_0.regf_0.rf[7][8] ),
    .S(_0938_),
    .X(_0941_));
 sky130_fd_sc_hd__clkbuf_1 _2493_ (.A(_0941_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2494_ (.A0(_0844_),
    .A1(\po_0.regf_0.rf[7][9] ),
    .S(_0938_),
    .X(_0942_));
 sky130_fd_sc_hd__clkbuf_1 _2495_ (.A(_0942_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2496_ (.A0(_0853_),
    .A1(\po_0.regf_0.rf[7][10] ),
    .S(_0938_),
    .X(_0943_));
 sky130_fd_sc_hd__clkbuf_1 _2497_ (.A(_0943_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _2498_ (.A0(_0862_),
    .A1(\po_0.regf_0.rf[7][11] ),
    .S(_0938_),
    .X(_0944_));
 sky130_fd_sc_hd__clkbuf_1 _2499_ (.A(_0944_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _2500_ (.A0(_0874_),
    .A1(\po_0.regf_0.rf[7][12] ),
    .S(_0930_),
    .X(_0945_));
 sky130_fd_sc_hd__clkbuf_1 _2501_ (.A(_0945_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _2502_ (.A0(_0883_),
    .A1(\po_0.regf_0.rf[7][13] ),
    .S(_0930_),
    .X(_0946_));
 sky130_fd_sc_hd__clkbuf_1 _2503_ (.A(_0946_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(_0896_),
    .A1(\po_0.regf_0.rf[7][14] ),
    .S(_0930_),
    .X(_0947_));
 sky130_fd_sc_hd__clkbuf_1 _2505_ (.A(_0947_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(_0904_),
    .A1(\po_0.regf_0.rf[7][15] ),
    .S(_0930_),
    .X(_0948_));
 sky130_fd_sc_hd__clkbuf_1 _2507_ (.A(_0948_),
    .X(_0063_));
 sky130_fd_sc_hd__clkbuf_2 _2508_ (.A(_0735_),
    .X(_0949_));
 sky130_fd_sc_hd__and4b_4 _2509_ (.A_N(_0742_),
    .B(_0927_),
    .C(_0906_),
    .D(_0741_),
    .X(_0950_));
 sky130_fd_sc_hd__buf_2 _2510_ (.A(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_1 _2511_ (.A0(\po_0.regf_0.rf[9][0] ),
    .A1(_0949_),
    .S(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__clkbuf_1 _2512_ (.A(_0952_),
    .X(_0064_));
 sky130_fd_sc_hd__clkbuf_2 _2513_ (.A(_0755_),
    .X(_0953_));
 sky130_fd_sc_hd__mux2_1 _2514_ (.A0(\po_0.regf_0.rf[9][1] ),
    .A1(_0953_),
    .S(_0951_),
    .X(_0954_));
 sky130_fd_sc_hd__clkbuf_1 _2515_ (.A(_0954_),
    .X(_0065_));
 sky130_fd_sc_hd__clkbuf_2 _2516_ (.A(_0767_),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(\po_0.regf_0.rf[9][2] ),
    .A1(_0955_),
    .S(_0951_),
    .X(_0956_));
 sky130_fd_sc_hd__clkbuf_1 _2518_ (.A(_0956_),
    .X(_0066_));
 sky130_fd_sc_hd__clkbuf_2 _2519_ (.A(_0777_),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(\po_0.regf_0.rf[9][3] ),
    .A1(_0957_),
    .S(_0951_),
    .X(_0958_));
 sky130_fd_sc_hd__clkbuf_1 _2521_ (.A(_0958_),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_2 _2522_ (.A(_0788_),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(\po_0.regf_0.rf[9][4] ),
    .A1(_0959_),
    .S(_0951_),
    .X(_0960_));
 sky130_fd_sc_hd__clkbuf_1 _2524_ (.A(_0960_),
    .X(_0068_));
 sky130_fd_sc_hd__clkbuf_2 _2525_ (.A(_0796_),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(\po_0.regf_0.rf[9][5] ),
    .A1(_0961_),
    .S(_0951_),
    .X(_0962_));
 sky130_fd_sc_hd__clkbuf_1 _2527_ (.A(_0962_),
    .X(_0069_));
 sky130_fd_sc_hd__clkbuf_2 _2528_ (.A(_0808_),
    .X(_0963_));
 sky130_fd_sc_hd__buf_2 _2529_ (.A(_0950_),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(\po_0.regf_0.rf[9][6] ),
    .A1(_0963_),
    .S(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__clkbuf_1 _2531_ (.A(_0965_),
    .X(_0070_));
 sky130_fd_sc_hd__clkbuf_2 _2532_ (.A(_0820_),
    .X(_0966_));
 sky130_fd_sc_hd__mux2_1 _2533_ (.A0(\po_0.regf_0.rf[9][7] ),
    .A1(_0966_),
    .S(_0964_),
    .X(_0967_));
 sky130_fd_sc_hd__clkbuf_1 _2534_ (.A(_0967_),
    .X(_0071_));
 sky130_fd_sc_hd__clkbuf_2 _2535_ (.A(_0835_),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_1 _2536_ (.A0(\po_0.regf_0.rf[9][8] ),
    .A1(_0968_),
    .S(_0964_),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_1 _2537_ (.A(_0969_),
    .X(_0072_));
 sky130_fd_sc_hd__clkbuf_2 _2538_ (.A(_0843_),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_1 _2539_ (.A0(\po_0.regf_0.rf[9][9] ),
    .A1(_0970_),
    .S(_0964_),
    .X(_0971_));
 sky130_fd_sc_hd__clkbuf_1 _2540_ (.A(_0971_),
    .X(_0073_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2541_ (.A(_0852_),
    .X(_0972_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(\po_0.regf_0.rf[9][10] ),
    .A1(_0972_),
    .S(_0964_),
    .X(_0973_));
 sky130_fd_sc_hd__clkbuf_1 _2543_ (.A(_0973_),
    .X(_0074_));
 sky130_fd_sc_hd__clkbuf_2 _2544_ (.A(_0861_),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_1 _2545_ (.A0(\po_0.regf_0.rf[9][11] ),
    .A1(_0974_),
    .S(_0964_),
    .X(_0975_));
 sky130_fd_sc_hd__clkbuf_1 _2546_ (.A(_0975_),
    .X(_0075_));
 sky130_fd_sc_hd__clkbuf_2 _2547_ (.A(_0873_),
    .X(_0976_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(\po_0.regf_0.rf[9][12] ),
    .A1(_0976_),
    .S(_0950_),
    .X(_0977_));
 sky130_fd_sc_hd__clkbuf_1 _2549_ (.A(_0977_),
    .X(_0076_));
 sky130_fd_sc_hd__clkbuf_2 _2550_ (.A(_0882_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(\po_0.regf_0.rf[9][13] ),
    .A1(_0978_),
    .S(_0950_),
    .X(_0979_));
 sky130_fd_sc_hd__clkbuf_1 _2552_ (.A(_0979_),
    .X(_0077_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2553_ (.A(_0895_),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_1 _2554_ (.A0(\po_0.regf_0.rf[9][14] ),
    .A1(_0980_),
    .S(_0950_),
    .X(_0981_));
 sky130_fd_sc_hd__clkbuf_1 _2555_ (.A(_0981_),
    .X(_0078_));
 sky130_fd_sc_hd__clkbuf_2 _2556_ (.A(_0903_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(\po_0.regf_0.rf[9][15] ),
    .A1(_0982_),
    .S(_0950_),
    .X(_0983_));
 sky130_fd_sc_hd__clkbuf_1 _2558_ (.A(_0983_),
    .X(_0079_));
 sky130_fd_sc_hd__and4bb_4 _2559_ (.A_N(_0929_),
    .B_N(\po_0.regf_0.w_addr[3] ),
    .C(_0906_),
    .D(_0741_),
    .X(_0984_));
 sky130_fd_sc_hd__clkbuf_4 _2560_ (.A(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(\po_0.regf_0.rf[1][0] ),
    .A1(_0949_),
    .S(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__clkbuf_1 _2562_ (.A(_0986_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2563_ (.A0(\po_0.regf_0.rf[1][1] ),
    .A1(_0953_),
    .S(_0985_),
    .X(_0987_));
 sky130_fd_sc_hd__clkbuf_1 _2564_ (.A(_0987_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(\po_0.regf_0.rf[1][2] ),
    .A1(_0955_),
    .S(_0985_),
    .X(_0988_));
 sky130_fd_sc_hd__clkbuf_1 _2566_ (.A(_0988_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(\po_0.regf_0.rf[1][3] ),
    .A1(_0957_),
    .S(_0985_),
    .X(_0989_));
 sky130_fd_sc_hd__clkbuf_1 _2568_ (.A(_0989_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(\po_0.regf_0.rf[1][4] ),
    .A1(_0959_),
    .S(_0985_),
    .X(_0990_));
 sky130_fd_sc_hd__clkbuf_1 _2570_ (.A(_0990_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2571_ (.A0(\po_0.regf_0.rf[1][5] ),
    .A1(_0961_),
    .S(_0985_),
    .X(_0991_));
 sky130_fd_sc_hd__clkbuf_1 _2572_ (.A(_0991_),
    .X(_0085_));
 sky130_fd_sc_hd__buf_2 _2573_ (.A(_0984_),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(\po_0.regf_0.rf[1][6] ),
    .A1(_0963_),
    .S(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__clkbuf_1 _2575_ (.A(_0993_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(\po_0.regf_0.rf[1][7] ),
    .A1(_0966_),
    .S(_0992_),
    .X(_0994_));
 sky130_fd_sc_hd__clkbuf_1 _2577_ (.A(_0994_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(\po_0.regf_0.rf[1][8] ),
    .A1(_0968_),
    .S(_0992_),
    .X(_0995_));
 sky130_fd_sc_hd__clkbuf_1 _2579_ (.A(_0995_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(\po_0.regf_0.rf[1][9] ),
    .A1(_0970_),
    .S(_0992_),
    .X(_0996_));
 sky130_fd_sc_hd__clkbuf_1 _2581_ (.A(_0996_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(\po_0.regf_0.rf[1][10] ),
    .A1(_0972_),
    .S(_0992_),
    .X(_0997_));
 sky130_fd_sc_hd__clkbuf_1 _2583_ (.A(_0997_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _2584_ (.A0(\po_0.regf_0.rf[1][11] ),
    .A1(_0974_),
    .S(_0992_),
    .X(_0998_));
 sky130_fd_sc_hd__clkbuf_1 _2585_ (.A(_0998_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _2586_ (.A0(\po_0.regf_0.rf[1][12] ),
    .A1(_0976_),
    .S(_0984_),
    .X(_0999_));
 sky130_fd_sc_hd__clkbuf_1 _2587_ (.A(_0999_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2588_ (.A0(\po_0.regf_0.rf[1][13] ),
    .A1(_0978_),
    .S(_0984_),
    .X(_1000_));
 sky130_fd_sc_hd__clkbuf_1 _2589_ (.A(_1000_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2590_ (.A0(\po_0.regf_0.rf[1][14] ),
    .A1(_0980_),
    .S(_0984_),
    .X(_1001_));
 sky130_fd_sc_hd__clkbuf_1 _2591_ (.A(_1001_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _2592_ (.A0(\po_0.regf_0.rf[1][15] ),
    .A1(_0982_),
    .S(_0984_),
    .X(_1002_));
 sky130_fd_sc_hd__clkbuf_1 _2593_ (.A(_1002_),
    .X(_0095_));
 sky130_fd_sc_hd__and4_4 _2594_ (.A(_0929_),
    .B(_0927_),
    .C(_0738_),
    .D(_0928_),
    .X(_1003_));
 sky130_fd_sc_hd__buf_2 _2595_ (.A(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_1 _2596_ (.A0(\po_0.regf_0.rf[15][0] ),
    .A1(_0949_),
    .S(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__clkbuf_1 _2597_ (.A(_1005_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _2598_ (.A0(\po_0.regf_0.rf[15][1] ),
    .A1(_0953_),
    .S(_1004_),
    .X(_1006_));
 sky130_fd_sc_hd__clkbuf_1 _2599_ (.A(_1006_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _2600_ (.A0(\po_0.regf_0.rf[15][2] ),
    .A1(_0955_),
    .S(_1004_),
    .X(_1007_));
 sky130_fd_sc_hd__clkbuf_1 _2601_ (.A(_1007_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _2602_ (.A0(\po_0.regf_0.rf[15][3] ),
    .A1(_0957_),
    .S(_1004_),
    .X(_1008_));
 sky130_fd_sc_hd__clkbuf_1 _2603_ (.A(_1008_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _2604_ (.A0(\po_0.regf_0.rf[15][4] ),
    .A1(_0959_),
    .S(_1004_),
    .X(_1009_));
 sky130_fd_sc_hd__clkbuf_1 _2605_ (.A(_1009_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2606_ (.A0(\po_0.regf_0.rf[15][5] ),
    .A1(_0961_),
    .S(_1004_),
    .X(_1010_));
 sky130_fd_sc_hd__clkbuf_1 _2607_ (.A(_1010_),
    .X(_0101_));
 sky130_fd_sc_hd__buf_2 _2608_ (.A(_1003_),
    .X(_1011_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(\po_0.regf_0.rf[15][6] ),
    .A1(_0963_),
    .S(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__clkbuf_1 _2610_ (.A(_1012_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(\po_0.regf_0.rf[15][7] ),
    .A1(_0966_),
    .S(_1011_),
    .X(_1013_));
 sky130_fd_sc_hd__clkbuf_1 _2612_ (.A(_1013_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _2613_ (.A0(\po_0.regf_0.rf[15][8] ),
    .A1(_0968_),
    .S(_1011_),
    .X(_1014_));
 sky130_fd_sc_hd__clkbuf_1 _2614_ (.A(_1014_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _2615_ (.A0(\po_0.regf_0.rf[15][9] ),
    .A1(_0970_),
    .S(_1011_),
    .X(_1015_));
 sky130_fd_sc_hd__clkbuf_1 _2616_ (.A(_1015_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2617_ (.A0(\po_0.regf_0.rf[15][10] ),
    .A1(_0972_),
    .S(_1011_),
    .X(_1016_));
 sky130_fd_sc_hd__clkbuf_1 _2618_ (.A(_1016_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _2619_ (.A0(\po_0.regf_0.rf[15][11] ),
    .A1(_0974_),
    .S(_1011_),
    .X(_1017_));
 sky130_fd_sc_hd__clkbuf_1 _2620_ (.A(_1017_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _2621_ (.A0(\po_0.regf_0.rf[15][12] ),
    .A1(_0976_),
    .S(_1003_),
    .X(_1018_));
 sky130_fd_sc_hd__clkbuf_1 _2622_ (.A(_1018_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _2623_ (.A0(\po_0.regf_0.rf[15][13] ),
    .A1(_0978_),
    .S(_1003_),
    .X(_1019_));
 sky130_fd_sc_hd__clkbuf_1 _2624_ (.A(_1019_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _2625_ (.A0(\po_0.regf_0.rf[15][14] ),
    .A1(_0980_),
    .S(_1003_),
    .X(_1020_));
 sky130_fd_sc_hd__clkbuf_1 _2626_ (.A(_1020_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _2627_ (.A0(\po_0.regf_0.rf[15][15] ),
    .A1(_0982_),
    .S(_1003_),
    .X(_1021_));
 sky130_fd_sc_hd__clkbuf_1 _2628_ (.A(_1021_),
    .X(_0111_));
 sky130_fd_sc_hd__nand3_1 _2629_ (.A(\po_0.regf_0.w_addr[2] ),
    .B(\po_0.regf_0.w_addr[3] ),
    .C(\po_0.regf_0.w_wr ),
    .Y(_1022_));
 sky130_fd_sc_hd__or3b_4 _2630_ (.A(_1022_),
    .B(_0740_),
    .C_N(_0739_),
    .X(_1023_));
 sky130_fd_sc_hd__buf_2 _2631_ (.A(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(_0736_),
    .A1(\po_0.regf_0.rf[14][0] ),
    .S(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__clkbuf_1 _2633_ (.A(_1025_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(_0756_),
    .A1(\po_0.regf_0.rf[14][1] ),
    .S(_1024_),
    .X(_1026_));
 sky130_fd_sc_hd__clkbuf_1 _2635_ (.A(_1026_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(_0768_),
    .A1(\po_0.regf_0.rf[14][2] ),
    .S(_1024_),
    .X(_1027_));
 sky130_fd_sc_hd__clkbuf_1 _2637_ (.A(_1027_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _2638_ (.A0(_0778_),
    .A1(\po_0.regf_0.rf[14][3] ),
    .S(_1024_),
    .X(_1028_));
 sky130_fd_sc_hd__clkbuf_1 _2639_ (.A(_1028_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _2640_ (.A0(_0789_),
    .A1(\po_0.regf_0.rf[14][4] ),
    .S(_1024_),
    .X(_1029_));
 sky130_fd_sc_hd__clkbuf_1 _2641_ (.A(_1029_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _2642_ (.A0(_0797_),
    .A1(\po_0.regf_0.rf[14][5] ),
    .S(_1024_),
    .X(_1030_));
 sky130_fd_sc_hd__clkbuf_1 _2643_ (.A(_1030_),
    .X(_0117_));
 sky130_fd_sc_hd__buf_2 _2644_ (.A(_1023_),
    .X(_1031_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(_0809_),
    .A1(\po_0.regf_0.rf[14][6] ),
    .S(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__clkbuf_1 _2646_ (.A(_1032_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _2647_ (.A0(_0821_),
    .A1(\po_0.regf_0.rf[14][7] ),
    .S(_1031_),
    .X(_1033_));
 sky130_fd_sc_hd__clkbuf_1 _2648_ (.A(_1033_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _2649_ (.A0(_0836_),
    .A1(\po_0.regf_0.rf[14][8] ),
    .S(_1031_),
    .X(_1034_));
 sky130_fd_sc_hd__clkbuf_1 _2650_ (.A(_1034_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _2651_ (.A0(_0844_),
    .A1(\po_0.regf_0.rf[14][9] ),
    .S(_1031_),
    .X(_1035_));
 sky130_fd_sc_hd__clkbuf_1 _2652_ (.A(_1035_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2653_ (.A0(_0853_),
    .A1(\po_0.regf_0.rf[14][10] ),
    .S(_1031_),
    .X(_1036_));
 sky130_fd_sc_hd__clkbuf_1 _2654_ (.A(_1036_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _2655_ (.A0(_0862_),
    .A1(\po_0.regf_0.rf[14][11] ),
    .S(_1031_),
    .X(_1037_));
 sky130_fd_sc_hd__clkbuf_1 _2656_ (.A(_1037_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _2657_ (.A0(_0874_),
    .A1(\po_0.regf_0.rf[14][12] ),
    .S(_1023_),
    .X(_1038_));
 sky130_fd_sc_hd__clkbuf_1 _2658_ (.A(_1038_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _2659_ (.A0(_0883_),
    .A1(\po_0.regf_0.rf[14][13] ),
    .S(_1023_),
    .X(_1039_));
 sky130_fd_sc_hd__clkbuf_1 _2660_ (.A(_1039_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2661_ (.A0(_0896_),
    .A1(\po_0.regf_0.rf[14][14] ),
    .S(_1023_),
    .X(_1040_));
 sky130_fd_sc_hd__clkbuf_1 _2662_ (.A(_1040_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _2663_ (.A0(_0904_),
    .A1(\po_0.regf_0.rf[14][15] ),
    .S(_1023_),
    .X(_1041_));
 sky130_fd_sc_hd__clkbuf_1 _2664_ (.A(_1041_),
    .X(_0127_));
 sky130_fd_sc_hd__or3b_4 _2665_ (.A(_0739_),
    .B(_1022_),
    .C_N(_0740_),
    .X(_1042_));
 sky130_fd_sc_hd__buf_2 _2666_ (.A(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__mux2_1 _2667_ (.A0(_0736_),
    .A1(\po_0.regf_0.rf[13][0] ),
    .S(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__clkbuf_1 _2668_ (.A(_1044_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _2669_ (.A0(_0756_),
    .A1(\po_0.regf_0.rf[13][1] ),
    .S(_1043_),
    .X(_1045_));
 sky130_fd_sc_hd__clkbuf_1 _2670_ (.A(_1045_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _2671_ (.A0(_0768_),
    .A1(\po_0.regf_0.rf[13][2] ),
    .S(_1043_),
    .X(_1046_));
 sky130_fd_sc_hd__clkbuf_1 _2672_ (.A(_1046_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _2673_ (.A0(_0778_),
    .A1(\po_0.regf_0.rf[13][3] ),
    .S(_1043_),
    .X(_1047_));
 sky130_fd_sc_hd__clkbuf_1 _2674_ (.A(_1047_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _2675_ (.A0(_0789_),
    .A1(\po_0.regf_0.rf[13][4] ),
    .S(_1043_),
    .X(_1048_));
 sky130_fd_sc_hd__clkbuf_1 _2676_ (.A(_1048_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2677_ (.A0(_0797_),
    .A1(\po_0.regf_0.rf[13][5] ),
    .S(_1043_),
    .X(_1049_));
 sky130_fd_sc_hd__clkbuf_1 _2678_ (.A(_1049_),
    .X(_0133_));
 sky130_fd_sc_hd__buf_2 _2679_ (.A(_1042_),
    .X(_1050_));
 sky130_fd_sc_hd__mux2_1 _2680_ (.A0(_0809_),
    .A1(\po_0.regf_0.rf[13][6] ),
    .S(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__clkbuf_1 _2681_ (.A(_1051_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _2682_ (.A0(_0821_),
    .A1(\po_0.regf_0.rf[13][7] ),
    .S(_1050_),
    .X(_1052_));
 sky130_fd_sc_hd__clkbuf_1 _2683_ (.A(_1052_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _2684_ (.A0(_0836_),
    .A1(\po_0.regf_0.rf[13][8] ),
    .S(_1050_),
    .X(_1053_));
 sky130_fd_sc_hd__clkbuf_1 _2685_ (.A(_1053_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _2686_ (.A0(_0844_),
    .A1(\po_0.regf_0.rf[13][9] ),
    .S(_1050_),
    .X(_1054_));
 sky130_fd_sc_hd__clkbuf_1 _2687_ (.A(_1054_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _2688_ (.A0(_0853_),
    .A1(\po_0.regf_0.rf[13][10] ),
    .S(_1050_),
    .X(_1055_));
 sky130_fd_sc_hd__clkbuf_1 _2689_ (.A(_1055_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _2690_ (.A0(_0862_),
    .A1(\po_0.regf_0.rf[13][11] ),
    .S(_1050_),
    .X(_1056_));
 sky130_fd_sc_hd__clkbuf_1 _2691_ (.A(_1056_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _2692_ (.A0(_0874_),
    .A1(\po_0.regf_0.rf[13][12] ),
    .S(_1042_),
    .X(_1057_));
 sky130_fd_sc_hd__clkbuf_1 _2693_ (.A(_1057_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(_0883_),
    .A1(\po_0.regf_0.rf[13][13] ),
    .S(_1042_),
    .X(_1058_));
 sky130_fd_sc_hd__clkbuf_1 _2695_ (.A(_1058_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2696_ (.A0(_0896_),
    .A1(\po_0.regf_0.rf[13][14] ),
    .S(_1042_),
    .X(_1059_));
 sky130_fd_sc_hd__clkbuf_1 _2697_ (.A(_1059_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _2698_ (.A0(_0904_),
    .A1(\po_0.regf_0.rf[13][15] ),
    .S(_1042_),
    .X(_1060_));
 sky130_fd_sc_hd__clkbuf_1 _2699_ (.A(_1060_),
    .X(_0143_));
 sky130_fd_sc_hd__nor2_1 _2700_ (.A(_0740_),
    .B(_0739_),
    .Y(_1061_));
 sky130_fd_sc_hd__and4_4 _2701_ (.A(_0929_),
    .B(_0927_),
    .C(_0738_),
    .D(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__buf_2 _2702_ (.A(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_1 _2703_ (.A0(\po_0.regf_0.rf[12][0] ),
    .A1(_0949_),
    .S(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__clkbuf_1 _2704_ (.A(_1064_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2705_ (.A0(\po_0.regf_0.rf[12][1] ),
    .A1(_0953_),
    .S(_1063_),
    .X(_1065_));
 sky130_fd_sc_hd__clkbuf_1 _2706_ (.A(_1065_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2707_ (.A0(\po_0.regf_0.rf[12][2] ),
    .A1(_0955_),
    .S(_1063_),
    .X(_1066_));
 sky130_fd_sc_hd__clkbuf_1 _2708_ (.A(_1066_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2709_ (.A0(\po_0.regf_0.rf[12][3] ),
    .A1(_0957_),
    .S(_1063_),
    .X(_1067_));
 sky130_fd_sc_hd__clkbuf_1 _2710_ (.A(_1067_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2711_ (.A0(\po_0.regf_0.rf[12][4] ),
    .A1(_0959_),
    .S(_1063_),
    .X(_1068_));
 sky130_fd_sc_hd__clkbuf_1 _2712_ (.A(_1068_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2713_ (.A0(\po_0.regf_0.rf[12][5] ),
    .A1(_0961_),
    .S(_1063_),
    .X(_1069_));
 sky130_fd_sc_hd__clkbuf_1 _2714_ (.A(_1069_),
    .X(_0149_));
 sky130_fd_sc_hd__buf_2 _2715_ (.A(_1062_),
    .X(_1070_));
 sky130_fd_sc_hd__mux2_1 _2716_ (.A0(\po_0.regf_0.rf[12][6] ),
    .A1(_0963_),
    .S(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__clkbuf_1 _2717_ (.A(_1071_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2718_ (.A0(\po_0.regf_0.rf[12][7] ),
    .A1(_0966_),
    .S(_1070_),
    .X(_1072_));
 sky130_fd_sc_hd__clkbuf_1 _2719_ (.A(_1072_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2720_ (.A0(\po_0.regf_0.rf[12][8] ),
    .A1(_0968_),
    .S(_1070_),
    .X(_1073_));
 sky130_fd_sc_hd__clkbuf_1 _2721_ (.A(_1073_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2722_ (.A0(\po_0.regf_0.rf[12][9] ),
    .A1(_0970_),
    .S(_1070_),
    .X(_1074_));
 sky130_fd_sc_hd__clkbuf_1 _2723_ (.A(_1074_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2724_ (.A0(\po_0.regf_0.rf[12][10] ),
    .A1(_0972_),
    .S(_1070_),
    .X(_1075_));
 sky130_fd_sc_hd__clkbuf_1 _2725_ (.A(_1075_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2726_ (.A0(\po_0.regf_0.rf[12][11] ),
    .A1(_0974_),
    .S(_1070_),
    .X(_1076_));
 sky130_fd_sc_hd__clkbuf_1 _2727_ (.A(_1076_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2728_ (.A0(\po_0.regf_0.rf[12][12] ),
    .A1(_0976_),
    .S(_1062_),
    .X(_1077_));
 sky130_fd_sc_hd__clkbuf_1 _2729_ (.A(_1077_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2730_ (.A0(\po_0.regf_0.rf[12][13] ),
    .A1(_0978_),
    .S(_1062_),
    .X(_1078_));
 sky130_fd_sc_hd__clkbuf_1 _2731_ (.A(_1078_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2732_ (.A0(\po_0.regf_0.rf[12][14] ),
    .A1(_0980_),
    .S(_1062_),
    .X(_1079_));
 sky130_fd_sc_hd__clkbuf_1 _2733_ (.A(_1079_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2734_ (.A0(\po_0.regf_0.rf[12][15] ),
    .A1(_0982_),
    .S(_1062_),
    .X(_1080_));
 sky130_fd_sc_hd__clkbuf_1 _2735_ (.A(_1080_),
    .X(_0159_));
 sky130_fd_sc_hd__and4b_4 _2736_ (.A_N(\po_0.regf_0.w_addr[2] ),
    .B(_0927_),
    .C(\po_0.regf_0.w_wr ),
    .D(_0928_),
    .X(_1081_));
 sky130_fd_sc_hd__clkbuf_4 _2737_ (.A(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__mux2_1 _2738_ (.A0(\po_0.regf_0.rf[11][0] ),
    .A1(_0949_),
    .S(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__clkbuf_1 _2739_ (.A(_1083_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2740_ (.A0(\po_0.regf_0.rf[11][1] ),
    .A1(_0953_),
    .S(_1082_),
    .X(_1084_));
 sky130_fd_sc_hd__clkbuf_1 _2741_ (.A(_1084_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2742_ (.A0(\po_0.regf_0.rf[11][2] ),
    .A1(_0955_),
    .S(_1082_),
    .X(_1085_));
 sky130_fd_sc_hd__clkbuf_1 _2743_ (.A(_1085_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2744_ (.A0(\po_0.regf_0.rf[11][3] ),
    .A1(_0957_),
    .S(_1082_),
    .X(_1086_));
 sky130_fd_sc_hd__clkbuf_1 _2745_ (.A(_1086_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2746_ (.A0(\po_0.regf_0.rf[11][4] ),
    .A1(_0959_),
    .S(_1082_),
    .X(_1087_));
 sky130_fd_sc_hd__clkbuf_1 _2747_ (.A(_1087_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(\po_0.regf_0.rf[11][5] ),
    .A1(_0961_),
    .S(_1082_),
    .X(_1088_));
 sky130_fd_sc_hd__clkbuf_1 _2749_ (.A(_1088_),
    .X(_0165_));
 sky130_fd_sc_hd__buf_2 _2750_ (.A(_1081_),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(\po_0.regf_0.rf[11][6] ),
    .A1(_0963_),
    .S(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__clkbuf_1 _2752_ (.A(_1090_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2753_ (.A0(\po_0.regf_0.rf[11][7] ),
    .A1(_0966_),
    .S(_1089_),
    .X(_1091_));
 sky130_fd_sc_hd__clkbuf_1 _2754_ (.A(_1091_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2755_ (.A0(\po_0.regf_0.rf[11][8] ),
    .A1(_0968_),
    .S(_1089_),
    .X(_1092_));
 sky130_fd_sc_hd__clkbuf_1 _2756_ (.A(_1092_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(\po_0.regf_0.rf[11][9] ),
    .A1(_0970_),
    .S(_1089_),
    .X(_1093_));
 sky130_fd_sc_hd__clkbuf_1 _2758_ (.A(_1093_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _2759_ (.A0(\po_0.regf_0.rf[11][10] ),
    .A1(_0972_),
    .S(_1089_),
    .X(_1094_));
 sky130_fd_sc_hd__clkbuf_1 _2760_ (.A(_1094_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2761_ (.A0(\po_0.regf_0.rf[11][11] ),
    .A1(_0974_),
    .S(_1089_),
    .X(_1095_));
 sky130_fd_sc_hd__clkbuf_1 _2762_ (.A(_1095_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _2763_ (.A0(\po_0.regf_0.rf[11][12] ),
    .A1(_0976_),
    .S(_1081_),
    .X(_1096_));
 sky130_fd_sc_hd__clkbuf_1 _2764_ (.A(_1096_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2765_ (.A0(\po_0.regf_0.rf[11][13] ),
    .A1(_0978_),
    .S(_1081_),
    .X(_1097_));
 sky130_fd_sc_hd__clkbuf_1 _2766_ (.A(_1097_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2767_ (.A0(\po_0.regf_0.rf[11][14] ),
    .A1(_0980_),
    .S(_1081_),
    .X(_1098_));
 sky130_fd_sc_hd__clkbuf_1 _2768_ (.A(_1098_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _2769_ (.A0(\po_0.regf_0.rf[11][15] ),
    .A1(_0982_),
    .S(_1081_),
    .X(_1099_));
 sky130_fd_sc_hd__clkbuf_1 _2770_ (.A(_1099_),
    .X(_0175_));
 sky130_fd_sc_hd__and4b_4 _2771_ (.A_N(\po_0.regf_0.w_addr[2] ),
    .B(_0737_),
    .C(\po_0.regf_0.w_wr ),
    .D(_0907_),
    .X(_1100_));
 sky130_fd_sc_hd__buf_2 _2772_ (.A(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__mux2_1 _2773_ (.A0(\po_0.regf_0.rf[10][0] ),
    .A1(_0949_),
    .S(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__clkbuf_1 _2774_ (.A(_1102_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2775_ (.A0(\po_0.regf_0.rf[10][1] ),
    .A1(_0953_),
    .S(_1101_),
    .X(_1103_));
 sky130_fd_sc_hd__clkbuf_1 _2776_ (.A(_1103_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2777_ (.A0(\po_0.regf_0.rf[10][2] ),
    .A1(_0955_),
    .S(_1101_),
    .X(_1104_));
 sky130_fd_sc_hd__clkbuf_1 _2778_ (.A(_1104_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2779_ (.A0(\po_0.regf_0.rf[10][3] ),
    .A1(_0957_),
    .S(_1101_),
    .X(_1105_));
 sky130_fd_sc_hd__clkbuf_1 _2780_ (.A(_1105_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _2781_ (.A0(\po_0.regf_0.rf[10][4] ),
    .A1(_0959_),
    .S(_1101_),
    .X(_1106_));
 sky130_fd_sc_hd__clkbuf_1 _2782_ (.A(_1106_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2783_ (.A0(\po_0.regf_0.rf[10][5] ),
    .A1(_0961_),
    .S(_1101_),
    .X(_1107_));
 sky130_fd_sc_hd__clkbuf_1 _2784_ (.A(_1107_),
    .X(_0181_));
 sky130_fd_sc_hd__buf_2 _2785_ (.A(_1100_),
    .X(_1108_));
 sky130_fd_sc_hd__mux2_1 _2786_ (.A0(\po_0.regf_0.rf[10][6] ),
    .A1(_0963_),
    .S(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__clkbuf_1 _2787_ (.A(_1109_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2788_ (.A0(\po_0.regf_0.rf[10][7] ),
    .A1(_0966_),
    .S(_1108_),
    .X(_1110_));
 sky130_fd_sc_hd__clkbuf_1 _2789_ (.A(_1110_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2790_ (.A0(\po_0.regf_0.rf[10][8] ),
    .A1(_0968_),
    .S(_1108_),
    .X(_1111_));
 sky130_fd_sc_hd__clkbuf_1 _2791_ (.A(_1111_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _2792_ (.A0(\po_0.regf_0.rf[10][9] ),
    .A1(_0970_),
    .S(_1108_),
    .X(_1112_));
 sky130_fd_sc_hd__clkbuf_1 _2793_ (.A(_1112_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _2794_ (.A0(\po_0.regf_0.rf[10][10] ),
    .A1(_0972_),
    .S(_1108_),
    .X(_1113_));
 sky130_fd_sc_hd__clkbuf_1 _2795_ (.A(_1113_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2796_ (.A0(\po_0.regf_0.rf[10][11] ),
    .A1(_0974_),
    .S(_1108_),
    .X(_1114_));
 sky130_fd_sc_hd__clkbuf_1 _2797_ (.A(_1114_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _2798_ (.A0(\po_0.regf_0.rf[10][12] ),
    .A1(_0976_),
    .S(_1100_),
    .X(_1115_));
 sky130_fd_sc_hd__clkbuf_1 _2799_ (.A(_1115_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _2800_ (.A0(\po_0.regf_0.rf[10][13] ),
    .A1(_0978_),
    .S(_1100_),
    .X(_1116_));
 sky130_fd_sc_hd__clkbuf_1 _2801_ (.A(_1116_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(\po_0.regf_0.rf[10][14] ),
    .A1(_0980_),
    .S(_1100_),
    .X(_1117_));
 sky130_fd_sc_hd__clkbuf_1 _2803_ (.A(_1117_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _2804_ (.A0(\po_0.regf_0.rf[10][15] ),
    .A1(_0982_),
    .S(_1100_),
    .X(_1118_));
 sky130_fd_sc_hd__clkbuf_1 _2805_ (.A(_1118_),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_2 _2806_ (.A(\uc_0._01_ ),
    .X(_1119_));
 sky130_fd_sc_hd__nor2_2 _2807_ (.A(\uc_0._00_ ),
    .B(\uc_0._02_ ),
    .Y(_1120_));
 sky130_fd_sc_hd__clkbuf_2 _2808_ (.A(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__clkbuf_2 _2809_ (.A(net61),
    .X(_1122_));
 sky130_fd_sc_hd__clkbuf_2 _2810_ (.A(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__clkbuf_2 _2811_ (.A(\uc_0._21_[0] ),
    .X(_1124_));
 sky130_fd_sc_hd__xnor2_1 _2812_ (.A(_1123_),
    .B(_1124_),
    .Y(_1125_));
 sky130_fd_sc_hd__clkbuf_2 _2813_ (.A(\uc_0._02_ ),
    .X(_1126_));
 sky130_fd_sc_hd__clkbuf_2 _2814_ (.A(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__clkbuf_2 _2815_ (.A(\uc_0._00_ ),
    .X(_1128_));
 sky130_fd_sc_hd__clkbuf_2 _2816_ (.A(\uc_0._02_ ),
    .X(_1129_));
 sky130_fd_sc_hd__nor3_2 _2817_ (.A(\uc_0._01_ ),
    .B(_1128_),
    .C(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__buf_2 _2818_ (.A(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__mux2_1 _2819_ (.A0(_1127_),
    .A1(_1131_),
    .S(_1123_),
    .X(_1132_));
 sky130_fd_sc_hd__a31o_1 _2820_ (.A1(_1119_),
    .A2(_1121_),
    .A3(_1125_),
    .B1(_1132_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_2 _2821_ (.A(net99),
    .X(_1133_));
 sky130_fd_sc_hd__or3_2 _2822_ (.A(_1119_),
    .B(_1128_),
    .C(_1126_),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_2 _2823_ (.A(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_2 _2824_ (.A(\uc_0._21_[1] ),
    .X(_1136_));
 sky130_fd_sc_hd__nor2_1 _2825_ (.A(net99),
    .B(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__and2_1 _2826_ (.A(net99),
    .B(\uc_0._21_[1] ),
    .X(_1138_));
 sky130_fd_sc_hd__or4_1 _2827_ (.A(_1122_),
    .B(_1124_),
    .C(_1137_),
    .D(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__o22ai_1 _2828_ (.A1(_1122_),
    .A2(\uc_0._21_[0] ),
    .B1(_1137_),
    .B2(_1138_),
    .Y(_1140_));
 sky130_fd_sc_hd__a21boi_1 _2829_ (.A1(_1122_),
    .A2(net99),
    .B1_N(_1129_),
    .Y(_1141_));
 sky130_fd_sc_hd__o22a_1 _2830_ (.A1(_1123_),
    .A2(_1133_),
    .B1(_1130_),
    .B2(_1141_),
    .X(_1142_));
 sky130_fd_sc_hd__a31o_1 _2831_ (.A1(_1139_),
    .A2(_1121_),
    .A3(_1140_),
    .B1(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__o21a_1 _2832_ (.A1(_1133_),
    .A2(_1135_),
    .B1(_1143_),
    .X(_0193_));
 sky130_fd_sc_hd__clkbuf_2 _2833_ (.A(net69),
    .X(_1144_));
 sky130_fd_sc_hd__a21o_1 _2834_ (.A1(_1123_),
    .A2(_1133_),
    .B1(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__nand3_1 _2835_ (.A(_1123_),
    .B(_1133_),
    .C(_1144_),
    .Y(_1146_));
 sky130_fd_sc_hd__clkbuf_2 _2836_ (.A(_1130_),
    .X(_1147_));
 sky130_fd_sc_hd__a31o_1 _2837_ (.A1(_1145_),
    .A2(_1146_),
    .A3(_1127_),
    .B1(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__o22a_1 _2838_ (.A1(net61),
    .A2(\uc_0._21_[0] ),
    .B1(_1137_),
    .B2(_1138_),
    .X(_1149_));
 sky130_fd_sc_hd__or2_1 _2839_ (.A(net69),
    .B(\uc_0._21_[2] ),
    .X(_1150_));
 sky130_fd_sc_hd__clkbuf_2 _2840_ (.A(\uc_0._21_[2] ),
    .X(_1151_));
 sky130_fd_sc_hd__nand2_1 _2841_ (.A(net69),
    .B(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__a2bb2o_1 _2842_ (.A1_N(net99),
    .A2_N(_1136_),
    .B1(_1150_),
    .B2(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__nand3_1 _2843_ (.A(_1150_),
    .B(_1152_),
    .C(_1137_),
    .Y(_1154_));
 sky130_fd_sc_hd__nand2_1 _2844_ (.A(_1153_),
    .B(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__buf_2 _2845_ (.A(_1128_),
    .X(_1156_));
 sky130_fd_sc_hd__clkbuf_2 _2846_ (.A(_1129_),
    .X(_1157_));
 sky130_fd_sc_hd__a211o_1 _2847_ (.A1(_1140_),
    .A2(_1155_),
    .B1(_1156_),
    .C1(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__a31oi_1 _2848_ (.A1(_1149_),
    .A2(_1153_),
    .A3(_1154_),
    .B1(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__o22a_1 _2849_ (.A1(_1144_),
    .A2(_1135_),
    .B1(_1148_),
    .B2(_1159_),
    .X(_0194_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2850_ (.A(net70),
    .X(_1160_));
 sky130_fd_sc_hd__clkbuf_2 _2851_ (.A(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__and2b_1 _2852_ (.A_N(net70),
    .B(\uc_0._21_[3] ),
    .X(_1162_));
 sky130_fd_sc_hd__clkbuf_2 _2853_ (.A(\uc_0._21_[3] ),
    .X(_1163_));
 sky130_fd_sc_hd__and2b_1 _2854_ (.A_N(_1163_),
    .B(_1160_),
    .X(_1164_));
 sky130_fd_sc_hd__nor2_1 _2855_ (.A(net69),
    .B(_1151_),
    .Y(_1165_));
 sky130_fd_sc_hd__o21ai_1 _2856_ (.A1(_1162_),
    .A2(_1164_),
    .B1(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__nor2_1 _2857_ (.A(_1160_),
    .B(_1163_),
    .Y(_1167_));
 sky130_fd_sc_hd__and2_1 _2858_ (.A(_1160_),
    .B(\uc_0._21_[3] ),
    .X(_1168_));
 sky130_fd_sc_hd__o21ai_1 _2859_ (.A1(_1167_),
    .A2(_1168_),
    .B1(_1150_),
    .Y(_1169_));
 sky130_fd_sc_hd__nand2_1 _2860_ (.A(_1166_),
    .B(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__a21oi_1 _2861_ (.A1(_1150_),
    .A2(_1152_),
    .B1(_1137_),
    .Y(_1171_));
 sky130_fd_sc_hd__a21oi_2 _2862_ (.A1(_1149_),
    .A2(_1154_),
    .B1(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__nor2_1 _2863_ (.A(_1170_),
    .B(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__a211o_1 _2864_ (.A1(_1172_),
    .A2(_1170_),
    .B1(_1128_),
    .C1(_1126_),
    .X(_1174_));
 sky130_fd_sc_hd__and3_1 _2865_ (.A(_1122_),
    .B(net68),
    .C(_1144_),
    .X(_1175_));
 sky130_fd_sc_hd__o21ai_1 _2866_ (.A1(_1161_),
    .A2(_1175_),
    .B1(_1126_),
    .Y(_1176_));
 sky130_fd_sc_hd__a41o_1 _2867_ (.A1(_1123_),
    .A2(_1133_),
    .A3(_1144_),
    .A4(_1161_),
    .B1(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__o211a_1 _2868_ (.A1(_1173_),
    .A2(_1174_),
    .B1(_1177_),
    .C1(_1134_),
    .X(_1178_));
 sky130_fd_sc_hd__o21ba_1 _2869_ (.A1(_1161_),
    .A2(_1135_),
    .B1_N(_1178_),
    .X(_0195_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2870_ (.A(net71),
    .X(_1179_));
 sky130_fd_sc_hd__nand3_1 _2871_ (.A(_1161_),
    .B(_1179_),
    .C(_1175_),
    .Y(_1180_));
 sky130_fd_sc_hd__a41o_1 _2872_ (.A1(_1122_),
    .A2(_1133_),
    .A3(_1144_),
    .A4(_1161_),
    .B1(_1179_),
    .X(_1181_));
 sky130_fd_sc_hd__a31o_1 _2873_ (.A1(_1180_),
    .A2(_1127_),
    .A3(_1181_),
    .B1(_1147_),
    .X(_1182_));
 sky130_fd_sc_hd__o32ai_4 _2874_ (.A1(_1165_),
    .A2(_1162_),
    .A3(_1164_),
    .B1(_1170_),
    .B2(_1172_),
    .Y(_1183_));
 sky130_fd_sc_hd__nand2_1 _2875_ (.A(\uc_0._21_[4] ),
    .B(net71),
    .Y(_1184_));
 sky130_fd_sc_hd__or2_1 _2876_ (.A(\uc_0._21_[4] ),
    .B(net71),
    .X(_1185_));
 sky130_fd_sc_hd__a21oi_2 _2877_ (.A1(_1184_),
    .A2(_1185_),
    .B1(_1167_),
    .Y(_1186_));
 sky130_fd_sc_hd__and3_1 _2878_ (.A(_1185_),
    .B(_1167_),
    .C(_1184_),
    .X(_1187_));
 sky130_fd_sc_hd__nor2_2 _2879_ (.A(_1186_),
    .B(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__and2_1 _2880_ (.A(_1183_),
    .B(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__or3_1 _2881_ (.A(_1128_),
    .B(_1126_),
    .C(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__o21ba_1 _2882_ (.A1(_1183_),
    .A2(_1188_),
    .B1_N(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__o22a_1 _2883_ (.A1(_1179_),
    .A2(_1135_),
    .B1(_1182_),
    .B2(_1191_),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _2884_ (.A(\uc_0._21_[5] ),
    .B(net72),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_2 _2885_ (.A(net72),
    .X(_1193_));
 sky130_fd_sc_hd__nand2_1 _2886_ (.A(\uc_0._21_[5] ),
    .B(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__nand2_1 _2887_ (.A(_1192_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__o21ai_1 _2888_ (.A1(\uc_0._21_[4] ),
    .A2(net71),
    .B1(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__nand3b_1 _2889_ (.A_N(_1185_),
    .B(_1192_),
    .C(_1194_),
    .Y(_1197_));
 sky130_fd_sc_hd__and2_1 _2890_ (.A(_1196_),
    .B(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__o21ai_1 _2891_ (.A1(_1186_),
    .A2(_1189_),
    .B1(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__a221o_1 _2892_ (.A1(_1196_),
    .A2(_1197_),
    .B1(_1183_),
    .B2(_1188_),
    .C1(_1186_),
    .X(_1200_));
 sky130_fd_sc_hd__and4_1 _2893_ (.A(_1160_),
    .B(_1179_),
    .C(_1193_),
    .D(_1175_),
    .X(_1201_));
 sky130_fd_sc_hd__a31o_1 _2894_ (.A1(_1160_),
    .A2(_1179_),
    .A3(_1175_),
    .B1(_1193_),
    .X(_1202_));
 sky130_fd_sc_hd__and3b_1 _2895_ (.A_N(_1201_),
    .B(_1202_),
    .C(_1129_),
    .X(_1203_));
 sky130_fd_sc_hd__a31o_1 _2896_ (.A1(_1199_),
    .A2(_1120_),
    .A3(_1200_),
    .B1(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__mux2_1 _2897_ (.A0(_1204_),
    .A1(_1193_),
    .S(_1131_),
    .X(_1205_));
 sky130_fd_sc_hd__clkbuf_1 _2898_ (.A(_1205_),
    .X(_0197_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2899_ (.A(net73),
    .X(_1206_));
 sky130_fd_sc_hd__nand2_1 _2900_ (.A(_1206_),
    .B(_1201_),
    .Y(_1207_));
 sky130_fd_sc_hd__a41o_1 _2901_ (.A1(_1161_),
    .A2(_1179_),
    .A3(_1193_),
    .A4(_1175_),
    .B1(_1206_),
    .X(_1208_));
 sky130_fd_sc_hd__a31o_1 _2902_ (.A1(_1207_),
    .A2(_1127_),
    .A3(_1208_),
    .B1(_1147_),
    .X(_1209_));
 sky130_fd_sc_hd__nand2_1 _2903_ (.A(\uc_0._21_[6] ),
    .B(net73),
    .Y(_1210_));
 sky130_fd_sc_hd__or2_1 _2904_ (.A(\uc_0._21_[6] ),
    .B(net73),
    .X(_1211_));
 sky130_fd_sc_hd__a21oi_1 _2905_ (.A1(_1210_),
    .A2(_1211_),
    .B1(_1192_),
    .Y(_1212_));
 sky130_fd_sc_hd__and3_1 _2906_ (.A(_1192_),
    .B(_1210_),
    .C(_1211_),
    .X(_1213_));
 sky130_fd_sc_hd__nor2_1 _2907_ (.A(_1212_),
    .B(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__o21a_1 _2908_ (.A1(_1549_),
    .A2(net71),
    .B1(_1195_),
    .X(_1215_));
 sky130_fd_sc_hd__o21a_1 _2909_ (.A1(_1186_),
    .A2(_1215_),
    .B1(_1197_),
    .X(_1216_));
 sky130_fd_sc_hd__a31oi_4 _2910_ (.A1(_1183_),
    .A2(_1188_),
    .A3(_1198_),
    .B1(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__nor2_1 _2911_ (.A(_1214_),
    .B(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__a211o_1 _2912_ (.A1(_1217_),
    .A2(_1214_),
    .B1(_1156_),
    .C1(_1127_),
    .X(_1219_));
 sky130_fd_sc_hd__nor2_1 _2913_ (.A(_1218_),
    .B(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__o22a_1 _2914_ (.A1(_1206_),
    .A2(_1134_),
    .B1(_1209_),
    .B2(_1220_),
    .X(_0198_));
 sky130_fd_sc_hd__nor2_1 _2915_ (.A(\uc_0._21_[7] ),
    .B(net74),
    .Y(_1221_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2916_ (.A(net74),
    .X(_1222_));
 sky130_fd_sc_hd__nand2_1 _2917_ (.A(_1559_),
    .B(_1222_),
    .Y(_1223_));
 sky130_fd_sc_hd__or4b_2 _2918_ (.A(\uc_0._21_[6] ),
    .B(net73),
    .C(_1221_),
    .D_N(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__or2_1 _2919_ (.A(\uc_0._21_[7] ),
    .B(_1222_),
    .X(_1225_));
 sky130_fd_sc_hd__a2bb2o_1 _2920_ (.A1_N(_1557_),
    .A2_N(net73),
    .B1(_1225_),
    .B2(_1223_),
    .X(_1226_));
 sky130_fd_sc_hd__a21boi_1 _2921_ (.A1(_1210_),
    .A2(_1211_),
    .B1_N(_1192_),
    .Y(_1227_));
 sky130_fd_sc_hd__a211oi_1 _2922_ (.A1(_1224_),
    .A2(_1226_),
    .B1(_1227_),
    .C1(_1218_),
    .Y(_1228_));
 sky130_fd_sc_hd__o211a_1 _2923_ (.A1(_1227_),
    .A2(_1218_),
    .B1(_1224_),
    .C1(_1226_),
    .X(_1229_));
 sky130_fd_sc_hd__and3_1 _2924_ (.A(_1206_),
    .B(_1222_),
    .C(_1201_),
    .X(_1230_));
 sky130_fd_sc_hd__a21oi_1 _2925_ (.A1(_1206_),
    .A2(_1201_),
    .B1(_1222_),
    .Y(_1231_));
 sky130_fd_sc_hd__or3b_1 _2926_ (.A(_1230_),
    .B(_1231_),
    .C_N(_1129_),
    .X(_1232_));
 sky130_fd_sc_hd__o41ai_1 _2927_ (.A1(_1128_),
    .A2(_1157_),
    .A3(_1228_),
    .A4(_1229_),
    .B1(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__mux2_1 _2928_ (.A0(_1233_),
    .A1(_1222_),
    .S(_1131_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _2929_ (.A(_1234_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_2 _2930_ (.A(net75),
    .X(_1235_));
 sky130_fd_sc_hd__o21ai_1 _2931_ (.A1(_1235_),
    .A2(_1230_),
    .B1(_1126_),
    .Y(_1236_));
 sky130_fd_sc_hd__and4_1 _2932_ (.A(_1206_),
    .B(_1222_),
    .C(net75),
    .D(_1201_),
    .X(_1237_));
 sky130_fd_sc_hd__o211ai_2 _2933_ (.A1(_1212_),
    .A2(_1213_),
    .B1(_1224_),
    .C1(_1226_),
    .Y(_1238_));
 sky130_fd_sc_hd__a2bb2o_1 _2934_ (.A1_N(_1555_),
    .A2_N(_1193_),
    .B1(_1210_),
    .B2(_1211_),
    .X(_1239_));
 sky130_fd_sc_hd__a21bo_1 _2935_ (.A1(_1239_),
    .A2(_1226_),
    .B1_N(_1224_),
    .X(_1240_));
 sky130_fd_sc_hd__o21ai_4 _2936_ (.A1(_1238_),
    .A2(_1217_),
    .B1(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__xor2_1 _2937_ (.A(net75),
    .B(_1221_),
    .X(_1242_));
 sky130_fd_sc_hd__nand2_1 _2938_ (.A(_1241_),
    .B(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__o21a_1 _2939_ (.A1(_1242_),
    .A2(_1241_),
    .B1(_1120_),
    .X(_1244_));
 sky130_fd_sc_hd__a2bb2o_1 _2940_ (.A1_N(_1236_),
    .A2_N(_1237_),
    .B1(_1243_),
    .B2(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_1 _2941_ (.A0(_1245_),
    .A1(_1235_),
    .S(_1131_),
    .X(_1246_));
 sky130_fd_sc_hd__clkbuf_1 _2942_ (.A(_1246_),
    .X(_0200_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2943_ (.A(net98),
    .X(_1247_));
 sky130_fd_sc_hd__buf_2 _2944_ (.A(_1157_),
    .X(_1248_));
 sky130_fd_sc_hd__and2_1 _2945_ (.A(net75),
    .B(net98),
    .X(_1249_));
 sky130_fd_sc_hd__o2bb2a_1 _2946_ (.A1_N(_1230_),
    .A2_N(_1249_),
    .B1(_1237_),
    .B2(_1247_),
    .X(_1250_));
 sky130_fd_sc_hd__a21o_1 _2947_ (.A1(_1248_),
    .A2(_1250_),
    .B1(_1147_),
    .X(_1251_));
 sky130_fd_sc_hd__o21a_1 _2948_ (.A1(_1235_),
    .A2(_1221_),
    .B1(_1243_),
    .X(_1252_));
 sky130_fd_sc_hd__nor2_1 _2949_ (.A(net75),
    .B(net98),
    .Y(_1253_));
 sky130_fd_sc_hd__nor2_1 _2950_ (.A(_1249_),
    .B(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__o21a_1 _2951_ (.A1(_1252_),
    .A2(_1254_),
    .B1(_1120_),
    .X(_1255_));
 sky130_fd_sc_hd__a21boi_1 _2952_ (.A1(_1252_),
    .A2(_1254_),
    .B1_N(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__o22a_1 _2953_ (.A1(_1247_),
    .A2(_1134_),
    .B1(_1251_),
    .B2(_1256_),
    .X(_0201_));
 sky130_fd_sc_hd__xnor2_1 _2954_ (.A(net98),
    .B(net62),
    .Y(_1257_));
 sky130_fd_sc_hd__o21a_1 _2955_ (.A1(_1249_),
    .A2(_1253_),
    .B1(_1242_),
    .X(_1258_));
 sky130_fd_sc_hd__nor2_1 _2956_ (.A(_1235_),
    .B(_1225_),
    .Y(_1259_));
 sky130_fd_sc_hd__o2bb2ai_1 _2957_ (.A1_N(_1258_),
    .A2_N(_1241_),
    .B1(_1247_),
    .B2(_1259_),
    .Y(_1260_));
 sky130_fd_sc_hd__or2_1 _2958_ (.A(_1257_),
    .B(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__nand2_1 _2959_ (.A(_1257_),
    .B(_1260_),
    .Y(_1262_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2960_ (.A(net62),
    .X(_1263_));
 sky130_fd_sc_hd__and3_2 _2961_ (.A(net98),
    .B(_1263_),
    .C(_1237_),
    .X(_1264_));
 sky130_fd_sc_hd__a31o_1 _2962_ (.A1(_1235_),
    .A2(_1247_),
    .A3(_1230_),
    .B1(_1263_),
    .X(_1265_));
 sky130_fd_sc_hd__and3b_1 _2963_ (.A_N(_1264_),
    .B(_1129_),
    .C(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__a31o_1 _2964_ (.A1(_1261_),
    .A2(_1120_),
    .A3(_1262_),
    .B1(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__mux2_1 _2965_ (.A0(_1267_),
    .A1(_1263_),
    .S(_1131_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_1 _2966_ (.A(_1268_),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_2 _2967_ (.A(net97),
    .X(_1269_));
 sky130_fd_sc_hd__or2b_1 _2968_ (.A(_1263_),
    .B_N(_1247_),
    .X(_1270_));
 sky130_fd_sc_hd__xnor2_1 _2969_ (.A(net62),
    .B(net97),
    .Y(_1271_));
 sky130_fd_sc_hd__a21bo_1 _2970_ (.A1(_1262_),
    .A2(_1270_),
    .B1_N(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__nand3b_1 _2971_ (.A_N(_1271_),
    .B(_1270_),
    .C(_1262_),
    .Y(_1273_));
 sky130_fd_sc_hd__and4_1 _2972_ (.A(_1247_),
    .B(_1263_),
    .C(_1269_),
    .D(_1237_),
    .X(_1274_));
 sky130_fd_sc_hd__o21ai_1 _2973_ (.A1(_1269_),
    .A2(_1264_),
    .B1(_1157_),
    .Y(_1275_));
 sky130_fd_sc_hd__o21ai_1 _2974_ (.A1(_1274_),
    .A2(_1275_),
    .B1(_1134_),
    .Y(_1276_));
 sky130_fd_sc_hd__a31o_1 _2975_ (.A1(_1272_),
    .A2(_1273_),
    .A3(_1121_),
    .B1(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__o41a_1 _2976_ (.A1(_1119_),
    .A2(_1156_),
    .A3(_1248_),
    .A4(_1269_),
    .B1(_1277_),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_2 _2977_ (.A(net96),
    .X(_1278_));
 sky130_fd_sc_hd__and3_1 _2978_ (.A(_1258_),
    .B(_1271_),
    .C(_1257_),
    .X(_1279_));
 sky130_fd_sc_hd__nor4_1 _2979_ (.A(_1235_),
    .B(net98),
    .C(_1263_),
    .D(_1225_),
    .Y(_1280_));
 sky130_fd_sc_hd__nor2_1 _2980_ (.A(net97),
    .B(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__nor2_1 _2981_ (.A(net97),
    .B(net96),
    .Y(_1282_));
 sky130_fd_sc_hd__and2_1 _2982_ (.A(net97),
    .B(net96),
    .X(_1283_));
 sky130_fd_sc_hd__a2111o_1 _2983_ (.A1(_1241_),
    .A2(_1279_),
    .B1(_1281_),
    .C1(_1282_),
    .D1(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__a21o_1 _2984_ (.A1(_1241_),
    .A2(_1279_),
    .B1(_1281_),
    .X(_1285_));
 sky130_fd_sc_hd__o21ai_1 _2985_ (.A1(_1283_),
    .A2(_1282_),
    .B1(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__nand2_1 _2986_ (.A(_1264_),
    .B(_1283_),
    .Y(_1287_));
 sky130_fd_sc_hd__o211a_1 _2987_ (.A1(_1278_),
    .A2(_1274_),
    .B1(_1157_),
    .C1(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__a311o_1 _2988_ (.A1(_1284_),
    .A2(_1286_),
    .A3(_1121_),
    .B1(_1288_),
    .C1(_1131_),
    .X(_1289_));
 sky130_fd_sc_hd__o41a_1 _2989_ (.A1(_1119_),
    .A2(_1156_),
    .A3(_1248_),
    .A4(_1278_),
    .B1(_1289_),
    .X(_0204_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2990_ (.A(net95),
    .X(_1290_));
 sky130_fd_sc_hd__or2b_1 _2991_ (.A(net96),
    .B_N(_1269_),
    .X(_1291_));
 sky130_fd_sc_hd__nand2_1 _2992_ (.A(net96),
    .B(net95),
    .Y(_1292_));
 sky130_fd_sc_hd__or2_1 _2993_ (.A(net64),
    .B(net95),
    .X(_1293_));
 sky130_fd_sc_hd__a22o_1 _2994_ (.A1(_1286_),
    .A2(_1291_),
    .B1(_1292_),
    .B2(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__nand4_1 _2995_ (.A(_1286_),
    .B(_1291_),
    .C(_1292_),
    .D(_1293_),
    .Y(_1295_));
 sky130_fd_sc_hd__a31o_1 _2996_ (.A1(_1269_),
    .A2(_1278_),
    .A3(_1264_),
    .B1(net95),
    .X(_1296_));
 sky130_fd_sc_hd__nand4_1 _2997_ (.A(_1269_),
    .B(_1278_),
    .C(_1290_),
    .D(_1264_),
    .Y(_1297_));
 sky130_fd_sc_hd__a31o_1 _2998_ (.A1(_1296_),
    .A2(_1297_),
    .A3(_1157_),
    .B1(_1130_),
    .X(_1298_));
 sky130_fd_sc_hd__a31o_1 _2999_ (.A1(_1294_),
    .A2(_1121_),
    .A3(_1295_),
    .B1(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__o41a_1 _3000_ (.A1(_1119_),
    .A2(_1156_),
    .A3(_1248_),
    .A4(_1290_),
    .B1(_1299_),
    .X(_0205_));
 sky130_fd_sc_hd__a31o_1 _3001_ (.A1(_1278_),
    .A2(_1290_),
    .A3(_1274_),
    .B1(net94),
    .X(_1300_));
 sky130_fd_sc_hd__nand4_1 _3002_ (.A(_1278_),
    .B(_1290_),
    .C(net94),
    .D(_1274_),
    .Y(_1301_));
 sky130_fd_sc_hd__a31oi_1 _3003_ (.A1(_1300_),
    .A2(_1301_),
    .A3(_1248_),
    .B1(_1147_),
    .Y(_1302_));
 sky130_fd_sc_hd__xnor2_1 _3004_ (.A(net65),
    .B(net94),
    .Y(_1303_));
 sky130_fd_sc_hd__a2bb2o_1 _3005_ (.A1_N(_1283_),
    .A2_N(_1282_),
    .B1(_1292_),
    .B2(_1293_),
    .X(_1304_));
 sky130_fd_sc_hd__a2bb2oi_1 _3006_ (.A1_N(net63),
    .A2_N(_1280_),
    .B1(_1279_),
    .B2(_1241_),
    .Y(_1305_));
 sky130_fd_sc_hd__o22ai_2 _3007_ (.A1(net95),
    .A2(_1282_),
    .B1(_1304_),
    .B2(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__o21a_1 _3008_ (.A1(_1303_),
    .A2(_1306_),
    .B1(_1120_),
    .X(_1307_));
 sky130_fd_sc_hd__nand2_1 _3009_ (.A(_1306_),
    .B(_1303_),
    .Y(_1308_));
 sky130_fd_sc_hd__nand2_1 _3010_ (.A(_1307_),
    .B(_1308_),
    .Y(_1309_));
 sky130_fd_sc_hd__o2bb2a_1 _3011_ (.A1_N(_1302_),
    .A2_N(_1309_),
    .B1(_1135_),
    .B2(net94),
    .X(_0206_));
 sky130_fd_sc_hd__xor2_1 _3012_ (.A(net94),
    .B(net67),
    .X(_1310_));
 sky130_fd_sc_hd__a31o_1 _3013_ (.A1(_1290_),
    .A2(_1264_),
    .A3(_1283_),
    .B1(net67),
    .X(_1311_));
 sky130_fd_sc_hd__o211a_1 _3014_ (.A1(_1297_),
    .A2(_1310_),
    .B1(_1127_),
    .C1(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__nor2_1 _3015_ (.A(_1147_),
    .B(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__or2b_1 _3016_ (.A(net66),
    .B_N(_1290_),
    .X(_1314_));
 sky130_fd_sc_hd__a21o_1 _3017_ (.A1(_1314_),
    .A2(_1308_),
    .B1(_1310_),
    .X(_1315_));
 sky130_fd_sc_hd__nand3_1 _3018_ (.A(_1314_),
    .B(_1308_),
    .C(_1310_),
    .Y(_1316_));
 sky130_fd_sc_hd__nand3_1 _3019_ (.A(_1315_),
    .B(_1121_),
    .C(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__a2bb2oi_1 _3020_ (.A1_N(net67),
    .A2_N(_1135_),
    .B1(_1313_),
    .B2(_1317_),
    .Y(_0207_));
 sky130_fd_sc_hd__and4b_4 _3021_ (.A_N(_0737_),
    .B(_0906_),
    .C(_1061_),
    .D(_0742_),
    .X(_1318_));
 sky130_fd_sc_hd__buf_2 _3022_ (.A(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__mux2_1 _3023_ (.A0(\po_0.regf_0.rf[4][0] ),
    .A1(_0735_),
    .S(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__clkbuf_1 _3024_ (.A(_1320_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _3025_ (.A0(\po_0.regf_0.rf[4][1] ),
    .A1(_0755_),
    .S(_1319_),
    .X(_1321_));
 sky130_fd_sc_hd__clkbuf_1 _3026_ (.A(_1321_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _3027_ (.A0(\po_0.regf_0.rf[4][2] ),
    .A1(_0767_),
    .S(_1319_),
    .X(_1322_));
 sky130_fd_sc_hd__clkbuf_1 _3028_ (.A(_1322_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _3029_ (.A0(\po_0.regf_0.rf[4][3] ),
    .A1(_0777_),
    .S(_1319_),
    .X(_1323_));
 sky130_fd_sc_hd__clkbuf_1 _3030_ (.A(_1323_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _3031_ (.A0(\po_0.regf_0.rf[4][4] ),
    .A1(_0788_),
    .S(_1319_),
    .X(_1324_));
 sky130_fd_sc_hd__clkbuf_1 _3032_ (.A(_1324_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _3033_ (.A0(\po_0.regf_0.rf[4][5] ),
    .A1(_0796_),
    .S(_1319_),
    .X(_1325_));
 sky130_fd_sc_hd__clkbuf_1 _3034_ (.A(_1325_),
    .X(_0213_));
 sky130_fd_sc_hd__buf_2 _3035_ (.A(_1318_),
    .X(_1326_));
 sky130_fd_sc_hd__mux2_1 _3036_ (.A0(\po_0.regf_0.rf[4][6] ),
    .A1(_0808_),
    .S(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__clkbuf_1 _3037_ (.A(_1327_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _3038_ (.A0(\po_0.regf_0.rf[4][7] ),
    .A1(_0820_),
    .S(_1326_),
    .X(_1328_));
 sky130_fd_sc_hd__clkbuf_1 _3039_ (.A(_1328_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _3040_ (.A0(\po_0.regf_0.rf[4][8] ),
    .A1(_0835_),
    .S(_1326_),
    .X(_1329_));
 sky130_fd_sc_hd__clkbuf_1 _3041_ (.A(_1329_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _3042_ (.A0(\po_0.regf_0.rf[4][9] ),
    .A1(_0843_),
    .S(_1326_),
    .X(_1330_));
 sky130_fd_sc_hd__clkbuf_1 _3043_ (.A(_1330_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _3044_ (.A0(\po_0.regf_0.rf[4][10] ),
    .A1(_0852_),
    .S(_1326_),
    .X(_1331_));
 sky130_fd_sc_hd__clkbuf_1 _3045_ (.A(_1331_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _3046_ (.A0(\po_0.regf_0.rf[4][11] ),
    .A1(_0861_),
    .S(_1326_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_1 _3047_ (.A(_1332_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _3048_ (.A0(\po_0.regf_0.rf[4][12] ),
    .A1(_0873_),
    .S(_1318_),
    .X(_1333_));
 sky130_fd_sc_hd__clkbuf_1 _3049_ (.A(_1333_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _3050_ (.A0(\po_0.regf_0.rf[4][13] ),
    .A1(_0882_),
    .S(_1318_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_1 _3051_ (.A(_1334_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(\po_0.regf_0.rf[4][14] ),
    .A1(_0895_),
    .S(_1318_),
    .X(_1335_));
 sky130_fd_sc_hd__clkbuf_1 _3053_ (.A(_1335_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _3054_ (.A0(\po_0.regf_0.rf[4][15] ),
    .A1(_0903_),
    .S(_1318_),
    .X(_1336_));
 sky130_fd_sc_hd__clkbuf_1 _3055_ (.A(_1336_),
    .X(_0223_));
 sky130_fd_sc_hd__buf_2 _3056_ (.A(\uc_0._03_ ),
    .X(_1337_));
 sky130_fd_sc_hd__mux2_1 _3057_ (.A0(_1124_),
    .A1(net17),
    .S(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__clkbuf_1 _3058_ (.A(_1338_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(_1136_),
    .A1(net24),
    .S(_1337_),
    .X(_1339_));
 sky130_fd_sc_hd__clkbuf_1 _3060_ (.A(_1339_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(_1151_),
    .A1(net25),
    .S(_1337_),
    .X(_1340_));
 sky130_fd_sc_hd__clkbuf_1 _3062_ (.A(_1340_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _3063_ (.A0(_1163_),
    .A1(net26),
    .S(_1337_),
    .X(_1341_));
 sky130_fd_sc_hd__clkbuf_1 _3064_ (.A(_1341_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _3065_ (.A0(_1549_),
    .A1(net27),
    .S(_1337_),
    .X(_1342_));
 sky130_fd_sc_hd__clkbuf_1 _3066_ (.A(_1342_),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_4 _3067_ (.A(\uc_0._03_ ),
    .X(_1343_));
 sky130_fd_sc_hd__buf_2 _3068_ (.A(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__mux2_1 _3069_ (.A0(_1555_),
    .A1(net28),
    .S(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__clkbuf_1 _3070_ (.A(_1345_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _3071_ (.A0(_1557_),
    .A1(net29),
    .S(_1344_),
    .X(_1346_));
 sky130_fd_sc_hd__clkbuf_1 _3072_ (.A(_1346_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _3073_ (.A0(_1559_),
    .A1(net30),
    .S(_1344_),
    .X(_1347_));
 sky130_fd_sc_hd__clkbuf_1 _3074_ (.A(_1347_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _3075_ (.A0(\uc_0._21_[8] ),
    .A1(net31),
    .S(_1344_),
    .X(_1348_));
 sky130_fd_sc_hd__clkbuf_1 _3076_ (.A(_1348_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _3077_ (.A0(\uc_0._21_[9] ),
    .A1(net32),
    .S(_1344_),
    .X(_1349_));
 sky130_fd_sc_hd__clkbuf_1 _3078_ (.A(_1349_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _3079_ (.A0(\uc_0._21_[10] ),
    .A1(net18),
    .S(_1344_),
    .X(_1350_));
 sky130_fd_sc_hd__clkbuf_1 _3080_ (.A(_1350_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _3081_ (.A0(\uc_0._21_[11] ),
    .A1(net19),
    .S(_1343_),
    .X(_1351_));
 sky130_fd_sc_hd__clkbuf_1 _3082_ (.A(_1351_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _3083_ (.A0(\uc_0._21_[12] ),
    .A1(net20),
    .S(_1343_),
    .X(_1352_));
 sky130_fd_sc_hd__clkbuf_1 _3084_ (.A(_1352_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _3085_ (.A0(\uc_0._21_[13] ),
    .A1(net21),
    .S(_1343_),
    .X(_1353_));
 sky130_fd_sc_hd__clkbuf_1 _3086_ (.A(_1353_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _3087_ (.A0(\uc_0._21_[14] ),
    .A1(net22),
    .S(_1343_),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_1 _3088_ (.A(_1354_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _3089_ (.A0(\uc_0._21_[15] ),
    .A1(net23),
    .S(_1343_),
    .X(_1355_));
 sky130_fd_sc_hd__clkbuf_1 _3090_ (.A(_1355_),
    .X(_0239_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3091_ (.A(_1517_),
    .X(_1356_));
 sky130_fd_sc_hd__nand3_1 _3092_ (.A(_1533_),
    .B(_1534_),
    .C(_1537_),
    .Y(_1357_));
 sky130_fd_sc_hd__or3_2 _3093_ (.A(_1356_),
    .B(_1357_),
    .C(_1546_),
    .X(_1358_));
 sky130_fd_sc_hd__o32a_1 _3094_ (.A1(\uc_0.bc_0._70_[2] ),
    .A2(\uc_0.bc_0._70_[3] ),
    .A3(_1358_),
    .B1(_1156_),
    .B2(_1356_),
    .X(_0240_));
 sky130_fd_sc_hd__and4bb_4 _3095_ (.A_N(_0742_),
    .B_N(\po_0.regf_0.w_addr[3] ),
    .C(_0906_),
    .D(_0928_),
    .X(_1359_));
 sky130_fd_sc_hd__clkbuf_4 _3096_ (.A(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__mux2_1 _3097_ (.A0(\po_0.regf_0.rf[3][0] ),
    .A1(_0735_),
    .S(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__clkbuf_1 _3098_ (.A(_1361_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _3099_ (.A0(\po_0.regf_0.rf[3][1] ),
    .A1(_0755_),
    .S(_1360_),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _3100_ (.A(_1362_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(\po_0.regf_0.rf[3][2] ),
    .A1(_0767_),
    .S(_1360_),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_1 _3102_ (.A(_1363_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(\po_0.regf_0.rf[3][3] ),
    .A1(_0777_),
    .S(_1360_),
    .X(_1364_));
 sky130_fd_sc_hd__clkbuf_1 _3104_ (.A(_1364_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _3105_ (.A0(\po_0.regf_0.rf[3][4] ),
    .A1(_0788_),
    .S(_1360_),
    .X(_1365_));
 sky130_fd_sc_hd__clkbuf_1 _3106_ (.A(_1365_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(\po_0.regf_0.rf[3][5] ),
    .A1(_0796_),
    .S(_1360_),
    .X(_1366_));
 sky130_fd_sc_hd__clkbuf_1 _3108_ (.A(_1366_),
    .X(_0246_));
 sky130_fd_sc_hd__buf_2 _3109_ (.A(_1359_),
    .X(_1367_));
 sky130_fd_sc_hd__mux2_1 _3110_ (.A0(\po_0.regf_0.rf[3][6] ),
    .A1(_0808_),
    .S(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__clkbuf_1 _3111_ (.A(_1368_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _3112_ (.A0(\po_0.regf_0.rf[3][7] ),
    .A1(_0820_),
    .S(_1367_),
    .X(_1369_));
 sky130_fd_sc_hd__clkbuf_1 _3113_ (.A(_1369_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _3114_ (.A0(\po_0.regf_0.rf[3][8] ),
    .A1(_0835_),
    .S(_1367_),
    .X(_1370_));
 sky130_fd_sc_hd__clkbuf_1 _3115_ (.A(_1370_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _3116_ (.A0(\po_0.regf_0.rf[3][9] ),
    .A1(_0843_),
    .S(_1367_),
    .X(_1371_));
 sky130_fd_sc_hd__clkbuf_1 _3117_ (.A(_1371_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _3118_ (.A0(\po_0.regf_0.rf[3][10] ),
    .A1(_0852_),
    .S(_1367_),
    .X(_1372_));
 sky130_fd_sc_hd__clkbuf_1 _3119_ (.A(_1372_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _3120_ (.A0(\po_0.regf_0.rf[3][11] ),
    .A1(_0861_),
    .S(_1367_),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_1 _3121_ (.A(_1373_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _3122_ (.A0(\po_0.regf_0.rf[3][12] ),
    .A1(_0873_),
    .S(_1359_),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_1 _3123_ (.A(_1374_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _3124_ (.A0(\po_0.regf_0.rf[3][13] ),
    .A1(_0882_),
    .S(_1359_),
    .X(_1375_));
 sky130_fd_sc_hd__clkbuf_1 _3125_ (.A(_1375_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _3126_ (.A0(\po_0.regf_0.rf[3][14] ),
    .A1(_0895_),
    .S(_1359_),
    .X(_1376_));
 sky130_fd_sc_hd__clkbuf_1 _3127_ (.A(_1376_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _3128_ (.A0(\po_0.regf_0.rf[3][15] ),
    .A1(_0903_),
    .S(_1359_),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_1 _3129_ (.A(_1377_),
    .X(_0256_));
 sky130_fd_sc_hd__or4bb_4 _3130_ (.A(_0929_),
    .B(_0737_),
    .C_N(_0738_),
    .D_N(_1061_),
    .X(_1378_));
 sky130_fd_sc_hd__buf_2 _3131_ (.A(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__mux2_1 _3132_ (.A0(_0736_),
    .A1(\po_0.regf_0.rf[0][0] ),
    .S(_1379_),
    .X(_1380_));
 sky130_fd_sc_hd__clkbuf_1 _3133_ (.A(_1380_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _3134_ (.A0(_0756_),
    .A1(\po_0.regf_0.rf[0][1] ),
    .S(_1379_),
    .X(_1381_));
 sky130_fd_sc_hd__clkbuf_1 _3135_ (.A(_1381_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _3136_ (.A0(_0768_),
    .A1(\po_0.regf_0.rf[0][2] ),
    .S(_1379_),
    .X(_1382_));
 sky130_fd_sc_hd__clkbuf_1 _3137_ (.A(_1382_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _3138_ (.A0(_0778_),
    .A1(\po_0.regf_0.rf[0][3] ),
    .S(_1379_),
    .X(_1383_));
 sky130_fd_sc_hd__clkbuf_1 _3139_ (.A(_1383_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _3140_ (.A0(_0789_),
    .A1(\po_0.regf_0.rf[0][4] ),
    .S(_1379_),
    .X(_1384_));
 sky130_fd_sc_hd__clkbuf_1 _3141_ (.A(_1384_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _3142_ (.A0(_0797_),
    .A1(\po_0.regf_0.rf[0][5] ),
    .S(_1379_),
    .X(_1385_));
 sky130_fd_sc_hd__clkbuf_1 _3143_ (.A(_1385_),
    .X(_0262_));
 sky130_fd_sc_hd__buf_2 _3144_ (.A(_1378_),
    .X(_1386_));
 sky130_fd_sc_hd__mux2_1 _3145_ (.A0(_0809_),
    .A1(\po_0.regf_0.rf[0][6] ),
    .S(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__clkbuf_1 _3146_ (.A(_1387_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _3147_ (.A0(_0821_),
    .A1(\po_0.regf_0.rf[0][7] ),
    .S(_1386_),
    .X(_1388_));
 sky130_fd_sc_hd__clkbuf_1 _3148_ (.A(_1388_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _3149_ (.A0(_0836_),
    .A1(\po_0.regf_0.rf[0][8] ),
    .S(_1386_),
    .X(_1389_));
 sky130_fd_sc_hd__clkbuf_1 _3150_ (.A(_1389_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _3151_ (.A0(_0844_),
    .A1(\po_0.regf_0.rf[0][9] ),
    .S(_1386_),
    .X(_1390_));
 sky130_fd_sc_hd__clkbuf_1 _3152_ (.A(_1390_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _3153_ (.A0(_0853_),
    .A1(\po_0.regf_0.rf[0][10] ),
    .S(_1386_),
    .X(_1391_));
 sky130_fd_sc_hd__clkbuf_1 _3154_ (.A(_1391_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _3155_ (.A0(_0862_),
    .A1(\po_0.regf_0.rf[0][11] ),
    .S(_1386_),
    .X(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _3156_ (.A(_1392_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _3157_ (.A0(_0874_),
    .A1(\po_0.regf_0.rf[0][12] ),
    .S(_1378_),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _3158_ (.A(_1393_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _3159_ (.A0(_0883_),
    .A1(\po_0.regf_0.rf[0][13] ),
    .S(_1378_),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _3160_ (.A(_1394_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _3161_ (.A0(_0896_),
    .A1(\po_0.regf_0.rf[0][14] ),
    .S(_1378_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_1 _3162_ (.A(_1395_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _3163_ (.A0(_0904_),
    .A1(\po_0.regf_0.rf[0][15] ),
    .S(_1378_),
    .X(_1396_));
 sky130_fd_sc_hd__clkbuf_1 _3164_ (.A(_1396_),
    .X(_0272_));
 sky130_fd_sc_hd__and4bb_4 _3165_ (.A_N(_0742_),
    .B_N(\po_0.regf_0.w_addr[3] ),
    .C(_0906_),
    .D(_0907_),
    .X(_1397_));
 sky130_fd_sc_hd__clkbuf_4 _3166_ (.A(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(\po_0.regf_0.rf[2][0] ),
    .A1(_0735_),
    .S(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_1 _3168_ (.A(_1399_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(\po_0.regf_0.rf[2][1] ),
    .A1(_0755_),
    .S(_1398_),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_1 _3170_ (.A(_1400_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _3171_ (.A0(\po_0.regf_0.rf[2][2] ),
    .A1(_0767_),
    .S(_1398_),
    .X(_1401_));
 sky130_fd_sc_hd__clkbuf_1 _3172_ (.A(_1401_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(\po_0.regf_0.rf[2][3] ),
    .A1(_0777_),
    .S(_1398_),
    .X(_1402_));
 sky130_fd_sc_hd__clkbuf_1 _3174_ (.A(_1402_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(\po_0.regf_0.rf[2][4] ),
    .A1(_0788_),
    .S(_1398_),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_1 _3176_ (.A(_1403_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _3177_ (.A0(\po_0.regf_0.rf[2][5] ),
    .A1(_0796_),
    .S(_1398_),
    .X(_1404_));
 sky130_fd_sc_hd__clkbuf_1 _3178_ (.A(_1404_),
    .X(_0278_));
 sky130_fd_sc_hd__buf_2 _3179_ (.A(_1397_),
    .X(_1405_));
 sky130_fd_sc_hd__mux2_1 _3180_ (.A0(\po_0.regf_0.rf[2][6] ),
    .A1(_0808_),
    .S(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _3181_ (.A(_1406_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _3182_ (.A0(\po_0.regf_0.rf[2][7] ),
    .A1(_0820_),
    .S(_1405_),
    .X(_1407_));
 sky130_fd_sc_hd__clkbuf_1 _3183_ (.A(_1407_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _3184_ (.A0(\po_0.regf_0.rf[2][8] ),
    .A1(_0835_),
    .S(_1405_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _3185_ (.A(_1408_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _3186_ (.A0(\po_0.regf_0.rf[2][9] ),
    .A1(_0843_),
    .S(_1405_),
    .X(_1409_));
 sky130_fd_sc_hd__clkbuf_1 _3187_ (.A(_1409_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _3188_ (.A0(\po_0.regf_0.rf[2][10] ),
    .A1(_0852_),
    .S(_1405_),
    .X(_1410_));
 sky130_fd_sc_hd__clkbuf_1 _3189_ (.A(_1410_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _3190_ (.A0(\po_0.regf_0.rf[2][11] ),
    .A1(_0861_),
    .S(_1405_),
    .X(_1411_));
 sky130_fd_sc_hd__clkbuf_1 _3191_ (.A(_1411_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _3192_ (.A0(\po_0.regf_0.rf[2][12] ),
    .A1(_0873_),
    .S(_1397_),
    .X(_1412_));
 sky130_fd_sc_hd__clkbuf_1 _3193_ (.A(_1412_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _3194_ (.A0(\po_0.regf_0.rf[2][13] ),
    .A1(_0882_),
    .S(_1397_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_1 _3195_ (.A(_1413_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _3196_ (.A0(\po_0.regf_0.rf[2][14] ),
    .A1(_0895_),
    .S(_1397_),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _3197_ (.A(_1414_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _3198_ (.A0(\po_0.regf_0.rf[2][15] ),
    .A1(_0903_),
    .S(_1397_),
    .X(_1415_));
 sky130_fd_sc_hd__clkbuf_1 _3199_ (.A(_1415_),
    .X(_0288_));
 sky130_fd_sc_hd__and4b_4 _3200_ (.A_N(\po_0.regf_0.w_addr[2] ),
    .B(_0737_),
    .C(\po_0.regf_0.w_wr ),
    .D(_1061_),
    .X(_1416_));
 sky130_fd_sc_hd__buf_2 _3201_ (.A(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(\po_0.regf_0.rf[8][0] ),
    .A1(_0735_),
    .S(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _3203_ (.A(_1418_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _3204_ (.A0(\po_0.regf_0.rf[8][1] ),
    .A1(_0755_),
    .S(_1417_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_1 _3205_ (.A(_1419_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _3206_ (.A0(\po_0.regf_0.rf[8][2] ),
    .A1(_0767_),
    .S(_1417_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _3207_ (.A(_1420_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _3208_ (.A0(\po_0.regf_0.rf[8][3] ),
    .A1(_0777_),
    .S(_1417_),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_1 _3209_ (.A(_1421_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _3210_ (.A0(\po_0.regf_0.rf[8][4] ),
    .A1(_0788_),
    .S(_1417_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_1 _3211_ (.A(_1422_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _3212_ (.A0(\po_0.regf_0.rf[8][5] ),
    .A1(_0796_),
    .S(_1417_),
    .X(_1423_));
 sky130_fd_sc_hd__clkbuf_1 _3213_ (.A(_1423_),
    .X(_0294_));
 sky130_fd_sc_hd__buf_2 _3214_ (.A(_1416_),
    .X(_1424_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(\po_0.regf_0.rf[8][6] ),
    .A1(_0808_),
    .S(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__clkbuf_1 _3216_ (.A(_1425_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _3217_ (.A0(\po_0.regf_0.rf[8][7] ),
    .A1(_0820_),
    .S(_1424_),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_1 _3218_ (.A(_1426_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _3219_ (.A0(\po_0.regf_0.rf[8][8] ),
    .A1(_0835_),
    .S(_1424_),
    .X(_1427_));
 sky130_fd_sc_hd__clkbuf_1 _3220_ (.A(_1427_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(\po_0.regf_0.rf[8][9] ),
    .A1(_0843_),
    .S(_1424_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_1 _3222_ (.A(_1428_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _3223_ (.A0(\po_0.regf_0.rf[8][10] ),
    .A1(_0852_),
    .S(_1424_),
    .X(_1429_));
 sky130_fd_sc_hd__clkbuf_1 _3224_ (.A(_1429_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _3225_ (.A0(\po_0.regf_0.rf[8][11] ),
    .A1(_0861_),
    .S(_1424_),
    .X(_1430_));
 sky130_fd_sc_hd__clkbuf_1 _3226_ (.A(_1430_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _3227_ (.A0(\po_0.regf_0.rf[8][12] ),
    .A1(_0873_),
    .S(_1416_),
    .X(_1431_));
 sky130_fd_sc_hd__clkbuf_1 _3228_ (.A(_1431_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _3229_ (.A0(\po_0.regf_0.rf[8][13] ),
    .A1(_0882_),
    .S(_1416_),
    .X(_1432_));
 sky130_fd_sc_hd__clkbuf_1 _3230_ (.A(_1432_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _3231_ (.A0(\po_0.regf_0.rf[8][14] ),
    .A1(_0895_),
    .S(_1416_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _3232_ (.A(_1433_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _3233_ (.A0(\po_0.regf_0.rf[8][15] ),
    .A1(_0903_),
    .S(_1416_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_1 _3234_ (.A(_1434_),
    .X(_0304_));
 sky130_fd_sc_hd__a21bo_1 _3235_ (.A1(_1551_),
    .A2(_0729_),
    .B1_N(_1550_),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_2 _3236_ (.A(_1546_),
    .X(_1435_));
 sky130_fd_sc_hd__and2_1 _3237_ (.A(_1550_),
    .B(_1551_),
    .X(_1436_));
 sky130_fd_sc_hd__a32o_1 _3238_ (.A1(_1520_),
    .A2(\uc_0.bc_0._70_[1] ),
    .A3(_1435_),
    .B1(_1436_),
    .B2(_1489_),
    .X(_0306_));
 sky130_fd_sc_hd__or4_1 _3239_ (.A(_1356_),
    .B(_1357_),
    .C(_1546_),
    .D(_0594_),
    .X(_1437_));
 sky130_fd_sc_hd__buf_2 _3240_ (.A(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__a21o_1 _3241_ (.A1(_1438_),
    .A2(net92),
    .B1(_1553_),
    .X(_0307_));
 sky130_fd_sc_hd__a21o_1 _3242_ (.A1(net88),
    .A2(_1358_),
    .B1(_0596_),
    .X(_0308_));
 sky130_fd_sc_hd__or3b_1 _3243_ (.A(_1357_),
    .B(_1517_),
    .C_N(_1520_),
    .X(_1439_));
 sky130_fd_sc_hd__inv_2 _3244_ (.A(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__and3_2 _3245_ (.A(_1520_),
    .B(\uc_0.bc_0._70_[0] ),
    .C(_1357_),
    .X(_1441_));
 sky130_fd_sc_hd__clkbuf_4 _3246_ (.A(_1552_),
    .X(_1442_));
 sky130_fd_sc_hd__a211oi_4 _3247_ (.A1(_1546_),
    .A2(_1440_),
    .B1(_1441_),
    .C1(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__a21bo_1 _3248_ (.A1(_0738_),
    .A2(_1438_),
    .B1_N(_1443_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _3249_ (.A0(\po_0.regf_0.rq_addr[0] ),
    .A1(_1549_),
    .S(_1553_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _3250_ (.A(_1444_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _3251_ (.A0(\po_0.regf_0.rq_addr[1] ),
    .A1(_1555_),
    .S(_1442_),
    .X(_1445_));
 sky130_fd_sc_hd__clkbuf_1 _3252_ (.A(_1445_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _3253_ (.A0(\po_0.regf_0.rq_addr[2] ),
    .A1(_1557_),
    .S(_1442_),
    .X(_1446_));
 sky130_fd_sc_hd__clkbuf_1 _3254_ (.A(_1446_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _3255_ (.A0(\po_0.regf_0.rq_addr[3] ),
    .A1(_1559_),
    .S(_1442_),
    .X(_1447_));
 sky130_fd_sc_hd__clkbuf_1 _3256_ (.A(_1447_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _3257_ (.A0(\po_0.regf_0.rp_addr[0] ),
    .A1(\uc_0._21_[8] ),
    .S(_0596_),
    .X(_1448_));
 sky130_fd_sc_hd__clkbuf_1 _3258_ (.A(_1448_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _3259_ (.A0(\po_0.regf_0.rp_addr[1] ),
    .A1(\uc_0._21_[9] ),
    .S(_0595_),
    .X(_1449_));
 sky130_fd_sc_hd__clkbuf_1 _3260_ (.A(_1449_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _3261_ (.A0(\po_0.regf_0.rp_addr[2] ),
    .A1(\uc_0._21_[10] ),
    .S(_0595_),
    .X(_1450_));
 sky130_fd_sc_hd__clkbuf_1 _3262_ (.A(_1450_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _3263_ (.A0(\po_0.regf_0.rp_addr[3] ),
    .A1(\uc_0._21_[11] ),
    .S(_0595_),
    .X(_1451_));
 sky130_fd_sc_hd__clkbuf_1 _3264_ (.A(_1451_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _3265_ (.A0(\uc_0._21_[8] ),
    .A1(_1124_),
    .S(_1442_),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_1 _3266_ (.A0(_1452_),
    .A1(_0740_),
    .S(_1443_),
    .X(_1453_));
 sky130_fd_sc_hd__clkbuf_1 _3267_ (.A(_1453_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _3268_ (.A0(\uc_0._21_[9] ),
    .A1(_1136_),
    .S(_1442_),
    .X(_1454_));
 sky130_fd_sc_hd__mux2_1 _3269_ (.A0(_1454_),
    .A1(_0739_),
    .S(_1443_),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_1 _3270_ (.A(_1455_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _3271_ (.A0(\uc_0._21_[10] ),
    .A1(_1151_),
    .S(_1552_),
    .X(_1456_));
 sky130_fd_sc_hd__mux2_1 _3272_ (.A0(_1456_),
    .A1(_0929_),
    .S(_1443_),
    .X(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _3273_ (.A(_1457_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _3274_ (.A0(\uc_0._21_[11] ),
    .A1(_1163_),
    .S(_1552_),
    .X(_1458_));
 sky130_fd_sc_hd__mux2_1 _3275_ (.A0(_1458_),
    .A1(_0927_),
    .S(_1443_),
    .X(_1459_));
 sky130_fd_sc_hd__clkbuf_1 _3276_ (.A(_1459_),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_2 _3277_ (.A(_1441_),
    .X(_1460_));
 sky130_fd_sc_hd__mux2_1 _3278_ (.A0(\po_0.muxf_0.rf_w_data[0] ),
    .A1(_1124_),
    .S(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__clkbuf_1 _3279_ (.A(_1461_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _3280_ (.A0(\po_0.muxf_0.rf_w_data[1] ),
    .A1(_1136_),
    .S(_1460_),
    .X(_1462_));
 sky130_fd_sc_hd__clkbuf_1 _3281_ (.A(_1462_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _3282_ (.A0(\po_0.muxf_0.rf_w_data[2] ),
    .A1(_1151_),
    .S(_1460_),
    .X(_1463_));
 sky130_fd_sc_hd__clkbuf_1 _3283_ (.A(_1463_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _3284_ (.A0(\po_0.muxf_0.rf_w_data[3] ),
    .A1(_1163_),
    .S(_1460_),
    .X(_1464_));
 sky130_fd_sc_hd__clkbuf_1 _3285_ (.A(_1464_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _3286_ (.A0(\po_0.muxf_0.rf_w_data[4] ),
    .A1(_1549_),
    .S(_1441_),
    .X(_1465_));
 sky130_fd_sc_hd__clkbuf_1 _3287_ (.A(_1465_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _3288_ (.A0(\po_0.muxf_0.rf_w_data[5] ),
    .A1(_1555_),
    .S(_1441_),
    .X(_1466_));
 sky130_fd_sc_hd__clkbuf_1 _3289_ (.A(_1466_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(\po_0.muxf_0.rf_w_data[6] ),
    .A1(_1557_),
    .S(_1441_),
    .X(_1467_));
 sky130_fd_sc_hd__clkbuf_1 _3291_ (.A(_1467_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _3292_ (.A0(\po_0.muxf_0.rf_w_data[7] ),
    .A1(_1559_),
    .S(_1441_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _3293_ (.A(_1468_),
    .X(_0329_));
 sky130_fd_sc_hd__a31o_1 _3294_ (.A1(\uc_0.bc_0._70_[2] ),
    .A2(_0593_),
    .A3(_1435_),
    .B1(\po_0.muxf_0.s0 ),
    .X(_1469_));
 sky130_fd_sc_hd__and3b_1 _3295_ (.A_N(_1460_),
    .B(_1469_),
    .C(_1436_),
    .X(_1470_));
 sky130_fd_sc_hd__clkbuf_1 _3296_ (.A(_1470_),
    .X(_0330_));
 sky130_fd_sc_hd__inv_2 _3297_ (.A(_1435_),
    .Y(_1471_));
 sky130_fd_sc_hd__clkbuf_4 _3298_ (.A(_1439_),
    .X(_1472_));
 sky130_fd_sc_hd__buf_2 _3299_ (.A(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__o221a_1 _3300_ (.A1(_1471_),
    .A2(_1473_),
    .B1(_1460_),
    .B2(\po_0.muxf_0.s1 ),
    .C1(_1436_),
    .X(_0331_));
 sky130_fd_sc_hd__a22o_1 _3301_ (.A1(\uc_0.bc_0._70_[0] ),
    .A2(_1440_),
    .B1(_1438_),
    .B2(net60),
    .X(_0332_));
 sky130_fd_sc_hd__a32o_1 _3302_ (.A1(\uc_0.bc_0._70_[2] ),
    .A2(_0593_),
    .A3(_1435_),
    .B1(_1438_),
    .B2(net59),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _3303_ (.A0(_1124_),
    .A1(net51),
    .S(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__clkbuf_1 _3304_ (.A(_1474_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _3305_ (.A0(_1136_),
    .A1(net52),
    .S(_1473_),
    .X(_1475_));
 sky130_fd_sc_hd__clkbuf_1 _3306_ (.A(_1475_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _3307_ (.A0(_1151_),
    .A1(net53),
    .S(_1473_),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_1 _3308_ (.A(_1476_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _3309_ (.A0(_1163_),
    .A1(net54),
    .S(_1472_),
    .X(_1477_));
 sky130_fd_sc_hd__clkbuf_1 _3310_ (.A(_1477_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _3311_ (.A0(_1549_),
    .A1(net55),
    .S(_1472_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_1 _3312_ (.A(_1478_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _3313_ (.A0(_1555_),
    .A1(net56),
    .S(_1472_),
    .X(_1479_));
 sky130_fd_sc_hd__clkbuf_1 _3314_ (.A(_1479_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _3315_ (.A0(_1557_),
    .A1(net57),
    .S(_1472_),
    .X(_1480_));
 sky130_fd_sc_hd__clkbuf_1 _3316_ (.A(_1480_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _3317_ (.A0(_1559_),
    .A1(net58),
    .S(_1472_),
    .X(_1481_));
 sky130_fd_sc_hd__clkbuf_1 _3318_ (.A(_1481_),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_1 _3319_ (.A(_0594_),
    .B(_1358_),
    .Y(_1482_));
 sky130_fd_sc_hd__o2bb2a_1 _3320_ (.A1_N(\uc_0.bc_0._70_[2] ),
    .A2_N(_0593_),
    .B1(_1482_),
    .B2(net77),
    .X(_0342_));
 sky130_fd_sc_hd__or3_1 _3321_ (.A(_1356_),
    .B(_0593_),
    .C(_1435_),
    .X(_1483_));
 sky130_fd_sc_hd__o221a_1 _3322_ (.A1(_0594_),
    .A2(_1483_),
    .B1(_1482_),
    .B2(_1337_),
    .C1(_1473_),
    .X(_0343_));
 sky130_fd_sc_hd__and3b_1 _3323_ (.A_N(_1535_),
    .B(_1519_),
    .C(_1539_),
    .X(_1484_));
 sky130_fd_sc_hd__o21ba_1 _3324_ (.A1(_1248_),
    .A2(_1484_),
    .B1_N(_1356_),
    .X(_1485_));
 sky130_fd_sc_hd__o311a_1 _3325_ (.A1(_1538_),
    .A2(_1435_),
    .A3(_0594_),
    .B1(_1473_),
    .C1(_1485_),
    .X(_0344_));
 sky130_fd_sc_hd__a311o_1 _3326_ (.A1(_1533_),
    .A2(_1534_),
    .A3(_1537_),
    .B1(_1356_),
    .C1(_1471_),
    .X(_1486_));
 sky130_fd_sc_hd__a2bb2o_1 _3327_ (.A1_N(_1548_),
    .A2_N(_1486_),
    .B1(_1119_),
    .B2(_1438_),
    .X(_0345_));
 sky130_fd_sc_hd__dfxtp_1 _3328_ (.CLK(net127),
    .D(_0016_),
    .Q(\po_0.regf_0.rf[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3329_ (.CLK(net129),
    .D(_0017_),
    .Q(\po_0.regf_0.rf[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3330_ (.CLK(net136),
    .D(_0018_),
    .Q(\po_0.regf_0.rf[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3331_ (.CLK(net129),
    .D(_0019_),
    .Q(\po_0.regf_0.rf[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3332_ (.CLK(net136),
    .D(_0020_),
    .Q(\po_0.regf_0.rf[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3333_ (.CLK(net134),
    .D(_0021_),
    .Q(\po_0.regf_0.rf[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3334_ (.CLK(net154),
    .D(_0022_),
    .Q(\po_0.regf_0.rf[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3335_ (.CLK(net154),
    .D(_0023_),
    .Q(\po_0.regf_0.rf[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3336_ (.CLK(net118),
    .D(_0024_),
    .Q(\po_0.regf_0.rf[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3337_ (.CLK(net115),
    .D(_0025_),
    .Q(\po_0.regf_0.rf[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3338_ (.CLK(net158),
    .D(_0026_),
    .Q(\po_0.regf_0.rf[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3339_ (.CLK(net118),
    .D(_0027_),
    .Q(\po_0.regf_0.rf[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3340_ (.CLK(net102),
    .D(_0028_),
    .Q(\po_0.regf_0.rf[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3341_ (.CLK(net109),
    .D(_0029_),
    .Q(\po_0.regf_0.rf[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3342_ (.CLK(net105),
    .D(_0030_),
    .Q(\po_0.regf_0.rf[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3343_ (.CLK(net100),
    .D(_0031_),
    .Q(\po_0.regf_0.rf[5][15] ));
 sky130_fd_sc_hd__dlxtp_1 _3344_ (.D(\po_0.regf_0._5_[0] ),
    .GATE(net93),
    .Q(\po_0._1_[0] ));
 sky130_fd_sc_hd__dlxtp_1 _3345_ (.D(\po_0.regf_0._5_[1] ),
    .GATE(net93),
    .Q(\po_0._1_[1] ));
 sky130_fd_sc_hd__dlxtp_1 _3346_ (.D(\po_0.regf_0._5_[2] ),
    .GATE(net93),
    .Q(\po_0._1_[2] ));
 sky130_fd_sc_hd__dlxtp_1 _3347_ (.D(\po_0.regf_0._5_[3] ),
    .GATE(net93),
    .Q(\po_0._1_[3] ));
 sky130_fd_sc_hd__dlxtp_1 _3348_ (.D(\po_0.regf_0._5_[4] ),
    .GATE(\po_0.regf_0.rq_rd ),
    .Q(\po_0._1_[4] ));
 sky130_fd_sc_hd__dlxtp_1 _3349_ (.D(\po_0.regf_0._5_[5] ),
    .GATE(\po_0.regf_0.rq_rd ),
    .Q(\po_0._1_[5] ));
 sky130_fd_sc_hd__dlxtp_1 _3350_ (.D(\po_0.regf_0._5_[6] ),
    .GATE(net91),
    .Q(\po_0._1_[6] ));
 sky130_fd_sc_hd__dlxtp_1 _3351_ (.D(\po_0.regf_0._5_[7] ),
    .GATE(net92),
    .Q(\po_0._1_[7] ));
 sky130_fd_sc_hd__dlxtp_1 _3352_ (.D(\po_0.regf_0._5_[8] ),
    .GATE(net92),
    .Q(\po_0._1_[8] ));
 sky130_fd_sc_hd__dlxtp_1 _3353_ (.D(\po_0.regf_0._5_[9] ),
    .GATE(net92),
    .Q(\po_0._1_[9] ));
 sky130_fd_sc_hd__dlxtp_1 _3354_ (.D(\po_0.regf_0._5_[10] ),
    .GATE(net92),
    .Q(\po_0._1_[10] ));
 sky130_fd_sc_hd__dlxtp_1 _3355_ (.D(\po_0.regf_0._5_[11] ),
    .GATE(net91),
    .Q(\po_0._1_[11] ));
 sky130_fd_sc_hd__dlxtp_1 _3356_ (.D(\po_0.regf_0._5_[12] ),
    .GATE(net91),
    .Q(\po_0._1_[12] ));
 sky130_fd_sc_hd__dlxtp_1 _3357_ (.D(\po_0.regf_0._5_[13] ),
    .GATE(net91),
    .Q(\po_0._1_[13] ));
 sky130_fd_sc_hd__dlxtp_1 _3358_ (.D(\po_0.regf_0._5_[14] ),
    .GATE(net91),
    .Q(\po_0._1_[14] ));
 sky130_fd_sc_hd__dlxtp_1 _3359_ (.D(\po_0.regf_0._5_[15] ),
    .GATE(net91),
    .Q(\po_0._1_[15] ));
 sky130_fd_sc_hd__dlxtp_1 _3360_ (.D(\po_0.regf_0._3_[0] ),
    .GATE(net89),
    .Q(net35));
 sky130_fd_sc_hd__dlxtp_1 _3361_ (.D(\po_0.regf_0._3_[1] ),
    .GATE(net89),
    .Q(net42));
 sky130_fd_sc_hd__dlxtp_1 _3362_ (.D(\po_0.regf_0._3_[2] ),
    .GATE(net90),
    .Q(net43));
 sky130_fd_sc_hd__dlxtp_1 _3363_ (.D(\po_0.regf_0._3_[3] ),
    .GATE(net89),
    .Q(net44));
 sky130_fd_sc_hd__dlxtp_1 _3364_ (.D(\po_0.regf_0._3_[4] ),
    .GATE(net90),
    .Q(net45));
 sky130_fd_sc_hd__dlxtp_1 _3365_ (.D(\po_0.regf_0._3_[5] ),
    .GATE(net90),
    .Q(net46));
 sky130_fd_sc_hd__dlxtp_1 _3366_ (.D(\po_0.regf_0._3_[6] ),
    .GATE(net89),
    .Q(net47));
 sky130_fd_sc_hd__dlxtp_1 _3367_ (.D(\po_0.regf_0._3_[7] ),
    .GATE(net88),
    .Q(net48));
 sky130_fd_sc_hd__dlxtp_1 _3368_ (.D(\po_0.regf_0._3_[8] ),
    .GATE(net88),
    .Q(net49));
 sky130_fd_sc_hd__dlxtp_1 _3369_ (.D(\po_0.regf_0._3_[9] ),
    .GATE(net89),
    .Q(net50));
 sky130_fd_sc_hd__dlxtp_1 _3370_ (.D(\po_0.regf_0._3_[10] ),
    .GATE(net88),
    .Q(net36));
 sky130_fd_sc_hd__dlxtp_1 _3371_ (.D(\po_0.regf_0._3_[11] ),
    .GATE(net88),
    .Q(net37));
 sky130_fd_sc_hd__dlxtp_1 _3372_ (.D(\po_0.regf_0._3_[12] ),
    .GATE(net90),
    .Q(net38));
 sky130_fd_sc_hd__dlxtp_1 _3373_ (.D(\po_0.regf_0._3_[13] ),
    .GATE(net90),
    .Q(net39));
 sky130_fd_sc_hd__dlxtp_1 _3374_ (.D(\po_0.regf_0._3_[14] ),
    .GATE(net88),
    .Q(net40));
 sky130_fd_sc_hd__dlxtp_1 _3375_ (.D(\po_0.regf_0._3_[15] ),
    .GATE(net90),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _3376_ (.CLK(net127),
    .D(_0032_),
    .Q(\po_0.regf_0.rf[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3377_ (.CLK(net129),
    .D(_0033_),
    .Q(\po_0.regf_0.rf[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3378_ (.CLK(net134),
    .D(_0034_),
    .Q(\po_0.regf_0.rf[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3379_ (.CLK(net129),
    .D(_0035_),
    .Q(\po_0.regf_0.rf[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3380_ (.CLK(net134),
    .D(_0036_),
    .Q(\po_0.regf_0.rf[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3381_ (.CLK(net135),
    .D(_0037_),
    .Q(\po_0.regf_0.rf[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3382_ (.CLK(net155),
    .D(_0038_),
    .Q(\po_0.regf_0.rf[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3383_ (.CLK(net154),
    .D(_0039_),
    .Q(\po_0.regf_0.rf[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3384_ (.CLK(net118),
    .D(_0040_),
    .Q(\po_0.regf_0.rf[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3385_ (.CLK(net115),
    .D(_0041_),
    .Q(\po_0.regf_0.rf[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3386_ (.CLK(net158),
    .D(_0042_),
    .Q(\po_0.regf_0.rf[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3387_ (.CLK(net115),
    .D(_0043_),
    .Q(\po_0.regf_0.rf[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3388_ (.CLK(net105),
    .D(_0044_),
    .Q(\po_0.regf_0.rf[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3389_ (.CLK(net109),
    .D(_0045_),
    .Q(\po_0.regf_0.rf[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3390_ (.CLK(net105),
    .D(_0046_),
    .Q(\po_0.regf_0.rf[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3391_ (.CLK(net101),
    .D(_0047_),
    .Q(\po_0.regf_0.rf[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3392_ (.CLK(net127),
    .D(_0048_),
    .Q(\po_0.regf_0.rf[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3393_ (.CLK(net129),
    .D(_0049_),
    .Q(\po_0.regf_0.rf[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3394_ (.CLK(net134),
    .D(_0050_),
    .Q(\po_0.regf_0.rf[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3395_ (.CLK(net129),
    .D(_0051_),
    .Q(\po_0.regf_0.rf[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3396_ (.CLK(net134),
    .D(_0052_),
    .Q(\po_0.regf_0.rf[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3397_ (.CLK(net134),
    .D(_0053_),
    .Q(\po_0.regf_0.rf[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3398_ (.CLK(net155),
    .D(_0054_),
    .Q(\po_0.regf_0.rf[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3399_ (.CLK(net154),
    .D(_0055_),
    .Q(\po_0.regf_0.rf[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3400_ (.CLK(net119),
    .D(_0056_),
    .Q(\po_0.regf_0.rf[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3401_ (.CLK(net115),
    .D(_0057_),
    .Q(\po_0.regf_0.rf[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3402_ (.CLK(net158),
    .D(_0058_),
    .Q(\po_0.regf_0.rf[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3403_ (.CLK(net115),
    .D(_0059_),
    .Q(\po_0.regf_0.rf[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3404_ (.CLK(net105),
    .D(_0060_),
    .Q(\po_0.regf_0.rf[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3405_ (.CLK(net109),
    .D(_0061_),
    .Q(\po_0.regf_0.rf[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3406_ (.CLK(net105),
    .D(_0062_),
    .Q(\po_0.regf_0.rf[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3407_ (.CLK(net100),
    .D(_0063_),
    .Q(\po_0.regf_0.rf[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3408_ (.CLK(net178),
    .D(_0008_),
    .Q(_0000_));
 sky130_fd_sc_hd__dfxtp_1 _3409_ (.CLK(net166),
    .D(_0009_),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_1 _3410_ (.CLK(net166),
    .D(_0010_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_2 _3411_ (.CLK(net164),
    .D(_0011_),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_1 _3412_ (.CLK(net145),
    .D(_0064_),
    .Q(\po_0.regf_0.rf[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3413_ (.CLK(net151),
    .D(_0065_),
    .Q(\po_0.regf_0.rf[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3414_ (.CLK(net150),
    .D(_0066_),
    .Q(\po_0.regf_0.rf[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3415_ (.CLK(net145),
    .D(_0067_),
    .Q(\po_0.regf_0.rf[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3416_ (.CLK(net149),
    .D(_0068_),
    .Q(\po_0.regf_0.rf[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3417_ (.CLK(net150),
    .D(_0069_),
    .Q(\po_0.regf_0.rf[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3418_ (.CLK(net166),
    .D(_0070_),
    .Q(\po_0.regf_0.rf[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3419_ (.CLK(net162),
    .D(_0071_),
    .Q(\po_0.regf_0.rf[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3420_ (.CLK(net122),
    .D(_0072_),
    .Q(\po_0.regf_0.rf[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3421_ (.CLK(net124),
    .D(_0073_),
    .Q(\po_0.regf_0.rf[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3422_ (.CLK(net164),
    .D(_0074_),
    .Q(\po_0.regf_0.rf[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3423_ (.CLK(net123),
    .D(_0075_),
    .Q(\po_0.regf_0.rf[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3424_ (.CLK(net109),
    .D(_0076_),
    .Q(\po_0.regf_0.rf[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3425_ (.CLK(net127),
    .D(_0077_),
    .Q(\po_0.regf_0.rf[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3426_ (.CLK(net112),
    .D(_0078_),
    .Q(\po_0.regf_0.rf[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3427_ (.CLK(net109),
    .D(_0079_),
    .Q(\po_0.regf_0.rf[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3428_ (.CLK(net143),
    .D(_0080_),
    .Q(\po_0.regf_0.rf[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3429_ (.CLK(net131),
    .D(_0081_),
    .Q(\po_0.regf_0.rf[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3430_ (.CLK(net149),
    .D(_0082_),
    .Q(\po_0.regf_0.rf[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3431_ (.CLK(net143),
    .D(_0083_),
    .Q(\po_0.regf_0.rf[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3432_ (.CLK(net140),
    .D(_0084_),
    .Q(\po_0.regf_0.rf[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3433_ (.CLK(net148),
    .D(_0085_),
    .Q(\po_0.regf_0.rf[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3434_ (.CLK(net159),
    .D(_0086_),
    .Q(\po_0.regf_0.rf[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3435_ (.CLK(net156),
    .D(_0087_),
    .Q(\po_0.regf_0.rf[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3436_ (.CLK(net120),
    .D(_0088_),
    .Q(\po_0.regf_0.rf[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3437_ (.CLK(net116),
    .D(_0089_),
    .Q(\po_0.regf_0.rf[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3438_ (.CLK(net159),
    .D(_0090_),
    .Q(\po_0.regf_0.rf[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3439_ (.CLK(net120),
    .D(_0091_),
    .Q(\po_0.regf_0.rf[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3440_ (.CLK(net112),
    .D(_0092_),
    .Q(\po_0.regf_0.rf[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3441_ (.CLK(net113),
    .D(_0093_),
    .Q(\po_0.regf_0.rf[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3442_ (.CLK(net103),
    .D(_0094_),
    .Q(\po_0.regf_0.rf[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3443_ (.CLK(net107),
    .D(_0095_),
    .Q(\po_0.regf_0.rf[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3444_ (.CLK(net132),
    .D(_0096_),
    .Q(\po_0.regf_0.rf[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3445_ (.CLK(net148),
    .D(_0097_),
    .Q(\po_0.regf_0.rf[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3446_ (.CLK(net149),
    .D(_0098_),
    .Q(\po_0.regf_0.rf[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3447_ (.CLK(net143),
    .D(_0099_),
    .Q(\po_0.regf_0.rf[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3448_ (.CLK(net140),
    .D(_0100_),
    .Q(\po_0.regf_0.rf[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3449_ (.CLK(net137),
    .D(_0101_),
    .Q(\po_0.regf_0.rf[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3450_ (.CLK(net164),
    .D(_0102_),
    .Q(\po_0.regf_0.rf[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3451_ (.CLK(net162),
    .D(_0103_),
    .Q(\po_0.regf_0.rf[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3452_ (.CLK(net122),
    .D(_0104_),
    .Q(\po_0.regf_0.rf[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3453_ (.CLK(net124),
    .D(_0105_),
    .Q(\po_0.regf_0.rf[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3454_ (.CLK(net164),
    .D(_0106_),
    .Q(\po_0.regf_0.rf[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3455_ (.CLK(net122),
    .D(_0107_),
    .Q(\po_0.regf_0.rf[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3456_ (.CLK(net107),
    .D(_0108_),
    .Q(\po_0.regf_0.rf[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3457_ (.CLK(net127),
    .D(_0109_),
    .Q(\po_0.regf_0.rf[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3458_ (.CLK(net112),
    .D(_0110_),
    .Q(\po_0.regf_0.rf[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3459_ (.CLK(net107),
    .D(_0111_),
    .Q(\po_0.regf_0.rf[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3460_ (.CLK(net132),
    .D(_0112_),
    .Q(\po_0.regf_0.rf[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3461_ (.CLK(net131),
    .D(_0113_),
    .Q(\po_0.regf_0.rf[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3462_ (.CLK(net139),
    .D(_0114_),
    .Q(\po_0.regf_0.rf[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3463_ (.CLK(net133),
    .D(_0115_),
    .Q(\po_0.regf_0.rf[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3464_ (.CLK(net139),
    .D(_0116_),
    .Q(\po_0.regf_0.rf[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3465_ (.CLK(net137),
    .D(_0117_),
    .Q(\po_0.regf_0.rf[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3466_ (.CLK(net162),
    .D(_0118_),
    .Q(\po_0.regf_0.rf[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3467_ (.CLK(net156),
    .D(_0119_),
    .Q(\po_0.regf_0.rf[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3468_ (.CLK(net120),
    .D(_0120_),
    .Q(\po_0.regf_0.rf[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3469_ (.CLK(net116),
    .D(_0121_),
    .Q(\po_0.regf_0.rf[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3470_ (.CLK(net159),
    .D(_0122_),
    .Q(\po_0.regf_0.rf[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3471_ (.CLK(net120),
    .D(_0123_),
    .Q(\po_0.regf_0.rf[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3472_ (.CLK(net100),
    .D(_0124_),
    .Q(\po_0.regf_0.rf[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3473_ (.CLK(net110),
    .D(_0125_),
    .Q(\po_0.regf_0.rf[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3474_ (.CLK(net103),
    .D(_0126_),
    .Q(\po_0.regf_0.rf[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3475_ (.CLK(net100),
    .D(_0127_),
    .Q(\po_0.regf_0.rf[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3476_ (.CLK(net132),
    .D(_0128_),
    .Q(\po_0.regf_0.rf[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3477_ (.CLK(net137),
    .D(_0129_),
    .Q(\po_0.regf_0.rf[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3478_ (.CLK(net139),
    .D(_0130_),
    .Q(\po_0.regf_0.rf[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3479_ (.CLK(net133),
    .D(_0131_),
    .Q(\po_0.regf_0.rf[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3480_ (.CLK(net139),
    .D(_0132_),
    .Q(\po_0.regf_0.rf[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3481_ (.CLK(net138),
    .D(_0133_),
    .Q(\po_0.regf_0.rf[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3482_ (.CLK(net156),
    .D(_0134_),
    .Q(\po_0.regf_0.rf[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3483_ (.CLK(net156),
    .D(_0135_),
    .Q(\po_0.regf_0.rf[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3484_ (.CLK(net120),
    .D(_0136_),
    .Q(\po_0.regf_0.rf[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3485_ (.CLK(net116),
    .D(_0137_),
    .Q(\po_0.regf_0.rf[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3486_ (.CLK(net159),
    .D(_0138_),
    .Q(\po_0.regf_0.rf[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3487_ (.CLK(net120),
    .D(_0139_),
    .Q(\po_0.regf_0.rf[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3488_ (.CLK(net100),
    .D(_0140_),
    .Q(\po_0.regf_0.rf[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3489_ (.CLK(net110),
    .D(_0141_),
    .Q(\po_0.regf_0.rf[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3490_ (.CLK(net104),
    .D(_0142_),
    .Q(\po_0.regf_0.rf[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3491_ (.CLK(net100),
    .D(_0143_),
    .Q(\po_0.regf_0.rf[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3492_ (.CLK(net132),
    .D(_0144_),
    .Q(\po_0.regf_0.rf[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3493_ (.CLK(net138),
    .D(_0145_),
    .Q(\po_0.regf_0.rf[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3494_ (.CLK(net149),
    .D(_0146_),
    .Q(\po_0.regf_0.rf[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3495_ (.CLK(net143),
    .D(_0147_),
    .Q(\po_0.regf_0.rf[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3496_ (.CLK(net140),
    .D(_0148_),
    .Q(\po_0.regf_0.rf[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3497_ (.CLK(net148),
    .D(_0149_),
    .Q(\po_0.regf_0.rf[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3498_ (.CLK(net165),
    .D(_0150_),
    .Q(\po_0.regf_0.rf[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3499_ (.CLK(net162),
    .D(_0151_),
    .Q(\po_0.regf_0.rf[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3500_ (.CLK(net123),
    .D(_0152_),
    .Q(\po_0.regf_0.rf[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3501_ (.CLK(net124),
    .D(_0153_),
    .Q(\po_0.regf_0.rf[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3502_ (.CLK(net164),
    .D(_0154_),
    .Q(\po_0.regf_0.rf[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3503_ (.CLK(net122),
    .D(_0155_),
    .Q(\po_0.regf_0.rf[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3504_ (.CLK(net107),
    .D(_0156_),
    .Q(\po_0.regf_0.rf[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3505_ (.CLK(net127),
    .D(_0157_),
    .Q(\po_0.regf_0.rf[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3506_ (.CLK(net112),
    .D(_0158_),
    .Q(\po_0.regf_0.rf[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3507_ (.CLK(net107),
    .D(_0159_),
    .Q(\po_0.regf_0.rf[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3508_ (.CLK(net145),
    .D(_0160_),
    .Q(\po_0.regf_0.rf[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3509_ (.CLK(net146),
    .D(_0161_),
    .Q(\po_0.regf_0.rf[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3510_ (.CLK(net150),
    .D(_0162_),
    .Q(\po_0.regf_0.rf[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3511_ (.CLK(net146),
    .D(_0163_),
    .Q(\po_0.regf_0.rf[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3512_ (.CLK(net150),
    .D(_0164_),
    .Q(\po_0.regf_0.rf[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3513_ (.CLK(net151),
    .D(_0165_),
    .Q(\po_0.regf_0.rf[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3514_ (.CLK(net166),
    .D(_0166_),
    .Q(\po_0.regf_0.rf[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3515_ (.CLK(net163),
    .D(_0167_),
    .Q(\po_0.regf_0.rf[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3516_ (.CLK(net162),
    .D(_0168_),
    .Q(\po_0.regf_0.rf[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3517_ (.CLK(net124),
    .D(_0169_),
    .Q(\po_0.regf_0.rf[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3518_ (.CLK(net164),
    .D(_0170_),
    .Q(\po_0.regf_0.rf[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3519_ (.CLK(net122),
    .D(_0171_),
    .Q(\po_0.regf_0.rf[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3520_ (.CLK(net110),
    .D(_0172_),
    .Q(\po_0.regf_0.rf[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3521_ (.CLK(net128),
    .D(_0173_),
    .Q(\po_0.regf_0.rf[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3522_ (.CLK(net112),
    .D(_0174_),
    .Q(\po_0.regf_0.rf[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3523_ (.CLK(net108),
    .D(_0175_),
    .Q(\po_0.regf_0.rf[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3524_ (.CLK(net145),
    .D(_0176_),
    .Q(\po_0.regf_0.rf[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3525_ (.CLK(net146),
    .D(_0177_),
    .Q(\po_0.regf_0.rf[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3526_ (.CLK(net150),
    .D(_0178_),
    .Q(\po_0.regf_0.rf[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3527_ (.CLK(net146),
    .D(_0179_),
    .Q(\po_0.regf_0.rf[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3528_ (.CLK(net150),
    .D(_0180_),
    .Q(\po_0.regf_0.rf[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3529_ (.CLK(net151),
    .D(_0181_),
    .Q(\po_0.regf_0.rf[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3530_ (.CLK(net166),
    .D(_0182_),
    .Q(\po_0.regf_0.rf[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3531_ (.CLK(net163),
    .D(_0183_),
    .Q(\po_0.regf_0.rf[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3532_ (.CLK(net162),
    .D(_0184_),
    .Q(\po_0.regf_0.rf[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3533_ (.CLK(net124),
    .D(_0185_),
    .Q(\po_0.regf_0.rf[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3534_ (.CLK(net165),
    .D(_0186_),
    .Q(\po_0.regf_0.rf[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3535_ (.CLK(net122),
    .D(_0187_),
    .Q(\po_0.regf_0.rf[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3536_ (.CLK(net109),
    .D(_0188_),
    .Q(\po_0.regf_0.rf[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3537_ (.CLK(net128),
    .D(_0189_),
    .Q(\po_0.regf_0.rf[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3538_ (.CLK(net112),
    .D(_0190_),
    .Q(\po_0.regf_0.rf[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3539_ (.CLK(net107),
    .D(_0191_),
    .Q(\po_0.regf_0.rf[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3540_ (.CLK(net181),
    .D(_0192_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _3541_ (.CLK(net183),
    .D(_0193_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_2 _3542_ (.CLK(net174),
    .D(_0194_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _3543_ (.CLK(net176),
    .D(_0195_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _3544_ (.CLK(net176),
    .D(_0196_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_2 _3545_ (.CLK(net171),
    .D(_0197_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_2 _3546_ (.CLK(net171),
    .D(_0198_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _3547_ (.CLK(net172),
    .D(_0199_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_2 _3548_ (.CLK(net173),
    .D(_0200_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _3549_ (.CLK(net173),
    .D(_0201_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_4 _3550_ (.CLK(net173),
    .D(_0202_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _3551_ (.CLK(net176),
    .D(_0203_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _3552_ (.CLK(net176),
    .D(_0204_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _3553_ (.CLK(net177),
    .D(_0205_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_1 _3554_ (.CLK(net181),
    .D(_0206_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_2 _3555_ (.CLK(net181),
    .D(_0207_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _3556_ (.CLK(net131),
    .D(_0208_),
    .Q(\po_0.regf_0.rf[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3557_ (.CLK(net135),
    .D(_0209_),
    .Q(\po_0.regf_0.rf[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3558_ (.CLK(net136),
    .D(_0210_),
    .Q(\po_0.regf_0.rf[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3559_ (.CLK(net130),
    .D(_0211_),
    .Q(\po_0.regf_0.rf[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3560_ (.CLK(net136),
    .D(_0212_),
    .Q(\po_0.regf_0.rf[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3561_ (.CLK(net135),
    .D(_0213_),
    .Q(\po_0.regf_0.rf[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3562_ (.CLK(net155),
    .D(_0214_),
    .Q(\po_0.regf_0.rf[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3563_ (.CLK(net154),
    .D(_0215_),
    .Q(\po_0.regf_0.rf[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3564_ (.CLK(net119),
    .D(_0216_),
    .Q(\po_0.regf_0.rf[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3565_ (.CLK(net115),
    .D(_0217_),
    .Q(\po_0.regf_0.rf[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3566_ (.CLK(net158),
    .D(_0218_),
    .Q(\po_0.regf_0.rf[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3567_ (.CLK(net118),
    .D(_0219_),
    .Q(\po_0.regf_0.rf[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3568_ (.CLK(net103),
    .D(_0220_),
    .Q(\po_0.regf_0.rf[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3569_ (.CLK(net110),
    .D(_0221_),
    .Q(\po_0.regf_0.rf[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3570_ (.CLK(net105),
    .D(_0222_),
    .Q(\po_0.regf_0.rf[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3571_ (.CLK(net101),
    .D(_0223_),
    .Q(\po_0.regf_0.rf[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3572_ (.CLK(net181),
    .D(_0224_),
    .Q(\uc_0._21_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3573_ (.CLK(net181),
    .D(_0225_),
    .Q(\uc_0._21_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3574_ (.CLK(net179),
    .D(_0226_),
    .Q(\uc_0._21_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3575_ (.CLK(net174),
    .D(_0227_),
    .Q(\uc_0._21_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3576_ (.CLK(net179),
    .D(_0228_),
    .Q(\uc_0._21_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3577_ (.CLK(net172),
    .D(_0229_),
    .Q(\uc_0._21_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3578_ (.CLK(net174),
    .D(_0230_),
    .Q(\uc_0._21_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3579_ (.CLK(net172),
    .D(_0231_),
    .Q(\uc_0._21_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3580_ (.CLK(net178),
    .D(_0232_),
    .Q(\uc_0._21_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3581_ (.CLK(net167),
    .D(_0233_),
    .Q(\uc_0._21_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3582_ (.CLK(net171),
    .D(_0234_),
    .Q(\uc_0._21_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3583_ (.CLK(net171),
    .D(_0235_),
    .Q(\uc_0._21_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3584_ (.CLK(net171),
    .D(_0236_),
    .Q(\uc_0._21_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3585_ (.CLK(net184),
    .D(_0237_),
    .Q(\uc_0._21_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3586_ (.CLK(net171),
    .D(_0238_),
    .Q(\uc_0._21_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3587_ (.CLK(net179),
    .D(_0239_),
    .Q(\uc_0._21_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3588_ (.CLK(net181),
    .D(_0240_),
    .Q(\uc_0._00_ ));
 sky130_fd_sc_hd__dfxtp_1 _3589_ (.CLK(net165),
    .D(_0012_),
    .Q(_0004_));
 sky130_fd_sc_hd__dfxtp_1 _3590_ (.CLK(net159),
    .D(_0013_),
    .Q(_0005_));
 sky130_fd_sc_hd__dfxtp_2 _3591_ (.CLK(net165),
    .D(_0014_),
    .Q(_0006_));
 sky130_fd_sc_hd__dfxtp_1 _3592_ (.CLK(net167),
    .D(_0015_),
    .Q(_0007_));
 sky130_fd_sc_hd__dfxtp_1 _3593_ (.CLK(net143),
    .D(_0241_),
    .Q(\po_0.regf_0.rf[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3594_ (.CLK(net131),
    .D(_0242_),
    .Q(\po_0.regf_0.rf[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3595_ (.CLK(net148),
    .D(_0243_),
    .Q(\po_0.regf_0.rf[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3596_ (.CLK(net144),
    .D(_0244_),
    .Q(\po_0.regf_0.rf[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3597_ (.CLK(net138),
    .D(_0245_),
    .Q(\po_0.regf_0.rf[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3598_ (.CLK(net144),
    .D(_0246_),
    .Q(\po_0.regf_0.rf[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3599_ (.CLK(net159),
    .D(_0247_),
    .Q(\po_0.regf_0.rf[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3600_ (.CLK(net156),
    .D(_0248_),
    .Q(\po_0.regf_0.rf[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3601_ (.CLK(net119),
    .D(_0249_),
    .Q(\po_0.regf_0.rf[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3602_ (.CLK(net117),
    .D(_0250_),
    .Q(\po_0.regf_0.rf[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3603_ (.CLK(net158),
    .D(_0251_),
    .Q(\po_0.regf_0.rf[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3604_ (.CLK(net118),
    .D(_0252_),
    .Q(\po_0.regf_0.rf[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3605_ (.CLK(net103),
    .D(_0253_),
    .Q(\po_0.regf_0.rf[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3606_ (.CLK(net113),
    .D(_0254_),
    .Q(\po_0.regf_0.rf[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3607_ (.CLK(net116),
    .D(_0255_),
    .Q(\po_0.regf_0.rf[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3608_ (.CLK(net108),
    .D(_0256_),
    .Q(\po_0.regf_0.rf[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3609_ (.CLK(net132),
    .D(_0257_),
    .Q(\po_0.regf_0.rf[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3610_ (.CLK(net137),
    .D(_0258_),
    .Q(\po_0.regf_0.rf[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3611_ (.CLK(net139),
    .D(_0259_),
    .Q(\po_0.regf_0.rf[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3612_ (.CLK(net131),
    .D(_0260_),
    .Q(\po_0.regf_0.rf[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3613_ (.CLK(net139),
    .D(_0261_),
    .Q(\po_0.regf_0.rf[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3614_ (.CLK(net137),
    .D(_0262_),
    .Q(\po_0.regf_0.rf[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3615_ (.CLK(net157),
    .D(_0263_),
    .Q(\po_0.regf_0.rf[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3616_ (.CLK(net156),
    .D(_0264_),
    .Q(\po_0.regf_0.rf[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3617_ (.CLK(net121),
    .D(_0265_),
    .Q(\po_0.regf_0.rf[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3618_ (.CLK(net116),
    .D(_0266_),
    .Q(\po_0.regf_0.rf[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3619_ (.CLK(net158),
    .D(_0267_),
    .Q(\po_0.regf_0.rf[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3620_ (.CLK(net116),
    .D(_0268_),
    .Q(\po_0.regf_0.rf[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3621_ (.CLK(net103),
    .D(_0269_),
    .Q(\po_0.regf_0.rf[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3622_ (.CLK(net128),
    .D(_0270_),
    .Q(\po_0.regf_0.rf[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3623_ (.CLK(net104),
    .D(_0271_),
    .Q(\po_0.regf_0.rf[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3624_ (.CLK(net108),
    .D(_0272_),
    .Q(\po_0.regf_0.rf[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3625_ (.CLK(net143),
    .D(_0273_),
    .Q(\po_0.regf_0.rf[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3626_ (.CLK(net131),
    .D(_0274_),
    .Q(\po_0.regf_0.rf[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3627_ (.CLK(net148),
    .D(_0275_),
    .Q(\po_0.regf_0.rf[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3628_ (.CLK(net144),
    .D(_0276_),
    .Q(\po_0.regf_0.rf[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3629_ (.CLK(net137),
    .D(_0277_),
    .Q(\po_0.regf_0.rf[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3630_ (.CLK(net148),
    .D(_0278_),
    .Q(\po_0.regf_0.rf[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3631_ (.CLK(net160),
    .D(_0279_),
    .Q(\po_0.regf_0.rf[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3632_ (.CLK(net154),
    .D(_0280_),
    .Q(\po_0.regf_0.rf[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3633_ (.CLK(net119),
    .D(_0281_),
    .Q(\po_0.regf_0.rf[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3634_ (.CLK(net117),
    .D(_0282_),
    .Q(\po_0.regf_0.rf[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3635_ (.CLK(net161),
    .D(_0283_),
    .Q(\po_0.regf_0.rf[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3636_ (.CLK(net118),
    .D(_0284_),
    .Q(\po_0.regf_0.rf[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3637_ (.CLK(net103),
    .D(_0285_),
    .Q(\po_0.regf_0.rf[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3638_ (.CLK(net113),
    .D(_0286_),
    .Q(\po_0.regf_0.rf[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3639_ (.CLK(net104),
    .D(_0287_),
    .Q(\po_0.regf_0.rf[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3640_ (.CLK(net101),
    .D(_0288_),
    .Q(\po_0.regf_0.rf[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3641_ (.CLK(net145),
    .D(_0289_),
    .Q(\po_0.regf_0.rf[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3642_ (.CLK(net151),
    .D(_0290_),
    .Q(\po_0.regf_0.rf[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3643_ (.CLK(net152),
    .D(_0291_),
    .Q(\po_0.regf_0.rf[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3644_ (.CLK(net146),
    .D(_0292_),
    .Q(\po_0.regf_0.rf[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3645_ (.CLK(net152),
    .D(_0293_),
    .Q(\po_0.regf_0.rf[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3646_ (.CLK(net151),
    .D(_0294_),
    .Q(\po_0.regf_0.rf[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3647_ (.CLK(net163),
    .D(_0295_),
    .Q(\po_0.regf_0.rf[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3648_ (.CLK(net163),
    .D(_0296_),
    .Q(\po_0.regf_0.rf[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3649_ (.CLK(net178),
    .D(_0297_),
    .Q(\po_0.regf_0.rf[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3650_ (.CLK(net123),
    .D(_0298_),
    .Q(\po_0.regf_0.rf[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3651_ (.CLK(net166),
    .D(_0299_),
    .Q(\po_0.regf_0.rf[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3652_ (.CLK(net123),
    .D(_0300_),
    .Q(\po_0.regf_0.rf[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3653_ (.CLK(net113),
    .D(_0301_),
    .Q(\po_0.regf_0.rf[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3654_ (.CLK(net128),
    .D(_0302_),
    .Q(\po_0.regf_0.rf[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3655_ (.CLK(net113),
    .D(_0303_),
    .Q(\po_0.regf_0.rf[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3656_ (.CLK(net110),
    .D(_0304_),
    .Q(\po_0.regf_0.rf[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _3657_ (.CLK(net179),
    .D(_0305_),
    .Q(\po_0.alu_0.s1 ));
 sky130_fd_sc_hd__dfxtp_1 _3658_ (.CLK(net180),
    .D(_0306_),
    .Q(\po_0.alu_0.s0 ));
 sky130_fd_sc_hd__dfxtp_1 _3659_ (.CLK(net178),
    .D(_0307_),
    .Q(\po_0.regf_0.rq_rd ));
 sky130_fd_sc_hd__dfxtp_1 _3660_ (.CLK(net189),
    .D(_0308_),
    .Q(\po_0.regf_0.rp_rd ));
 sky130_fd_sc_hd__dfxtp_1 _3661_ (.CLK(net145),
    .D(_0309_),
    .Q(\po_0.regf_0.w_wr ));
 sky130_fd_sc_hd__dfxtp_1 _3662_ (.CLK(net174),
    .D(_0310_),
    .Q(\po_0.regf_0.rq_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3663_ (.CLK(net172),
    .D(_0311_),
    .Q(\po_0.regf_0.rq_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3664_ (.CLK(net160),
    .D(_0312_),
    .Q(\po_0.regf_0.rq_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3665_ (.CLK(net165),
    .D(_0313_),
    .Q(\po_0.regf_0.rq_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3666_ (.CLK(net179),
    .D(_0314_),
    .Q(\po_0.regf_0.rp_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3667_ (.CLK(net167),
    .D(_0315_),
    .Q(\po_0.regf_0.rp_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3668_ (.CLK(net174),
    .D(_0316_),
    .Q(\po_0.regf_0.rp_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3669_ (.CLK(net175),
    .D(_0317_),
    .Q(\po_0.regf_0.rp_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3670_ (.CLK(net178),
    .D(_0318_),
    .Q(\po_0.regf_0.w_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3671_ (.CLK(net178),
    .D(_0319_),
    .Q(\po_0.regf_0.w_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3672_ (.CLK(net123),
    .D(_0320_),
    .Q(\po_0.regf_0.w_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3673_ (.CLK(net125),
    .D(_0321_),
    .Q(\po_0.regf_0.w_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3674_ (.CLK(net180),
    .D(_0322_),
    .Q(\po_0.muxf_0.rf_w_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3675_ (.CLK(net187),
    .D(_0323_),
    .Q(\po_0.muxf_0.rf_w_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3676_ (.CLK(net187),
    .D(_0324_),
    .Q(\po_0.muxf_0.rf_w_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3677_ (.CLK(net180),
    .D(_0325_),
    .Q(\po_0.muxf_0.rf_w_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3678_ (.CLK(net187),
    .D(_0326_),
    .Q(\po_0.muxf_0.rf_w_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3679_ (.CLK(net180),
    .D(_0327_),
    .Q(\po_0.muxf_0.rf_w_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3680_ (.CLK(net179),
    .D(_0328_),
    .Q(\po_0.muxf_0.rf_w_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3681_ (.CLK(net187),
    .D(_0329_),
    .Q(\po_0.muxf_0.rf_w_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3682_ (.CLK(net187),
    .D(_0330_),
    .Q(\po_0.muxf_0.s0 ));
 sky130_fd_sc_hd__dfxtp_1 _3683_ (.CLK(net188),
    .D(_0331_),
    .Q(\po_0.muxf_0.s1 ));
 sky130_fd_sc_hd__dfxtp_1 _3684_ (.CLK(net184),
    .D(_0332_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_2 _3685_ (.CLK(net184),
    .D(_0333_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_2 _3686_ (.CLK(net175),
    .D(_0334_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _3687_ (.CLK(net182),
    .D(_0335_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _3688_ (.CLK(net175),
    .D(_0336_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _3689_ (.CLK(net180),
    .D(_0337_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _3690_ (.CLK(net187),
    .D(_0338_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _3691_ (.CLK(net174),
    .D(_0339_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _3692_ (.CLK(net160),
    .D(_0340_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _3693_ (.CLK(net160),
    .D(_0341_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _3694_ (.CLK(net184),
    .D(_0342_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _3695_ (.CLK(net185),
    .D(_0343_),
    .Q(\uc_0._03_ ));
 sky130_fd_sc_hd__dfxtp_1 _3696_ (.CLK(net183),
    .D(_0344_),
    .Q(\uc_0._02_ ));
 sky130_fd_sc_hd__dfxtp_1 _3697_ (.CLK(net183),
    .D(_0345_),
    .Q(\uc_0._01_ ));
 sky130_fd_sc_hd__dfxtp_1 _3698_ (.CLK(net184),
    .D(\uc_0.bc_0._70_[0] ),
    .Q(\uc_0.bc_0._05_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3699_ (.CLK(net184),
    .D(\uc_0.bc_0._70_[1] ),
    .Q(\uc_0.bc_0._05_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3700_ (.CLK(net182),
    .D(\uc_0.bc_0._70_[2] ),
    .Q(\uc_0.bc_0._05_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3701_ (.CLK(net182),
    .D(\uc_0.bc_0._70_[3] ),
    .Q(\uc_0.bc_0._05_[3] ));
 sky130_fd_sc_hd__clkbuf_1 _3702_ (.A(net173),
    .X(net78));
 sky130_fd_sc_hd__ebufn_1 _3703_ (.A(\po_0.alu_0._10_[0] ),
    .TE_B(_1624_),
    .Z(\po_0.alu_0._11_[0] ));
 sky130_fd_sc_hd__ebufn_1 _3704_ (.A(\po_0.alu_0._10_[1] ),
    .TE_B(_1625_),
    .Z(\po_0.alu_0._11_[1] ));
 sky130_fd_sc_hd__ebufn_1 _3705_ (.A(\po_0.alu_0._10_[2] ),
    .TE_B(_1626_),
    .Z(\po_0.alu_0._11_[2] ));
 sky130_fd_sc_hd__ebufn_1 _3706_ (.A(\po_0.alu_0._10_[3] ),
    .TE_B(_1627_),
    .Z(\po_0.alu_0._11_[3] ));
 sky130_fd_sc_hd__ebufn_1 _3707_ (.A(\po_0.alu_0._10_[4] ),
    .TE_B(_1628_),
    .Z(\po_0.alu_0._11_[4] ));
 sky130_fd_sc_hd__ebufn_1 _3708_ (.A(\po_0.alu_0._10_[5] ),
    .TE_B(_1629_),
    .Z(\po_0.alu_0._11_[5] ));
 sky130_fd_sc_hd__ebufn_1 _3709_ (.A(\po_0.alu_0._10_[6] ),
    .TE_B(_1630_),
    .Z(\po_0.alu_0._11_[6] ));
 sky130_fd_sc_hd__ebufn_1 _3710_ (.A(\po_0.alu_0._10_[7] ),
    .TE_B(_1631_),
    .Z(\po_0.alu_0._11_[7] ));
 sky130_fd_sc_hd__ebufn_1 _3711_ (.A(\po_0.alu_0._10_[8] ),
    .TE_B(_1632_),
    .Z(\po_0.alu_0._11_[8] ));
 sky130_fd_sc_hd__ebufn_1 _3712_ (.A(\po_0.alu_0._10_[9] ),
    .TE_B(_1633_),
    .Z(\po_0.alu_0._11_[9] ));
 sky130_fd_sc_hd__ebufn_1 _3713_ (.A(\po_0.alu_0._10_[10] ),
    .TE_B(_1634_),
    .Z(\po_0.alu_0._11_[10] ));
 sky130_fd_sc_hd__ebufn_1 _3714_ (.A(\po_0.alu_0._10_[11] ),
    .TE_B(_1635_),
    .Z(\po_0.alu_0._11_[11] ));
 sky130_fd_sc_hd__ebufn_1 _3715_ (.A(\po_0.alu_0._10_[12] ),
    .TE_B(_1636_),
    .Z(\po_0.alu_0._11_[12] ));
 sky130_fd_sc_hd__ebufn_1 _3716_ (.A(\po_0.alu_0._10_[13] ),
    .TE_B(_1637_),
    .Z(\po_0.alu_0._11_[13] ));
 sky130_fd_sc_hd__ebufn_1 _3717_ (.A(\po_0.alu_0._10_[14] ),
    .TE_B(_1638_),
    .Z(\po_0.alu_0._11_[14] ));
 sky130_fd_sc_hd__ebufn_1 _3718_ (.A(\po_0.alu_0._10_[15] ),
    .TE_B(_1639_),
    .Z(\po_0.alu_0._11_[15] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout100 (.A(net102),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 fanout101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 fanout102 (.A(net106),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 fanout103 (.A(net106),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 fanout104 (.A(net106),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout106 (.A(net126),
    .X(net106));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout107 (.A(net111),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 fanout108 (.A(net111),
    .X(net108));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 fanout111 (.A(net114),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 fanout112 (.A(net114),
    .X(net112));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 fanout114 (.A(net126),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 fanout115 (.A(net117),
    .X(net115));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout117 (.A(net125),
    .X(net117));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout118 (.A(net121),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 fanout119 (.A(net121),
    .X(net119));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout121 (.A(net125),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout126 (.A(net191),
    .X(net126));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout127 (.A(net130),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 fanout128 (.A(net130),
    .X(net128));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 fanout130 (.A(net133),
    .X(net130));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout133 (.A(net142),
    .X(net133));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout134 (.A(net136),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 fanout136 (.A(net142),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 fanout137 (.A(net141),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 fanout138 (.A(net141),
    .X(net138));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout139 (.A(net141),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 fanout140 (.A(net141),
    .X(net140));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 fanout142 (.A(net153),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 fanout143 (.A(net147),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 fanout144 (.A(net147),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 fanout145 (.A(net147),
    .X(net145));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 fanout147 (.A(net153),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 fanout148 (.A(net152),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 fanout149 (.A(net152),
    .X(net149));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 fanout151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout153 (.A(net191),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 fanout154 (.A(net157),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 fanout155 (.A(net157),
    .X(net155));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout157 (.A(net170),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 fanout158 (.A(net161),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 fanout159 (.A(net161),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout161 (.A(net170),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 fanout162 (.A(net169),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 fanout163 (.A(net169),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 fanout164 (.A(net168),
    .X(net164));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout165 (.A(net168),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 fanout166 (.A(net168),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout170 (.A(net190),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 fanout171 (.A(net173),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 fanout173 (.A(net177),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 fanout174 (.A(net176),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout177 (.A(net190),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 fanout178 (.A(net189),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 fanout179 (.A(net186),
    .X(net179));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout180 (.A(net186),
    .X(net180));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout181 (.A(net183),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout183 (.A(net185),
    .X(net183));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 fanout186 (.A(net188),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 fanout191 (.A(net33),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 fanout83 (.A(net39),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 fanout84 (.A(net38),
    .X(net84));
 sky130_fd_sc_hd__buf_2 fanout85 (.A(net37),
    .X(net85));
 sky130_fd_sc_hd__buf_2 fanout86 (.A(net49),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 fanout87 (.A(net42),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 fanout88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 fanout89 (.A(\po_0.regf_0.rp_rd ),
    .X(net89));
 sky130_fd_sc_hd__buf_2 fanout90 (.A(\po_0.regf_0.rp_rd ),
    .X(net90));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout91 (.A(net93),
    .X(net91));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 fanout93 (.A(\po_0.regf_0.rq_rd ),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(net66),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 fanout95 (.A(net65),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(net64),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 fanout97 (.A(net63),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 fanout98 (.A(net76),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 fanout99 (.A(net68),
    .X(net99));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(D_R_data[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(D_R_data[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(D_R_data[4]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(D_R_data[5]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(D_R_data[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(D_R_data[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(D_R_data[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(D_R_data[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(I_data[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(I_data[10]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(I_data[11]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(D_R_data[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(I_data[12]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(I_data[13]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(I_data[14]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(I_data[15]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(I_data[1]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(I_data[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(I_data[3]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(I_data[4]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(I_data[5]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(I_data[6]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(D_R_data[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(I_data[7]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(I_data[8]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(I_data[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(clock),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(reset),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(D_R_data[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(D_R_data[13]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(D_R_data[14]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(D_R_data[15]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(D_R_data[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(D_R_data[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(D_W_data[0]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(D_W_data[10]));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net37),
    .X(D_W_data[11]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net84),
    .X(D_W_data[12]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(D_W_data[13]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(D_W_data[14]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(D_W_data[15]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(D_W_data[1]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(D_W_data[2]));
 sky130_fd_sc_hd__clkbuf_4 output44 (.A(net44),
    .X(D_W_data[3]));
 sky130_fd_sc_hd__clkbuf_4 output45 (.A(net45),
    .X(D_W_data[4]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(D_W_data[5]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(D_W_data[6]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(D_W_data[7]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net86),
    .X(D_W_data[8]));
 sky130_fd_sc_hd__clkbuf_4 output50 (.A(net50),
    .X(D_W_data[9]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(D_addr[0]));
 sky130_fd_sc_hd__clkbuf_4 output52 (.A(net52),
    .X(D_addr[1]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(D_addr[2]));
 sky130_fd_sc_hd__clkbuf_4 output54 (.A(net54),
    .X(D_addr[3]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(D_addr[4]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(D_addr[5]));
 sky130_fd_sc_hd__clkbuf_4 output57 (.A(net57),
    .X(D_addr[6]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(D_addr[7]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(D_rd));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(D_wr));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(I_addr[0]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(I_addr[10]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net97),
    .X(I_addr[11]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net96),
    .X(I_addr[12]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net95),
    .X(I_addr[13]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net94),
    .X(I_addr[14]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(I_addr[15]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net99),
    .X(I_addr[1]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(I_addr[2]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(I_addr[3]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(I_addr[4]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(I_addr[5]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(I_addr[6]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(I_addr[7]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(I_addr[8]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(I_addr[9]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(I_rd));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net78),
    .X(led_clock));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(leds[0]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(leds[1]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(leds[2]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(leds[3]));
endmodule

